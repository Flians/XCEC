//
// Conformal-LEC Version 20.10-d213 (02-Sep-2020)
//
module top(RIbe28de0_41,RIbe27b98_2,RIbe29920_65,RIbe28c78_38,RIbe28318_18,RIbe29038_46,RIbe29650_59,RIbe296c8_60,RIbe290b0_47,
        RIbe29a88_68,RIbe27d78_6,RIbe286d8_26,RIbe27ee0_9,RIbe28e58_42,RIbe27c10_3,RIbe284f8_22,RIbe28750_27,RIbe28c00_37,RIbe27d00_5,
        RIbe28840_29,RIbe28570_23,RIbe28fc0_45,RIbe29380_53,RIbe28048_12,RIbe29308_52,RIbe280c0_13,RIbe281b0_15,RIbe28228_16,RIbe29560_57,
        RIbe28930_31,RIbe29830_63,RIbe29470_55,RIbe294e8_56,RIbe288b8_30,RIbe28a98_34,RIbe28138_14,RIbe282a0_17,RIbe289a8_32,RIbe28a20_33,
        RIbe293f8_54,RIbe29740_61,RIbe297b8_62,RIbe28b88_36,RIbe29290_51,RIbe295d8_58,RIbe29a10_67,RIbe29b00_69,RIbe298a8_64,RIbe29998_66,
        RIbe27e68_8,RIbe27f58_10,RIbe27fd0_11,RIbe28480_21,RIbe287c8_28,RIbe285e8_24,RIbe28b10_35,RIbe28390_19,RIbe27c88_4,RIbe27df0_7,
        RIbe27b20_1,RIbe28660_25,RIbe28408_20,RIbe28cf0_39,RIbe28d68_40,RIbe28ed0_43,RIbe28f48_44,RIbe29128_48,RIbe291a0_49,RIbe29218_50,
        RIbe29bf0_71,RIbe29c68_72,RIbe29b78_70,RIbe29ce0_73,RIbe29d58_74,RIbe29dd0_75,RIbe29e48_76,RIbe29ec0_77,RIbe2a028_80,RIbe29fb0_79,
        RIbe29f38_78,RIbe2b6a8_128,RIbe2aa78_102,RIbe2a2f8_86,RIbe2acd0_107,RIbe2aa00_101,RIbe2a370_87,RIbe2a3e8_88,RIbe2a898_98,RIbe2a910_99,
        RIbe2b5b8_126,RIbe2a820_97,RIbe2a118_82,RIbe2a0a0_81,RIbe2a550_91,RIbe2a988_100,RIbe2b360_121,RIbe2a190_83,RIbe2a5c8_92,RIbe2adc0_109,
        RIbe2a460_89,RIbe2a4d8_90,RIbe2b2e8_120,RIbe2b540_125,RIbe2a280_85,RIbe2a208_84,RIbe2ad48_108,RIbe2b108_116,RIbe2b090_115,RIbe2b4c8_124,
        RIbe2a6b8_94,RIbe2b180_117,RIbe2b270_119,RIbe2afa0_113,RIbe2b018_114,RIbe2af28_112,RIbe2abe0_105,RIbe2ac58_106,RIbe2b1f8_118,RIbe2a640_93,
        RIbe2a730_95,RIbe2a7a8_96,RIbe2aaf0_103,RIbe2b630_127,RIbe2b450_123,RIbe2b3d8_122,RIbe2aeb0_111,RIbe2ae38_110,RIbe2ab68_104,R_81_9fc6f08,
        R_82_9fc5ea0,R_83_90f04e0,R_84_90effa0,R_85_90e8ad0,R_86_90e3e08,R_87_90f1a88,R_88_90e8638,R_89_90f1200,R_8a_90f12a8,R_8b_90f0cc0,
        R_8c_90ef088,R_8d_90f1158,R_8e_90e49d8,R_8f_90e3eb0,R_90_9fc69c8,R_91_90e9c88,R_92_90f0588,R_93_90eacf0,R_94_90ebb60,R_95_90e66b8,
        R_96_9fc6d10,R_97_90ead98,R_98_90e90b8,R_99_90eb038,R_9a_90e9d30,R_9b_90e7bb8,R_9c_9fc7b80,R_9d_90ebd58,R_9e_90e9a90,R_9f_90efb08,
        R_a0_90e6e98,R_a1_90f0780,R_a2_90e2da0,R_a3_90f0240,R_a4_9fc7ad8,R_a5_9fc73a0,R_a6_9fc6680,R_a7_90e4f18,R_a8_90e3388,R_a9_9fc67d0,
        R_aa_90f17e8,R_ab_90e4888,R_ac_90e9010,R_ad_90eee90,R_ae_90e53b0,R_af_90ebc08,R_b0_90e8440,R_b1_90ea900,R_b2_90e9400,R_b3_9fc6bc0,
        R_b4_90e4690,R_b5_90e3778,R_b6_90e9160,R_b7_90e29b0,R_b8_90e2278,R_b9_9fc6a70,R_ba_90ebf50,R_bb_90f0e10,R_bc_9fc7640,R_bd_90f1dd0,
        R_be_90f0630,R_bf_90f0eb8,R_c0_90e34d8,R_c1_90e9f28,R_c2_90f0d68,R_c3_90ea7b0,R_c4_9fc7448,R_c5_90eb428,R_c6_90e81a0,R_c7_90f0a20,
        R_c8_90efda8,R_c9_90e2c50,R_ca_90e88d8,R_cb_9fc6530,R_cc_90f06d8,R_cd_90efa60,R_ce_90e2b00,R_cf_9fc6920,R_d0_90f1f20,R_d1_90e7678,
        R_d2_90efd00,R_d3_90e7e58,R_d4_90e7d08,R_d5_90eaa50,R_d6_90e3040,R_d7_90efe50,R_d8_90f1350,R_d9_9fc71a8,R_da_9fc9cf8,R_db_90ef9b8,
        R_dc_90e4540,R_dd_90f0ac8,R_de_90e30e8,R_df_9fc6290,R_e0_9fc78e0,R_e1_90e5500,R_e2_90e68b0,R_e3_90eede8,R_e4_90e64c0,R_e5_9fc7100,
        R_e6_90e2470,R_e7_90ebea8,R_e8_90e4a80,R_e9_90ef910,R_ea_9fc7c28,R_eb_90eb4d0,R_ec_90f14a0,R_ed_90ef5c8,R_ee_90e4498,R_ef_90e4000,
        R_f0_90f0048,R_f1_90ea3c0,R_f2_90f1e78,R_f3_90f00f0);
input RIbe28de0_41,RIbe27b98_2,RIbe29920_65,RIbe28c78_38,RIbe28318_18,RIbe29038_46,RIbe29650_59,RIbe296c8_60,RIbe290b0_47,
        RIbe29a88_68,RIbe27d78_6,RIbe286d8_26,RIbe27ee0_9,RIbe28e58_42,RIbe27c10_3,RIbe284f8_22,RIbe28750_27,RIbe28c00_37,RIbe27d00_5,
        RIbe28840_29,RIbe28570_23,RIbe28fc0_45,RIbe29380_53,RIbe28048_12,RIbe29308_52,RIbe280c0_13,RIbe281b0_15,RIbe28228_16,RIbe29560_57,
        RIbe28930_31,RIbe29830_63,RIbe29470_55,RIbe294e8_56,RIbe288b8_30,RIbe28a98_34,RIbe28138_14,RIbe282a0_17,RIbe289a8_32,RIbe28a20_33,
        RIbe293f8_54,RIbe29740_61,RIbe297b8_62,RIbe28b88_36,RIbe29290_51,RIbe295d8_58,RIbe29a10_67,RIbe29b00_69,RIbe298a8_64,RIbe29998_66,
        RIbe27e68_8,RIbe27f58_10,RIbe27fd0_11,RIbe28480_21,RIbe287c8_28,RIbe285e8_24,RIbe28b10_35,RIbe28390_19,RIbe27c88_4,RIbe27df0_7,
        RIbe27b20_1,RIbe28660_25,RIbe28408_20,RIbe28cf0_39,RIbe28d68_40,RIbe28ed0_43,RIbe28f48_44,RIbe29128_48,RIbe291a0_49,RIbe29218_50,
        RIbe29bf0_71,RIbe29c68_72,RIbe29b78_70,RIbe29ce0_73,RIbe29d58_74,RIbe29dd0_75,RIbe29e48_76,RIbe29ec0_77,RIbe2a028_80,RIbe29fb0_79,
        RIbe29f38_78,RIbe2b6a8_128,RIbe2aa78_102,RIbe2a2f8_86,RIbe2acd0_107,RIbe2aa00_101,RIbe2a370_87,RIbe2a3e8_88,RIbe2a898_98,RIbe2a910_99,
        RIbe2b5b8_126,RIbe2a820_97,RIbe2a118_82,RIbe2a0a0_81,RIbe2a550_91,RIbe2a988_100,RIbe2b360_121,RIbe2a190_83,RIbe2a5c8_92,RIbe2adc0_109,
        RIbe2a460_89,RIbe2a4d8_90,RIbe2b2e8_120,RIbe2b540_125,RIbe2a280_85,RIbe2a208_84,RIbe2ad48_108,RIbe2b108_116,RIbe2b090_115,RIbe2b4c8_124,
        RIbe2a6b8_94,RIbe2b180_117,RIbe2b270_119,RIbe2afa0_113,RIbe2b018_114,RIbe2af28_112,RIbe2abe0_105,RIbe2ac58_106,RIbe2b1f8_118,RIbe2a640_93,
        RIbe2a730_95,RIbe2a7a8_96,RIbe2aaf0_103,RIbe2b630_127,RIbe2b450_123,RIbe2b3d8_122,RIbe2aeb0_111,RIbe2ae38_110,RIbe2ab68_104;
output R_81_9fc6f08,R_82_9fc5ea0,R_83_90f04e0,R_84_90effa0,R_85_90e8ad0,R_86_90e3e08,R_87_90f1a88,R_88_90e8638,R_89_90f1200,
        R_8a_90f12a8,R_8b_90f0cc0,R_8c_90ef088,R_8d_90f1158,R_8e_90e49d8,R_8f_90e3eb0,R_90_9fc69c8,R_91_90e9c88,R_92_90f0588,R_93_90eacf0,
        R_94_90ebb60,R_95_90e66b8,R_96_9fc6d10,R_97_90ead98,R_98_90e90b8,R_99_90eb038,R_9a_90e9d30,R_9b_90e7bb8,R_9c_9fc7b80,R_9d_90ebd58,
        R_9e_90e9a90,R_9f_90efb08,R_a0_90e6e98,R_a1_90f0780,R_a2_90e2da0,R_a3_90f0240,R_a4_9fc7ad8,R_a5_9fc73a0,R_a6_9fc6680,R_a7_90e4f18,
        R_a8_90e3388,R_a9_9fc67d0,R_aa_90f17e8,R_ab_90e4888,R_ac_90e9010,R_ad_90eee90,R_ae_90e53b0,R_af_90ebc08,R_b0_90e8440,R_b1_90ea900,
        R_b2_90e9400,R_b3_9fc6bc0,R_b4_90e4690,R_b5_90e3778,R_b6_90e9160,R_b7_90e29b0,R_b8_90e2278,R_b9_9fc6a70,R_ba_90ebf50,R_bb_90f0e10,
        R_bc_9fc7640,R_bd_90f1dd0,R_be_90f0630,R_bf_90f0eb8,R_c0_90e34d8,R_c1_90e9f28,R_c2_90f0d68,R_c3_90ea7b0,R_c4_9fc7448,R_c5_90eb428,
        R_c6_90e81a0,R_c7_90f0a20,R_c8_90efda8,R_c9_90e2c50,R_ca_90e88d8,R_cb_9fc6530,R_cc_90f06d8,R_cd_90efa60,R_ce_90e2b00,R_cf_9fc6920,
        R_d0_90f1f20,R_d1_90e7678,R_d2_90efd00,R_d3_90e7e58,R_d4_90e7d08,R_d5_90eaa50,R_d6_90e3040,R_d7_90efe50,R_d8_90f1350,R_d9_9fc71a8,
        R_da_9fc9cf8,R_db_90ef9b8,R_dc_90e4540,R_dd_90f0ac8,R_de_90e30e8,R_df_9fc6290,R_e0_9fc78e0,R_e1_90e5500,R_e2_90e68b0,R_e3_90eede8,
        R_e4_90e64c0,R_e5_9fc7100,R_e6_90e2470,R_e7_90ebea8,R_e8_90e4a80,R_e9_90ef910,R_ea_9fc7c28,R_eb_90eb4d0,R_ec_90f14a0,R_ed_90ef5c8,
        R_ee_90e4498,R_ef_90e4000,R_f0_90f0048,R_f1_90ea3c0,R_f2_90f1e78,R_f3_90f00f0;

wire \244 , \245_N$1 , \246_ZERO , \247_ONE , \248 , \249 , \250 , \251 , \252 ,
         \253 , \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 , \262 ,
         \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 , \272 ,
         \273 , \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 , \282 ,
         \283 , \284 , \285 , \286 , \287 , \288 , \289 , \290 , \291 , \292 ,
         \293 , \294 , \295 , \296 , \297 , \298 , \299 , \300 , \301 , \302 ,
         \303 , \304 , \305 , \306 , \307 , \308 , \309 , \310 , \311 , \312 ,
         \313 , \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321 , \322 ,
         \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331 , \332 ,
         \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 , \342 ,
         \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 , \351 , \352 ,
         \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 , \362 ,
         \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 ,
         \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 ,
         \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 ,
         \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 ,
         \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 ,
         \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 ,
         \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 ,
         \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 ,
         \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 ,
         \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 ,
         \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 ,
         \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 ,
         \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 ,
         \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 ,
         \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 ,
         \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 ,
         \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 ,
         \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 ,
         \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 ,
         \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 ,
         \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 ,
         \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 ,
         \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 ,
         \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 ,
         \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 ,
         \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 ,
         \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 ,
         \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 ,
         \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 ,
         \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 ,
         \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 ,
         \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 ,
         \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 ,
         \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 ,
         \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 ,
         \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 ,
         \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 ,
         \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 ,
         \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 ,
         \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 ,
         \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 ,
         \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 ,
         \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 ,
         \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 ,
         \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 ,
         \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 ,
         \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 ,
         \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 ,
         \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 ,
         \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 ,
         \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 ,
         \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 ,
         \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 ,
         \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 ,
         \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 ,
         \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 ,
         \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 ,
         \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 ,
         \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 ,
         \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 ,
         \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 ,
         \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 ,
         \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 ,
         \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 ,
         \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 ,
         \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 ,
         \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 ,
         \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 ,
         \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 ,
         \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 ,
         \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 ,
         \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 ,
         \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 ,
         \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 ,
         \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 ,
         \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 ,
         \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 ,
         \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
         \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 ,
         \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 ,
         \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 ,
         \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 ,
         \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 ,
         \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 ,
         \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 ,
         \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 ,
         \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 ,
         \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 ,
         \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 ,
         \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 ,
         \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 ,
         \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 ,
         \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 ,
         \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 ,
         \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 ,
         \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 ,
         \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
         \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 ,
         \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 ,
         \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 ,
         \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 ,
         \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 ,
         \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 ,
         \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 ,
         \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 ,
         \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 ,
         \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 ,
         \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 ,
         \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 ,
         \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 ,
         \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 ,
         \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 ,
         \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 ,
         \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 ,
         \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 ,
         \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 ,
         \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 ,
         \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 ,
         \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 ,
         \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 ,
         \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 ,
         \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 ,
         \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 ,
         \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 ,
         \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 ,
         \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 ,
         \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 ,
         \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 ,
         \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 ,
         \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 ,
         \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 ,
         \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 ,
         \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 ,
         \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 ,
         \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 ,
         \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 ,
         \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 ,
         \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 ,
         \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 ,
         \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 ,
         \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 ,
         \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 ,
         \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 ,
         \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 ,
         \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 ,
         \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 ,
         \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 ,
         \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 ,
         \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 ,
         \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 ,
         \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 ,
         \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 ,
         \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 ,
         \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 ,
         \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 ,
         \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 ,
         \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 ,
         \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 ,
         \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 ,
         \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 ,
         \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 ,
         \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 ,
         \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 ,
         \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 ,
         \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 ,
         \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 ,
         \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 ,
         \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 ,
         \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 ,
         \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 ,
         \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 ,
         \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 ,
         \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 ,
         \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 ,
         \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 ,
         \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 ,
         \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 ,
         \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 ,
         \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 ,
         \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 ,
         \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 ,
         \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 ,
         \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 ,
         \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 ,
         \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 ,
         \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 ,
         \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 ,
         \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 ,
         \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 ,
         \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 ,
         \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 ,
         \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 ,
         \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 ,
         \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 ,
         \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 ,
         \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 ,
         \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 ,
         \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 ,
         \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 ,
         \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 ,
         \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 ,
         \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 ,
         \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 ,
         \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 ,
         \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 ,
         \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 ,
         \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 ,
         \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 ,
         \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 ,
         \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 ,
         \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 ,
         \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 ,
         \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 ,
         \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 ,
         \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 ,
         \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 ,
         \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 ,
         \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 ,
         \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 ,
         \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 ,
         \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 ,
         \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 ,
         \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 ,
         \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 ,
         \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 ,
         \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 ,
         \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 ,
         \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 ,
         \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 ,
         \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 ,
         \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 ,
         \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 ,
         \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 ,
         \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 ,
         \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 ,
         \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 ,
         \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 ,
         \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 ,
         \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 ,
         \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 ,
         \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 ,
         \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 ,
         \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 ,
         \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 ,
         \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 ,
         \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 ,
         \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 ,
         \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 ,
         \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 ,
         \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 ,
         \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 ,
         \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 ,
         \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 ,
         \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 ,
         \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 ,
         \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 ,
         \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 ,
         \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 ,
         \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 ,
         \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 ,
         \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 ,
         \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 ,
         \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 ,
         \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 ,
         \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 ,
         \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 ,
         \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 ,
         \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 ,
         \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 ,
         \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 ,
         \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 ,
         \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 ,
         \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 ,
         \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 ,
         \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 ,
         \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 ,
         \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 ,
         \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 ,
         \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 ,
         \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 ,
         \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 ,
         \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 ,
         \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 ,
         \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 ,
         \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 ,
         \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 ,
         \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 ,
         \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 ,
         \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 ,
         \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 ,
         \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 ,
         \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 ,
         \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 ,
         \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 ,
         \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 ,
         \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 ,
         \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 ,
         \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 ,
         \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 ,
         \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 ,
         \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 ,
         \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 ,
         \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 ,
         \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 ,
         \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 ,
         \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 ,
         \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 ,
         \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 ,
         \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 ,
         \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 ,
         \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 ,
         \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 ,
         \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 ,
         \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 ,
         \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 ,
         \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 ,
         \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 ,
         \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 ,
         \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 ,
         \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 ,
         \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 ,
         \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 ,
         \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 ,
         \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 ,
         \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 ,
         \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 ,
         \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 ,
         \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 ,
         \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 ,
         \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 ,
         \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 ,
         \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 ,
         \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 ,
         \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 ,
         \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 ,
         \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 ,
         \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 ,
         \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 ,
         \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 ,
         \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 ,
         \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 ,
         \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 ,
         \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 ,
         \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 ,
         \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 ,
         \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 ,
         \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 ,
         \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 ,
         \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 ,
         \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 ,
         \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 ,
         \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 ,
         \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 ,
         \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 ,
         \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 ,
         \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 ,
         \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 ,
         \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 ,
         \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 ,
         \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 ,
         \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 ,
         \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 ,
         \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 ,
         \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 ,
         \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 ,
         \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 ,
         \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 ,
         \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 ,
         \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 ,
         \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 ,
         \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 ,
         \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 ,
         \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 ,
         \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 ,
         \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 ,
         \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 ,
         \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 ,
         \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 ,
         \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 ,
         \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 ,
         \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 ,
         \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 ,
         \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 ,
         \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 ,
         \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 ,
         \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 ,
         \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 ,
         \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 ,
         \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 ,
         \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 ,
         \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 ,
         \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 ,
         \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 ,
         \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 ,
         \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 ,
         \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 ,
         \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 ,
         \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 ,
         \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 ,
         \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 ,
         \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 ,
         \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 ,
         \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 ,
         \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 ,
         \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 ,
         \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 ,
         \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 ,
         \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 ,
         \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 ,
         \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 ,
         \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 ,
         \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 ,
         \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 ,
         \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 ,
         \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 ,
         \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 ,
         \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 ,
         \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 ,
         \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 ,
         \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 ,
         \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 ,
         \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 ,
         \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 ,
         \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 ,
         \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 ,
         \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 ,
         \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 ,
         \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 ,
         \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 ,
         \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 ,
         \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 ,
         \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 ,
         \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 ,
         \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 ,
         \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 ,
         \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 ,
         \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 ,
         \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 ,
         \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 ,
         \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 ,
         \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 ,
         \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 ,
         \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 ,
         \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 ,
         \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 ,
         \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 ,
         \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 ,
         \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 ,
         \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 ,
         \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 ,
         \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 ,
         \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 ,
         \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 ,
         \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 ,
         \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 ,
         \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 ,
         \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 ,
         \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 ,
         \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 ,
         \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 ,
         \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 ,
         \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 ,
         \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 ,
         \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 ,
         \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 ,
         \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 ,
         \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 ,
         \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 ,
         \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 ,
         \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 ,
         \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 ,
         \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 ,
         \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 ,
         \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 ,
         \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 ,
         \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 ,
         \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 ,
         \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 ,
         \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 ,
         \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 ,
         \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 ,
         \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 ,
         \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 ,
         \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 ,
         \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 ,
         \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 ,
         \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 ,
         \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 ,
         \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 ,
         \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 ,
         \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 ,
         \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 ,
         \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 ,
         \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 ,
         \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 ,
         \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 ,
         \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 ,
         \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 ,
         \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 ,
         \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 ,
         \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 ,
         \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 ,
         \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 ,
         \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 ,
         \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 ,
         \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 ,
         \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 ,
         \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 ,
         \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 ,
         \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 ,
         \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 ,
         \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 ,
         \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 ,
         \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 ,
         \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 ,
         \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 ,
         \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 ,
         \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 ,
         \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 ,
         \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 ,
         \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 ,
         \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 ,
         \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 ,
         \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 ,
         \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 ,
         \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 ,
         \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 ,
         \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 ,
         \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 ,
         \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 ,
         \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 ,
         \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 ,
         \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 ,
         \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 ,
         \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 ,
         \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 ,
         \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 ,
         \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 ,
         \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 ,
         \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 ,
         \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 ,
         \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 ,
         \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 ,
         \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 ,
         \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 ,
         \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 ,
         \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 ,
         \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 ,
         \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 ,
         \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 ,
         \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 ,
         \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 ,
         \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 ,
         \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 ,
         \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 ,
         \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 ,
         \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 ,
         \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 ,
         \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 ,
         \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 ,
         \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 ,
         \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 ,
         \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 ,
         \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 ,
         \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 ,
         \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 ,
         \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 ,
         \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 ,
         \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 ,
         \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 ,
         \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 ,
         \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 ,
         \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 ,
         \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 ,
         \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 ,
         \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 ,
         \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 ,
         \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 ,
         \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 ,
         \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 ,
         \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 ,
         \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 ,
         \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 ,
         \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 ,
         \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 ,
         \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 ,
         \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 ,
         \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 ,
         \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 ,
         \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 ,
         \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 ,
         \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 ,
         \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 ,
         \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 ,
         \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 ,
         \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 ,
         \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 ,
         \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 ,
         \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 ,
         \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 ,
         \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 ,
         \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 ,
         \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 ,
         \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 ,
         \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 ,
         \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 ,
         \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 ,
         \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 ,
         \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 ,
         \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 ,
         \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 ,
         \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 ,
         \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 ,
         \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 ,
         \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 ,
         \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 ,
         \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 ,
         \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 ,
         \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 ,
         \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 ,
         \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 ,
         \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 ,
         \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 ,
         \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 ,
         \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 ,
         \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 ,
         \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 ,
         \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 ,
         \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 ,
         \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 ,
         \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 ,
         \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 ,
         \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 ,
         \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 ,
         \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 ,
         \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 ,
         \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 ,
         \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 ,
         \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 ,
         \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 ,
         \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 ,
         \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 ,
         \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 ,
         \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 ,
         \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 ,
         \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 ,
         \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 ,
         \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 ,
         \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 ,
         \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 ,
         \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 ,
         \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 ,
         \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 ,
         \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 ,
         \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 ,
         \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 ,
         \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 ,
         \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 ,
         \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 ,
         \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 ,
         \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 ,
         \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 ,
         \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 ,
         \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 ,
         \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 ,
         \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 ,
         \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 ,
         \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 ,
         \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 ,
         \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 ,
         \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 ,
         \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 ,
         \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 ,
         \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 ,
         \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 ,
         \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 ,
         \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 ,
         \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 ,
         \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 ,
         \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 ,
         \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 ,
         \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 ,
         \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 ,
         \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 ,
         \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 ,
         \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 ,
         \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 ,
         \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 ,
         \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 ,
         \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 ,
         \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 ,
         \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 ,
         \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 ,
         \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 ,
         \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 ,
         \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 ,
         \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 ,
         \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 ,
         \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 ,
         \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 ,
         \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 ,
         \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 ,
         \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 ,
         \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 ,
         \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 ,
         \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 ,
         \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 ,
         \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 ,
         \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 ,
         \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 ,
         \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 ,
         \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 ,
         \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 ,
         \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 ,
         \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 ,
         \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 ,
         \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 ,
         \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 ,
         \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 ,
         \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 ,
         \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 ,
         \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 ,
         \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 ,
         \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 ,
         \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 ,
         \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 ,
         \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 ,
         \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 ,
         \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 ,
         \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 ,
         \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 ,
         \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 ,
         \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 ,
         \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 ,
         \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 ,
         \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 ,
         \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 ,
         \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 ,
         \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 ,
         \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 ,
         \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 ,
         \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 ,
         \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 ,
         \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 ,
         \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 ,
         \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 ,
         \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 ,
         \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 ,
         \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 ,
         \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 ,
         \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 ,
         \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 ,
         \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 ,
         \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 ,
         \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 ,
         \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 ,
         \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 ,
         \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 ,
         \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 ,
         \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 ,
         \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 ,
         \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 ,
         \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 ,
         \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 ,
         \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 ,
         \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 ,
         \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 ,
         \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 ,
         \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 ,
         \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 ,
         \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 ,
         \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 ,
         \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 ,
         \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 ,
         \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 ,
         \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 ,
         \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 ,
         \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 ,
         \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 ,
         \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 ,
         \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 ,
         \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 ,
         \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 ,
         \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 ,
         \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 ,
         \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 ,
         \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 ,
         \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 ,
         \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 ,
         \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 ,
         \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 ,
         \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 ,
         \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 ,
         \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 ,
         \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 ,
         \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 ,
         \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 ,
         \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 ,
         \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 ,
         \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 ,
         \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 ,
         \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 ,
         \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 ,
         \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 ,
         \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 ,
         \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 ,
         \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 ,
         \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 ,
         \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 ,
         \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 ,
         \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 ,
         \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 ,
         \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 ,
         \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 ,
         \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 ,
         \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 ,
         \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 ,
         \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 ,
         \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 ,
         \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 ,
         \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 ,
         \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 ,
         \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 ,
         \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 ,
         \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 ,
         \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 ,
         \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 ,
         \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 ,
         \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 ,
         \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 ,
         \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 ,
         \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 ,
         \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 ,
         \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 ,
         \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 ,
         \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 ,
         \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 ,
         \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 ,
         \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 ,
         \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 ,
         \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 ,
         \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 ,
         \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 ,
         \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 ,
         \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 ,
         \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 ,
         \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 ,
         \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 ,
         \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 ,
         \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 ,
         \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 ,
         \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 ,
         \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 ,
         \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 ,
         \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 ,
         \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 ,
         \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 ,
         \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 ,
         \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 ,
         \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 ,
         \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 ,
         \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 ,
         \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 ,
         \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 ,
         \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 ,
         \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 ,
         \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 ,
         \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 ,
         \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 ,
         \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 ,
         \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 ,
         \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 ,
         \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 ,
         \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 ,
         \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 ,
         \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 ,
         \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 ,
         \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 ,
         \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 ,
         \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 ,
         \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 ,
         \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 ,
         \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 ,
         \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 ,
         \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 ,
         \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 ,
         \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 ,
         \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 ,
         \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 ,
         \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 ,
         \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 ,
         \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 ,
         \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 ,
         \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 ,
         \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 ,
         \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 ,
         \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 ,
         \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 ,
         \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 ,
         \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 ,
         \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 ,
         \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 ,
         \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 ,
         \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 ,
         \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 ,
         \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 ,
         \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 ,
         \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 ,
         \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 ,
         \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 ,
         \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 ,
         \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 ,
         \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 ,
         \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 ,
         \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 ,
         \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 ,
         \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 ,
         \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 ,
         \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 ,
         \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 ,
         \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 ,
         \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 ,
         \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 ,
         \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 ,
         \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 ,
         \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 ,
         \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 ,
         \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 ,
         \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 ,
         \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 ,
         \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 ,
         \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 ,
         \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 ,
         \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 ,
         \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 ,
         \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 ,
         \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 ,
         \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 ,
         \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 ,
         \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 ,
         \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 ,
         \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 ,
         \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 ,
         \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 ,
         \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 ,
         \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 ,
         \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 ,
         \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 ,
         \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 ,
         \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 ,
         \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 ,
         \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 ,
         \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 ,
         \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 ,
         \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 ,
         \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 ,
         \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 ,
         \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 ,
         \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 ,
         \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 ,
         \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 ,
         \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 ,
         \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 ,
         \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 ,
         \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 ,
         \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 ,
         \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 ,
         \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 ,
         \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 ,
         \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 ,
         \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 ,
         \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 ,
         \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 ,
         \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 ,
         \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 ,
         \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 ,
         \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 ,
         \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 ,
         \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 ,
         \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 ,
         \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 ,
         \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 ,
         \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 ,
         \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 ,
         \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 ,
         \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 ,
         \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 ,
         \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 ,
         \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 ,
         \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 ,
         \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 ,
         \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 ,
         \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 ,
         \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 ,
         \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 ,
         \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 ,
         \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 ,
         \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 ,
         \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 ,
         \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 ,
         \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 ,
         \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 ,
         \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 ,
         \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 ,
         \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 ,
         \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 ,
         \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 ,
         \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 ,
         \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 ,
         \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 ,
         \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 ,
         \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 ,
         \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 ,
         \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 ,
         \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 ,
         \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 ,
         \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 ,
         \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 ,
         \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 ,
         \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 ,
         \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 ,
         \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 ,
         \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 ,
         \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 ,
         \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 ,
         \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 ,
         \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 ,
         \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 ,
         \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 ,
         \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 ,
         \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 ,
         \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 ,
         \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 ,
         \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 ,
         \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 ,
         \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 ,
         \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 ,
         \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 ,
         \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 ,
         \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 ,
         \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 ,
         \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 ,
         \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 ,
         \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 ,
         \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 ,
         \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 ,
         \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 ,
         \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 ,
         \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 ,
         \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 ,
         \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 ,
         \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 ,
         \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 ,
         \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 ,
         \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 ,
         \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 ,
         \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 ,
         \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 , \10941 , \10942 ,
         \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 , \10951 , \10952 ,
         \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 , \10961 , \10962 ,
         \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 , \10971 , \10972 ,
         \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 , \10981 , \10982 ,
         \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 , \10991 , \10992 ,
         \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 , \11001 , \11002 ,
         \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 , \11011 , \11012 ,
         \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 , \11021 , \11022 ,
         \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 , \11031 , \11032 ,
         \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 , \11041 , \11042 ,
         \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 , \11051 , \11052 ,
         \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 , \11061 , \11062 ,
         \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 , \11071 , \11072 ,
         \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 , \11081 , \11082 ,
         \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 , \11091 , \11092 ,
         \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 , \11101 , \11102 ,
         \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 , \11111 , \11112 ,
         \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 , \11121 , \11122 ,
         \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 , \11131 , \11132 ,
         \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 , \11141 , \11142 ,
         \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 , \11151 , \11152 ,
         \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 , \11161 , \11162 ,
         \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 , \11171 , \11172 ,
         \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 , \11181 , \11182 ,
         \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 , \11191 , \11192 ,
         \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 , \11201 , \11202 ,
         \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 , \11211 , \11212 ,
         \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 , \11221 , \11222 ,
         \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 , \11231 , \11232 ,
         \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 , \11241 , \11242 ,
         \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 , \11251 , \11252 ,
         \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 , \11261 , \11262 ,
         \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 , \11271 , \11272 ,
         \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 , \11281 , \11282 ,
         \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 , \11291 , \11292 ,
         \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 , \11301 , \11302 ,
         \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 , \11311 , \11312 ,
         \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 , \11321 , \11322 ,
         \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 , \11331 , \11332 ,
         \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 , \11341 , \11342 ,
         \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 , \11351 , \11352 ,
         \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 , \11361 , \11362 ,
         \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 , \11371 , \11372 ,
         \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 , \11381 , \11382 ,
         \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 , \11391 , \11392 ,
         \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 , \11401 , \11402 ,
         \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 , \11411 , \11412 ,
         \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 , \11421 , \11422 ,
         \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 , \11431 , \11432 ,
         \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 , \11441 , \11442 ,
         \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 , \11451 , \11452 ,
         \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 , \11461 , \11462 ,
         \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 , \11471 , \11472 ,
         \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 , \11481 , \11482 ,
         \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 , \11491 , \11492 ,
         \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 , \11501 , \11502 ,
         \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 , \11511 , \11512 ,
         \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 , \11521 , \11522 ,
         \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 , \11531 , \11532 ,
         \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 , \11541 , \11542 ,
         \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 , \11551 , \11552 ,
         \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 , \11561 , \11562 ,
         \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 , \11571 , \11572 ,
         \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 , \11581 , \11582 ,
         \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 , \11591 , \11592 ,
         \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 , \11601 , \11602 ,
         \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 , \11611 , \11612 ,
         \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 , \11621 , \11622 ,
         \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 , \11631 , \11632 ,
         \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 , \11641 , \11642 ,
         \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 , \11651 , \11652 ,
         \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 , \11661 , \11662 ,
         \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 , \11671 , \11672 ,
         \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 , \11681 , \11682 ,
         \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 , \11691 , \11692 ,
         \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 , \11701 , \11702 ,
         \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 , \11711 , \11712 ,
         \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 , \11721 , \11722 ,
         \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 , \11731 , \11732 ,
         \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 , \11741 , \11742 ,
         \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 , \11751 , \11752 ,
         \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 , \11761 , \11762 ,
         \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 , \11771 , \11772 ,
         \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 , \11781 , \11782 ,
         \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 , \11791 , \11792 ,
         \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 , \11801 , \11802 ,
         \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 , \11811 , \11812 ,
         \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 , \11821 , \11822 ,
         \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 , \11831 , \11832 ,
         \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 , \11841 , \11842 ,
         \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 , \11851 , \11852 ,
         \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 , \11861 , \11862 ,
         \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 , \11871 , \11872 ,
         \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 , \11881 , \11882 ,
         \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 , \11891 , \11892 ,
         \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 , \11901 , \11902 ,
         \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 , \11911 , \11912 ,
         \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 , \11921 , \11922 ,
         \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 , \11931 , \11932 ,
         \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 , \11941 , \11942 ,
         \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 , \11951 , \11952 ,
         \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 , \11961 , \11962 ,
         \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 , \11971 , \11972 ,
         \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 , \11981 , \11982 ,
         \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 , \11991 , \11992 ,
         \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 , \12001 , \12002 ,
         \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 , \12011 , \12012 ,
         \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 , \12021 , \12022 ,
         \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 , \12031 , \12032 ,
         \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 , \12041 , \12042 ,
         \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 , \12051 , \12052 ,
         \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 , \12061 , \12062 ,
         \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 , \12071 , \12072 ,
         \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 , \12081 , \12082 ,
         \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 , \12091 , \12092 ,
         \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 , \12101 , \12102 ,
         \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 , \12111 , \12112 ,
         \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 , \12121 , \12122 ,
         \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 , \12131 , \12132 ,
         \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 , \12141 , \12142 ,
         \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 , \12151 , \12152 ,
         \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 , \12161 , \12162 ,
         \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 , \12171 , \12172 ,
         \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 , \12181 , \12182 ,
         \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 , \12191 , \12192 ,
         \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 , \12201 , \12202 ,
         \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 , \12211 , \12212 ,
         \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 , \12221 , \12222 ,
         \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 , \12231 , \12232 ,
         \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 , \12241 , \12242 ,
         \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 , \12251 , \12252 ,
         \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 , \12261 , \12262 ,
         \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 , \12271 , \12272 ,
         \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 , \12281 , \12282 ,
         \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 , \12291 , \12292 ,
         \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 , \12301 , \12302 ,
         \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 , \12311 , \12312 ,
         \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 , \12321 , \12322 ,
         \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 , \12331 , \12332 ,
         \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 , \12341 , \12342 ,
         \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 , \12351 , \12352 ,
         \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 , \12361 , \12362 ,
         \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 , \12371 , \12372 ,
         \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 , \12381 , \12382 ,
         \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 , \12391 , \12392 ,
         \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 , \12401 , \12402 ,
         \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 , \12411 , \12412 ,
         \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 , \12421 , \12422 ,
         \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 , \12431 , \12432 ,
         \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 , \12441 , \12442 ,
         \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 , \12451 , \12452 ,
         \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 , \12461 , \12462 ,
         \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 , \12471 , \12472 ,
         \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 , \12481 , \12482 ,
         \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 , \12491 , \12492 ,
         \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 , \12501 , \12502 ,
         \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 , \12511 , \12512 ,
         \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 , \12521 , \12522 ,
         \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 , \12531 , \12532 ,
         \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 , \12541 , \12542 ,
         \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 , \12551 , \12552 ,
         \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 , \12561 , \12562 ,
         \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 , \12571 , \12572 ,
         \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 , \12581 , \12582 ,
         \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 , \12591 , \12592 ,
         \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 , \12601 , \12602 ,
         \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 , \12611 , \12612 ,
         \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 , \12621 , \12622 ,
         \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 , \12631 , \12632 ,
         \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 , \12641 , \12642 ,
         \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 , \12651 , \12652 ,
         \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 , \12661 , \12662 ,
         \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 , \12671 , \12672 ,
         \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 , \12681 , \12682 ,
         \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 , \12691 , \12692 ,
         \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 , \12701 , \12702 ,
         \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 , \12711 , \12712 ,
         \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 , \12721 , \12722 ,
         \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 , \12731 , \12732 ,
         \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 , \12741 , \12742 ,
         \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 , \12751 , \12752 ,
         \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 , \12761 , \12762 ,
         \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 , \12771 , \12772 ,
         \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 , \12781 , \12782 ,
         \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 , \12791 , \12792 ,
         \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 , \12801 , \12802 ,
         \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 , \12811 , \12812 ,
         \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 , \12821 , \12822 ,
         \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 , \12831 , \12832 ,
         \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 , \12841 , \12842 ,
         \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 , \12851 , \12852 ,
         \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 , \12861 , \12862 ,
         \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 , \12871 , \12872 ,
         \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 , \12881 , \12882 ,
         \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 , \12891 , \12892 ,
         \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 , \12901 , \12902 ,
         \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 , \12911 , \12912 ,
         \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 , \12921 , \12922 ,
         \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 , \12931 , \12932 ,
         \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 , \12941 , \12942 ,
         \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 , \12951 , \12952 ,
         \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 , \12961 , \12962 ,
         \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 , \12971 , \12972 ,
         \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 , \12981 , \12982 ,
         \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 , \12991 , \12992 ,
         \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 , \13001 , \13002 ,
         \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 , \13011 , \13012 ,
         \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 , \13021 , \13022 ,
         \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 , \13031 , \13032 ,
         \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 , \13041 , \13042 ,
         \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 , \13051 , \13052 ,
         \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 , \13061 , \13062 ,
         \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 , \13071 , \13072 ,
         \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 , \13081 , \13082 ,
         \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 , \13091 , \13092 ,
         \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 , \13101 , \13102 ,
         \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 , \13111 , \13112 ,
         \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 , \13121 , \13122 ,
         \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 , \13131 , \13132 ,
         \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 , \13141 , \13142 ,
         \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 , \13151 , \13152 ,
         \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 , \13161 , \13162 ,
         \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 , \13171 , \13172 ,
         \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 , \13181 , \13182 ,
         \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 , \13191 , \13192 ,
         \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 , \13201 , \13202 ,
         \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 , \13211 , \13212 ,
         \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 , \13221 , \13222 ,
         \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 , \13231 , \13232 ,
         \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 , \13241 , \13242 ,
         \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 , \13251 , \13252 ,
         \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 , \13261 , \13262 ,
         \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 , \13271 , \13272 ,
         \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 , \13281 , \13282 ,
         \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 , \13291 , \13292 ,
         \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 , \13301 , \13302 ,
         \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 , \13311 , \13312 ,
         \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 , \13321 , \13322 ,
         \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 , \13331 , \13332 ,
         \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 , \13341 , \13342 ,
         \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 , \13351 , \13352 ,
         \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 , \13361 , \13362 ,
         \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 , \13371 , \13372 ,
         \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 , \13381 , \13382 ,
         \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 , \13391 , \13392 ,
         \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 , \13401 , \13402 ,
         \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 , \13411 , \13412 ,
         \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 , \13421 , \13422 ,
         \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 , \13431 , \13432 ,
         \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 , \13441 , \13442 ,
         \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 , \13451 , \13452 ,
         \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 , \13461 , \13462 ,
         \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 , \13471 , \13472 ,
         \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 , \13481 , \13482 ,
         \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 , \13491 , \13492 ,
         \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 , \13501 , \13502 ,
         \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 , \13511 , \13512 ,
         \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 , \13521 , \13522 ,
         \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 , \13531 , \13532 ,
         \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 , \13541 , \13542 ,
         \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 , \13551 , \13552 ,
         \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 , \13561 , \13562 ,
         \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 , \13571 , \13572 ,
         \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 , \13581 , \13582 ,
         \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 , \13591 , \13592 ,
         \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 , \13601 , \13602 ,
         \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 , \13611 , \13612 ,
         \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 , \13621 , \13622 ,
         \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 , \13631 , \13632 ,
         \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 , \13641 , \13642 ,
         \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 , \13651 , \13652 ,
         \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 , \13661 , \13662 ,
         \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 , \13671 , \13672 ,
         \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 , \13681 , \13682 ,
         \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 , \13691 , \13692 ,
         \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 , \13701 , \13702 ,
         \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 , \13711 , \13712 ,
         \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 , \13721 , \13722 ,
         \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 , \13731 , \13732 ,
         \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 , \13741 , \13742 ,
         \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 , \13751 , \13752 ,
         \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 , \13761 , \13762 ,
         \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 , \13771 , \13772 ,
         \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 , \13781 , \13782 ,
         \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 , \13791 , \13792 ,
         \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 , \13801 , \13802 ,
         \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 , \13811 , \13812 ,
         \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 , \13821 , \13822 ,
         \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 , \13831 , \13832 ,
         \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 , \13841 , \13842 ,
         \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 , \13851 , \13852 ,
         \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 , \13861 , \13862 ,
         \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 , \13871 , \13872 ,
         \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 , \13881 , \13882 ,
         \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 , \13891 , \13892 ,
         \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 , \13901 , \13902 ,
         \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 , \13911 , \13912 ,
         \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 , \13921 , \13922 ,
         \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 , \13931 , \13932 ,
         \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 , \13941 , \13942 ,
         \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 , \13951 , \13952 ,
         \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 , \13961 , \13962 ,
         \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 , \13971 , \13972 ,
         \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 , \13981 , \13982 ,
         \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 , \13991 , \13992 ,
         \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 , \14001 , \14002 ,
         \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 , \14011 , \14012 ,
         \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 , \14021 , \14022 ,
         \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 , \14031 , \14032 ,
         \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 , \14041 , \14042 ,
         \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 , \14051 , \14052 ,
         \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 , \14061 , \14062 ,
         \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 , \14071 , \14072 ,
         \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 , \14081 , \14082 ,
         \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 , \14091 , \14092 ,
         \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 , \14101 , \14102 ,
         \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 , \14111 , \14112 ,
         \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 , \14121 , \14122 ,
         \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 , \14131 , \14132 ,
         \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 , \14141 , \14142 ,
         \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 , \14151 , \14152 ,
         \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 , \14161 , \14162 ,
         \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 , \14171 , \14172 ,
         \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 , \14181 , \14182 ,
         \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 , \14191 , \14192 ,
         \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 , \14201 , \14202 ,
         \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 , \14211 , \14212 ,
         \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 , \14221 , \14222 ,
         \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 , \14231 , \14232 ,
         \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 , \14241 , \14242 ,
         \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 , \14251 , \14252 ,
         \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 , \14261 , \14262 ,
         \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 , \14271 , \14272 ,
         \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 , \14281 , \14282 ,
         \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 , \14291 , \14292 ,
         \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 , \14301 , \14302 ,
         \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 , \14311 , \14312 ,
         \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 , \14321 , \14322 ,
         \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 , \14331 , \14332 ,
         \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 , \14341 , \14342 ,
         \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 , \14351 , \14352 ,
         \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 , \14361 , \14362 ,
         \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 , \14371 , \14372 ,
         \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 , \14381 , \14382 ,
         \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 , \14391 , \14392 ,
         \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 , \14401 , \14402 ,
         \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 , \14411 , \14412 ,
         \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 , \14421 , \14422 ,
         \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 , \14431 , \14432 ,
         \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 , \14441 , \14442 ,
         \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 , \14451 , \14452 ,
         \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 , \14461 , \14462 ,
         \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 , \14471 , \14472 ,
         \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 , \14481 , \14482 ,
         \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 , \14491 , \14492 ,
         \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 , \14501 , \14502 ,
         \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 , \14511 , \14512 ,
         \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 , \14521 , \14522 ,
         \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 , \14531 , \14532 ,
         \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 , \14541 , \14542 ,
         \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 , \14551 , \14552 ,
         \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 , \14561 , \14562 ,
         \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 , \14571 , \14572 ,
         \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 , \14581 , \14582 ,
         \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 , \14591 , \14592 ,
         \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 , \14601 , \14602 ,
         \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 , \14611 , \14612 ,
         \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 , \14621 , \14622 ,
         \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 , \14631 , \14632 ,
         \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 , \14641 , \14642 ,
         \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 , \14651 , \14652 ,
         \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 , \14661 , \14662 ,
         \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 , \14671 , \14672 ,
         \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 , \14681 , \14682 ,
         \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 , \14691 , \14692 ,
         \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 , \14701 , \14702 ,
         \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 , \14711 , \14712 ,
         \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 , \14721 , \14722 ,
         \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 , \14731 , \14732 ,
         \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 , \14741 , \14742 ,
         \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 , \14751 , \14752 ,
         \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 , \14761 , \14762 ,
         \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 , \14771 , \14772 ,
         \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 , \14781 , \14782 ,
         \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 , \14791 , \14792 ,
         \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 , \14801 , \14802 ,
         \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 , \14811 , \14812 ,
         \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 , \14821 , \14822 ,
         \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 , \14831 , \14832 ,
         \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 , \14841 , \14842 ,
         \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 , \14851 , \14852 ,
         \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 , \14861 , \14862 ,
         \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 , \14871 , \14872 ,
         \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 , \14881 , \14882 ,
         \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 , \14891 , \14892 ,
         \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 , \14901 , \14902 ,
         \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 , \14911 , \14912 ,
         \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 , \14921 , \14922 ,
         \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 , \14931 , \14932 ,
         \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 , \14941 , \14942 ,
         \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 , \14951 , \14952 ,
         \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 , \14961 , \14962 ,
         \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 , \14971 , \14972 ,
         \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 , \14981 , \14982 ,
         \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 , \14991 , \14992 ,
         \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 , \15001 , \15002 ,
         \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 , \15011 , \15012 ,
         \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 , \15021 , \15022 ,
         \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 , \15031 , \15032 ,
         \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 , \15041 , \15042 ,
         \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 , \15051 , \15052 ,
         \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 , \15061 , \15062 ,
         \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 , \15071 , \15072 ,
         \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 , \15081 , \15082 ,
         \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 , \15091 , \15092 ,
         \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 , \15101 , \15102 ,
         \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 , \15111 , \15112 ,
         \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 , \15121 , \15122 ,
         \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 , \15131 , \15132 ,
         \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 , \15141 , \15142 ,
         \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 , \15151 , \15152 ,
         \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 , \15161 , \15162 ,
         \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 , \15171 , \15172 ,
         \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 , \15181 , \15182 ,
         \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 , \15191 , \15192 ,
         \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 , \15201 , \15202 ,
         \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 , \15211 , \15212 ,
         \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 , \15221 , \15222 ,
         \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 , \15231 , \15232 ,
         \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 , \15241 , \15242 ,
         \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 , \15251 , \15252 ,
         \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 , \15261 , \15262 ,
         \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 , \15271 , \15272 ,
         \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 , \15281 , \15282 ,
         \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 , \15291 , \15292 ,
         \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 , \15301 , \15302 ,
         \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 , \15311 , \15312 ,
         \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 , \15321 , \15322 ,
         \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 , \15331 , \15332 ,
         \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 , \15341 , \15342 ,
         \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 , \15351 , \15352 ,
         \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 , \15361 , \15362 ,
         \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 , \15371 , \15372 ,
         \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 , \15381 , \15382 ,
         \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 , \15391 , \15392 ,
         \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 , \15401 , \15402 ,
         \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 , \15411 , \15412 ,
         \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 , \15421 , \15422 ,
         \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 , \15431 , \15432 ,
         \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 , \15441 , \15442 ,
         \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 , \15451 , \15452 ,
         \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 , \15461 , \15462 ,
         \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 , \15471 , \15472 ,
         \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 , \15481 , \15482 ,
         \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 , \15491 , \15492 ,
         \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 , \15501 , \15502 ,
         \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 , \15511 , \15512 ,
         \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 , \15521 , \15522 ,
         \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 , \15531 , \15532 ,
         \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 , \15541 , \15542 ,
         \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 , \15551 , \15552 ,
         \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 , \15561 , \15562 ,
         \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 , \15571 , \15572 ,
         \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 , \15581 , \15582 ,
         \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 , \15591 , \15592 ,
         \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 , \15601 , \15602 ,
         \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 , \15611 , \15612 ,
         \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 , \15621 , \15622 ,
         \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 , \15631 , \15632 ,
         \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 , \15641 , \15642 ,
         \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 , \15651 , \15652 ,
         \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 , \15661 , \15662 ,
         \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 , \15671 , \15672 ,
         \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 , \15681 , \15682 ,
         \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 , \15691 , \15692 ,
         \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 , \15701 , \15702 ,
         \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 , \15711 , \15712 ,
         \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 , \15721 , \15722 ,
         \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 , \15731 , \15732 ,
         \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 , \15741 , \15742 ,
         \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 , \15751 , \15752 ,
         \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 , \15761 , \15762 ,
         \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 , \15771 , \15772 ,
         \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 , \15781 , \15782 ,
         \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 , \15791 , \15792 ,
         \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 , \15801 , \15802 ,
         \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 , \15811 , \15812 ,
         \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 , \15821 , \15822 ,
         \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 , \15831 , \15832 ,
         \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 , \15841 , \15842 ,
         \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 , \15851 , \15852 ,
         \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 , \15861 , \15862 ,
         \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 , \15871 , \15872 ,
         \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 , \15881 , \15882 ,
         \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 , \15891 , \15892 ,
         \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 , \15901 , \15902 ,
         \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 , \15911 , \15912 ,
         \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 , \15921 , \15922 ,
         \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 , \15931 , \15932 ,
         \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 , \15941 , \15942 ,
         \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 , \15951 , \15952 ,
         \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 , \15961 , \15962 ,
         \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 , \15971 , \15972 ,
         \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 , \15981 , \15982 ,
         \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 , \15991 , \15992 ,
         \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 , \16001 , \16002 ,
         \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 , \16011 , \16012 ,
         \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 , \16021 , \16022 ,
         \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 , \16031 , \16032 ,
         \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 , \16041 , \16042 ,
         \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 , \16051 , \16052 ,
         \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 , \16061 , \16062 ,
         \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 , \16071 , \16072 ,
         \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 , \16081 , \16082 ,
         \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 , \16091 , \16092 ,
         \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 , \16101 , \16102 ,
         \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 , \16111 , \16112 ,
         \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 , \16121 , \16122 ,
         \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 , \16131 , \16132 ,
         \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 , \16141 , \16142 ,
         \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 , \16151 , \16152 ,
         \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 , \16161 , \16162 ,
         \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 , \16171 , \16172 ,
         \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 , \16181 , \16182 ,
         \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 , \16191 , \16192 ,
         \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 , \16201 , \16202 ,
         \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 , \16211 , \16212 ,
         \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 , \16221 , \16222 ,
         \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 , \16231 , \16232 ,
         \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 , \16241 , \16242 ,
         \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 , \16251 , \16252 ,
         \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 , \16261 , \16262 ,
         \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 , \16271 , \16272 ,
         \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 , \16281 , \16282 ,
         \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 , \16291 , \16292 ,
         \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 , \16301 , \16302 ,
         \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 , \16311 , \16312 ,
         \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 , \16321 , \16322 ,
         \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 , \16331 , \16332 ,
         \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 , \16341 , \16342 ,
         \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 , \16351 , \16352 ,
         \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 , \16361 , \16362 ,
         \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 , \16371 , \16372 ,
         \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 , \16381 , \16382 ,
         \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 , \16391 , \16392 ,
         \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 , \16401 , \16402 ,
         \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 , \16411 , \16412 ,
         \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 , \16421 , \16422 ,
         \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 , \16431 , \16432 ,
         \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 , \16441 , \16442 ,
         \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 , \16451 , \16452 ,
         \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 , \16461 , \16462 ,
         \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 , \16471 , \16472 ,
         \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 , \16481 , \16482 ,
         \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 , \16491 , \16492 ,
         \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 , \16501 , \16502 ,
         \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 , \16511 , \16512 ,
         \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 , \16521 , \16522 ,
         \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 , \16531 , \16532 ,
         \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 , \16541 , \16542 ,
         \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 , \16551 , \16552 ,
         \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 , \16561 , \16562 ,
         \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 , \16571 , \16572 ,
         \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 , \16581 , \16582 ,
         \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 , \16591 , \16592 ,
         \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 , \16601 , \16602 ,
         \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 , \16611 , \16612 ,
         \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 , \16621 , \16622 ,
         \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 , \16631 , \16632 ,
         \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 , \16641 , \16642 ,
         \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 , \16651 , \16652 ,
         \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 , \16661 , \16662 ,
         \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 , \16671 , \16672 ,
         \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 , \16681 , \16682 ,
         \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 , \16691 , \16692 ,
         \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 , \16701 , \16702 ,
         \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 , \16711 , \16712 ,
         \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 , \16721 , \16722 ,
         \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 , \16731 , \16732 ,
         \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 , \16741 , \16742 ,
         \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 , \16751 , \16752 ,
         \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 , \16761 , \16762 ,
         \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 , \16771 , \16772 ,
         \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 , \16781 , \16782 ,
         \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 , \16791 , \16792 ,
         \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 , \16801 , \16802 ,
         \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 , \16811 , \16812 ,
         \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 , \16821 , \16822 ,
         \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 , \16831 , \16832 ,
         \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 , \16841 , \16842 ,
         \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 , \16851 , \16852 ,
         \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 , \16861 , \16862 ,
         \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 , \16871 , \16872 ,
         \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 , \16881 , \16882 ,
         \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 , \16891 , \16892 ,
         \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 , \16901 , \16902 ,
         \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 , \16911 , \16912 ,
         \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 , \16921 , \16922 ,
         \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 , \16931 , \16932 ,
         \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 , \16941 , \16942 ,
         \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 , \16951 , \16952 ,
         \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 , \16961 , \16962 ,
         \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 , \16971 , \16972 ,
         \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 , \16981 , \16982 ,
         \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 , \16991 , \16992 ,
         \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 , \17001 , \17002 ,
         \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 , \17011 , \17012 ,
         \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 , \17021 , \17022 ,
         \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 , \17031 , \17032 ,
         \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 , \17041 , \17042 ,
         \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 , \17051 , \17052 ,
         \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 , \17061 , \17062 ,
         \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 , \17071 , \17072 ,
         \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 , \17081 , \17082 ,
         \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 , \17091 , \17092 ,
         \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 , \17101 , \17102 ,
         \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 , \17111 , \17112 ,
         \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 , \17121 , \17122 ,
         \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 , \17131 , \17132 ,
         \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 , \17141 , \17142 ,
         \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 , \17151 , \17152 ,
         \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 , \17161 , \17162 ,
         \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 , \17171 , \17172 ,
         \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 , \17181 , \17182 ,
         \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 , \17191 , \17192 ,
         \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 , \17201 , \17202 ,
         \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 , \17211 , \17212 ,
         \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 , \17221 , \17222 ,
         \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 , \17231 , \17232 ,
         \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 , \17241 , \17242 ,
         \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 , \17251 , \17252 ,
         \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 , \17261 , \17262 ,
         \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 , \17271 , \17272 ,
         \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 , \17281 , \17282 ,
         \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 , \17291 , \17292 ,
         \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 , \17301 , \17302 ,
         \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 , \17311 , \17312 ,
         \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 , \17321 , \17322 ,
         \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 , \17331 , \17332 ,
         \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 , \17341 , \17342 ,
         \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 , \17351 , \17352 ,
         \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 , \17361 , \17362 ,
         \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 , \17371 , \17372 ,
         \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 , \17381 , \17382 ,
         \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 , \17391 , \17392 ,
         \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 , \17401 , \17402 ,
         \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 , \17411 , \17412 ,
         \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 , \17421 , \17422 ,
         \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 , \17431 , \17432 ,
         \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 , \17441 , \17442 ,
         \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 , \17451 , \17452 ,
         \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 , \17461 , \17462 ,
         \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 , \17471 , \17472 ,
         \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 , \17481 , \17482 ,
         \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 , \17491 , \17492 ,
         \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 , \17501 , \17502 ,
         \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 , \17511 , \17512 ,
         \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 , \17521 , \17522 ,
         \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 , \17531 , \17532 ,
         \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 , \17541 , \17542 ,
         \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 , \17551 , \17552 ,
         \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 , \17561 , \17562 ,
         \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 , \17571 , \17572 ,
         \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 , \17581 , \17582 ,
         \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 , \17591 , \17592 ,
         \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 , \17601 , \17602 ,
         \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 , \17611 , \17612 ,
         \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 , \17621 , \17622 ,
         \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 , \17631 , \17632 ,
         \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 , \17641 , \17642 ,
         \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 , \17651 , \17652 ,
         \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 , \17661 , \17662 ,
         \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 , \17671 , \17672 ,
         \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 , \17681 , \17682 ,
         \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 , \17691 , \17692 ,
         \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 , \17701 , \17702 ,
         \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 , \17711 , \17712 ,
         \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 , \17721 , \17722 ,
         \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 , \17731 , \17732 ,
         \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 , \17741 , \17742 ,
         \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 , \17751 , \17752 ,
         \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 , \17761 , \17762 ,
         \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 , \17771 , \17772 ,
         \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 , \17781 , \17782 ,
         \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 , \17791 , \17792 ,
         \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 , \17801 , \17802 ,
         \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 , \17811 , \17812 ,
         \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 , \17821 , \17822 ,
         \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 , \17831 , \17832 ,
         \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 , \17841 , \17842 ,
         \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 , \17851 , \17852 ,
         \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 , \17861 , \17862 ,
         \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 , \17871 , \17872 ,
         \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 , \17881 , \17882 ,
         \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 , \17891 , \17892 ,
         \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 , \17901 , \17902 ,
         \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 , \17911 , \17912 ,
         \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 , \17921 , \17922 ,
         \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 , \17931 , \17932 ,
         \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 , \17941 , \17942 ,
         \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 , \17951 , \17952 ,
         \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 , \17961 , \17962 ,
         \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 , \17971 , \17972 ,
         \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 , \17981 , \17982 ,
         \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 , \17991 , \17992 ,
         \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 , \18001 , \18002 ,
         \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 , \18011 , \18012 ,
         \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 , \18021 , \18022 ,
         \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 , \18031 , \18032 ,
         \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 , \18041 , \18042 ,
         \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 , \18051 , \18052 ,
         \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 , \18061 , \18062 ,
         \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 , \18071 , \18072 ,
         \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 , \18081 , \18082 ,
         \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 , \18091 , \18092 ,
         \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 , \18101 , \18102 ,
         \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 , \18111 , \18112 ,
         \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 , \18121 , \18122 ,
         \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 , \18131 , \18132 ,
         \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 , \18141 , \18142 ,
         \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 , \18151 , \18152 ,
         \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 , \18161 , \18162 ,
         \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 , \18171 , \18172 ,
         \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 , \18181 , \18182 ,
         \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 , \18191 , \18192 ,
         \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 , \18201 , \18202 ,
         \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 , \18211 , \18212 ,
         \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 , \18221 , \18222 ,
         \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 , \18231 , \18232 ,
         \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 , \18241 , \18242 ,
         \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 , \18251 , \18252 ,
         \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 , \18261 , \18262 ,
         \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 , \18271 , \18272 ,
         \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 , \18281 , \18282 ,
         \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 , \18291 , \18292 ,
         \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 , \18301 , \18302 ,
         \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 , \18311 , \18312 ,
         \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 , \18321 , \18322 ,
         \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 , \18331 , \18332 ,
         \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 , \18341 , \18342 ,
         \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 , \18351 , \18352 ,
         \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 , \18361 , \18362 ,
         \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 , \18371 , \18372 ,
         \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 , \18381 , \18382 ,
         \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 , \18391 , \18392 ,
         \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 , \18401 , \18402 ,
         \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 , \18411 , \18412 ,
         \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 , \18421 , \18422 ,
         \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 , \18431 , \18432 ,
         \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 , \18441 , \18442 ,
         \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 , \18451 , \18452 ,
         \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 , \18461 , \18462 ,
         \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 , \18471 , \18472 ,
         \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 , \18481 , \18482 ,
         \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 , \18491 , \18492 ,
         \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 , \18501 , \18502 ,
         \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 , \18511 , \18512 ,
         \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 , \18521 , \18522 ,
         \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 , \18531 , \18532 ,
         \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 , \18541 , \18542 ,
         \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 , \18551 , \18552 ,
         \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 , \18561 , \18562 ,
         \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 , \18571 , \18572 ,
         \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 , \18581 , \18582 ,
         \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 , \18591 , \18592 ,
         \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 , \18601 , \18602 ,
         \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 , \18611 , \18612 ,
         \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 , \18621 , \18622 ,
         \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 , \18631 , \18632 ,
         \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 , \18641 , \18642 ,
         \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 , \18651 , \18652 ,
         \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 , \18661 , \18662 ,
         \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 , \18671 , \18672 ,
         \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 , \18681 , \18682 ,
         \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 , \18691 , \18692 ,
         \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 , \18701 , \18702 ,
         \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 , \18711 , \18712 ,
         \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 , \18721 , \18722 ,
         \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 , \18731 , \18732 ,
         \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 , \18741 , \18742 ,
         \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 , \18751 , \18752 ,
         \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 , \18761 , \18762 ,
         \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 , \18771 , \18772 ,
         \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 , \18781 , \18782 ,
         \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 , \18791 , \18792 ,
         \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 , \18801 , \18802 ,
         \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 , \18811 , \18812 ,
         \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 , \18821 , \18822 ,
         \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 , \18831 , \18832 ,
         \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 , \18841 , \18842 ,
         \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 , \18851 , \18852 ,
         \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 , \18861 , \18862 ,
         \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 , \18871 , \18872 ,
         \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 , \18881 , \18882 ,
         \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 , \18891 , \18892 ,
         \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 , \18901 , \18902 ,
         \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 , \18911 , \18912 ,
         \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 , \18921 , \18922 ,
         \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 , \18931 , \18932 ,
         \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 , \18941 , \18942 ,
         \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 , \18951 , \18952 ,
         \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 , \18961 , \18962 ,
         \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 , \18971 , \18972 ,
         \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 , \18981 , \18982 ,
         \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 , \18991 , \18992 ,
         \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 , \19001 , \19002 ,
         \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 , \19011 , \19012 ,
         \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 , \19021 , \19022 ,
         \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 , \19031 , \19032 ,
         \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 , \19041 , \19042 ,
         \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 , \19051 , \19052 ,
         \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 , \19061 , \19062 ,
         \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 , \19071 , \19072 ,
         \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 , \19081 , \19082 ,
         \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 , \19091 , \19092 ,
         \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 , \19101 , \19102 ,
         \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 , \19111 , \19112 ,
         \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 , \19121 , \19122 ,
         \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 , \19131 , \19132 ,
         \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 , \19141 , \19142 ,
         \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 , \19151 , \19152 ,
         \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 , \19161 , \19162 ,
         \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 , \19171 , \19172 ,
         \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 , \19181 , \19182 ,
         \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 , \19191 , \19192 ,
         \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 , \19201 , \19202 ,
         \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 , \19211 , \19212 ,
         \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 , \19221 , \19222 ,
         \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 , \19231 , \19232 ,
         \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 , \19241 , \19242 ,
         \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 , \19251 , \19252 ,
         \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 , \19261 , \19262 ,
         \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 , \19271 , \19272 ,
         \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 , \19281 , \19282 ,
         \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 , \19291 , \19292 ,
         \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 , \19301 , \19302 ,
         \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 , \19311 , \19312 ,
         \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 , \19321 , \19322 ,
         \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 , \19331 , \19332 ,
         \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 , \19341 , \19342 ,
         \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 , \19351 , \19352 ,
         \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 , \19361 , \19362 ,
         \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 , \19371 , \19372 ,
         \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 , \19381 , \19382 ,
         \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 , \19391 , \19392 ,
         \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 , \19401 , \19402 ,
         \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 , \19411 , \19412 ,
         \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 , \19421 , \19422 ,
         \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 , \19431 , \19432 ,
         \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 , \19441 , \19442 ,
         \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 , \19451 , \19452 ,
         \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 , \19461 , \19462 ,
         \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 , \19471 , \19472 ,
         \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 , \19481 , \19482 ,
         \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 , \19491 , \19492 ,
         \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 , \19501 , \19502 ,
         \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 , \19511 , \19512 ,
         \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 , \19521 , \19522 ,
         \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 , \19531 , \19532 ,
         \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 , \19541 , \19542 ,
         \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 , \19551 , \19552 ,
         \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 , \19561 , \19562 ,
         \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 , \19571 , \19572 ,
         \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 , \19581 , \19582 ,
         \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 , \19591 , \19592 ,
         \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 , \19601 , \19602 ,
         \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 , \19611 , \19612 ,
         \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 , \19621 , \19622 ,
         \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 , \19631 , \19632 ,
         \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 , \19641 , \19642 ,
         \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 , \19651 , \19652 ,
         \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 , \19661 , \19662 ,
         \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 , \19671 , \19672 ,
         \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 , \19681 , \19682 ,
         \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 , \19691 , \19692 ,
         \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 , \19701 , \19702 ,
         \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 , \19711 , \19712 ,
         \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 , \19721 , \19722 ,
         \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 , \19731 , \19732 ,
         \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 , \19741 , \19742 ,
         \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 , \19751 , \19752 ,
         \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 , \19761 , \19762 ,
         \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 , \19771 , \19772 ,
         \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 , \19781 , \19782 ,
         \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 , \19791 , \19792 ,
         \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 , \19801 , \19802 ,
         \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 , \19811 , \19812 ,
         \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 , \19821 , \19822 ,
         \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 , \19831 , \19832 ,
         \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 , \19841 , \19842 ,
         \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 , \19851 , \19852 ,
         \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 , \19861 , \19862 ,
         \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 , \19871 , \19872 ,
         \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 , \19881 , \19882 ,
         \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 , \19891 , \19892 ,
         \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 , \19901 , \19902 ,
         \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 , \19911 , \19912 ,
         \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 , \19921 , \19922 ,
         \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 , \19931 , \19932 ,
         \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 , \19941 , \19942 ,
         \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 , \19951 , \19952 ,
         \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 , \19961 , \19962 ,
         \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 , \19971 , \19972 ,
         \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 , \19981 , \19982 ,
         \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 , \19991 , \19992 ,
         \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 , \20001 , \20002 ,
         \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 , \20011 , \20012 ,
         \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 , \20021 , \20022 ,
         \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 , \20031 , \20032 ,
         \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 , \20041 , \20042 ,
         \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 , \20051 , \20052 ,
         \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 , \20061 , \20062 ,
         \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 , \20071 , \20072 ,
         \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 , \20081 , \20082 ,
         \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 , \20091 , \20092 ,
         \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 , \20101 , \20102 ,
         \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 , \20111 , \20112 ,
         \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 , \20121 , \20122 ,
         \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 , \20131 , \20132 ,
         \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 , \20141 , \20142 ,
         \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 , \20151 , \20152 ,
         \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 , \20161 , \20162 ,
         \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 , \20171 , \20172 ,
         \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 , \20181 , \20182 ,
         \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 , \20191 , \20192 ,
         \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 , \20201 , \20202 ,
         \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 , \20211 , \20212 ,
         \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 , \20221 , \20222 ,
         \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 , \20231 , \20232 ,
         \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 , \20241 , \20242 ,
         \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 , \20251 , \20252 ,
         \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 , \20261 , \20262 ,
         \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 , \20271 , \20272 ,
         \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 , \20281 , \20282 ,
         \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 , \20291 , \20292 ,
         \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 , \20301 , \20302 ,
         \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 , \20311 , \20312 ,
         \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 , \20321 , \20322 ,
         \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 , \20331 , \20332 ,
         \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 , \20341 , \20342 ,
         \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 , \20351 , \20352 ,
         \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 , \20361 , \20362 ,
         \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 , \20371 , \20372 ,
         \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 , \20381 , \20382 ,
         \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 , \20391 , \20392 ,
         \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 , \20401 , \20402 ,
         \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 , \20411 , \20412 ,
         \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 , \20421 , \20422 ,
         \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 , \20431 , \20432 ,
         \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 , \20441 , \20442 ,
         \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 , \20451 , \20452 ,
         \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 , \20461 , \20462 ,
         \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 , \20471 , \20472 ,
         \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 , \20481 , \20482 ,
         \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 , \20491 , \20492 ,
         \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 , \20501 , \20502 ,
         \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 , \20511 , \20512 ,
         \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 , \20521 , \20522 ,
         \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 , \20531 , \20532 ,
         \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 , \20541 , \20542 ,
         \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 , \20551 , \20552 ,
         \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 , \20561 , \20562 ,
         \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 , \20571 , \20572 ,
         \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 , \20581 , \20582 ,
         \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 , \20591 , \20592 ,
         \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 , \20601 , \20602 ,
         \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 , \20611 , \20612 ,
         \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 , \20621 , \20622 ,
         \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 , \20631 , \20632 ,
         \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 , \20641 , \20642 ,
         \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 , \20651 , \20652 ,
         \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 , \20661 , \20662 ,
         \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 , \20671 , \20672 ,
         \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 , \20681 , \20682 ,
         \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 , \20691 , \20692 ,
         \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 , \20701 , \20702 ,
         \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 , \20711 , \20712 ,
         \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 , \20721 , \20722 ,
         \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 , \20731 , \20732 ,
         \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 , \20741 , \20742 ,
         \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 , \20751 , \20752 ,
         \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 , \20761 , \20762 ,
         \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 , \20771 , \20772 ,
         \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 , \20781 , \20782 ,
         \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 , \20791 , \20792 ,
         \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 , \20801 , \20802 ,
         \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 , \20811 , \20812 ,
         \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 , \20821 , \20822 ,
         \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 , \20831 , \20832 ,
         \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 , \20841 , \20842 ,
         \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 , \20851 , \20852 ,
         \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 , \20861 , \20862 ,
         \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 , \20871 , \20872 ,
         \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 , \20881 , \20882 ,
         \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 , \20891 , \20892 ,
         \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 , \20901 , \20902 ,
         \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 , \20911 , \20912 ,
         \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 , \20921 , \20922 ,
         \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 , \20931 , \20932 ,
         \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 , \20941 , \20942 ,
         \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 , \20951 , \20952 ,
         \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 , \20961 , \20962 ,
         \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 , \20971 , \20972 ,
         \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 , \20981 , \20982 ,
         \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 , \20991 , \20992 ,
         \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 , \21001 , \21002 ,
         \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 , \21011 , \21012 ,
         \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 , \21021 , \21022 ,
         \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 , \21031 , \21032 ,
         \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 , \21041 , \21042 ,
         \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 , \21051 , \21052 ,
         \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 , \21061 , \21062 ,
         \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 , \21071 , \21072 ,
         \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 , \21081 , \21082 ,
         \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 , \21091 , \21092 ,
         \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 , \21101 , \21102 ,
         \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 , \21111 , \21112 ,
         \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 , \21121 , \21122 ,
         \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 , \21131 , \21132 ,
         \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 , \21141 , \21142 ,
         \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 , \21151 , \21152 ,
         \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 , \21161 , \21162 ,
         \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 , \21171 , \21172 ,
         \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 , \21181 , \21182 ,
         \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 , \21191 , \21192 ,
         \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 , \21201 , \21202 ,
         \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 , \21211 , \21212 ,
         \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 , \21221 , \21222 ,
         \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 , \21231 , \21232 ,
         \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 , \21241 , \21242 ,
         \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 , \21251 , \21252 ,
         \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 , \21261 , \21262 ,
         \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 , \21271 , \21272 ,
         \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 , \21281 , \21282 ,
         \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 , \21291 , \21292 ,
         \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 , \21301 , \21302 ,
         \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 , \21311 , \21312 ,
         \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 , \21321 , \21322 ,
         \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 , \21331 , \21332 ,
         \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 , \21341 , \21342 ,
         \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 , \21351 , \21352 ,
         \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 , \21361 , \21362 ,
         \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370 , \21371 , \21372 ,
         \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 , \21381 , \21382 ,
         \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 , \21391 , \21392 ,
         \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 , \21401 , \21402 ,
         \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 , \21411 , \21412 ,
         \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 , \21421 , \21422 ,
         \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 , \21431 , \21432 ,
         \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 , \21441 , \21442 ,
         \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 , \21451 , \21452 ,
         \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 , \21461 , \21462 ,
         \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 , \21471 , \21472 ,
         \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 , \21481 , \21482 ,
         \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 , \21491 , \21492 ,
         \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 , \21501 , \21502 ,
         \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 , \21511 , \21512 ,
         \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 , \21521 , \21522 ,
         \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 , \21531 , \21532 ,
         \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 , \21541 , \21542 ,
         \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 , \21551 , \21552 ,
         \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 , \21561 , \21562 ,
         \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 , \21571 , \21572 ,
         \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 , \21581 , \21582 ,
         \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 , \21591 , \21592 ,
         \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 , \21601 , \21602 ,
         \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 , \21611 , \21612 ,
         \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 , \21621 , \21622 ,
         \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 , \21631 , \21632 ,
         \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 , \21641 , \21642 ,
         \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 , \21651 , \21652 ,
         \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 , \21661 , \21662 ,
         \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 , \21671 , \21672 ,
         \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 , \21681 , \21682 ,
         \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 , \21691 , \21692 ,
         \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 , \21701 , \21702 ,
         \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 , \21711 , \21712 ,
         \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 , \21721 , \21722 ,
         \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 , \21731 , \21732 ,
         \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 , \21741 , \21742 ,
         \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 , \21751 , \21752 ,
         \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 , \21761 , \21762 ,
         \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 , \21771 , \21772 ,
         \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 , \21781 , \21782 ,
         \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 , \21791 , \21792 ,
         \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 , \21801 , \21802 ,
         \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 , \21811 , \21812 ,
         \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 , \21821 , \21822 ,
         \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 , \21831 , \21832 ,
         \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 , \21841 , \21842 ,
         \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 , \21851 , \21852 ,
         \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 , \21861 , \21862 ,
         \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 , \21871 , \21872 ,
         \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 , \21881 , \21882 ,
         \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 , \21891 , \21892 ,
         \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 , \21901 , \21902 ,
         \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 , \21911 , \21912 ,
         \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 , \21921 , \21922 ,
         \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 , \21931 , \21932 ,
         \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 , \21941 , \21942 ,
         \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 , \21951 , \21952 ,
         \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 , \21961 , \21962 ,
         \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 , \21971 , \21972 ,
         \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 , \21981 , \21982 ,
         \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 , \21991 , \21992 ,
         \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 , \22001 , \22002 ,
         \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 , \22011 , \22012 ,
         \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 , \22021 , \22022 ,
         \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 , \22031 , \22032 ,
         \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 , \22041 , \22042 ,
         \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 , \22051 , \22052 ,
         \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 , \22061 , \22062 ,
         \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 , \22071 , \22072 ,
         \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 , \22081 , \22082 ,
         \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 , \22091 , \22092 ,
         \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 , \22101 , \22102 ,
         \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 , \22111 , \22112 ,
         \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 , \22121 , \22122 ,
         \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 , \22131 , \22132 ,
         \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 , \22141 , \22142 ,
         \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 , \22151 , \22152 ,
         \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 , \22161 , \22162 ,
         \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 , \22171 , \22172 ,
         \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 , \22181 , \22182 ,
         \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 , \22191 , \22192 ,
         \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 , \22201 , \22202 ,
         \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 , \22211 , \22212 ,
         \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 , \22221 , \22222 ,
         \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 , \22231 , \22232 ,
         \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 , \22241 , \22242 ,
         \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 , \22251 , \22252 ,
         \22253 , \22254 , \22255 , \22256 , \22257 , \22258 , \22259 , \22260 , \22261 , \22262 ,
         \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , \22269 , \22270 , \22271 , \22272 ,
         \22273 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 , \22281 , \22282 ,
         \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 , \22291 , \22292 ,
         \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 , \22301 , \22302 ,
         \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 , \22311 , \22312 ,
         \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 , \22321 , \22322 ,
         \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 , \22331 , \22332 ,
         \22333 , \22334 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 , \22341 , \22342 ,
         \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 , \22351 , \22352 ,
         \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 , \22361 , \22362 ,
         \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 , \22371 , \22372 ,
         \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 , \22381 , \22382 ,
         \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 , \22391 , \22392 ,
         \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 , \22401 , \22402 ,
         \22403 , \22404 , \22405 , \22406 , \22407 , \22408 , \22409 , \22410 , \22411 , \22412 ,
         \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 , \22421 , \22422 ,
         \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 , \22431 , \22432 ,
         \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 , \22441 , \22442 ,
         \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 , \22451 , \22452 ,
         \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 , \22461 , \22462 ,
         \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 , \22470 , \22471 , \22472 ,
         \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 , \22481 , \22482 ,
         \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 , \22491 , \22492 ,
         \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 , \22501 , \22502 ,
         \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 , \22511 , \22512 ,
         \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 , \22521 , \22522 ,
         \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 , \22531 , \22532 ,
         \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 , \22541 , \22542 ,
         \22543 , \22544 , \22545 , \22546 , \22547 , \22548 , \22549 , \22550 , \22551 , \22552 ,
         \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 , \22561 , \22562 ,
         \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 , \22571 , \22572 ,
         \22573 , \22574 , \22575 , \22576 , \22577 , \22578 , \22579 , \22580 , \22581 , \22582 ,
         \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 , \22591 , \22592 ,
         \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 , \22601 , \22602 ,
         \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 , \22611 , \22612 ,
         \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 , \22621 , \22622 ,
         \22623 , \22624 , \22625 , \22626 , \22627 , \22628 , \22629 , \22630 , \22631 , \22632 ,
         \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 , \22641 , \22642 ,
         \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 , \22651 , \22652 ,
         \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 , \22661 , \22662 ,
         \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 , \22671 , \22672 ,
         \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 , \22681 , \22682 ,
         \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 , \22691 , \22692 ,
         \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 , \22701 , \22702 ,
         \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 , \22711 , \22712 ,
         \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 , \22721 , \22722 ,
         \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 , \22731 , \22732 ,
         \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 , \22741 , \22742 ,
         \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 , \22751 , \22752 ,
         \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 , \22761 , \22762 ,
         \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 , \22771 , \22772 ,
         \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 , \22781 , \22782 ,
         \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 , \22791 , \22792 ,
         \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 , \22801 , \22802 ,
         \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 , \22811 , \22812 ,
         \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 , \22821 , \22822 ,
         \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 , \22831 , \22832 ,
         \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 , \22841 , \22842 ,
         \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 , \22851 , \22852 ,
         \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 , \22861 , \22862 ,
         \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 , \22871 , \22872 ,
         \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 , \22881 , \22882 ,
         \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 , \22891 , \22892 ,
         \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 , \22901 , \22902 ,
         \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 , \22911 , \22912 ,
         \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 , \22921 , \22922 ,
         \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 , \22931 , \22932 ,
         \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 , \22941 , \22942 ,
         \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 , \22951 , \22952 ,
         \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 , \22961 , \22962 ,
         \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 , \22971 , \22972 ,
         \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 , \22981 , \22982 ,
         \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 , \22991 , \22992 ,
         \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 , \23001 , \23002 ,
         \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 , \23011 , \23012 ,
         \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 , \23021 , \23022 ,
         \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 , \23031 , \23032 ,
         \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 , \23041 , \23042 ,
         \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 , \23051 , \23052 ,
         \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 , \23061 , \23062 ,
         \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 , \23071 , \23072 ,
         \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 , \23081 , \23082 ,
         \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 , \23091 , \23092 ,
         \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 , \23101 , \23102 ,
         \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 , \23111 , \23112 ,
         \23113 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 , \23121 , \23122 ,
         \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 , \23131 , \23132 ,
         \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 , \23141 , \23142 ,
         \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 , \23151 , \23152 ,
         \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 , \23161 , \23162 ,
         \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 , \23171 , \23172 ,
         \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 , \23181 , \23182 ,
         \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 , \23191 , \23192 ,
         \23193 , \23194 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 , \23201 , \23202 ,
         \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 , \23211 , \23212 ,
         \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 , \23220 , \23221 , \23222 ,
         \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 , \23231 , \23232 ,
         \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 , \23241 , \23242 ,
         \23243 , \23244 , \23245 , \23246 , \23247 , \23248 , \23249 , \23250 , \23251 , \23252 ,
         \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 , \23261 , \23262 ,
         \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 , \23271 , \23272 ,
         \23273 , \23274 , \23275 , \23276 , \23277 , \23278 , \23279 , \23280 , \23281 , \23282 ,
         \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 , \23291 , \23292 ,
         \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 , \23301 , \23302 ,
         \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 , \23311 , \23312 ,
         \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 , \23321 , \23322 ,
         \23323 , \23324 , \23325 , \23326 , \23327 , \23328 , \23329 , \23330 , \23331 , \23332 ,
         \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 , \23341 , \23342 ,
         \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 , \23351 , \23352 ,
         \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 , \23361 , \23362 ,
         \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 , \23371 , \23372 ,
         \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 , \23381 , \23382 ,
         \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 , \23391 , \23392 ,
         \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 , \23401 , \23402 ,
         \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 , \23411 , \23412 ,
         \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 , \23421 , \23422 ,
         \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 , \23431 , \23432 ,
         \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 , \23441 , \23442 ,
         \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 , \23451 , \23452 ,
         \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 , \23461 , \23462 ,
         \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 , \23471 , \23472 ,
         \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 , \23481 , \23482 ,
         \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 , \23491 , \23492 ,
         \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 , \23501 , \23502 ,
         \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 , \23511 , \23512 ,
         \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 , \23521 , \23522 ,
         \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 , \23531 , \23532 ,
         \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 , \23541 , \23542 ,
         \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 , \23551 , \23552 ,
         \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 , \23561 , \23562 ,
         \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 , \23571 , \23572 ,
         \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 , \23581 , \23582 ,
         \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 , \23591 , \23592 ,
         \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 , \23601 , \23602 ,
         \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 , \23611 , \23612 ,
         \23613 , \23614 , \23615 , \23616 , \23617 , \23618 , \23619 , \23620 , \23621 , \23622 ,
         \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 , \23631 , \23632 ,
         \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 , \23641 , \23642 ,
         \23643 , \23644 , \23645 , \23646 , \23647 , \23648 , \23649 , \23650 , \23651 , \23652 ,
         \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 , \23661 , \23662 ,
         \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 , \23671 , \23672 ,
         \23673 , \23674 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 , \23681 , \23682 ,
         \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 , \23691 , \23692 ,
         \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 , \23700 , \23701 , \23702 ,
         \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 , \23711 , \23712 ,
         \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 , \23721 , \23722 ,
         \23723 , \23724 , \23725 , \23726 , \23727 , \23728 , \23729 , \23730 , \23731 , \23732 ,
         \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 , \23741 , \23742 ,
         \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 , \23751 , \23752 ,
         \23753 , \23754 , \23755 , \23756 , \23757 , \23758 , \23759 , \23760 , \23761 , \23762 ,
         \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 , \23771 , \23772 ,
         \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 , \23781 , \23782 ,
         \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 , \23791 , \23792 ,
         \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 , \23801 , \23802 ,
         \23803 , \23804 , \23805 , \23806 , \23807 , \23808 , \23809 , \23810 , \23811 , \23812 ,
         \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 , \23821 , \23822 ,
         \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 , \23831 , \23832 ,
         \23833 , \23834 , \23835 , \23836 , \23837 , \23838 , \23839 , \23840 , \23841 , \23842 ,
         \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 , \23851 , \23852 ,
         \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 , \23861 , \23862 ,
         \23863 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 , \23871 , \23872 ,
         \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 , \23881 , \23882 ,
         \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 , \23891 , \23892 ,
         \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 , \23901 , \23902 ,
         \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 , \23911 , \23912 ,
         \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 , \23921 , \23922 ,
         \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 , \23931 , \23932 ,
         \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 , \23941 , \23942 ,
         \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 , \23951 , \23952 ,
         \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 , \23961 , \23962 ,
         \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 , \23971 , \23972 ,
         \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 , \23981 , \23982 ,
         \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 , \23991 , \23992 ,
         \23993 , \23994 , \23995 , \23996 , \23997 , \23998 , \23999 , \24000 , \24001 , \24002 ,
         \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 , \24011 , \24012 ,
         \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 , \24021 , \24022 ,
         \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 , \24031 , \24032 ,
         \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 , \24041 , \24042 ,
         \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 , \24051 , \24052 ,
         \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 , \24061 , \24062 ,
         \24063 , \24064 , \24065 , \24066 , \24067 , \24068 , \24069 , \24070 , \24071 , \24072 ,
         \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 , \24081 , \24082 ,
         \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 , \24091 , \24092 ,
         \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 , \24101 , \24102 ,
         \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 , \24111 , \24112 ,
         \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 , \24121 , \24122 ,
         \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 , \24131 , \24132 ,
         \24133 , \24134 , \24135 , \24136 , \24137 , \24138 , \24139 , \24140 , \24141 , \24142 ,
         \24143 , \24144 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 , \24151 , \24152 ,
         \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 , \24161 , \24162 ,
         \24163 , \24164 , \24165 , \24166 , \24167 , \24168 , \24169 , \24170 , \24171 , \24172 ,
         \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 , \24181 , \24182 ,
         \24183 , \24184 , \24185 , \24186 , \24187 , \24188 , \24189 , \24190 , \24191 , \24192 ,
         \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 , \24201 , \24202 ,
         \24203 , \24204 , \24205 , \24206 , \24207 , \24208 , \24209 , \24210 , \24211 , \24212 ,
         \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 , \24221 , \24222 ,
         \24223 , \24224 , \24225 , \24226 , \24227 , \24228 , \24229 , \24230 , \24231 , \24232 ,
         \24233 , \24234 , \24235 , \24236 , \24237 , \24238 , \24239 , \24240 , \24241 , \24242 ,
         \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 , \24251 , \24252 ,
         \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 , \24261 , \24262 ,
         \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 , \24271 , \24272 ,
         \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 , \24281 , \24282 ,
         \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 , \24291 , \24292 ,
         \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 , \24301 , \24302 ,
         \24303 , \24304 , \24305 , \24306 , \24307 , \24308 , \24309 , \24310 , \24311 , \24312 ,
         \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 , \24321 , \24322 ,
         \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 , \24331 , \24332 ,
         \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 , \24341 , \24342 ,
         \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 , \24351 , \24352 ,
         \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 , \24361 , \24362 ,
         \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 , \24370 , \24371 , \24372 ,
         \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 , \24381 , \24382 ,
         \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 , \24391 , \24392 ,
         \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 , \24401 , \24402 ,
         \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 , \24411 , \24412 ,
         \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 , \24421 , \24422 ,
         \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 , \24431 , \24432 ,
         \24433 , \24434 , \24435 , \24436 , \24437 , \24438 , \24439 , \24440 , \24441 , \24442 ,
         \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 , \24451 , \24452 ,
         \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 , \24461 , \24462 ,
         \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 , \24471 , \24472 ,
         \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 , \24481 , \24482 ,
         \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 , \24491 , \24492 ,
         \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 , \24501 , \24502 ,
         \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , \24509 , \24510 , \24511 , \24512 ,
         \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 , \24521 , \24522 ,
         \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 , \24531 , \24532 ,
         \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 , \24541 , \24542 ,
         \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 , \24551 , \24552 ,
         \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 , \24561 , \24562 ,
         \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 , \24571 , \24572 ,
         \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 , \24581 , \24582 ,
         \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 , \24591 , \24592 ,
         \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 , \24601 , \24602 ,
         \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 , \24611 , \24612 ,
         \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 , \24621 , \24622 ,
         \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 , \24631 , \24632 ,
         \24633 , \24634 , \24635 , \24636 , \24637 , \24638 , \24639 , \24640 , \24641 , \24642 ,
         \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 , \24651 , \24652 ,
         \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 , \24661 , \24662 ,
         \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 , \24671 , \24672 ,
         \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 , \24681 , \24682 ,
         \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 , \24691 , \24692 ,
         \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 , \24701 , \24702 ,
         \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 , \24711 , \24712 ,
         \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 , \24721 , \24722 ,
         \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 , \24731 , \24732 ,
         \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 , \24741 , \24742 ,
         \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 , \24751 , \24752 ,
         \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 , \24761 , \24762 ,
         \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 , \24771 , \24772 ,
         \24773 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 , \24781 , \24782 ,
         \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 , \24791 , \24792 ,
         \24793 , \24794 , \24795 , \24796 , \24797 , \24798 , \24799 , \24800 , \24801 , \24802 ,
         \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 , \24811 , \24812 ,
         \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 , \24821 , \24822 ,
         \24823 , \24824 , \24825 , \24826 , \24827 , \24828 , \24829 , \24830 , \24831 , \24832 ,
         \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 , \24841 , \24842 ,
         \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 , \24851 , \24852 ,
         \24853 , \24854 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 , \24861 , \24862 ,
         \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 , \24871 , \24872 ,
         \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 , \24880 , \24881 , \24882 ,
         \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 , \24891 , \24892 ,
         \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 , \24901 , \24902 ,
         \24903 , \24904 , \24905 , \24906 , \24907 , \24908 , \24909 , \24910 , \24911 , \24912 ,
         \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 , \24921 , \24922 ,
         \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 , \24931 , \24932 ,
         \24933 , \24934 , \24935 , \24936 , \24937 , \24938 , \24939 , \24940 , \24941 , \24942 ,
         \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 , \24951 , \24952 ,
         \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 , \24961 , \24962 ,
         \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 , \24971 , \24972 ,
         \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 , \24981 , \24982 ,
         \24983 , \24984 , \24985 , \24986 , \24987 , \24988 , \24989 , \24990 , \24991 , \24992 ,
         \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 , \25001 , \25002 ,
         \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 , \25011 , \25012 ,
         \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 , \25021 , \25022 ,
         \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 , \25031 , \25032 ,
         \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 , \25041 , \25042 ,
         \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 , \25051 , \25052 ,
         \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 , \25061 , \25062 ,
         \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 , \25071 , \25072 ,
         \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 , \25081 , \25082 ,
         \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 , \25091 , \25092 ,
         \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 , \25101 , \25102 ,
         \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 , \25111 , \25112 ,
         \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 , \25121 , \25122 ,
         \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 , \25131 , \25132 ,
         \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 , \25141 , \25142 ,
         \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 , \25151 , \25152 ,
         \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 , \25161 , \25162 ,
         \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 , \25171 , \25172 ,
         \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 , \25181 , \25182 ,
         \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 , \25191 , \25192 ,
         \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 , \25201 , \25202 ,
         \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 , \25211 , \25212 ,
         \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 , \25221 , \25222 ,
         \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 , \25231 , \25232 ,
         \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 , \25241 , \25242 ,
         \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 , \25251 , \25252 ,
         \25253 , \25254 , \25255 , \25256 , \25257 , \25258 , \25259 , \25260 , \25261 , \25262 ,
         \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 , \25271 , \25272 ,
         \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 , \25281 , \25282 ,
         \25283 , \25284 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 , \25291 , \25292 ,
         \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 , \25301 , \25302 ,
         \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 , \25310 , \25311 , \25312 ,
         \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 , \25321 , \25322 ,
         \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 , \25331 , \25332 ,
         \25333 , \25334 , \25335 , \25336 , \25337 , \25338 , \25339 , \25340 , \25341 , \25342 ,
         \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 , \25351 , \25352 ,
         \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 , \25361 , \25362 ,
         \25363 , \25364 , \25365 , \25366 , \25367 , \25368 , \25369 , \25370 , \25371 , \25372 ,
         \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 , \25381 , \25382 ,
         \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 , \25391 , \25392 ,
         \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 , \25401 , \25402 ,
         \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 , \25411 , \25412 ,
         \25413 , \25414 , \25415 , \25416 , \25417 , \25418 , \25419 , \25420 , \25421 , \25422 ,
         \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 , \25431 , \25432 ,
         \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 , \25441 , \25442 ,
         \25443 , \25444 , \25445 , \25446 , \25447 , \25448 , \25449 , \25450 , \25451 , \25452 ,
         \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 , \25461 , \25462 ,
         \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 , \25471 , \25472 ,
         \25473 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 , \25481 , \25482 ,
         \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 , \25491 , \25492 ,
         \25493 , \25494 , \25495 , \25496 , \25497 , \25498 , \25499 , \25500 , \25501 , \25502 ,
         \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 , \25511 , \25512 ,
         \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 , \25521 , \25522 ,
         \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 , \25531 , \25532 ,
         \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 , \25541 , \25542 ,
         \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 , \25551 , \25552 ,
         \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 , \25561 , \25562 ,
         \25563 , \25564 , \25565 , \25566 , \25567 , \25568 , \25569 , \25570 , \25571 , \25572 ,
         \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 , \25581 , \25582 ,
         \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 , \25591 , \25592 ,
         \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 , \25601 , \25602 ,
         \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 , \25611 , \25612 ,
         \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 , \25621 , \25622 ,
         \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 , \25631 , \25632 ,
         \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 , \25641 , \25642 ,
         \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 , \25651 , \25652 ,
         \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 , \25661 , \25662 ,
         \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 , \25671 , \25672 ,
         \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 , \25681 , \25682 ,
         \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 , \25691 , \25692 ,
         \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 , \25701 , \25702 ,
         \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 , \25711 , \25712 ,
         \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 , \25721 , \25722 ,
         \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 , \25731 , \25732 ,
         \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 , \25741 , \25742 ,
         \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 , \25751 , \25752 ,
         \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 , \25761 , \25762 ,
         \25763 , \25764 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 , \25771 , \25772 ,
         \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 , \25781 , \25782 ,
         \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 , \25790 , \25791 , \25792 ,
         \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 , \25801 , \25802 ,
         \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 , \25811 , \25812 ,
         \25813 , \25814 , \25815 , \25816 , \25817 , \25818 , \25819 , \25820 , \25821 , \25822 ,
         \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 , \25831 , \25832 ,
         \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 , \25841 , \25842 ,
         \25843 , \25844 , \25845 , \25846 , \25847 , \25848 , \25849 , \25850 , \25851 , \25852 ,
         \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 , \25861 , \25862 ,
         \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 , \25871 , \25872 ,
         \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 , \25881 , \25882 ,
         \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 , \25891 , \25892 ,
         \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 , \25901 , \25902 ,
         \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 , \25911 , \25912 ,
         \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 , \25921 , \25922 ,
         \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 , \25931 , \25932 ,
         \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 , \25941 , \25942 ,
         \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 , \25951 , \25952 ,
         \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 , \25961 , \25962 ,
         \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 , \25971 , \25972 ,
         \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 , \25981 , \25982 ,
         \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 , \25991 , \25992 ,
         \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 , \26001 , \26002 ,
         \26003 , \26004 , \26005 , \26006 , \26007 , \26008 , \26009 , \26010 , \26011 , \26012 ,
         \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 , \26021 , \26022 ,
         \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 , \26031 , \26032 ,
         \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 , \26041 , \26042 ,
         \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 , \26051 , \26052 ,
         \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 , \26061 , \26062 ,
         \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 , \26071 , \26072 ,
         \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 , \26081 , \26082 ,
         \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 , \26091 , \26092 ,
         \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 , \26101 , \26102 ,
         \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 , \26111 , \26112 ,
         \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 , \26121 , \26122 ,
         \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 , \26131 , \26132 ,
         \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 , \26141 , \26142 ,
         \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 , \26151 , \26152 ,
         \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 , \26161 , \26162 ,
         \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 , \26171 , \26172 ,
         \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 , \26181 , \26182 ,
         \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 , \26191 , \26192 ,
         \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 , \26201 , \26202 ,
         \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 , \26211 , \26212 ,
         \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 , \26221 , \26222 ,
         \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 , \26231 , \26232 ,
         \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 , \26241 , \26242 ,
         \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 , \26251 , \26252 ,
         \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 , \26261 , \26262 ,
         \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 , \26271 , \26272 ,
         \26273 , \26274 , \26275 , \26276 , \26277 , \26278 , \26279 , \26280 , \26281 , \26282 ,
         \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 , \26291 , \26292 ,
         \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 , \26301 , \26302 ,
         \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 , \26311 , \26312 ,
         \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 , \26321 , \26322 ,
         \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 , \26331 , \26332 ,
         \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 , \26341 , \26342 ,
         \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 , \26351 , \26352 ,
         \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 , \26361 , \26362 ,
         \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 , \26371 , \26372 ,
         \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 , \26381 , \26382 ,
         \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 , \26391 , \26392 ,
         \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 , \26401 , \26402 ,
         \26403 , \26404 , \26405 , \26406 , \26407 , \26408 , \26409 , \26410 , \26411 , \26412 ,
         \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 , \26421 , \26422 ,
         \26423 , \26424 , \26425 , \26426 , \26427 , \26428 , \26429 , \26430 , \26431 , \26432 ,
         \26433 , \26434 , \26435 , \26436 , \26437 , \26438 , \26439 , \26440 , \26441 , \26442 ,
         \26443 , \26444 , \26445 , \26446 , \26447 , \26448 , \26449 , \26450 , \26451 , \26452 ,
         \26453 , \26454 , \26455 , \26456 , \26457 , \26458 , \26459 , \26460 , \26461 , \26462 ,
         \26463 , \26464 , \26465 , \26466 , \26467 , \26468 , \26469 , \26470 , \26471 , \26472 ,
         \26473 , \26474 , \26475 , \26476 , \26477 , \26478 , \26479 , \26480 , \26481 , \26482 ,
         \26483 , \26484 , \26485 , \26486 , \26487 , \26488 , \26489 , \26490 , \26491 , \26492 ,
         \26493 , \26494 , \26495 , \26496 , \26497 , \26498 , \26499 , \26500 , \26501 , \26502 ,
         \26503 , \26504 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 , \26511 , \26512 ,
         \26513 , \26514 , \26515 , \26516 , \26517 , \26518 , \26519 , \26520 , \26521 , \26522 ,
         \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 , \26531 , \26532 ,
         \26533 , \26534 , \26535 , \26536 , \26537 , \26538 , \26539 , \26540 , \26541 , \26542 ,
         \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 , \26551 , \26552 ,
         \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 , \26561 , \26562 ,
         \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 , \26571 , \26572 ,
         \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 , \26581 , \26582 ,
         \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 , \26591 , \26592 ,
         \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 , \26601 , \26602 ,
         \26603 , \26604 , \26605 , \26606 , \26607 , \26608 , \26609 , \26610 , \26611 , \26612 ,
         \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 , \26621 , \26622 ,
         \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 , \26631 , \26632 ,
         \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 , \26641 , \26642 ,
         \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 , \26651 , \26652 ,
         \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 , \26661 , \26662 ,
         \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 , \26670 , \26671 , \26672 ,
         \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 , \26681 , \26682 ,
         \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 , \26691 , \26692 ,
         \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 , \26701 , \26702 ,
         \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 , \26711 , \26712 ,
         \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 , \26721 , \26722 ,
         \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 , \26731 , \26732 ,
         \26733 , \26734 , \26735 , \26736 , \26737 , \26738 , \26739 , \26740 , \26741 , \26742 ,
         \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 , \26751 , \26752 ,
         \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 , \26761 , \26762 ,
         \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 , \26771 , \26772 ,
         \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 , \26781 , \26782 ,
         \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 , \26791 , \26792 ,
         \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 , \26801 , \26802 ,
         \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 , \26811 , \26812 ,
         \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 , \26820 , \26821 , \26822 ,
         \26823 , \26824 , \26825 , \26826 , \26827 , \26828 , \26829 , \26830 , \26831 , \26832 ,
         \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 , \26841 , \26842 ,
         \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 , \26851 , \26852 ,
         \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 , \26861 , \26862 ,
         \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 , \26871 , \26872 ,
         \26873 , \26874 , \26875 , \26876 , \26877 , \26878 , \26879 , \26880 , \26881 , \26882 ,
         \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 , \26891 , \26892 ,
         \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 , \26901 , \26902 ,
         \26903 , \26904 , \26905 , \26906 , \26907 , \26908 , \26909 , \26910 , \26911 , \26912 ,
         \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 , \26921 , \26922 ,
         \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 , \26931 , \26932 ,
         \26933 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 , \26941 , \26942 ,
         \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 , \26951 , \26952 ,
         \26953 , \26954 , \26955 , \26956 , \26957 , \26958 , \26959 , \26960 , \26961 , \26962 ,
         \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 , \26971 , \26972 ,
         \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 , \26981 , \26982 ,
         \26983 , \26984 , \26985 , \26986 , \26987 , \26988 , \26989 , \26990 , \26991 , \26992 ,
         \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 , \27001 , \27002 ,
         \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 , \27011 , \27012 ,
         \27013 , \27014 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 , \27021 , \27022 ,
         \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 , \27031 , \27032 ,
         \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 , \27041 , \27042 ,
         \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 , \27051 , \27052 ,
         \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 , \27061 , \27062 ,
         \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 , \27071 , \27072 ,
         \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 , \27081 , \27082 ,
         \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 , \27091 , \27092 ,
         \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 , \27101 , \27102 ,
         \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 , \27111 , \27112 ,
         \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 , \27121 , \27122 ,
         \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 , \27131 , \27132 ,
         \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 , \27141 , \27142 ,
         \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 , \27151 , \27152 ,
         \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 , \27161 , \27162 ,
         \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 , \27171 , \27172 ,
         \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 , \27181 , \27182 ,
         \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 , \27191 , \27192 ,
         \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 , \27201 , \27202 ,
         \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 , \27211 , \27212 ,
         \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 , \27221 , \27222 ,
         \27223 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 , \27231 , \27232 ,
         \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 , \27241 , \27242 ,
         \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 , \27251 , \27252 ,
         \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 , \27261 , \27262 ,
         \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 , \27271 , \27272 ,
         \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 , \27281 , \27282 ,
         \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 , \27291 , \27292 ,
         \27293 , \27294 , \27295 , \27296 , \27297 , \27298 , \27299 , \27300 , \27301 , \27302 ,
         \27303 , \27304 , \27305 , \27306 , \27307 , \27308 , \27309 , \27310 , \27311 , \27312 ,
         \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 , \27321 , \27322 ,
         \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 , \27331 , \27332 ,
         \27333 , \27334 , \27335 , \27336 , \27337 , \27338 , \27339 , \27340 , \27341 , \27342 ,
         \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 , \27351 , \27352 ,
         \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 , \27361 , \27362 ,
         \27363 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 , \27371 , \27372 ,
         \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 , \27381 , \27382 ,
         \27383 , \27384 , \27385 , \27386 , \27387 , \27388 , \27389 , \27390 , \27391 , \27392 ,
         \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 , \27401 , \27402 ,
         \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 , \27411 , \27412 ,
         \27413 , \27414 , \27415 , \27416 , \27417 , \27418 , \27419 , \27420 , \27421 , \27422 ,
         \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 , \27431 , \27432 ,
         \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 , \27441 , \27442 ,
         \27443 , \27444 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 , \27451 , \27452 ,
         \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 , \27461 , \27462 ,
         \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 , \27470 , \27471 , \27472 ,
         \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 , \27481 , \27482 ,
         \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 , \27491 , \27492 ,
         \27493 , \27494 , \27495 , \27496 , \27497 , \27498 , \27499 , \27500 , \27501 , \27502 ,
         \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 , \27511 , \27512 ,
         \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 , \27521 , \27522 ,
         \27523 , \27524 , \27525 , \27526 , \27527 , \27528 , \27529 , \27530 , \27531 , \27532 ,
         \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 , \27541 , \27542 ,
         \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 , \27551 , \27552 ,
         \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 , \27561 , \27562 ,
         \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 , \27571 , \27572 ,
         \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 , \27581 , \27582 ,
         \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 , \27591 , \27592 ,
         \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 , \27601 , \27602 ,
         \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 , \27611 , \27612 ,
         \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 , \27621 , \27622 ,
         \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 , \27631 , \27632 ,
         \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 , \27641 , \27642 ,
         \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 , \27651 , \27652 ,
         \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 , \27661 , \27662 ,
         \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 , \27671 , \27672 ,
         \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 , \27681 , \27682 ,
         \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 , \27691 , \27692 ,
         \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 , \27701 , \27702 ,
         \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 , \27711 , \27712 ,
         \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 , \27721 , \27722 ,
         \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 , \27731 , \27732 ,
         \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 , \27741 , \27742 ,
         \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 , \27751 , \27752 ,
         \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 , \27761 , \27762 ,
         \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 , \27771 , \27772 ,
         \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 , \27781 , \27782 ,
         \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 , \27791 , \27792 ,
         \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 , \27801 , \27802 ,
         \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 , \27811 , \27812 ,
         \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 , \27821 , \27822 ,
         \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 , \27831 , \27832 ,
         \27833 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 , \27841 , \27842 ,
         \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 , \27851 , \27852 ,
         \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 , \27861 , \27862 ,
         \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 , \27871 , \27872 ,
         \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 , \27881 , \27882 ,
         \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 , \27891 , \27892 ,
         \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 , \27901 , \27902 ,
         \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 , \27911 , \27912 ,
         \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 , \27921 , \27922 ,
         \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 , \27931 , \27932 ,
         \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 , \27941 , \27942 ,
         \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 , \27951 , \27952 ,
         \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 , \27961 , \27962 ,
         \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 , \27970 , \27971 , \27972 ,
         \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 , \27981 , \27982 ,
         \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 , \27991 , \27992 ,
         \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 , \28001 , \28002 ,
         \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 , \28011 , \28012 ,
         \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 , \28021 , \28022 ,
         \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 , \28031 , \28032 ,
         \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 , \28041 , \28042 ,
         \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 , \28051 , \28052 ,
         \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 , \28061 , \28062 ,
         \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 , \28071 , \28072 ,
         \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 , \28081 , \28082 ,
         \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 , \28091 , \28092 ,
         \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 , \28101 , \28102 ,
         \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 , \28111 , \28112 ,
         \28113 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 , \28121 , \28122 ,
         \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 , \28131 , \28132 ,
         \28133 , \28134 , \28135 , \28136 , \28137 , \28138 , \28139 , \28140 , \28141 , \28142 ,
         \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 , \28151 , \28152 ,
         \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 , \28161 , \28162 ,
         \28163 , \28164 , \28165 , \28166 , \28167 , \28168 , \28169 , \28170 , \28171 , \28172 ,
         \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 , \28181 , \28182 ,
         \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 , \28191 , \28192 ,
         \28193 , \28194 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 , \28201 , \28202 ,
         \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 , \28211 , \28212 ,
         \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 , \28220 , \28221 , \28222 ,
         \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 , \28231 , \28232 ,
         \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 , \28241 , \28242 ,
         \28243 , \28244 , \28245 , \28246 , \28247 , \28248 , \28249 , \28250 , \28251 , \28252 ,
         \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 , \28261 , \28262 ,
         \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 , \28271 , \28272 ,
         \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 , \28281 , \28282 ,
         \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 , \28291 , \28292 ,
         \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 , \28301 , \28302 ,
         \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 , \28311 , \28312 ,
         \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 , \28321 , \28322 ,
         \28323 , \28324 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 , \28331 , \28332 ,
         \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 , \28341 , \28342 ,
         \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 , \28351 , \28352 ,
         \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 , \28361 , \28362 ,
         \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 , \28371 , \28372 ,
         \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 , \28381 , \28382 ,
         \28383 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 , \28391 , \28392 ,
         \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 , \28401 , \28402 ,
         \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 , \28411 , \28412 ,
         \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 , \28421 , \28422 ,
         \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 , \28431 , \28432 ,
         \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 , \28441 , \28442 ,
         \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 , \28451 , \28452 ,
         \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 , \28461 , \28462 ,
         \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 , \28471 , \28472 ,
         \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 , \28481 , \28482 ,
         \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 , \28491 , \28492 ,
         \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 , \28501 , \28502 ,
         \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 , \28511 , \28512 ,
         \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 , \28521 , \28522 ,
         \28523 , \28524 , \28525 , \28526 , \28527 , \28528 , \28529 , \28530 , \28531 , \28532 ,
         \28533 , \28534 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 , \28541 , \28542 ,
         \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 , \28551 , \28552 ,
         \28553 , \28554 , \28555 , \28556 , \28557 , \28558 , \28559 , \28560 , \28561 , \28562 ,
         \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 , \28571 , \28572 ,
         \28573 , \28574 , \28575 , \28576 , \28577 , \28578 , \28579 , \28580 , \28581 , \28582 ,
         \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 , \28591 , \28592 ,
         \28593 , \28594 , \28595 , \28596 , \28597 , \28598 , \28599 , \28600 , \28601 , \28602 ,
         \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 , \28611 , \28612 ,
         \28613 , \28614 , \28615 , \28616 , \28617 , \28618 , \28619 , \28620 , \28621 , \28622 ,
         \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 , \28631 , \28632 ,
         \28633 , \28634 , \28635 , \28636 , \28637 , \28638 , \28639 , \28640 , \28641 , \28642 ,
         \28643 , \28644 , \28645 , \28646 , \28647 , \28648 , \28649 , \28650 , \28651 , \28652 ,
         \28653 , \28654 , \28655 , \28656 , \28657 , \28658 , \28659 , \28660 , \28661 , \28662 ,
         \28663 , \28664 , \28665 , \28666 , \28667 , \28668 , \28669 , \28670 , \28671 , \28672 ,
         \28673 , \28674 , \28675 , \28676 , \28677 , \28678 , \28679 , \28680 , \28681 , \28682 ,
         \28683 , \28684 , \28685 , \28686 , \28687 , \28688 , \28689 , \28690 , \28691 , \28692 ,
         \28693 , \28694 , \28695 , \28696 , \28697 , \28698 , \28699 , \28700 , \28701 , \28702 ,
         \28703 , \28704 , \28705 , \28706 , \28707 , \28708 , \28709 , \28710 , \28711 , \28712 ,
         \28713 , \28714 , \28715 , \28716 , \28717 , \28718 , \28719 , \28720 , \28721 , \28722 ,
         \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 , \28731 , \28732 ,
         \28733 , \28734 , \28735 , \28736 , \28737 , \28738 , \28739 , \28740 , \28741 , \28742 ,
         \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 , \28751 , \28752 ,
         \28753 , \28754 , \28755 , \28756 , \28757 , \28758 , \28759 , \28760 , \28761 , \28762 ,
         \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , \28770 , \28771 , \28772 ,
         \28773 , \28774 , \28775 , \28776 , \28777 , \28778 , \28779 , \28780 , \28781 , \28782 ,
         \28783 , \28784 , \28785 , \28786 , \28787 , \28788 , \28789 , \28790 , \28791 , \28792 ,
         \28793 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 , \28801 , \28802 ,
         \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 , \28811 , \28812 ,
         \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 , \28821 , \28822 ,
         \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 , \28831 , \28832 ,
         \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 , \28841 , \28842 ,
         \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 , \28851 , \28852 ,
         \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 , \28861 , \28862 ,
         \28863 , \28864 , \28865 , \28866 , \28867 , \28868 , \28869 , \28870 , \28871 , \28872 ,
         \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 , \28881 , \28882 ,
         \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 , \28891 , \28892 ,
         \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 , \28901 , \28902 ,
         \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 , \28911 , \28912 ,
         \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 , \28921 , \28922 ,
         \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 , \28931 , \28932 ,
         \28933 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 , \28941 , \28942 ,
         \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 , \28951 , \28952 ,
         \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 , \28961 , \28962 ,
         \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 , \28971 , \28972 ,
         \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 , \28981 , \28982 ,
         \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 , \28991 , \28992 ,
         \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 , \29001 , \29002 ,
         \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 , \29011 , \29012 ,
         \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 , \29021 , \29022 ,
         \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 , \29031 , \29032 ,
         \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 , \29041 , \29042 ,
         \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 , \29051 , \29052 ,
         \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 , \29061 , \29062 ,
         \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 , \29071 , \29072 ,
         \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 , \29081 , \29082 ,
         \29083 , \29084 , \29085 , \29086 , \29087 , \29088 , \29089 , \29090 , \29091 , \29092 ,
         \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 , \29101 , \29102 ,
         \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 , \29111 , \29112 ,
         \29113 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 , \29121 , \29122 ,
         \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 , \29131 , \29132 ,
         \29133 , \29134 , \29135 , \29136 , \29137 , \29138 , \29139 , \29140 , \29141 , \29142 ,
         \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 , \29151 , \29152 ,
         \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 , \29161 , \29162 ,
         \29163 , \29164 , \29165 , \29166 , \29167 , \29168 , \29169 , \29170 , \29171 , \29172 ,
         \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 , \29181 , \29182 ,
         \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 , \29191 , \29192 ,
         \29193 , \29194 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 , \29201 , \29202 ,
         \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 , \29211 , \29212 ,
         \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 , \29220 , \29221 , \29222 ,
         \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 , \29231 , \29232 ,
         \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 , \29241 , \29242 ,
         \29243 , \29244 , \29245 , \29246 , \29247 , \29248 , \29249 , \29250 , \29251 , \29252 ,
         \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 , \29261 , \29262 ,
         \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 , \29271 , \29272 ,
         \29273 , \29274 , \29275 , \29276 , \29277 , \29278 , \29279 , \29280 , \29281 , \29282 ,
         \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 , \29291 , \29292 ,
         \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 , \29301 , \29302 ,
         \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 , \29311 , \29312 ,
         \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 , \29321 , \29322 ,
         \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 , \29331 , \29332 ,
         \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 , \29341 , \29342 ,
         \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 , \29351 , \29352 ,
         \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 , \29361 , \29362 ,
         \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 , \29371 , \29372 ,
         \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 , \29381 , \29382 ,
         \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 , \29391 , \29392 ,
         \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 , \29401 , \29402 ,
         \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 , \29411 , \29412 ,
         \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 , \29421 , \29422 ,
         \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 , \29431 , \29432 ,
         \29433 , \29434 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 , \29441 , \29442 ,
         \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 , \29451 , \29452 ,
         \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 , \29461 , \29462 ,
         \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 , \29471 , \29472 ,
         \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 , \29481 , \29482 ,
         \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 , \29491 , \29492 ,
         \29493 , \29494 , \29495 , \29496 , \29497 , \29498 , \29499 , \29500 , \29501 , \29502 ,
         \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 , \29511 , \29512 ,
         \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 , \29521 , \29522 ,
         \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 , \29531 , \29532 ,
         \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 , \29541 , \29542 ,
         \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 , \29551 , \29552 ,
         \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 , \29561 , \29562 ,
         \29563 , \29564 , \29565 , \29566 , \29567 , \29568 , \29569 , \29570 , \29571 , \29572 ,
         \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 , \29581 , \29582 ,
         \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 , \29591 , \29592 ,
         \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 , \29601 , \29602 ,
         \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 , \29611 , \29612 ,
         \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 , \29621 , \29622 ,
         \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 , \29631 , \29632 ,
         \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 , \29641 , \29642 ,
         \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 , \29651 , \29652 ,
         \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 , \29661 , \29662 ,
         \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 , \29671 , \29672 ,
         \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 , \29681 , \29682 ,
         \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 , \29691 , \29692 ,
         \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 , \29701 , \29702 ,
         \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 , \29711 , \29712 ,
         \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 , \29721 , \29722 ,
         \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 , \29731 , \29732 ,
         \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 , \29741 , \29742 ,
         \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 , \29751 , \29752 ,
         \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 , \29761 , \29762 ,
         \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 , \29771 , \29772 ,
         \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 , \29781 , \29782 ,
         \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 , \29791 , \29792 ,
         \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 , \29801 , \29802 ,
         \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 , \29811 , \29812 ,
         \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 , \29821 , \29822 ,
         \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 , \29831 , \29832 ,
         \29833 , \29834 , \29835 , \29836 , \29837 , \29838 , \29839 , \29840 , \29841 , \29842 ,
         \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 , \29851 , \29852 ,
         \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 , \29861 , \29862 ,
         \29863 , \29864 , \29865 , \29866 , \29867 , \29868 , \29869 , \29870 , \29871 , \29872 ,
         \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 , \29881 , \29882 ,
         \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 , \29891 , \29892 ,
         \29893 , \29894 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 , \29901 , \29902 ,
         \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 , \29911 , \29912 ,
         \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 , \29920 , \29921 , \29922 ,
         \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 , \29931 , \29932 ,
         \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 , \29941 , \29942 ,
         \29943 , \29944 , \29945 , \29946 , \29947 , \29948 , \29949 , \29950 , \29951 , \29952 ,
         \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 , \29961 , \29962 ,
         \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 , \29971 , \29972 ,
         \29973 , \29974 , \29975 , \29976 , \29977 , \29978 , \29979 , \29980 , \29981 , \29982 ,
         \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 , \29991 , \29992 ,
         \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 , \30001 , \30002 ,
         \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 , \30011 , \30012 ,
         \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 , \30021 , \30022 ,
         \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 , \30031 , \30032 ,
         \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 , \30041 , \30042 ,
         \30043 , \30044 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 , \30051 , \30052 ,
         \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 , \30061 , \30062 ,
         \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 , \30071 , \30072 ,
         \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 , \30081 , \30082 ,
         \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 , \30091 , \30092 ,
         \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 , \30101 , \30102 ,
         \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 , \30111 , \30112 ,
         \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 , \30121 , \30122 ,
         \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 , \30131 , \30132 ,
         \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 , \30141 , \30142 ,
         \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 , \30151 , \30152 ,
         \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 , \30161 , \30162 ,
         \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 , \30171 , \30172 ,
         \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 , \30181 , \30182 ,
         \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 , \30191 , \30192 ,
         \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 , \30201 , \30202 ,
         \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 , \30211 , \30212 ,
         \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 , \30221 , \30222 ,
         \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 , \30231 , \30232 ,
         \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 , \30241 , \30242 ,
         \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 , \30251 , \30252 ,
         \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 , \30261 , \30262 ,
         \30263 , \30264 , \30265 , \30266 , \30267 , \30268 , \30269 , \30270 , \30271 , \30272 ,
         \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 , \30281 , \30282 ,
         \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 , \30291 , \30292 ,
         \30293 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 , \30301 , \30302 ,
         \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 , \30311 , \30312 ,
         \30313 , \30314 , \30315 , \30316 , \30317 , \30318 , \30319 , \30320 , \30321 , \30322 ,
         \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 , \30331 , \30332 ,
         \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 , \30341 , \30342 ,
         \30343 , \30344 , \30345 , \30346 , \30347 , \30348 , \30349 , \30350 , \30351 , \30352 ,
         \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 , \30361 , \30362 ,
         \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 , \30371 , \30372 ,
         \30373 , \30374 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 , \30381 , \30382 ,
         \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 , \30391 , \30392 ,
         \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 , \30400 , \30401 , \30402 ,
         \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 , \30411 , \30412 ,
         \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 , \30421 , \30422 ,
         \30423 , \30424 , \30425 , \30426 , \30427 , \30428 , \30429 , \30430 , \30431 , \30432 ,
         \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 , \30441 , \30442 ,
         \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 , \30451 , \30452 ,
         \30453 , \30454 , \30455 , \30456 , \30457 , \30458 , \30459 , \30460 , \30461 , \30462 ,
         \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 , \30471 , \30472 ,
         \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 , \30481 , \30482 ,
         \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 , \30491 , \30492 ,
         \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 , \30501 , \30502 ,
         \30503 , \30504 , \30505 , \30506 , \30507 , \30508 , \30509 , \30510 , \30511 , \30512 ,
         \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 , \30521 , \30522 ,
         \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 , \30531 , \30532 ,
         \30533 , \30534 , \30535 , \30536 , \30537 , \30538 , \30539 , \30540 , \30541 , \30542 ,
         \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 , \30551 , \30552 ,
         \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 , \30561 , \30562 ,
         \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 , \30571 , \30572 ,
         \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 , \30581 , \30582 ,
         \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 , \30591 , \30592 ,
         \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 , \30601 , \30602 ,
         \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 , \30611 , \30612 ,
         \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 , \30621 , \30622 ,
         \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 , \30631 , \30632 ,
         \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 , \30641 , \30642 ,
         \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 , \30651 , \30652 ,
         \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 , \30661 , \30662 ,
         \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 , \30671 , \30672 ,
         \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 , \30681 , \30682 ,
         \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 , \30691 , \30692 ,
         \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 , \30701 , \30702 ,
         \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 , \30711 , \30712 ,
         \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 , \30721 , \30722 ,
         \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 , \30731 , \30732 ,
         \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 , \30741 , \30742 ,
         \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 , \30751 , \30752 ,
         \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 , \30761 , \30762 ,
         \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 , \30771 , \30772 ,
         \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 , \30781 , \30782 ,
         \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 , \30791 , \30792 ,
         \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 , \30801 , \30802 ,
         \30803 , \30804 , \30805 , \30806 , \30807 , \30808 , \30809 , \30810 , \30811 , \30812 ,
         \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 , \30821 , \30822 ,
         \30823 , \30824 , \30825 , \30826 , \30827 , \30828 , \30829 , \30830 , \30831 , \30832 ,
         \30833 , \30834 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 , \30841 , \30842 ,
         \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 , \30851 , \30852 ,
         \30853 , \30854 , \30855 , \30856 , \30857 , \30858 , \30859 , \30860 , \30861 , \30862 ,
         \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 , \30871 , \30872 ,
         \30873 , \30874 , \30875 , \30876 , \30877 , \30878 , \30879 , \30880 , \30881 , \30882 ,
         \30883 , \30884 , \30885 , \30886 , \30887 , \30888 , \30889 , \30890 , \30891 , \30892 ,
         \30893 , \30894 , \30895 , \30896 , \30897 , \30898 , \30899 , \30900 , \30901 , \30902 ,
         \30903 , \30904 , \30905 , \30906 , \30907 , \30908 , \30909 , \30910 , \30911 , \30912 ,
         \30913 , \30914 , \30915 , \30916 , \30917 , \30918 , \30919 , \30920 , \30921 , \30922 ,
         \30923 , \30924 , \30925 , \30926 , \30927 , \30928 , \30929 , \30930 , \30931 , \30932 ,
         \30933 , \30934 , \30935 , \30936 , \30937 , \30938 , \30939 , \30940 , \30941 , \30942 ,
         \30943 , \30944 , \30945 , \30946 , \30947 , \30948 , \30949 , \30950 , \30951 , \30952 ,
         \30953 , \30954 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 , \30961 , \30962 ,
         \30963 , \30964 , \30965 , \30966 , \30967 , \30968 , \30969 , \30970 , \30971 , \30972 ,
         \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 , \30981 , \30982 ,
         \30983 , \30984 , \30985 , \30986 , \30987 , \30988 , \30989 , \30990 , \30991 , \30992 ,
         \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 , \31001 , \31002 ,
         \31003 , \31004 , \31005 , \31006 , \31007 , \31008 , \31009 , \31010 , \31011 , \31012 ,
         \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 , \31021 , \31022 ,
         \31023 , \31024 , \31025 , \31026 , \31027 , \31028 , \31029 , \31030 , \31031 , \31032 ,
         \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 , \31041 , \31042 ,
         \31043 , \31044 , \31045 , \31046 , \31047 , \31048 , \31049 , \31050 , \31051 , \31052 ,
         \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 , \31061 , \31062 ,
         \31063 , \31064 , \31065 , \31066 , \31067 , \31068 , \31069 , \31070 , \31071 , \31072 ,
         \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 , \31081 , \31082 ,
         \31083 , \31084 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 , \31091 , \31092 ,
         \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 , \31101 , \31102 ,
         \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 , \31111 , \31112 ,
         \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 , \31121 , \31122 ,
         \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 , \31131 , \31132 ,
         \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 , \31141 , \31142 ,
         \31143 , \31144 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 , \31151 , \31152 ,
         \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 , \31161 , \31162 ,
         \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 , \31171 , \31172 ,
         \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 , \31181 , \31182 ,
         \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 , \31191 , \31192 ,
         \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 , \31201 , \31202 ,
         \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 , \31211 , \31212 ,
         \31213 , \31214 , \31215 , \31216 , \31217 , \31218 , \31219 , \31220 , \31221 , \31222 ,
         \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 , \31231 , \31232 ,
         \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 , \31241 , \31242 ,
         \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 , \31251 , \31252 ,
         \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 , \31261 , \31262 ,
         \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 , \31271 , \31272 ,
         \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 , \31281 , \31282 ,
         \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 , \31291 , \31292 ,
         \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 , \31301 , \31302 ,
         \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 , \31311 , \31312 ,
         \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 , \31321 , \31322 ,
         \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 , \31331 , \31332 ,
         \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 , \31341 , \31342 ,
         \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 , \31351 , \31352 ,
         \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 , \31361 , \31362 ,
         \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 , \31371 , \31372 ,
         \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 , \31381 , \31382 ,
         \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 , \31391 , \31392 ,
         \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 , \31401 , \31402 ,
         \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 , \31411 , \31412 ,
         \31413 , \31414 , \31415 , \31416 , \31417 , \31418 , \31419 , \31420 , \31421 , \31422 ,
         \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 , \31431 , \31432 ,
         \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 , \31441 , \31442 ,
         \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 , \31451 , \31452 ,
         \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 , \31461 , \31462 ,
         \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 , \31471 , \31472 ,
         \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 , \31481 , \31482 ,
         \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 , \31491 , \31492 ,
         \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 , \31501 , \31502 ,
         \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 , \31511 , \31512 ,
         \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 , \31521 , \31522 ,
         \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 , \31531 , \31532 ,
         \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 , \31541 , \31542 ,
         \31543 , \31544 , \31545 , \31546 , \31547 , \31548 , \31549 , \31550 , \31551 , \31552 ,
         \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 , \31561 , \31562 ,
         \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 , \31571 , \31572 ,
         \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 , \31581 , \31582 ,
         \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 , \31591 , \31592 ,
         \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 , \31601 , \31602 ,
         \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 , \31611 , \31612 ,
         \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 , \31621 , \31622 ,
         \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 , \31630 , \31631 , \31632 ,
         \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 , \31641 , \31642 ,
         \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 , \31651 , \31652 ,
         \31653 , \31654 , \31655 , \31656 , \31657 , \31658 , \31659 , \31660 , \31661 , \31662 ,
         \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 , \31671 , \31672 ,
         \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 , \31681 , \31682 ,
         \31683 , \31684 , \31685 , \31686 , \31687 , \31688 , \31689 , \31690 , \31691 , \31692 ,
         \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 , \31701 , \31702 ,
         \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 , \31711 , \31712 ,
         \31713 , \31714 , \31715 , \31716 , \31717 , \31718 , \31719 , \31720 , \31721 , \31722 ,
         \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 , \31731 , \31732 ,
         \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 , \31741 , \31742 ,
         \31743 , \31744 , \31745 , \31746 , \31747 , \31748 , \31749 , \31750 , \31751 , \31752 ,
         \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 , \31761 , \31762 ,
         \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 , \31771 , \31772 ,
         \31773 , \31774 , \31775 , \31776 , \31777 , \31778 , \31779 , \31780 , \31781 , \31782 ,
         \31783 , \31784 , \31785 , \31786 , \31787 , \31788 , \31789 , \31790 , \31791 , \31792 ,
         \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 , \31801 , \31802 ,
         \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 , \31811 , \31812 ,
         \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 , \31821 , \31822 ,
         \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 , \31831 , \31832 ,
         \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 , \31841 , \31842 ,
         \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 , \31851 , \31852 ,
         \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 , \31861 , \31862 ,
         \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 , \31871 , \31872 ,
         \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 , \31881 , \31882 ,
         \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 , \31891 , \31892 ,
         \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 , \31901 , \31902 ,
         \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 , \31911 , \31912 ,
         \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 , \31921 , \31922 ,
         \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 , \31931 , \31932 ,
         \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 , \31941 , \31942 ,
         \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 , \31951 , \31952 ,
         \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 , \31961 , \31962 ,
         \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 , \31971 , \31972 ,
         \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 , \31981 , \31982 ,
         \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 , \31991 , \31992 ,
         \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 , \32001 , \32002 ,
         \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 , \32011 , \32012 ,
         \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 , \32021 , \32022 ,
         \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 , \32031 , \32032 ,
         \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 , \32041 , \32042 ,
         \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 , \32051 , \32052 ,
         \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 , \32060 , \32061 , \32062 ,
         \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 , \32071 , \32072 ,
         \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 , \32081 , \32082 ,
         \32083 , \32084 , \32085 , \32086 , \32087 , \32088 , \32089 , \32090 , \32091 , \32092 ,
         \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 , \32101 , \32102 ,
         \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 , \32111 , \32112 ,
         \32113 , \32114 , \32115 , \32116 , \32117 , \32118 , \32119 , \32120 , \32121 , \32122 ,
         \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 , \32131 , \32132 ,
         \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 , \32141 , \32142 ,
         \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 , \32151 , \32152 ,
         \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 , \32161 , \32162 ,
         \32163 , \32164 , \32165 , \32166 , \32167 , \32168 , \32169 , \32170 , \32171 , \32172 ,
         \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 , \32181 , \32182 ,
         \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 , \32191 , \32192 ,
         \32193 , \32194 , \32195 , \32196 , \32197 , \32198 , \32199 , \32200 , \32201 , \32202 ,
         \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 , \32211 , \32212 ,
         \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 , \32221 , \32222 ,
         \32223 , \32224 , \32225 , \32226 , \32227 , \32228 , \32229 , \32230 , \32231 , \32232 ,
         \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 , \32241 , \32242 ,
         \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 , \32251 , \32252 ,
         \32253 , \32254 , \32255 , \32256 , \32257 , \32258 , \32259 , \32260 , \32261 , \32262 ,
         \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 , \32271 , \32272 ,
         \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 , \32281 , \32282 ,
         \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32289 , \32290 , \32291 , \32292 ,
         \32293 , \32294 , \32295 , \32296 , \32297 , \32298 , \32299 , \32300 , \32301 , \32302 ,
         \32303 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 , \32311 , \32312 ,
         \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 , \32320 , \32321 , \32322 ,
         \32323 , \32324 , \32325 , \32326 , \32327 , \32328 , \32329 , \32330 , \32331 , \32332 ,
         \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 , \32341 , \32342 ,
         \32343 , \32344 , \32345 , \32346 , \32347 , \32348 , \32349 , \32350 , \32351 , \32352 ,
         \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 , \32361 , \32362 ,
         \32363 , \32364 , \32365 , \32366 , \32367 , \32368 , \32369 , \32370 , \32371 , \32372 ,
         \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 , \32381 , \32382 ,
         \32383 , \32384 , \32385 , \32386 , \32387 , \32388 , \32389 , \32390 , \32391 , \32392 ,
         \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 , \32401 , \32402 ,
         \32403 , \32404 , \32405 , \32406 , \32407 , \32408 , \32409 , \32410 , \32411 , \32412 ,
         \32413 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 , \32421 , \32422 ,
         \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 , \32430 , \32431 , \32432 ,
         \32433 , \32434 , \32435 , \32436 , \32437 , \32438 , \32439 , \32440 , \32441 , \32442 ,
         \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 , \32451 , \32452 ,
         \32453 , \32454 , \32455 , \32456 , \32457 , \32458 , \32459 , \32460 , \32461 , \32462 ,
         \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 , \32471 , \32472 ,
         \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 , \32481 , \32482 ,
         \32483 , \32484 , \32485 , \32486 , \32487 , \32488 , \32489 , \32490 , \32491 , \32492 ,
         \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 , \32501 , \32502 ,
         \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 , \32511 , \32512 ,
         \32513 , \32514 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 , \32521 , \32522 ,
         \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 , \32531 , \32532 ,
         \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 , \32541 , \32542 ,
         \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 , \32551 , \32552 ,
         \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 , \32561 , \32562 ,
         \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 , \32571 , \32572 ,
         \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 , \32581 , \32582 ,
         \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 , \32591 , \32592 ,
         \32593 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 , \32601 , \32602 ,
         \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 , \32611 , \32612 ,
         \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 , \32621 , \32622 ,
         \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 , \32631 , \32632 ,
         \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 , \32641 , \32642 ,
         \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 , \32651 , \32652 ,
         \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 , \32661 , \32662 ,
         \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 , \32671 , \32672 ,
         \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 , \32681 , \32682 ,
         \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 , \32691 , \32692 ,
         \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 , \32701 , \32702 ,
         \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 , \32711 , \32712 ,
         \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 , \32721 , \32722 ,
         \32723 , \32724 , \32725 , \32726 , \32727 , \32728 , \32729 , \32730 , \32731 , \32732 ,
         \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 , \32741 , \32742 ,
         \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 , \32751 , \32752 ,
         \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 , \32761 , \32762 ,
         \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 , \32771 , \32772 ,
         \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 , \32781 , \32782 ,
         \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 , \32791 , \32792 ,
         \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 , \32801 , \32802 ,
         \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 , \32810 , \32811 , \32812 ,
         \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 , \32821 , \32822 ,
         \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 , \32831 , \32832 ,
         \32833 , \32834 , \32835 , \32836 , \32837 , \32838 , \32839 , \32840 , \32841 , \32842 ,
         \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 , \32851 , \32852 ,
         \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 , \32861 , \32862 ,
         \32863 , \32864 , \32865 , \32866 , \32867 , \32868 , \32869 , \32870 , \32871 , \32872 ,
         \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 , \32881 , \32882 ,
         \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 , \32891 , \32892 ,
         \32893 , \32894 , \32895 , \32896 , \32897 , \32898 , \32899 , \32900 , \32901 , \32902 ,
         \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 , \32911 , \32912 ,
         \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 , \32921 , \32922 ,
         \32923 , \32924 , \32925 , \32926 , \32927 , \32928 , \32929 , \32930 , \32931 , \32932 ,
         \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 , \32941 , \32942 ,
         \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 , \32951 , \32952 ,
         \32953 , \32954 , \32955 , \32956 , \32957 , \32958 , \32959 , \32960 , \32961 , \32962 ,
         \32963 , \32964 , \32965 , \32966 , \32967 , \32968 , \32969 , \32970 , \32971 , \32972 ,
         \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 , \32981 , \32982 ,
         \32983 , \32984 , \32985 , \32986 , \32987 , \32988 , \32989 , \32990 , \32991 , \32992 ,
         \32993 , \32994 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 , \33001 , \33002 ,
         \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 , \33011 , \33012 ,
         \33013 , \33014 , \33015 , \33016 , \33017 , \33018 , \33019 , \33020 , \33021 , \33022 ,
         \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 , \33031 , \33032 ,
         \33033 , \33034 , \33035 , \33036 , \33037 , \33038 , \33039 , \33040 , \33041 , \33042 ,
         \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 , \33051 , \33052 ,
         \33053 , \33054 , \33055 , \33056 , \33057 , \33058 , \33059 , \33060 , \33061 , \33062 ,
         \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 , \33071 , \33072 ,
         \33073 , \33074 , \33075 , \33076 , \33077 , \33078 , \33079 , \33080 , \33081 , \33082 ,
         \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 , \33091 , \33092 ,
         \33093 , \33094 , \33095 , \33096 , \33097 , \33098 , \33099 , \33100 , \33101 , \33102 ,
         \33103 , \33104 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 , \33111 , \33112 ,
         \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 , \33121 , \33122 ,
         \33123 , \33124 , \33125 , \33126 , \33127 , \33128 , \33129 , \33130 , \33131 , \33132 ,
         \33133 , \33134 , \33135 , \33136 , \33137 , \33138 , \33139 , \33140 , \33141 , \33142 ,
         \33143 , \33144 , \33145 , \33146 , \33147 , \33148 , \33149 , \33150 , \33151 , \33152 ,
         \33153 , \33154 , \33155 , \33156 , \33157 , \33158 , \33159 , \33160 , \33161 , \33162 ,
         \33163 , \33164 , \33165 , \33166 , \33167 , \33168 , \33169 , \33170 , \33171 , \33172 ,
         \33173 , \33174 , \33175 , \33176 , \33177 , \33178 , \33179 , \33180 , \33181 , \33182 ,
         \33183 , \33184 , \33185 , \33186 , \33187 , \33188 , \33189 , \33190 , \33191 , \33192 ,
         \33193 , \33194 , \33195 , \33196 , \33197 , \33198 , \33199 , \33200 , \33201 , \33202 ,
         \33203 , \33204 , \33205 , \33206 , \33207 , \33208 , \33209 , \33210 , \33211 , \33212 ,
         \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 , \33221 , \33222 ,
         \33223 , \33224 , \33225 , \33226 , \33227 , \33228 , \33229 , \33230 , \33231 , \33232 ,
         \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 , \33241 , \33242 ,
         \33243 , \33244 , \33245 , \33246 , \33247 , \33248 , \33249 , \33250 , \33251 , \33252 ,
         \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 , \33261 , \33262 ,
         \33263 , \33264 , \33265 , \33266 , \33267 , \33268 , \33269 , \33270 , \33271 , \33272 ,
         \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 , \33281 , \33282 ,
         \33283 , \33284 , \33285 , \33286 , \33287 , \33288 , \33289 , \33290 , \33291 , \33292 ,
         \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 , \33301 , \33302 ,
         \33303 , \33304 , \33305 , \33306 , \33307 , \33308 , \33309 , \33310 , \33311 , \33312 ,
         \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 , \33321 , \33322 ,
         \33323 , \33324 , \33325 , \33326 , \33327 , \33328 , \33329 , \33330 , \33331 , \33332 ,
         \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 , \33341 , \33342 ,
         \33343 , \33344 , \33345 , \33346 , \33347 , \33348 , \33349 , \33350 , \33351 , \33352 ,
         \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 , \33361 , \33362 ,
         \33363 , \33364 , \33365 , \33366 , \33367 , \33368 , \33369 , \33370 , \33371 , \33372 ,
         \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 , \33381 , \33382 ,
         \33383 , \33384 , \33385 , \33386 , \33387 , \33388 , \33389 , \33390 , \33391 , \33392 ,
         \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 , \33401 , \33402 ,
         \33403 , \33404 , \33405 , \33406 , \33407 , \33408 , \33409 , \33410 , \33411 , \33412 ,
         \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 , \33421 , \33422 ,
         \33423 , \33424 , \33425 , \33426 , \33427 , \33428 , \33429 , \33430 , \33431 , \33432 ,
         \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 , \33441 , \33442 ,
         \33443 , \33444 , \33445 , \33446 , \33447 , \33448 , \33449 , \33450 , \33451 , \33452 ,
         \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 , \33461 , \33462 ,
         \33463 , \33464 , \33465 , \33466 , \33467 , \33468 , \33469 , \33470 , \33471 , \33472 ,
         \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 , \33481 , \33482 ,
         \33483 , \33484 , \33485 , \33486 , \33487 , \33488 , \33489 , \33490 , \33491 , \33492 ,
         \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 , \33501 , \33502 ,
         \33503 , \33504 , \33505 , \33506 , \33507 , \33508 , \33509 , \33510 , \33511 , \33512 ,
         \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 , \33521 , \33522 ,
         \33523 , \33524 , \33525 , \33526 , \33527 , \33528 , \33529 , \33530 , \33531 , \33532 ,
         \33533 , \33534 , \33535 , \33536 , \33537 , \33538 , \33539 , \33540 , \33541 , \33542 ,
         \33543 , \33544 , \33545 , \33546 , \33547 , \33548 , \33549 , \33550 , \33551 , \33552 ,
         \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 , \33561 , \33562 ,
         \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 , \33571 , \33572 ,
         \33573 , \33574 , \33575 , \33576 , \33577 , \33578 , \33579 , \33580 , \33581 , \33582 ,
         \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 , \33591 , \33592 ,
         \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 , \33601 , \33602 ,
         \33603 , \33604 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 , \33611 , \33612 ,
         \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 , \33621 , \33622 ,
         \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 , \33630 , \33631 , \33632 ,
         \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 , \33641 , \33642 ,
         \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 , \33651 , \33652 ,
         \33653 , \33654 , \33655 , \33656 , \33657 , \33658 , \33659 , \33660 , \33661 , \33662 ,
         \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 , \33671 , \33672 ,
         \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 , \33681 , \33682 ,
         \33683 , \33684 , \33685 , \33686 , \33687 , \33688 , \33689 , \33690 , \33691 , \33692 ,
         \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 , \33701 , \33702 ,
         \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 , \33711 , \33712 ,
         \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 , \33721 , \33722 ,
         \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 , \33731 , \33732 ,
         \33733 , \33734 , \33735 , \33736 , \33737 , \33738 , \33739 , \33740 , \33741 , \33742 ,
         \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 , \33751 , \33752 ,
         \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 , \33761 , \33762 ,
         \33763 , \33764 , \33765 , \33766 , \33767 , \33768 , \33769 , \33770 , \33771 , \33772 ,
         \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 , \33781 , \33782 ,
         \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 , \33791 , \33792 ,
         \33793 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 , \33801 , \33802 ,
         \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 , \33811 , \33812 ,
         \33813 , \33814 , \33815 , \33816 , \33817 , \33818 , \33819 , \33820 , \33821 , \33822 ,
         \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 , \33831 , \33832 ,
         \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 , \33841 , \33842 ,
         \33843 , \33844 , \33845 , \33846 , \33847 , \33848 , \33849 , \33850 , \33851 , \33852 ,
         \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 , \33861 , \33862 ,
         \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 , \33871 , \33872 ,
         \33873 , \33874 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 , \33881 , \33882 ,
         \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 , \33891 , \33892 ,
         \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 , \33900 , \33901 , \33902 ,
         \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 , \33911 , \33912 ,
         \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 , \33921 , \33922 ,
         \33923 , \33924 , \33925 , \33926 , \33927 , \33928 , \33929 , \33930 , \33931 , \33932 ,
         \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 , \33941 , \33942 ,
         \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 , \33951 , \33952 ,
         \33953 , \33954 , \33955 , \33956 , \33957 , \33958 , \33959 , \33960 , \33961 , \33962 ,
         \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 , \33971 , \33972 ,
         \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 , \33981 , \33982 ,
         \33983 , \33984 , \33985 , \33986 , \33987 , \33988 , \33989 , \33990 , \33991 , \33992 ,
         \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 , \34001 , \34002 ,
         \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 , \34011 , \34012 ,
         \34013 , \34014 , \34015 , \34016 , \34017 , \34018 , \34019 , \34020 , \34021 , \34022 ,
         \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 , \34031 , \34032 ,
         \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 , \34041 , \34042 ,
         \34043 , \34044 , \34045 , \34046 , \34047 , \34048 , \34049 , \34050 , \34051 , \34052 ,
         \34053 , \34054 , \34055 , \34056 , \34057 , \34058 , \34059 , \34060 , \34061 , \34062 ,
         \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 , \34071 , \34072 ,
         \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 , \34081 , \34082 ,
         \34083 , \34084 , \34085 , \34086 , \34087 , \34088 , \34089 , \34090 , \34091 , \34092 ,
         \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 , \34101 , \34102 ,
         \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 , \34111 , \34112 ,
         \34113 , \34114 , \34115 , \34116 , \34117 , \34118 , \34119 , \34120 , \34121 , \34122 ,
         \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 , \34131 , \34132 ,
         \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 , \34141 , \34142 ,
         \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 , \34151 , \34152 ,
         \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 , \34161 , \34162 ,
         \34163 , \34164 , \34165 , \34166 , \34167 , \34168 , \34169 , \34170 , \34171 , \34172 ,
         \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 , \34181 , \34182 ,
         \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 , \34191 , \34192 ,
         \34193 , \34194 , \34195 , \34196 , \34197 , \34198 , \34199 , \34200 , \34201 , \34202 ,
         \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 , \34211 , \34212 ,
         \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 , \34221 , \34222 ,
         \34223 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 , \34231 , \34232 ,
         \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 , \34241 , \34242 ,
         \34243 , \34244 , \34245 , \34246 , \34247 , \34248 , \34249 , \34250 , \34251 , \34252 ,
         \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 , \34261 , \34262 ,
         \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 , \34271 , \34272 ,
         \34273 , \34274 , \34275 , \34276 , \34277 , \34278 , \34279 , \34280 , \34281 , \34282 ,
         \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 , \34291 , \34292 ,
         \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 , \34301 , \34302 ,
         \34303 , \34304 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 , \34311 , \34312 ,
         \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 , \34321 , \34322 ,
         \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 , \34330 , \34331 , \34332 ,
         \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 , \34341 , \34342 ,
         \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 , \34351 , \34352 ,
         \34353 , \34354 , \34355 , \34356 , \34357 , \34358 , \34359 , \34360 , \34361 , \34362 ,
         \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 , \34371 , \34372 ,
         \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 , \34381 , \34382 ,
         \34383 , \34384 , \34385 , \34386 , \34387 , \34388 , \34389 , \34390 , \34391 , \34392 ,
         \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 , \34401 , \34402 ,
         \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 , \34411 , \34412 ,
         \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 , \34421 , \34422 ,
         \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 , \34431 , \34432 ,
         \34433 , \34434 , \34435 , \34436 , \34437 , \34438 , \34439 , \34440 , \34441 , \34442 ,
         \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 , \34451 , \34452 ,
         \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 , \34461 , \34462 ,
         \34463 , \34464 , \34465 , \34466 , \34467 , \34468 , \34469 , \34470 , \34471 , \34472 ,
         \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 , \34481 , \34482 ,
         \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 , \34491 , \34492 ,
         \34493 , \34494 , \34495 , \34496 , \34497 , \34498 , \34499 , \34500 , \34501 , \34502 ,
         \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 , \34511 , \34512 ,
         \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 , \34521 , \34522 ,
         \34523 , \34524 , \34525 , \34526 , \34527 , \34528 , \34529 , \34530 , \34531 , \34532 ,
         \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 , \34541 , \34542 ,
         \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 , \34551 , \34552 ,
         \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34559 , \34560 , \34561 , \34562 ,
         \34563 , \34564 , \34565 , \34566 , \34567 , \34568 , \34569 , \34570 , \34571 , \34572 ,
         \34573 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 , \34581 , \34582 ,
         \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 , \34590 , \34591 , \34592 ,
         \34593 , \34594 , \34595 , \34596 , \34597 , \34598 , \34599 , \34600 , \34601 , \34602 ,
         \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 , \34611 , \34612 ,
         \34613 , \34614 , \34615 , \34616 , \34617 , \34618 , \34619 , \34620 , \34621 , \34622 ,
         \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 , \34631 , \34632 ,
         \34633 , \34634 , \34635 , \34636 , \34637 , \34638 , \34639 , \34640 , \34641 , \34642 ,
         \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 , \34651 , \34652 ,
         \34653 , \34654 , \34655 , \34656 , \34657 , \34658 , \34659 , \34660 , \34661 , \34662 ,
         \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 , \34671 , \34672 ,
         \34673 , \34674 , \34675 , \34676 , \34677 , \34678 , \34679 , \34680 , \34681 , \34682 ,
         \34683 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 , \34691 , \34692 ,
         \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 , \34700 , \34701 , \34702 ,
         \34703 , \34704 , \34705 , \34706 , \34707 , \34708 , \34709 , \34710 , \34711 , \34712 ,
         \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 , \34721 , \34722 ,
         \34723 , \34724 , \34725 , \34726 , \34727 , \34728 , \34729 , \34730 , \34731 , \34732 ,
         \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 , \34741 , \34742 ,
         \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 , \34751 , \34752 ,
         \34753 , \34754 , \34755 , \34756 , \34757 , \34758 , \34759 , \34760 , \34761 , \34762 ,
         \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 , \34771 , \34772 ,
         \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 , \34781 , \34782 ,
         \34783 , \34784 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 , \34791 , \34792 ,
         \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 , \34801 , \34802 ,
         \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 , \34810 , \34811 , \34812 ,
         \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 , \34821 , \34822 ,
         \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 , \34831 , \34832 ,
         \34833 , \34834 , \34835 , \34836 , \34837 , \34838 , \34839 , \34840 , \34841 , \34842 ,
         \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 , \34851 , \34852 ,
         \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 , \34861 , \34862 ,
         \34863 , \34864 , \34865 , \34866 , \34867 , \34868 , \34869 , \34870 , \34871 , \34872 ,
         \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 , \34881 , \34882 ,
         \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 , \34891 , \34892 ,
         \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 , \34901 , \34902 ,
         \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 , \34911 , \34912 ,
         \34913 , \34914 , \34915 , \34916 , \34917 , \34918 , \34919 , \34920 , \34921 , \34922 ,
         \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 , \34931 , \34932 ,
         \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 , \34941 , \34942 ,
         \34943 , \34944 , \34945 , \34946 , \34947 , \34948 , \34949 , \34950 , \34951 , \34952 ,
         \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 , \34961 , \34962 ,
         \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 , \34971 , \34972 ,
         \34973 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 , \34981 , \34982 ,
         \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 , \34991 , \34992 ,
         \34993 , \34994 , \34995 , \34996 , \34997 , \34998 , \34999 , \35000 , \35001 , \35002 ,
         \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 , \35011 , \35012 ,
         \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 , \35021 , \35022 ,
         \35023 , \35024 , \35025 , \35026 , \35027 , \35028 , \35029 , \35030 , \35031 , \35032 ,
         \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 , \35041 , \35042 ,
         \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 , \35051 , \35052 ,
         \35053 , \35054 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 , \35061 , \35062 ,
         \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 , \35071 , \35072 ,
         \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 , \35080 , \35081 , \35082 ,
         \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 , \35091 , \35092 ,
         \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 , \35101 , \35102 ,
         \35103 , \35104 , \35105 , \35106 , \35107 , \35108 , \35109 , \35110 , \35111 , \35112 ,
         \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 , \35121 , \35122 ,
         \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 , \35131 , \35132 ,
         \35133 , \35134 , \35135 , \35136 , \35137 , \35138 , \35139 , \35140 , \35141 , \35142 ,
         \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 , \35151 , \35152 ,
         \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 , \35161 , \35162 ,
         \35163 , \35164 , \35165 , \35166 , \35167 , \35168 , \35169 , \35170 , \35171 , \35172 ,
         \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 , \35181 , \35182 ,
         \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 , \35191 , \35192 ,
         \35193 , \35194 , \35195 , \35196 , \35197 , \35198 , \35199 , \35200 , \35201 , \35202 ,
         \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 , \35211 , \35212 ,
         \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 , \35221 , \35222 ,
         \35223 , \35224 , \35225 , \35226 , \35227 , \35228 , \35229 , \35230 , \35231 , \35232 ,
         \35233 , \35234 , \35235 , \35236 , \35237 , \35238 , \35239 , \35240 , \35241 , \35242 ,
         \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 , \35251 , \35252 ,
         \35253 , \35254 , \35255 , \35256 , \35257 , \35258 , \35259 , \35260 , \35261 , \35262 ,
         \35263 , \35264 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 , \35271 , \35272 ,
         \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 , \35281 , \35282 ,
         \35283 , \35284 , \35285 , \35286 , \35287 , \35288 , \35289 , \35290 , \35291 , \35292 ,
         \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 , \35301 , \35302 ,
         \35303 , \35304 , \35305 , \35306 , \35307 , \35308 , \35309 , \35310 , \35311 , \35312 ,
         \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 , \35321 , \35322 ,
         \35323 , \35324 , \35325 , \35326 , \35327 , \35328 , \35329 , \35330 , \35331 , \35332 ,
         \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 , \35341 , \35342 ,
         \35343 , \35344 , \35345 , \35346 , \35347 , \35348 , \35349 , \35350 , \35351 , \35352 ,
         \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 , \35361 , \35362 ,
         \35363 , \35364 , \35365 , \35366 , \35367 , \35368 , \35369 , \35370 , \35371 , \35372 ,
         \35373 , \35374 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 , \35381 , \35382 ,
         \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 , \35391 , \35392 ,
         \35393 , \35394 , \35395 , \35396 , \35397 , \35398 , \35399 , \35400 , \35401 , \35402 ,
         \35403 , \35404 , \35405 , \35406 , \35407 , \35408 , \35409 , \35410 , \35411 , \35412 ,
         \35413 , \35414 , \35415 , \35416 , \35417 , \35418 , \35419 , \35420 , \35421 , \35422 ,
         \35423 , \35424 , \35425 , \35426 , \35427 , \35428 , \35429 , \35430 , \35431 , \35432 ,
         \35433 , \35434 , \35435 , \35436 , \35437 , \35438 , \35439 , \35440 , \35441 , \35442 ,
         \35443 , \35444 , \35445 , \35446 , \35447 , \35448 , \35449 , \35450 , \35451 , \35452 ,
         \35453 , \35454 , \35455 , \35456 , \35457 , \35458 , \35459 , \35460 , \35461 , \35462 ,
         \35463 , \35464 , \35465 , \35466 , \35467 , \35468 , \35469 , \35470 , \35471 , \35472 ,
         \35473 , \35474 , \35475 , \35476 , \35477 , \35478 , \35479 , \35480 , \35481 , \35482 ,
         \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 , \35491 , \35492 ,
         \35493 , \35494 , \35495 , \35496 , \35497 , \35498 , \35499 , \35500 , \35501 , \35502 ,
         \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 , \35511 , \35512 ,
         \35513 , \35514 , \35515 , \35516 , \35517 , \35518 , \35519 , \35520 , \35521 , \35522 ,
         \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 , \35531 , \35532 ,
         \35533 , \35534 , \35535 , \35536 , \35537 , \35538 , \35539 , \35540 , \35541 , \35542 ,
         \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 , \35551 , \35552 ,
         \35553 , \35554 , \35555 , \35556 , \35557 , \35558 , \35559 , \35560 , \35561 , \35562 ,
         \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 , \35571 , \35572 ,
         \35573 , \35574 , \35575 , \35576 , \35577 , \35578 , \35579 , \35580 , \35581 , \35582 ,
         \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 , \35591 , \35592 ,
         \35593 , \35594 , \35595 , \35596 , \35597 , \35598 , \35599 , \35600 , \35601 , \35602 ,
         \35603 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 , \35611 , \35612 ,
         \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , \35619 , \35620 , \35621 , \35622 ,
         \35623 , \35624 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 , \35631 , \35632 ,
         \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , \35640 , \35641 , \35642 ,
         \35643 , \35644 , \35645 , \35646 , \35647 , \35648 , \35649 , \35650 , \35651 , \35652 ,
         \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 , \35661 , \35662 ,
         \35663 , \35664 , \35665 , \35666 , \35667 , \35668 , \35669 , \35670 , \35671 , \35672 ,
         \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 , \35681 , \35682 ,
         \35683 , \35684 , \35685 , \35686 , \35687 , \35688 , \35689 , \35690 , \35691 , \35692 ,
         \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 , \35701 , \35702 ,
         \35703 , \35704 , \35705 , \35706 , \35707 , \35708 , \35709 , \35710 , \35711 , \35712 ,
         \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 , \35721 , \35722 ,
         \35723 , \35724 , \35725 , \35726 , \35727 , \35728 , \35729 , \35730 , \35731 , \35732 ,
         \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 , \35741 , \35742 ,
         \35743 , \35744 , \35745 , \35746 , \35747 , \35748 , \35749 , \35750 , \35751 , \35752 ,
         \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 , \35761 , \35762 ,
         \35763 , \35764 , \35765 , \35766 , \35767 , \35768 , \35769 , \35770 , \35771 , \35772 ,
         \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 , \35781 , \35782 ,
         \35783 , \35784 , \35785 , \35786 , \35787 , \35788 , \35789 , \35790 , \35791 , \35792 ,
         \35793 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 , \35801 , \35802 ,
         \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , \35809 , \35810 , \35811 , \35812 ,
         \35813 , \35814 , \35815 , \35816 , \35817 , \35818 , \35819 , \35820 , \35821 , \35822 ,
         \35823 , \35824 , \35825 , \35826 , \35827 , \35828 , \35829 , \35830 , \35831 , \35832 ,
         \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 , \35841 , \35842 ,
         \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 , \35851 , \35852 ,
         \35853 , \35854 , \35855 , \35856 , \35857 , \35858 , \35859 , \35860 , \35861 , \35862 ,
         \35863 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 , \35871 , \35872 ,
         \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 , \35881 , \35882 ,
         \35883 , \35884 , \35885 , \35886 , \35887 , \35888 , \35889 , \35890 , \35891 , \35892 ,
         \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 , \35901 , \35902 ,
         \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 , \35911 , \35912 ,
         \35913 , \35914 , \35915 , \35916 , \35917 , \35918 , \35919 , \35920 , \35921 , \35922 ,
         \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 , \35931 , \35932 ,
         \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 , \35941 , \35942 ,
         \35943 , \35944 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 , \35951 , \35952 ,
         \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 , \35961 , \35962 ,
         \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 , \35970 , \35971 , \35972 ,
         \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 , \35981 , \35982 ,
         \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 , \35991 , \35992 ,
         \35993 , \35994 , \35995 , \35996 , \35997 , \35998 , \35999 , \36000 , \36001 , \36002 ,
         \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 , \36011 , \36012 ,
         \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 , \36021 , \36022 ,
         \36023 , \36024 , \36025 , \36026 , \36027 , \36028 , \36029 , \36030 , \36031 , \36032 ,
         \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 , \36041 , \36042 ,
         \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 , \36051 , \36052 ,
         \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 , \36061 , \36062 ,
         \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 , \36071 , \36072 ,
         \36073 , \36074 , \36075 , \36076 , \36077 , \36078 , \36079 , \36080 , \36081 , \36082 ,
         \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 , \36091 , \36092 ,
         \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 , \36101 , \36102 ,
         \36103 , \36104 , \36105 , \36106 , \36107 , \36108 , \36109 , \36110 , \36111 , \36112 ,
         \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 , \36121 , \36122 ,
         \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 , \36131 , \36132 ,
         \36133 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 , \36141 , \36142 ,
         \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 , \36151 , \36152 ,
         \36153 , \36154 , \36155 , \36156 , \36157 , \36158 , \36159 , \36160 , \36161 , \36162 ,
         \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 , \36171 , \36172 ,
         \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 , \36181 , \36182 ,
         \36183 , \36184 , \36185 , \36186 , \36187 , \36188 , \36189 , \36190 , \36191 , \36192 ,
         \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 , \36201 , \36202 ,
         \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 , \36211 , \36212 ,
         \36213 , \36214 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 , \36221 , \36222 ,
         \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 , \36231 , \36232 ,
         \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 , \36240 , \36241 , \36242 ,
         \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 , \36251 , \36252 ,
         \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 , \36261 , \36262 ,
         \36263 , \36264 , \36265 , \36266 , \36267 , \36268 , \36269 , \36270 , \36271 , \36272 ,
         \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 , \36281 , \36282 ,
         \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 , \36291 , \36292 ,
         \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 , \36301 , \36302 ,
         \36303 , \36304 , \36305 , \36306 , \36307 , \36308 , \36309 , \36310 , \36311 , \36312 ,
         \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 , \36321 , \36322 ,
         \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 , \36331 , \36332 ,
         \36333 , \36334 , \36335 , \36336 , \36337 , \36338 , \36339 , \36340 , \36341 , \36342 ,
         \36343 , \36344 , \36345 , \36346 , \36347 , \36348 , \36349 , \36350 , \36351 , \36352 ,
         \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 , \36361 , \36362 ,
         \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 , \36371 , \36372 ,
         \36373 , \36374 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 , \36381 , \36382 ,
         \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 , \36391 , \36392 ,
         \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 , \36400 , \36401 , \36402 ,
         \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 , \36411 , \36412 ,
         \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 , \36421 , \36422 ,
         \36423 , \36424 , \36425 , \36426 , \36427 , \36428 , \36429 , \36430 , \36431 , \36432 ,
         \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 , \36441 , \36442 ,
         \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 , \36451 , \36452 ,
         \36453 , \36454 , \36455 , \36456 , \36457 , \36458 , \36459 , \36460 , \36461 , \36462 ,
         \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 , \36471 , \36472 ,
         \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 , \36481 , \36482 ,
         \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 , \36491 , \36492 ,
         \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 , \36501 , \36502 ,
         \36503 , \36504 , \36505 , \36506 , \36507 , \36508 , \36509 , \36510 , \36511 , \36512 ,
         \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 , \36521 , \36522 ,
         \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 , \36531 , \36532 ,
         \36533 , \36534 , \36535 , \36536 , \36537 , \36538 , \36539 , \36540 , \36541 , \36542 ,
         \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 , \36551 , \36552 ,
         \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 , \36561 , \36562 ,
         \36563 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 , \36571 , \36572 ,
         \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 , \36581 , \36582 ,
         \36583 , \36584 , \36585 , \36586 , \36587 , \36588 , \36589 , \36590 , \36591 , \36592 ,
         \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 , \36601 , \36602 ,
         \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 , \36611 , \36612 ,
         \36613 , \36614 , \36615 , \36616 , \36617 , \36618 , \36619 , \36620 , \36621 , \36622 ,
         \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 , \36631 , \36632 ,
         \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 , \36641 , \36642 ,
         \36643 , \36644 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 , \36651 , \36652 ,
         \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 , \36661 , \36662 ,
         \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 , \36670 , \36671 , \36672 ,
         \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 , \36681 , \36682 ,
         \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 , \36691 , \36692 ,
         \36693 , \36694 , \36695 , \36696 , \36697 , \36698 , \36699 , \36700 , \36701 , \36702 ,
         \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 , \36711 , \36712 ,
         \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 , \36721 , \36722 ,
         \36723 , \36724 , \36725 , \36726 , \36727 , \36728 , \36729 , \36730 , \36731 , \36732 ,
         \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 , \36741 , \36742 ,
         \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 , \36751 , \36752 ,
         \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 , \36761 , \36762 ,
         \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 , \36771 , \36772 ,
         \36773 , \36774 , \36775 , \36776 , \36777 , \36778 , \36779 , \36780 , \36781 , \36782 ,
         \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 , \36791 , \36792 ,
         \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 , \36801 , \36802 ,
         \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 , \36811 , \36812 ,
         \36813 , \36814 , \36815 , \36816 , \36817 , \36818 , \36819 , \36820 , \36821 , \36822 ,
         \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 , \36831 , \36832 ,
         \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 , \36841 , \36842 ,
         \36843 , \36844 , \36845 , \36846 , \36847 , \36848 , \36849 , \36850 , \36851 , \36852 ,
         \36853 , \36854 , \36855 , \36856 , \36857 , \36858 , \36859 , \36860 , \36861 , \36862 ,
         \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 , \36871 , \36872 ,
         \36873 , \36874 , \36875 , \36876 , \36877 , \36878 , \36879 , \36880 , \36881 , \36882 ,
         \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 , \36891 , \36892 ,
         \36893 , \36894 , \36895 , \36896 , \36897 , \36898 , \36899 , \36900 , \36901 , \36902 ,
         \36903 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 , \36911 , \36912 ,
         \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 , \36920 , \36921 , \36922 ,
         \36923 , \36924 , \36925 , \36926 , \36927 , \36928 , \36929 , \36930 , \36931 , \36932 ,
         \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 , \36941 , \36942 ,
         \36943 , \36944 , \36945 , \36946 , \36947 , \36948 , \36949 , \36950 , \36951 , \36952 ,
         \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 , \36961 , \36962 ,
         \36963 , \36964 , \36965 , \36966 , \36967 , \36968 , \36969 , \36970 , \36971 , \36972 ,
         \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 , \36981 , \36982 ,
         \36983 , \36984 , \36985 , \36986 , \36987 , \36988 , \36989 , \36990 , \36991 , \36992 ,
         \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 , \37001 , \37002 ,
         \37003 , \37004 , \37005 , \37006 , \37007 , \37008 , \37009 , \37010 , \37011 , \37012 ,
         \37013 , \37014 , \37015 , \37016 , \37017 , \37018 , \37019 , \37020 , \37021 , \37022 ,
         \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 , \37031 , \37032 ,
         \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 , \37041 , \37042 ,
         \37043 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 , \37051 , \37052 ,
         \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 , \37061 , \37062 ,
         \37063 , \37064 , \37065 , \37066 , \37067 , \37068 , \37069 , \37070 , \37071 , \37072 ,
         \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 , \37081 , \37082 ,
         \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 , \37091 , \37092 ,
         \37093 , \37094 , \37095 , \37096 , \37097 , \37098 , \37099 , \37100 , \37101 , \37102 ,
         \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 , \37111 , \37112 ,
         \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 , \37121 , \37122 ,
         \37123 , \37124 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 , \37131 , \37132 ,
         \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 , \37141 , \37142 ,
         \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 , \37150 , \37151 , \37152 ,
         \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 , \37161 , \37162 ,
         \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 , \37171 , \37172 ,
         \37173 , \37174 , \37175 , \37176 , \37177 , \37178 , \37179 , \37180 , \37181 , \37182 ,
         \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 , \37191 , \37192 ,
         \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 , \37201 , \37202 ,
         \37203 , \37204 , \37205 , \37206 , \37207 , \37208 , \37209 , \37210 , \37211 , \37212 ,
         \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 , \37221 , \37222 ,
         \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 , \37231 , \37232 ,
         \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 , \37241 , \37242 ,
         \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 , \37251 , \37252 ,
         \37253 , \37254 , \37255 , \37256 , \37257 , \37258 , \37259 , \37260 , \37261 , \37262 ,
         \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 , \37271 , \37272 ,
         \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 , \37281 , \37282 ,
         \37283 , \37284 , \37285 , \37286 , \37287 , \37288 , \37289 , \37290 , \37291 , \37292 ,
         \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 , \37301 , \37302 ,
         \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 , \37311 , \37312 ,
         \37313 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 , \37321 , \37322 ,
         \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 , \37331 , \37332 ,
         \37333 , \37334 , \37335 , \37336 , \37337 , \37338 , \37339 , \37340 , \37341 , \37342 ,
         \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 , \37351 , \37352 ,
         \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 , \37361 , \37362 ,
         \37363 , \37364 , \37365 , \37366 , \37367 , \37368 , \37369 , \37370 , \37371 , \37372 ,
         \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 , \37381 , \37382 ,
         \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 , \37391 , \37392 ,
         \37393 , \37394 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 , \37401 , \37402 ,
         \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 , \37411 , \37412 ,
         \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 , \37420 , \37421 , \37422 ,
         \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 , \37431 , \37432 ,
         \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 , \37441 , \37442 ,
         \37443 , \37444 , \37445 , \37446 , \37447 , \37448 , \37449 , \37450 , \37451 , \37452 ,
         \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 , \37461 , \37462 ,
         \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 , \37471 , \37472 ,
         \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 , \37481 , \37482 ,
         \37483 , \37484 , \37485 , \37486 , \37487 , \37488 , \37489 , \37490 , \37491 , \37492 ,
         \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 , \37501 , \37502 ,
         \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 , \37511 , \37512 ,
         \37513 , \37514 , \37515 , \37516 , \37517 , \37518 , \37519 , \37520 , \37521 , \37522 ,
         \37523 , \37524 , \37525 , \37526 , \37527 , \37528 , \37529 , \37530 , \37531 , \37532 ,
         \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 , \37541 , \37542 ,
         \37543 , \37544 , \37545 , \37546 , \37547 , \37548 , \37549 , \37550 , \37551 , \37552 ,
         \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 , \37561 , \37562 ,
         \37563 , \37564 , \37565 , \37566 , \37567 , \37568 , \37569 , \37570 , \37571 , \37572 ,
         \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 , \37581 , \37582 ,
         \37583 , \37584 , \37585 , \37586 , \37587 , \37588 , \37589 , \37590 , \37591 , \37592 ,
         \37593 , \37594 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 , \37601 , \37602 ,
         \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 , \37611 , \37612 ,
         \37613 , \37614 , \37615 , \37616 , \37617 , \37618 , \37619 , \37620 , \37621 , \37622 ,
         \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 , \37631 , \37632 ,
         \37633 , \37634 , \37635 , \37636 , \37637 , \37638 , \37639 , \37640 , \37641 , \37642 ,
         \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 , \37651 , \37652 ,
         \37653 , \37654 , \37655 , \37656 , \37657 , \37658 , \37659 , \37660 , \37661 , \37662 ,
         \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 , \37671 , \37672 ,
         \37673 , \37674 , \37675 , \37676 , \37677 , \37678 , \37679 , \37680 , \37681 , \37682 ,
         \37683 , \37684 , \37685 , \37686 , \37687 , \37688 , \37689 , \37690 , \37691 , \37692 ,
         \37693 , \37694 , \37695 , \37696 , \37697 , \37698 , \37699 , \37700 , \37701 , \37702 ,
         \37703 , \37704 , \37705 , \37706 , \37707 , \37708 , \37709 , \37710 , \37711 , \37712 ,
         \37713 , \37714 , \37715 , \37716 , \37717 , \37718 , \37719 , \37720 , \37721 , \37722 ,
         \37723 , \37724 , \37725 , \37726 , \37727 , \37728 , \37729 , \37730 , \37731 , \37732 ,
         \37733 , \37734 , \37735 , \37736 , \37737 , \37738 , \37739 , \37740 , \37741 , \37742 ,
         \37743 , \37744 , \37745 , \37746 , \37747 , \37748 , \37749 , \37750 , \37751 , \37752 ,
         \37753 , \37754 , \37755 , \37756 , \37757 , \37758 , \37759 , \37760 , \37761 , \37762 ,
         \37763 , \37764 , \37765 , \37766 , \37767 , \37768 , \37769 , \37770 , \37771 , \37772 ,
         \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 , \37781 , \37782 ,
         \37783 , \37784 , \37785 , \37786 , \37787 , \37788 , \37789 , \37790 , \37791 , \37792 ,
         \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 , \37801 , \37802 ,
         \37803 , \37804 , \37805 , \37806 , \37807 , \37808 , \37809 , \37810 , \37811 , \37812 ,
         \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 , \37821 , \37822 ,
         \37823 , \37824 , \37825 , \37826 , \37827 , \37828 , \37829 , \37830 , \37831 , \37832 ,
         \37833 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 , \37841 , \37842 ,
         \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 , \37850 , \37851 , \37852 ,
         \37853 , \37854 , \37855 , \37856 , \37857 , \37858 , \37859 , \37860 , \37861 , \37862 ,
         \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 , \37871 , \37872 ,
         \37873 , \37874 , \37875 , \37876 , \37877 , \37878 , \37879 , \37880 , \37881 , \37882 ,
         \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 , \37891 , \37892 ,
         \37893 , \37894 , \37895 , \37896 , \37897 , \37898 , \37899 , \37900 , \37901 , \37902 ,
         \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 , \37911 , \37912 ,
         \37913 , \37914 , \37915 , \37916 , \37917 , \37918 , \37919 , \37920 , \37921 , \37922 ,
         \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 , \37931 , \37932 ,
         \37933 , \37934 , \37935 , \37936 , \37937 , \37938 , \37939 , \37940 , \37941 , \37942 ,
         \37943 , \37944 , \37945 , \37946 , \37947 , \37948 , \37949 , \37950 , \37951 , \37952 ,
         \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 , \37961 , \37962 ,
         \37963 , \37964 , \37965 , \37966 , \37967 , \37968 , \37969 , \37970 , \37971 , \37972 ,
         \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 , \37981 , \37982 ,
         \37983 , \37984 , \37985 , \37986 , \37987 , \37988 , \37989 , \37990 , \37991 , \37992 ,
         \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 , \38001 , \38002 ,
         \38003 , \38004 , \38005 , \38006 , \38007 , \38008 , \38009 , \38010 , \38011 , \38012 ,
         \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 , \38021 , \38022 ,
         \38023 , \38024 , \38025 , \38026 , \38027 , \38028 , \38029 , \38030 , \38031 , \38032 ,
         \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 , \38041 , \38042 ,
         \38043 , \38044 , \38045 , \38046 , \38047 , \38048 , \38049 , \38050 , \38051 , \38052 ,
         \38053 , \38054 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 , \38061 , \38062 ,
         \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 , \38071 , \38072 ,
         \38073 , \38074 , \38075 , \38076 , \38077 , \38078 , \38079 , \38080 , \38081 , \38082 ,
         \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 , \38091 , \38092 ,
         \38093 , \38094 , \38095 , \38096 , \38097 , \38098 , \38099 , \38100 , \38101 , \38102 ,
         \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 , \38111 , \38112 ,
         \38113 , \38114 , \38115 , \38116 , \38117 , \38118 , \38119 , \38120 , \38121 , \38122 ,
         \38123 , \38124 , \38125 , \38126 , \38127 , \38128 , \38129 , \38130 , \38131 , \38132 ,
         \38133 , \38134 , \38135 , \38136 , \38137 , \38138 , \38139 , \38140 , \38141 , \38142 ,
         \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 , \38151 , \38152 ,
         \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 , \38161 , \38162 ,
         \38163 , \38164 , \38165 , \38166 , \38167 , \38168 , \38169 , \38170 , \38171 , \38172 ,
         \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 , \38181 , \38182 ,
         \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 , \38191 , \38192 ,
         \38193 , \38194 , \38195 , \38196 , \38197 , \38198 , \38199 , \38200 , \38201 , \38202 ,
         \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 , \38211 , \38212 ,
         \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 , \38221 , \38222 ,
         \38223 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 , \38231 , \38232 ,
         \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 , \38241 , \38242 ,
         \38243 , \38244 , \38245 , \38246 , \38247 , \38248 , \38249 , \38250 , \38251 , \38252 ,
         \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 , \38261 , \38262 ,
         \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 , \38271 , \38272 ,
         \38273 , \38274 , \38275 , \38276 , \38277 , \38278 , \38279 , \38280 , \38281 , \38282 ,
         \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 , \38291 , \38292 ,
         \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 , \38301 , \38302 ,
         \38303 , \38304 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 , \38311 , \38312 ,
         \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 , \38321 , \38322 ,
         \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 , \38330 , \38331 , \38332 ,
         \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 , \38341 , \38342 ,
         \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 , \38351 , \38352 ,
         \38353 , \38354 , \38355 , \38356 , \38357 , \38358 , \38359 , \38360 , \38361 , \38362 ,
         \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 , \38371 , \38372 ,
         \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 , \38381 , \38382 ,
         \38383 , \38384 , \38385 , \38386 , \38387 , \38388 , \38389 , \38390 , \38391 , \38392 ,
         \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 , \38401 , \38402 ,
         \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 , \38411 , \38412 ,
         \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 , \38421 , \38422 ,
         \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 , \38431 , \38432 ,
         \38433 , \38434 , \38435 , \38436 , \38437 , \38438 , \38439 , \38440 , \38441 , \38442 ,
         \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 , \38451 , \38452 ,
         \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 , \38461 , \38462 ,
         \38463 , \38464 , \38465 , \38466 , \38467 , \38468 , \38469 , \38470 , \38471 , \38472 ,
         \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 , \38481 , \38482 ,
         \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 , \38491 , \38492 ,
         \38493 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 , \38501 , \38502 ,
         \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 , \38511 , \38512 ,
         \38513 , \38514 , \38515 , \38516 , \38517 , \38518 , \38519 , \38520 , \38521 , \38522 ,
         \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 , \38531 , \38532 ,
         \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 , \38541 , \38542 ,
         \38543 , \38544 , \38545 , \38546 , \38547 , \38548 , \38549 , \38550 , \38551 , \38552 ,
         \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 , \38561 , \38562 ,
         \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 , \38571 , \38572 ,
         \38573 , \38574 , \38575 , \38576 , \38577 , \38578 , \38579 , \38580 , \38581 , \38582 ,
         \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 , \38591 , \38592 ,
         \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 , \38601 , \38602 ,
         \38603 , \38604 , \38605 , \38606 , \38607 , \38608 , \38609 , \38610 , \38611 , \38612 ,
         \38613 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 , \38621 , \38622 ,
         \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 , \38631 , \38632 ,
         \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38640 , \38641 , \38642 ,
         \38643 , \38644 , \38645 , \38646 , \38647 , \38648 , \38649 , \38650 , \38651 , \38652 ,
         \38653 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 , \38661 , \38662 ,
         \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 , \38671 , \38672 ,
         \38673 , \38674 , \38675 , \38676 , \38677 , \38678 , \38679 , \38680 , \38681 , \38682 ,
         \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 , \38691 , \38692 ,
         \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 , \38701 , \38702 ,
         \38703 , \38704 , \38705 , \38706 , \38707 , \38708 , \38709 , \38710 , \38711 , \38712 ,
         \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 , \38721 , \38722 ,
         \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 , \38731 , \38732 ,
         \38733 , \38734 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 , \38741 , \38742 ,
         \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 , \38751 , \38752 ,
         \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 , \38760 , \38761 , \38762 ,
         \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 , \38771 , \38772 ,
         \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 , \38781 , \38782 ,
         \38783 , \38784 , \38785 , \38786 , \38787 , \38788 , \38789 , \38790 , \38791 , \38792 ,
         \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 , \38801 , \38802 ,
         \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 , \38811 , \38812 ,
         \38813 , \38814 , \38815 , \38816 , \38817 , \38818 , \38819 , \38820 , \38821 , \38822 ,
         \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 , \38831 , \38832 ,
         \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 , \38841 , \38842 ,
         \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 , \38851 , \38852 ,
         \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 , \38861 , \38862 ,
         \38863 , \38864 , \38865 , \38866 , \38867 , \38868 , \38869 , \38870 , \38871 , \38872 ,
         \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 , \38881 , \38882 ,
         \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 , \38891 , \38892 ,
         \38893 , \38894 , \38895 , \38896 , \38897 , \38898 , \38899 , \38900 , \38901 , \38902 ,
         \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 , \38911 , \38912 ,
         \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 , \38921 , \38922 ,
         \38923 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 , \38931 , \38932 ,
         \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 , \38941 , \38942 ,
         \38943 , \38944 , \38945 , \38946 , \38947 , \38948 , \38949 , \38950 , \38951 , \38952 ,
         \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 , \38961 , \38962 ,
         \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 , \38971 , \38972 ,
         \38973 , \38974 , \38975 , \38976 , \38977 , \38978 , \38979 , \38980 , \38981 , \38982 ,
         \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 , \38991 , \38992 ,
         \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 , \39001 , \39002 ,
         \39003 , \39004 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 , \39011 , \39012 ,
         \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 , \39021 , \39022 ,
         \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 , \39030 , \39031 , \39032 ,
         \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 , \39041 , \39042 ,
         \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 , \39051 , \39052 ,
         \39053 , \39054 , \39055 , \39056 , \39057 , \39058 , \39059 , \39060 , \39061 , \39062 ,
         \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 , \39071 , \39072 ,
         \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 , \39081 , \39082 ,
         \39083 , \39084 , \39085 , \39086 , \39087 , \39088 , \39089 , \39090 , \39091 , \39092 ,
         \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 , \39101 , \39102 ,
         \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 , \39111 , \39112 ,
         \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 , \39120 , \39121 , \39122 ,
         \39123 , \39124 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 , \39131 , \39132 ,
         \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 , \39141 , \39142 ,
         \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 , \39151 , \39152 ,
         \39153 , \39154 , \39155 , \39156 , \39157 , \39158 , \39159 , \39160 , \39161 , \39162 ,
         \39163 , \39164 , \39165 , \39166 , \39167 , \39168 , \39169 , \39170 , \39171 , \39172 ,
         \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 , \39181 , \39182 ,
         \39183 , \39184 , \39185 , \39186 , \39187 , \39188 , \39189 , \39190 , \39191 , \39192 ,
         \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 , \39201 , \39202 ,
         \39203 , \39204 , \39205 , \39206 , \39207 , \39208 , \39209 , \39210 , \39211 , \39212 ,
         \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 , \39221 , \39222 ,
         \39223 , \39224 , \39225 , \39226 , \39227 , \39228 , \39229 , \39230 , \39231 , \39232 ,
         \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 , \39241 , \39242 ,
         \39243 , \39244 , \39245 , \39246 , \39247 , \39248 , \39249 , \39250 , \39251 , \39252 ,
         \39253 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 , \39261 , \39262 ,
         \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 , \39270 , \39271 , \39272 ,
         \39273 , \39274 , \39275 , \39276 , \39277 , \39278 , \39279 , \39280 , \39281 , \39282 ,
         \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 , \39291 , \39292 ,
         \39293 , \39294 , \39295 , \39296 , \39297 , \39298 , \39299 , \39300 , \39301 , \39302 ,
         \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 , \39311 , \39312 ,
         \39313 , \39314 , \39315 , \39316 , \39317 , \39318 , \39319 , \39320 , \39321 , \39322 ,
         \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 , \39331 , \39332 ,
         \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 , \39341 , \39342 ,
         \39343 , \39344 , \39345 , \39346 , \39347 , \39348 , \39349 , \39350 , \39351 , \39352 ,
         \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 , \39361 , \39362 ,
         \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 , \39371 , \39372 ,
         \39373 , \39374 , \39375 , \39376 , \39377 , \39378 , \39379 , \39380 , \39381 ;
buf \U$labajz3969 ( R_81_9fc6f08, \37902 );
buf \U$labajz3970 ( R_82_9fc5ea0, \37934 );
buf \U$labajz3971 ( R_83_90f04e0, \37947 );
buf \U$labajz3972 ( R_84_90effa0, \37960 );
buf \U$labajz3973 ( R_85_90e8ad0, \37975 );
buf \U$labajz3974 ( R_86_90e3e08, \37987 );
buf \U$labajz3975 ( R_87_90f1a88, \37999 );
buf \U$labajz3976 ( R_88_90e8638, \38002 );
buf \U$labajz3977 ( R_89_90f1200, \38022 );
buf \U$labajz3978 ( R_8a_90f12a8, \38036 );
buf \U$labajz3979 ( R_8b_90f0cc0, \38050 );
buf \U$labajz3980 ( R_8c_90ef088, \38057 );
buf \U$labajz3981 ( R_8d_90f1158, \38087 );
buf \U$labajz3982 ( R_8e_90e49d8, \38100 );
buf \U$labajz3983 ( R_8f_90e3eb0, \38112 );
buf \U$labajz3984 ( R_90_9fc69c8, \38119 );
buf \U$labajz3985 ( R_91_90e9c88, \38130 );
buf \U$labajz3986 ( R_92_90f0588, \38151 );
buf \U$labajz3987 ( R_93_90eacf0, \38166 );
buf \U$labajz3988 ( R_94_90ebb60, \38179 );
buf \U$labajz3989 ( R_95_90e66b8, \38205 );
buf \U$labajz3990 ( R_96_9fc6d10, \38217 );
buf \U$labajz3991 ( R_97_90ead98, \38230 );
buf \U$labajz3992 ( R_98_90e90b8, \38242 );
buf \U$labajz3993 ( R_99_90eb038, \38285 );
buf \U$labajz3994 ( R_9a_90e9d30, \38292 );
buf \U$labajz3995 ( R_9b_90e7bb8, \38314 );
buf \U$labajz3996 ( R_9c_9fc7b80, \38321 );
buf \U$labajz3997 ( R_9d_90ebd58, \38335 );
buf \U$labajz3998 ( R_9e_90e9a90, \38347 );
buf \U$labajz3999 ( R_9f_90efb08, \38359 );
buf \U$labajz4000 ( R_a0_90e6e98, \38367 );
buf \U$labajz4001 ( R_a1_90f0780, \38407 );
buf \U$labajz4002 ( R_a2_90e2da0, \38430 );
buf \U$labajz4003 ( R_a3_90f0240, \38441 );
buf \U$labajz4004 ( R_a4_9fc7ad8, \38448 );
buf \U$labajz4005 ( R_a5_9fc73a0, \38474 );
buf \U$labajz4006 ( R_a6_9fc6680, \38482 );
buf \U$labajz4007 ( R_a7_90e4f18, \38494 );
buf \U$labajz4008 ( R_a8_90e3388, \38501 );
buf \U$labajz4009 ( R_a9_9fc67d0, \38524 );
buf \U$labajz4010 ( R_aa_90f17e8, \38532 );
buf \U$labajz4011 ( R_ab_90e4888, \38544 );
buf \U$labajz4012 ( R_ac_90e9010, \38551 );
buf \U$labajz4013 ( R_ad_90eee90, \38565 );
buf \U$labajz4014 ( R_ae_90e53b0, \38577 );
buf \U$labajz4015 ( R_af_90ebc08, \38588 );
buf \U$labajz4016 ( R_b0_90e8440, \38595 );
buf \U$labajz4017 ( R_b1_90ea900, \38620 );
buf \U$labajz4018 ( R_b2_90e9400, \38629 );
buf \U$labajz4019 ( R_b3_9fc6bc0, \38642 );
buf \U$labajz4020 ( R_b4_90e4690, \38649 );
buf \U$labajz4021 ( R_b5_90e3778, \38663 );
buf \U$labajz4022 ( R_b6_90e9160, \38681 );
buf \U$labajz4023 ( R_b7_90e29b0, \38693 );
buf \U$labajz4024 ( R_b8_90e2278, \38701 );
buf \U$labajz4025 ( R_b9_9fc6a70, \38727 );
buf \U$labajz4026 ( R_ba_90ebf50, \38734 );
buf \U$labajz4027 ( R_bb_90f0e10, \38746 );
buf \U$labajz4028 ( R_bc_9fc7640, \38753 );
buf \U$labajz4029 ( R_bd_90f1dd0, \38773 );
buf \U$labajz4030 ( R_be_90f0630, \38781 );
buf \U$labajz4031 ( R_bf_90f0eb8, \38793 );
buf \U$labajz4032 ( R_c0_90e34d8, \38800 );
buf \U$labajz4033 ( R_c1_90e9f28, \38829 );
buf \U$labajz4034 ( R_c2_90f0d68, \38836 );
buf \U$labajz4035 ( R_c3_90ea7b0, \38844 );
buf \U$labajz4036 ( R_c4_9fc7448, \38851 );
buf \U$labajz4037 ( R_c5_90eb428, \38870 );
buf \U$labajz4038 ( R_c6_90e81a0, \38877 );
buf \U$labajz4039 ( R_c7_90f0a20, \38891 );
buf \U$labajz4040 ( R_c8_90efda8, \38898 );
buf \U$labajz4041 ( R_c9_90e2c50, \38921 );
buf \U$labajz4042 ( R_ca_90e88d8, \38928 );
buf \U$labajz4043 ( R_cb_9fc6530, \38940 );
buf \U$labajz4044 ( R_cc_90f06d8, \38947 );
buf \U$labajz4045 ( R_cd_90efa60, \38965 );
buf \U$labajz4046 ( R_ce_90e2b00, \38972 );
buf \U$labajz4047 ( R_cf_9fc6920, \38980 );
buf \U$labajz4048 ( R_d0_90f1f20, \38987 );
buf \U$labajz4049 ( R_d1_90e7678, \39014 );
buf \U$labajz4050 ( R_d2_90efd00, \39021 );
buf \U$labajz4051 ( R_d3_90e7e58, \39033 );
buf \U$labajz4052 ( R_d4_90e7d08, \39040 );
buf \U$labajz4053 ( R_d5_90eaa50, \39061 );
buf \U$labajz4054 ( R_d6_90e3040, \39068 );
buf \U$labajz4055 ( R_d7_90efe50, \39075 );
buf \U$labajz4056 ( R_d8_90f1350, \39083 );
buf \U$labajz4057 ( R_d9_9fc71a8, \39108 );
buf \U$labajz4058 ( R_da_9fc9cf8, \39115 );
buf \U$labajz4059 ( R_db_90ef9b8, \39124 );
buf \U$labajz4060 ( R_dc_90e4540, \39131 );
buf \U$labajz4061 ( R_dd_90f0ac8, \39151 );
buf \U$labajz4062 ( R_de_90e30e8, \39158 );
buf \U$labajz4063 ( R_df_9fc6290, \39167 );
buf \U$labajz4064 ( R_e0_9fc78e0, \39174 );
buf \U$labajz4065 ( R_e1_90e5500, \39197 );
buf \U$labajz4066 ( R_e2_90e68b0, \39204 );
buf \U$labajz4067 ( R_e3_90eede8, \39215 );
buf \U$labajz4068 ( R_e4_90e64c0, \39222 );
buf \U$labajz4069 ( R_e5_9fc7100, \39241 );
buf \U$labajz4070 ( R_e6_90e2470, \39248 );
buf \U$labajz4071 ( R_e7_90ebea8, \39256 );
buf \U$labajz4072 ( R_e8_90e4a80, \39263 );
buf \U$labajz4073 ( R_e9_90ef910, \39282 );
buf \U$labajz4074 ( R_ea_9fc7c28, \39289 );
buf \U$labajz4075 ( R_eb_90eb4d0, \39299 );
buf \U$labajz4076 ( R_ec_90f14a0, \39302 );
buf \U$labajz4077 ( R_ed_90ef5c8, \39321 );
buf \U$labajz4078 ( R_ee_90e4498, \39328 );
buf \U$labajz4079 ( R_ef_90e4000, \39341 );
buf \U$labajz4080 ( R_f0_90f0048, \39348 );
buf \U$labajz4081 ( R_f1_90ea3c0, \39361 );
buf \U$labajz4082 ( R_f2_90f1e78, \39368 );
buf \U$labajz4083 ( R_f3_90f00f0, \39381 );
not \U$1 ( \248 , RIbe28de0_41);
not \U$2 ( \249 , RIbe27b98_2);
nand \U$3 ( \250 , \248 , \249 );
not \U$4 ( \251 , RIbe29920_65);
nand \U$5 ( \252 , \251 , RIbe28de0_41);
nand \U$6 ( \253 , RIbe27b98_2, RIbe29920_65);
nand \U$7 ( \254 , \250 , \252 , \253 );
buf \U$8 ( \255 , \254 );
not \U$9 ( \256 , \255 );
not \U$10 ( \257 , \256 );
not \U$11 ( \258 , \257 );
not \U$12 ( \259 , \258 );
not \U$13 ( \260 , \259 );
or \U$14 ( \261 , RIbe27b98_2, RIbe28c78_38);
nand \U$15 ( \262 , RIbe27b98_2, RIbe28c78_38);
nand \U$16 ( \263 , \261 , \262 );
not \U$17 ( \264 , \263 );
and \U$18 ( \265 , \260 , \264 );
xor \U$19 ( \266 , RIbe28de0_41, RIbe29920_65);
buf \U$20 ( \267 , \266 );
not \U$21 ( \268 , \267 );
not \U$22 ( \269 , \268 );
nand \U$23 ( \270 , RIbe27b98_2, RIbe28318_18);
not \U$24 ( \271 , \270 );
nor \U$25 ( \272 , RIbe27b98_2, RIbe28318_18);
nor \U$26 ( \273 , \271 , \272 );
and \U$27 ( \274 , \269 , \273 );
nor \U$28 ( \275 , \265 , \274 );
xor \U$29 ( \276 , RIbe29038_46, RIbe29650_59);
xor \U$30 ( \277 , RIbe29650_59, RIbe296c8_60);
not \U$31 ( \278 , \277 );
nand \U$32 ( \279 , \276 , \278 );
not \U$33 ( \280 , \279 );
buf \U$34 ( \281 , \280 );
buf \U$35 ( \282 , \281 );
not \U$36 ( \283 , \282 );
buf \U$37 ( \284 , \277 );
not \U$38 ( \285 , \284 );
not \U$39 ( \286 , \285 );
buf \U$40 ( \287 , \286 );
not \U$41 ( \288 , \287 );
and \U$42 ( \289 , \283 , \288 );
not \U$43 ( \290 , RIbe29038_46);
nor \U$44 ( \291 , \289 , \290 );
xnor \U$45 ( \292 , \275 , \291 );
and \U$46 ( \293 , RIbe290b0_47, RIbe29a88_68);
not \U$47 ( \294 , RIbe290b0_47);
and \U$48 ( \295 , \294 , RIbe27d78_6);
nor \U$49 ( \296 , \293 , \295 );
not \U$50 ( \297 , \296 );
nand \U$51 ( \298 , RIbe27d78_6, RIbe29a88_68);
nand \U$52 ( \299 , \297 , \298 );
buf \U$53 ( \300 , \299 );
buf \U$54 ( \301 , \300 );
not \U$55 ( \302 , \301 );
not \U$56 ( \303 , RIbe27d78_6);
not \U$57 ( \304 , RIbe286d8_26);
and \U$58 ( \305 , \303 , \304 );
and \U$59 ( \306 , RIbe27d78_6, RIbe286d8_26);
nor \U$60 ( \307 , \305 , \306 );
and \U$61 ( \308 , \302 , \307 );
not \U$62 ( \309 , RIbe290b0_47);
not \U$63 ( \310 , RIbe29a88_68);
and \U$64 ( \311 , \309 , \310 );
and \U$65 ( \312 , RIbe290b0_47, RIbe29a88_68);
nor \U$66 ( \313 , \311 , \312 );
buf \U$67 ( \314 , \313 );
buf \U$68 ( \315 , \314 );
or \U$69 ( \316 , \303 , RIbe27ee0_9);
not \U$70 ( \317 , RIbe27ee0_9);
or \U$71 ( \318 , \317 , RIbe27d78_6);
nand \U$72 ( \319 , \316 , \318 );
and \U$73 ( \320 , \315 , \319 );
nor \U$74 ( \321 , \308 , \320 );
or \U$75 ( \322 , \292 , \321 );
or \U$76 ( \323 , \275 , \291 );
nand \U$77 ( \324 , \322 , \323 );
or \U$78 ( \325 , RIbe28de0_41, RIbe28e58_42);
nand \U$79 ( \326 , RIbe27c10_3, RIbe28de0_41);
nand \U$80 ( \327 , \325 , \326 );
not \U$81 ( \328 , RIbe28e58_42);
nor \U$82 ( \329 , \328 , RIbe27c10_3);
nor \U$83 ( \330 , \327 , \329 );
buf \U$84 ( \331 , \330 );
buf \U$85 ( \332 , \331 );
not \U$86 ( \333 , \332 );
not \U$87 ( \334 , \333 );
not \U$88 ( \335 , RIbe284f8_22);
not \U$89 ( \336 , RIbe28de0_41);
and \U$90 ( \337 , \335 , \336 );
and \U$91 ( \338 , RIbe284f8_22, RIbe28de0_41);
nor \U$92 ( \339 , \337 , \338 );
and \U$93 ( \340 , \334 , \339 );
not \U$94 ( \341 , RIbe27c10_3);
not \U$95 ( \342 , RIbe28e58_42);
and \U$96 ( \343 , \341 , \342 );
and \U$97 ( \344 , RIbe27c10_3, RIbe28e58_42);
nor \U$98 ( \345 , \343 , \344 );
buf \U$99 ( \346 , \345 );
buf \U$100 ( \347 , \346 );
not \U$101 ( \348 , \347 );
not \U$102 ( \349 , \348 );
xor \U$103 ( \350 , RIbe28750_27, RIbe28de0_41);
and \U$104 ( \351 , \349 , \350 );
nor \U$105 ( \352 , \340 , \351 );
nand \U$106 ( \353 , RIbe27b98_2, RIbe28c00_37);
xnor \U$107 ( \354 , \352 , \353 );
xor \U$108 ( \355 , RIbe27d00_5, RIbe27d78_6);
not \U$109 ( \356 , \355 );
xor \U$110 ( \357 , RIbe27c10_3, RIbe27d00_5);
nand \U$111 ( \358 , \356 , \357 );
buf \U$112 ( \359 , \358 );
buf \U$113 ( \360 , \359 );
not \U$114 ( \361 , \360 );
buf \U$115 ( \362 , \361 );
not \U$116 ( \363 , RIbe27c10_3);
not \U$117 ( \364 , RIbe28840_29);
and \U$118 ( \365 , \363 , \364 );
and \U$119 ( \366 , RIbe27c10_3, RIbe28840_29);
nor \U$120 ( \367 , \365 , \366 );
and \U$121 ( \368 , \362 , \367 );
not \U$122 ( \369 , \356 );
buf \U$123 ( \370 , \369 );
not \U$124 ( \371 , RIbe28570_23);
and \U$125 ( \372 , \363 , \371 );
and \U$126 ( \373 , RIbe27c10_3, RIbe28570_23);
nor \U$127 ( \374 , \372 , \373 );
and \U$128 ( \375 , \370 , \374 );
nor \U$129 ( \376 , \368 , \375 );
or \U$130 ( \377 , \354 , \376 );
or \U$131 ( \378 , \352 , \353 );
nand \U$132 ( \379 , \377 , \378 );
xor \U$133 ( \380 , \324 , \379 );
xnor \U$134 ( \381 , RIbe28fc0_45, RIbe29038_46);
xor \U$135 ( \382 , RIbe28fc0_45, RIbe290b0_47);
nand \U$136 ( \383 , \381 , \382 );
buf \U$137 ( \384 , \383 );
buf \U$138 ( \385 , \384 );
not \U$139 ( \386 , \385 );
not \U$140 ( \387 , RIbe290b0_47);
not \U$141 ( \388 , RIbe29380_53);
and \U$142 ( \389 , \387 , \388 );
and \U$143 ( \390 , RIbe290b0_47, RIbe29380_53);
nor \U$144 ( \391 , \389 , \390 );
and \U$145 ( \392 , \386 , \391 );
and \U$146 ( \393 , RIbe28fc0_45, RIbe29038_46);
not \U$147 ( \394 , RIbe28fc0_45);
not \U$148 ( \395 , RIbe29038_46);
and \U$149 ( \396 , \394 , \395 );
nor \U$150 ( \397 , \393 , \396 );
buf \U$151 ( \398 , \397 );
buf \U$152 ( \399 , \398 );
and \U$153 ( \400 , \399 , RIbe290b0_47);
nor \U$154 ( \401 , \392 , \400 );
xnor \U$155 ( \402 , \401 , \262 );
and \U$156 ( \403 , \362 , \374 );
and \U$157 ( \404 , \363 , \304 );
and \U$158 ( \405 , RIbe27c10_3, RIbe286d8_26);
nor \U$159 ( \406 , \404 , \405 );
and \U$160 ( \407 , \370 , \406 );
nor \U$161 ( \408 , \403 , \407 );
xor \U$162 ( \409 , \402 , \408 );
and \U$163 ( \410 , \380 , \409 );
and \U$164 ( \411 , \324 , \379 );
nor \U$165 ( \412 , \410 , \411 );
not \U$166 ( \413 , \259 );
and \U$167 ( \414 , \413 , \273 );
xor \U$168 ( \415 , RIbe284f8_22, RIbe27b98_2);
and \U$169 ( \416 , \269 , \415 );
nor \U$170 ( \417 , \414 , \416 );
not \U$171 ( \418 , \417 );
buf \U$172 ( \419 , \334 );
and \U$173 ( \420 , \419 , \350 );
not \U$174 ( \421 , RIbe28de0_41);
and \U$175 ( \422 , \364 , \421 );
and \U$176 ( \423 , RIbe28840_29, RIbe28de0_41);
nor \U$177 ( \424 , \422 , \423 );
and \U$178 ( \425 , \349 , \424 );
nor \U$179 ( \426 , \420 , \425 );
not \U$180 ( \427 , \426 );
and \U$181 ( \428 , \418 , \427 );
xor \U$182 ( \429 , \417 , \426 );
and \U$183 ( \430 , \302 , \319 );
not \U$184 ( \431 , RIbe28048_12);
and \U$185 ( \432 , \431 , \303 );
and \U$186 ( \433 , RIbe27d78_6, RIbe28048_12);
nor \U$187 ( \434 , \432 , \433 );
and \U$188 ( \435 , \315 , \434 );
nor \U$189 ( \436 , \430 , \435 );
and \U$190 ( \437 , \429 , \436 );
nor \U$191 ( \438 , \428 , \437 );
and \U$192 ( \439 , \419 , \424 );
and \U$193 ( \440 , \421 , \371 );
and \U$194 ( \441 , RIbe28570_23, RIbe28de0_41);
nor \U$195 ( \442 , \440 , \441 );
and \U$196 ( \443 , \349 , \442 );
nor \U$197 ( \444 , \439 , \443 );
xor \U$198 ( \445 , \444 , \270 );
buf \U$199 ( \446 , \269 );
not \U$200 ( \447 , \446 );
not \U$201 ( \448 , \447 );
or \U$202 ( \449 , RIbe27b98_2, RIbe28750_27);
nand \U$203 ( \450 , RIbe27b98_2, RIbe28750_27);
nand \U$204 ( \451 , \449 , \450 );
not \U$205 ( \452 , \451 );
and \U$206 ( \453 , \448 , \452 );
and \U$207 ( \454 , \413 , \415 );
nor \U$208 ( \455 , \453 , \454 );
xor \U$209 ( \456 , \445 , \455 );
xor \U$210 ( \457 , \438 , \456 );
or \U$211 ( \458 , \402 , \408 );
or \U$212 ( \459 , \401 , \262 );
nand \U$213 ( \460 , \458 , \459 );
not \U$214 ( \461 , \436 );
and \U$215 ( \462 , \460 , \461 );
not \U$216 ( \463 , \460 );
and \U$217 ( \464 , \463 , \436 );
nor \U$218 ( \465 , \462 , \464 );
buf \U$219 ( \466 , \386 );
not \U$220 ( \467 , \466 );
not \U$221 ( \468 , \398 );
not \U$222 ( \469 , \468 );
not \U$223 ( \470 , \469 );
and \U$224 ( \471 , \467 , \470 );
nor \U$225 ( \472 , \471 , \387 );
and \U$226 ( \473 , \302 , \434 );
and \U$227 ( \474 , \303 , \388 );
and \U$228 ( \475 , RIbe27d78_6, RIbe29380_53);
nor \U$229 ( \476 , \474 , \475 );
and \U$230 ( \477 , \315 , \476 );
nor \U$231 ( \478 , \473 , \477 );
xnor \U$232 ( \479 , \472 , \478 );
and \U$233 ( \480 , \362 , \406 );
and \U$234 ( \481 , \363 , \317 );
and \U$235 ( \482 , RIbe27c10_3, RIbe27ee0_9);
nor \U$236 ( \483 , \481 , \482 );
and \U$237 ( \484 , \370 , \483 );
nor \U$238 ( \485 , \480 , \484 );
xor \U$239 ( \486 , \479 , \485 );
xnor \U$240 ( \487 , \465 , \486 );
xor \U$241 ( \488 , \457 , \487 );
xor \U$242 ( \489 , \412 , \488 );
and \U$243 ( \490 , \290 , \388 );
and \U$244 ( \491 , RIbe29038_46, RIbe29380_53);
nor \U$245 ( \492 , \490 , \491 );
not \U$246 ( \493 , \492 );
not \U$247 ( \494 , \282 );
or \U$248 ( \495 , \493 , \494 );
nand \U$249 ( \496 , \287 , RIbe29038_46);
nand \U$250 ( \497 , \495 , \496 );
not \U$251 ( \498 , \497 );
and \U$252 ( \499 , \431 , \387 );
and \U$253 ( \500 , RIbe28048_12, RIbe290b0_47);
nor \U$254 ( \501 , \499 , \500 );
and \U$255 ( \502 , \466 , \501 );
and \U$256 ( \503 , \469 , \391 );
nor \U$257 ( \504 , \502 , \503 );
not \U$258 ( \505 , \504 );
or \U$259 ( \506 , \498 , \505 );
or \U$260 ( \507 , \504 , \497 );
nand \U$261 ( \508 , \506 , \507 );
not \U$262 ( \509 , \508 );
xor \U$263 ( \510 , RIbe28318_18, RIbe28de0_41);
not \U$264 ( \511 , \510 );
not \U$265 ( \512 , \334 );
or \U$266 ( \513 , \511 , \512 );
buf \U$267 ( \514 , \346 );
nand \U$268 ( \515 , \514 , \339 );
nand \U$269 ( \516 , \513 , \515 );
not \U$270 ( \517 , \516 );
nand \U$271 ( \518 , RIbe27b98_2, RIbe29308_52);
not \U$272 ( \519 , \518 );
and \U$273 ( \520 , \517 , \519 );
and \U$274 ( \521 , \516 , \518 );
nor \U$275 ( \522 , \520 , \521 );
not \U$276 ( \523 , \384 );
not \U$277 ( \524 , \523 );
not \U$278 ( \525 , \524 );
xor \U$279 ( \526 , RIbe27ee0_9, RIbe290b0_47);
and \U$280 ( \527 , \525 , \526 );
and \U$281 ( \528 , \399 , \501 );
nor \U$282 ( \529 , \527 , \528 );
or \U$283 ( \530 , \522 , \529 );
not \U$284 ( \531 , \516 );
or \U$285 ( \532 , \531 , \518 );
nand \U$286 ( \533 , \530 , \532 );
not \U$287 ( \534 , \533 );
or \U$288 ( \535 , \509 , \534 );
not \U$289 ( \536 , \497 );
or \U$290 ( \537 , \536 , \504 );
nand \U$291 ( \538 , \535 , \537 );
xor \U$292 ( \539 , \417 , \426 );
xor \U$293 ( \540 , \539 , \436 );
and \U$294 ( \541 , \538 , \540 );
not \U$295 ( \542 , \269 );
not \U$296 ( \543 , \542 );
not \U$297 ( \544 , \263 );
and \U$298 ( \545 , \543 , \544 );
not \U$299 ( \546 , \257 );
not \U$300 ( \547 , \353 );
nor \U$301 ( \548 , RIbe27b98_2, RIbe28c00_37);
nor \U$302 ( \549 , \547 , \548 );
and \U$303 ( \550 , \546 , \549 );
nor \U$304 ( \551 , \545 , \550 );
and \U$305 ( \552 , \303 , \371 );
and \U$306 ( \553 , RIbe27d78_6, RIbe28570_23);
nor \U$307 ( \554 , \552 , \553 );
and \U$308 ( \555 , \302 , \554 );
and \U$309 ( \556 , \315 , \307 );
nor \U$310 ( \557 , \555 , \556 );
xor \U$311 ( \558 , \551 , \557 );
not \U$312 ( \559 , RIbe27c10_3);
not \U$313 ( \560 , RIbe28750_27);
and \U$314 ( \561 , \559 , \560 );
and \U$315 ( \562 , RIbe27c10_3, RIbe28750_27);
nor \U$316 ( \563 , \561 , \562 );
and \U$317 ( \564 , \362 , \563 );
and \U$318 ( \565 , \370 , \367 );
nor \U$319 ( \566 , \564 , \565 );
and \U$320 ( \567 , \558 , \566 );
and \U$321 ( \568 , \551 , \557 );
nor \U$322 ( \569 , \567 , \568 );
xor \U$323 ( \570 , \376 , \354 );
xor \U$324 ( \571 , \569 , \570 );
xor \U$325 ( \572 , \292 , \321 );
and \U$326 ( \573 , \571 , \572 );
and \U$327 ( \574 , \569 , \570 );
or \U$328 ( \575 , \573 , \574 );
xor \U$329 ( \576 , \417 , \426 );
xor \U$330 ( \577 , \576 , \436 );
and \U$331 ( \578 , \575 , \577 );
and \U$332 ( \579 , \538 , \575 );
or \U$333 ( \580 , \541 , \578 , \579 );
not \U$334 ( \581 , \580 );
and \U$335 ( \582 , \489 , \581 );
and \U$336 ( \583 , \412 , \488 );
or \U$337 ( \584 , \582 , \583 );
not \U$338 ( \585 , \584 );
not \U$339 ( \586 , \585 );
not \U$340 ( \587 , \259 );
not \U$341 ( \588 , \451 );
and \U$342 ( \589 , \587 , \588 );
nand \U$343 ( \590 , RIbe27b98_2, RIbe28840_29);
not \U$344 ( \591 , \590 );
nor \U$345 ( \592 , RIbe27b98_2, RIbe28840_29);
nor \U$346 ( \593 , \591 , \592 );
and \U$347 ( \594 , \269 , \593 );
nor \U$348 ( \595 , \589 , \594 );
and \U$349 ( \596 , \419 , \442 );
and \U$350 ( \597 , \421 , \304 );
and \U$351 ( \598 , RIbe286d8_26, RIbe28de0_41);
nor \U$352 ( \599 , \597 , \598 );
and \U$353 ( \600 , \349 , \599 );
nor \U$354 ( \601 , \596 , \600 );
xnor \U$355 ( \602 , \595 , \601 );
and \U$356 ( \603 , \362 , \483 );
and \U$357 ( \604 , \431 , \363 );
and \U$358 ( \605 , RIbe27c10_3, RIbe28048_12);
nor \U$359 ( \606 , \604 , \605 );
and \U$360 ( \607 , \370 , \606 );
nor \U$361 ( \608 , \603 , \607 );
xor \U$362 ( \609 , \602 , \608 );
xor \U$363 ( \610 , \444 , \270 );
and \U$364 ( \611 , \610 , \455 );
and \U$365 ( \612 , \444 , \270 );
nor \U$366 ( \613 , \611 , \612 );
xor \U$367 ( \614 , \609 , \613 );
or \U$368 ( \615 , \479 , \485 );
or \U$369 ( \616 , \472 , \478 );
nand \U$370 ( \617 , \615 , \616 );
and \U$371 ( \618 , RIbe284f8_22, RIbe27b98_2);
not \U$372 ( \619 , \618 );
and \U$373 ( \620 , \302 , \476 );
and \U$374 ( \621 , \315 , RIbe27d78_6);
nor \U$375 ( \622 , \620 , \621 );
not \U$376 ( \623 , \622 );
not \U$377 ( \624 , \623 );
or \U$378 ( \625 , \619 , \624 );
or \U$379 ( \626 , \623 , \618 );
nand \U$380 ( \627 , \625 , \626 );
xor \U$381 ( \628 , \617 , \627 );
xnor \U$382 ( \629 , \614 , \628 );
and \U$383 ( \630 , \465 , \486 );
and \U$384 ( \631 , \460 , \461 );
nor \U$385 ( \632 , \630 , \631 );
xor \U$386 ( \633 , \629 , \632 );
xor \U$387 ( \634 , \438 , \456 );
and \U$388 ( \635 , \634 , \487 );
and \U$389 ( \636 , \438 , \456 );
or \U$390 ( \637 , \635 , \636 );
xor \U$391 ( \638 , \633 , \637 );
nand \U$392 ( \639 , \586 , \638 );
xor \U$393 ( \640 , \629 , \632 );
and \U$394 ( \641 , \640 , \637 );
and \U$395 ( \642 , \629 , \632 );
or \U$396 ( \643 , \641 , \642 );
and \U$397 ( \644 , \614 , \628 );
and \U$398 ( \645 , \609 , \613 );
nor \U$399 ( \646 , \644 , \645 );
and \U$400 ( \647 , \617 , \627 );
and \U$401 ( \648 , \622 , \618 );
nor \U$402 ( \649 , \647 , \648 );
xor \U$403 ( \650 , \646 , \649 );
and \U$404 ( \651 , \419 , \599 );
and \U$405 ( \652 , \317 , \421 );
and \U$406 ( \653 , RIbe27ee0_9, RIbe28de0_41);
nor \U$407 ( \654 , \652 , \653 );
and \U$408 ( \655 , \349 , \654 );
nor \U$409 ( \656 , \651 , \655 );
xnor \U$410 ( \657 , \656 , \450 );
and \U$411 ( \658 , \413 , \593 );
and \U$412 ( \659 , \249 , \371 );
nand \U$413 ( \660 , RIbe27b98_2, RIbe28570_23);
not \U$414 ( \661 , \660 );
nor \U$415 ( \662 , \659 , \661 );
and \U$416 ( \663 , \446 , \662 );
nor \U$417 ( \664 , \658 , \663 );
xor \U$418 ( \665 , \657 , \664 );
or \U$419 ( \666 , \602 , \608 );
or \U$420 ( \667 , \595 , \601 );
nand \U$421 ( \668 , \666 , \667 );
xor \U$422 ( \669 , \665 , \668 );
not \U$423 ( \670 , \315 );
and \U$424 ( \671 , \301 , \670 );
nor \U$425 ( \672 , \671 , \303 );
and \U$426 ( \673 , \672 , \623 );
not \U$427 ( \674 , \672 );
and \U$428 ( \675 , \674 , \622 );
nor \U$429 ( \676 , \673 , \675 );
and \U$430 ( \677 , \362 , \606 );
and \U$431 ( \678 , \363 , \388 );
and \U$432 ( \679 , RIbe27c10_3, RIbe29380_53);
nor \U$433 ( \680 , \678 , \679 );
and \U$434 ( \681 , \370 , \680 );
nor \U$435 ( \682 , \677 , \681 );
xor \U$436 ( \683 , \676 , \682 );
xnor \U$437 ( \684 , \669 , \683 );
xor \U$438 ( \685 , \650 , \684 );
nand \U$439 ( \686 , \643 , \685 );
and \U$440 ( \687 , \639 , \686 );
not \U$441 ( \688 , \687 );
xor \U$442 ( \689 , \646 , \649 );
and \U$443 ( \690 , \689 , \684 );
and \U$444 ( \691 , \646 , \649 );
or \U$445 ( \692 , \690 , \691 );
not \U$446 ( \693 , \692 );
or \U$447 ( \694 , \657 , \664 );
or \U$448 ( \695 , \656 , \450 );
nand \U$449 ( \696 , \694 , \695 );
and \U$450 ( \697 , \362 , \680 );
and \U$451 ( \698 , \370 , RIbe27c10_3);
nor \U$452 ( \699 , \697 , \698 );
and \U$453 ( \700 , \696 , \699 );
not \U$454 ( \701 , \696 );
not \U$455 ( \702 , \699 );
and \U$456 ( \703 , \701 , \702 );
nor \U$457 ( \704 , \700 , \703 );
and \U$458 ( \705 , \419 , \654 );
and \U$459 ( \706 , \431 , \421 );
and \U$460 ( \707 , RIbe28048_12, RIbe28de0_41);
nor \U$461 ( \708 , \706 , \707 );
and \U$462 ( \709 , \349 , \708 );
nor \U$463 ( \710 , \705 , \709 );
xnor \U$464 ( \711 , \710 , \590 );
and \U$465 ( \712 , \413 , \662 );
not \U$466 ( \713 , RIbe27b98_2);
and \U$467 ( \714 , \713 , \304 );
nor \U$468 ( \715 , \304 , \249 );
nor \U$469 ( \716 , \714 , \715 );
and \U$470 ( \717 , \446 , \716 );
nor \U$471 ( \718 , \712 , \717 );
xor \U$472 ( \719 , \711 , \718 );
xor \U$473 ( \720 , \704 , \719 );
not \U$474 ( \721 , \720 );
and \U$475 ( \722 , \669 , \683 );
and \U$476 ( \723 , \668 , \665 );
nor \U$477 ( \724 , \722 , \723 );
not \U$478 ( \725 , \724 );
or \U$479 ( \726 , \676 , \682 );
or \U$480 ( \727 , \672 , \622 );
nand \U$481 ( \728 , \726 , \727 );
not \U$482 ( \729 , \728 );
and \U$483 ( \730 , \725 , \729 );
and \U$484 ( \731 , \724 , \728 );
nor \U$485 ( \732 , \730 , \731 );
not \U$486 ( \733 , \732 );
or \U$487 ( \734 , \721 , \733 );
or \U$488 ( \735 , \732 , \720 );
nand \U$489 ( \736 , \734 , \735 );
nor \U$490 ( \737 , \693 , \736 );
nor \U$491 ( \738 , \688 , \737 );
and \U$492 ( \739 , \720 , \728 );
not \U$493 ( \740 , \720 );
not \U$494 ( \741 , \728 );
and \U$495 ( \742 , \740 , \741 );
nor \U$496 ( \743 , \742 , \724 );
nor \U$497 ( \744 , \739 , \743 );
or \U$498 ( \745 , \711 , \718 );
or \U$499 ( \746 , \710 , \590 );
nand \U$500 ( \747 , \745 , \746 );
or \U$501 ( \748 , \362 , \370 );
nand \U$502 ( \749 , \748 , RIbe27c10_3);
and \U$503 ( \750 , \749 , \702 );
not \U$504 ( \751 , \749 );
and \U$505 ( \752 , \751 , \699 );
nor \U$506 ( \753 , \750 , \752 );
xnor \U$507 ( \754 , \747 , \753 );
and \U$508 ( \755 , \419 , \708 );
and \U$509 ( \756 , \421 , \388 );
and \U$510 ( \757 , RIbe28de0_41, RIbe29380_53);
nor \U$511 ( \758 , \756 , \757 );
and \U$512 ( \759 , \349 , \758 );
nor \U$513 ( \760 , \755 , \759 );
xor \U$514 ( \761 , \760 , \660 );
and \U$515 ( \762 , \413 , \716 );
and \U$516 ( \763 , \713 , \317 );
nor \U$517 ( \764 , \317 , \249 );
nor \U$518 ( \765 , \763 , \764 );
and \U$519 ( \766 , \446 , \765 );
nor \U$520 ( \767 , \762 , \766 );
xor \U$521 ( \768 , \761 , \767 );
xor \U$522 ( \769 , \754 , \768 );
and \U$523 ( \770 , \704 , \719 );
and \U$524 ( \771 , \696 , \699 );
nor \U$525 ( \772 , \770 , \771 );
xor \U$526 ( \773 , \769 , \772 );
nand \U$527 ( \774 , \744 , \773 );
and \U$528 ( \775 , \738 , \774 );
and \U$529 ( \776 , \747 , \753 );
and \U$530 ( \777 , \702 , \749 );
nor \U$531 ( \778 , \776 , \777 );
not \U$532 ( \779 , \778 );
and \U$533 ( \780 , \413 , \765 );
and \U$534 ( \781 , \713 , \431 );
nand \U$535 ( \782 , RIbe27b98_2, RIbe28048_12);
not \U$536 ( \783 , \782 );
nor \U$537 ( \784 , \781 , \783 );
and \U$538 ( \785 , \446 , \784 );
nor \U$539 ( \786 , \780 , \785 );
not \U$540 ( \787 , \715 );
and \U$541 ( \788 , \786 , \787 );
not \U$542 ( \789 , \786 );
and \U$543 ( \790 , \789 , \715 );
nor \U$544 ( \791 , \788 , \790 );
and \U$545 ( \792 , \419 , \758 );
and \U$546 ( \793 , \349 , RIbe28de0_41);
nor \U$547 ( \794 , \792 , \793 );
xor \U$548 ( \795 , \791 , \794 );
xor \U$549 ( \796 , \760 , \660 );
and \U$550 ( \797 , \796 , \767 );
and \U$551 ( \798 , \760 , \660 );
nor \U$552 ( \799 , \797 , \798 );
xor \U$553 ( \800 , \795 , \799 );
not \U$554 ( \801 , \800 );
or \U$555 ( \802 , \779 , \801 );
or \U$556 ( \803 , \778 , \800 );
nand \U$557 ( \804 , \802 , \803 );
not \U$558 ( \805 , \804 );
xor \U$559 ( \806 , \754 , \768 );
and \U$560 ( \807 , \806 , \772 );
and \U$561 ( \808 , \754 , \768 );
or \U$562 ( \809 , \807 , \808 );
nand \U$563 ( \810 , \805 , \809 );
or \U$564 ( \811 , \791 , \794 );
or \U$565 ( \812 , \786 , \715 );
nand \U$566 ( \813 , \811 , \812 );
or \U$567 ( \814 , \813 , \787 );
nand \U$568 ( \815 , \813 , \787 );
nand \U$569 ( \816 , \814 , \815 );
or \U$570 ( \817 , \419 , \349 );
nand \U$571 ( \818 , \817 , RIbe28de0_41);
xor \U$572 ( \819 , \818 , \764 );
not \U$573 ( \820 , \784 );
not \U$574 ( \821 , \413 );
or \U$575 ( \822 , \820 , \821 );
or \U$576 ( \823 , RIbe27b98_2, RIbe29380_53);
nand \U$577 ( \824 , RIbe27b98_2, RIbe29380_53);
nand \U$578 ( \825 , \823 , \824 );
or \U$579 ( \826 , \447 , \825 );
nand \U$580 ( \827 , \822 , \826 );
xor \U$581 ( \828 , \819 , \827 );
xnor \U$582 ( \829 , \816 , \828 );
and \U$583 ( \830 , \795 , \799 );
not \U$584 ( \831 , \795 );
not \U$585 ( \832 , \799 );
and \U$586 ( \833 , \831 , \832 );
nor \U$587 ( \834 , \833 , \778 );
nor \U$588 ( \835 , \830 , \834 );
nand \U$589 ( \836 , \829 , \835 );
and \U$590 ( \837 , \810 , \836 );
and \U$591 ( \838 , \816 , \828 );
and \U$592 ( \839 , \813 , \715 );
nor \U$593 ( \840 , \838 , \839 );
and \U$594 ( \841 , \819 , \827 );
and \U$595 ( \842 , \818 , \764 );
nor \U$596 ( \843 , \841 , \842 );
not \U$597 ( \844 , \259 );
not \U$598 ( \845 , \825 );
and \U$599 ( \846 , \844 , \845 );
and \U$600 ( \847 , \446 , RIbe27b98_2);
nor \U$601 ( \848 , \846 , \847 );
and \U$602 ( \849 , \848 , \782 );
nor \U$603 ( \850 , \848 , \782 );
nor \U$604 ( \851 , \849 , \850 );
xnor \U$605 ( \852 , \843 , \851 );
nand \U$606 ( \853 , \840 , \852 );
and \U$607 ( \854 , \775 , \837 , \853 );
not \U$608 ( \855 , \854 );
xnor \U$609 ( \856 , RIbe280c0_13, RIbe281b0_15);
xor \U$610 ( \857 , RIbe281b0_15, RIbe28228_16);
nor \U$611 ( \858 , \856 , \857 );
not \U$612 ( \859 , \858 );
not \U$613 ( \860 , \859 );
buf \U$614 ( \861 , \860 );
buf \U$615 ( \862 , \861 );
not \U$616 ( \863 , \862 );
not \U$617 ( \864 , \863 );
xnor \U$618 ( \865 , RIbe280c0_13, RIbe28570_23);
not \U$619 ( \866 , \865 );
and \U$620 ( \867 , \864 , \866 );
buf \U$621 ( \868 , \857 );
buf \U$622 ( \869 , \868 );
and \U$623 ( \870 , RIbe280c0_13, RIbe286d8_26);
not \U$624 ( \871 , RIbe280c0_13);
and \U$625 ( \872 , \871 , \304 );
nor \U$626 ( \873 , \870 , \872 );
and \U$627 ( \874 , \869 , \873 );
nor \U$628 ( \875 , \867 , \874 );
xnor \U$629 ( \876 , RIbe28228_16, RIbe29560_57);
xor \U$630 ( \877 , RIbe28930_31, RIbe29560_57);
nor \U$631 ( \878 , \876 , \877 );
buf \U$632 ( \879 , \878 );
not \U$633 ( \880 , \879 );
not \U$634 ( \881 , \880 );
xnor \U$635 ( \882 , RIbe27ee0_9, RIbe28228_16);
not \U$636 ( \883 , \882 );
and \U$637 ( \884 , \881 , \883 );
buf \U$638 ( \885 , \877 );
not \U$639 ( \886 , \885 );
not \U$640 ( \887 , \886 );
not \U$641 ( \888 , RIbe28228_16);
and \U$642 ( \889 , \888 , \431 );
and \U$643 ( \890 , RIbe28048_12, RIbe28228_16);
nor \U$644 ( \891 , \889 , \890 );
and \U$645 ( \892 , \887 , \891 );
nor \U$646 ( \893 , \884 , \892 );
xor \U$647 ( \894 , \875 , \893 );
xor \U$648 ( \895 , RIbe280c0_13, RIbe29830_63);
not \U$649 ( \896 , \895 );
xor \U$650 ( \897 , RIbe296c8_60, RIbe29830_63);
nand \U$651 ( \898 , \896 , \897 );
buf \U$652 ( \899 , \898 );
not \U$653 ( \900 , \899 );
not \U$654 ( \901 , RIbe296c8_60);
not \U$655 ( \902 , RIbe28750_27);
and \U$656 ( \903 , \901 , \902 );
and \U$657 ( \904 , RIbe28750_27, RIbe296c8_60);
nor \U$658 ( \905 , \903 , \904 );
and \U$659 ( \906 , \900 , \905 );
buf \U$660 ( \907 , \895 );
buf \U$661 ( \908 , \907 );
xor \U$662 ( \909 , RIbe28840_29, RIbe296c8_60);
and \U$663 ( \910 , \908 , \909 );
nor \U$664 ( \911 , \906 , \910 );
and \U$665 ( \912 , \894 , \911 );
and \U$666 ( \913 , \875 , \893 );
or \U$667 ( \914 , \912 , \913 );
not \U$668 ( \915 , \914 );
not \U$669 ( \916 , \915 );
and \U$670 ( \917 , RIbe28de0_41, RIbe29470_55);
not \U$671 ( \918 , RIbe28de0_41);
not \U$672 ( \919 , RIbe29470_55);
and \U$673 ( \920 , \918 , \919 );
nor \U$674 ( \921 , \917 , \920 );
not \U$675 ( \922 , \921 );
buf \U$676 ( \923 , \330 );
buf \U$677 ( \924 , \923 );
buf \U$678 ( \925 , \924 );
not \U$679 ( \926 , \925 );
or \U$680 ( \927 , \922 , \926 );
xor \U$681 ( \928 , RIbe28de0_41, RIbe294e8_56);
nand \U$682 ( \929 , \514 , \928 );
nand \U$683 ( \930 , \927 , \929 );
not \U$684 ( \931 , RIbe288b8_30);
and \U$685 ( \932 , \363 , \931 );
and \U$686 ( \933 , RIbe27c10_3, RIbe288b8_30);
nor \U$687 ( \934 , \932 , \933 );
not \U$688 ( \935 , \934 );
not \U$689 ( \936 , \359 );
not \U$690 ( \937 , \936 );
or \U$691 ( \938 , \935 , \937 );
or \U$692 ( \939 , \363 , RIbe28a98_34);
not \U$693 ( \940 , RIbe28a98_34);
or \U$694 ( \941 , \940 , RIbe27c10_3);
nand \U$695 ( \942 , \939 , \941 );
nand \U$696 ( \943 , \370 , \942 );
nand \U$697 ( \944 , \938 , \943 );
xor \U$698 ( \945 , \930 , \944 );
not \U$699 ( \946 , \546 );
or \U$700 ( \947 , RIbe27b98_2, RIbe28138_14);
nand \U$701 ( \948 , RIbe27b98_2, RIbe28138_14);
nand \U$702 ( \949 , \947 , \948 );
or \U$703 ( \950 , \946 , \949 );
not \U$704 ( \951 , RIbe282a0_17);
and \U$705 ( \952 , RIbe27b98_2, \951 );
not \U$706 ( \953 , RIbe27b98_2);
and \U$707 ( \954 , \953 , RIbe282a0_17);
nor \U$708 ( \955 , \952 , \954 );
or \U$709 ( \956 , \542 , \955 );
nand \U$710 ( \957 , \950 , \956 );
and \U$711 ( \958 , \945 , \957 );
and \U$712 ( \959 , \930 , \944 );
or \U$713 ( \960 , \958 , \959 );
xor \U$714 ( \961 , RIbe28930_31, RIbe289a8_32);
not \U$715 ( \962 , \961 );
xor \U$716 ( \963 , RIbe289a8_32, RIbe28a20_33);
nor \U$717 ( \964 , \962 , \963 );
buf \U$718 ( \965 , \964 );
buf \U$719 ( \966 , \965 );
not \U$720 ( \967 , \966 );
xnor \U$721 ( \968 , RIbe28930_31, RIbe29380_53);
or \U$722 ( \969 , \967 , \968 );
buf \U$723 ( \970 , \963 );
buf \U$724 ( \971 , \970 );
not \U$725 ( \972 , \971 );
not \U$726 ( \973 , RIbe28930_31);
or \U$727 ( \974 , \972 , \973 );
nand \U$728 ( \975 , \969 , \974 );
not \U$729 ( \976 , \975 );
xor \U$730 ( \977 , RIbe28318_18, RIbe29038_46);
not \U$731 ( \978 , \977 );
buf \U$732 ( \979 , \281 );
not \U$733 ( \980 , \979 );
or \U$734 ( \981 , \978 , \980 );
xor \U$735 ( \982 , RIbe284f8_22, RIbe29038_46);
nand \U$736 ( \983 , \287 , \982 );
nand \U$737 ( \984 , \981 , \983 );
xor \U$738 ( \985 , RIbe28c00_37, RIbe290b0_47);
not \U$739 ( \986 , \985 );
not \U$740 ( \987 , \466 );
or \U$741 ( \988 , \986 , \987 );
not \U$742 ( \989 , RIbe28c78_38);
not \U$743 ( \990 , RIbe290b0_47);
and \U$744 ( \991 , \989 , \990 );
and \U$745 ( \992 , RIbe28c78_38, RIbe290b0_47);
nor \U$746 ( \993 , \991 , \992 );
nand \U$747 ( \994 , \399 , \993 );
nand \U$748 ( \995 , \988 , \994 );
xor \U$749 ( \996 , \984 , \995 );
not \U$750 ( \997 , \996 );
or \U$751 ( \998 , \976 , \997 );
nand \U$752 ( \999 , \984 , \995 );
nand \U$753 ( \1000 , \998 , \999 );
xor \U$754 ( \1001 , \960 , \1000 );
not \U$755 ( \1002 , \1001 );
or \U$756 ( \1003 , \916 , \1002 );
nand \U$757 ( \1004 , \1000 , \960 );
nand \U$758 ( \1005 , \1003 , \1004 );
xnor \U$759 ( \1006 , RIbe28750_27, RIbe29038_46);
or \U$760 ( \1007 , \283 , \1006 );
not \U$761 ( \1008 , RIbe28840_29);
not \U$762 ( \1009 , RIbe29038_46);
and \U$763 ( \1010 , \1008 , \1009 );
and \U$764 ( \1011 , RIbe28840_29, RIbe29038_46);
nor \U$765 ( \1012 , \1010 , \1011 );
not \U$766 ( \1013 , \1012 );
or \U$767 ( \1014 , \288 , \1013 );
nand \U$768 ( \1015 , \1007 , \1014 );
xor \U$769 ( \1016 , RIbe28318_18, RIbe290b0_47);
not \U$770 ( \1017 , \1016 );
not \U$771 ( \1018 , \466 );
or \U$772 ( \1019 , \1017 , \1018 );
and \U$773 ( \1020 , RIbe284f8_22, RIbe290b0_47);
nor \U$774 ( \1021 , RIbe284f8_22, RIbe290b0_47);
nor \U$775 ( \1022 , \1020 , \1021 );
nand \U$776 ( \1023 , \399 , \1022 );
nand \U$777 ( \1024 , \1019 , \1023 );
not \U$778 ( \1025 , \1024 );
nand \U$779 ( \1026 , RIbe27b98_2, RIbe282a0_17);
not \U$780 ( \1027 , \1026 );
and \U$781 ( \1028 , \1025 , \1027 );
and \U$782 ( \1029 , \1024 , \1026 );
nor \U$783 ( \1030 , \1028 , \1029 );
and \U$784 ( \1031 , \1015 , \1030 );
not \U$785 ( \1032 , \1015 );
not \U$786 ( \1033 , \1030 );
and \U$787 ( \1034 , \1032 , \1033 );
or \U$788 ( \1035 , \1031 , \1034 );
not \U$789 ( \1036 , \670 );
xor \U$790 ( \1037 , RIbe27d78_6, RIbe29308_52);
not \U$791 ( \1038 , \1037 );
not \U$792 ( \1039 , \1038 );
and \U$793 ( \1040 , \1036 , \1039 );
not \U$794 ( \1041 , \296 );
nand \U$795 ( \1042 , \1041 , \298 );
not \U$796 ( \1043 , \1042 );
buf \U$797 ( \1044 , \1043 );
not \U$798 ( \1045 , RIbe27d78_6);
not \U$799 ( \1046 , RIbe293f8_54);
and \U$800 ( \1047 , \1045 , \1046 );
and \U$801 ( \1048 , RIbe27d78_6, RIbe293f8_54);
nor \U$802 ( \1049 , \1047 , \1048 );
and \U$803 ( \1050 , \1044 , \1049 );
nor \U$804 ( \1051 , \1040 , \1050 );
not \U$805 ( \1052 , \873 );
not \U$806 ( \1053 , \859 );
buf \U$807 ( \1054 , \1053 );
not \U$808 ( \1055 , \1054 );
or \U$809 ( \1056 , \1052 , \1055 );
xor \U$810 ( \1057 , RIbe27ee0_9, RIbe280c0_13);
nand \U$811 ( \1058 , \869 , \1057 );
nand \U$812 ( \1059 , \1056 , \1058 );
xor \U$813 ( \1060 , \1051 , \1059 );
buf \U$814 ( \1061 , \879 );
and \U$815 ( \1062 , \1061 , \891 );
and \U$816 ( \1063 , \888 , \388 );
and \U$817 ( \1064 , RIbe28228_16, RIbe29380_53);
nor \U$818 ( \1065 , \1063 , \1064 );
and \U$819 ( \1066 , \887 , \1065 );
nor \U$820 ( \1067 , \1062 , \1066 );
or \U$821 ( \1068 , \1060 , \1067 );
not \U$822 ( \1069 , \1059 );
or \U$823 ( \1070 , \1069 , \1051 );
nand \U$824 ( \1071 , \1068 , \1070 );
xor \U$825 ( \1072 , \1035 , \1071 );
and \U$826 ( \1073 , \1005 , \1072 );
and \U$827 ( \1074 , \1035 , \1071 );
nor \U$828 ( \1075 , \1073 , \1074 );
not \U$829 ( \1076 , \1015 );
not \U$830 ( \1077 , \1033 );
or \U$831 ( \1078 , \1076 , \1077 );
not \U$832 ( \1079 , \1026 );
nand \U$833 ( \1080 , \1079 , \1024 );
nand \U$834 ( \1081 , \1078 , \1080 );
not \U$835 ( \1082 , \886 );
not \U$836 ( \1083 , \880 );
or \U$837 ( \1084 , \1082 , \1083 );
nand \U$838 ( \1085 , \1084 , RIbe28228_16);
not \U$839 ( \1086 , \301 );
not \U$840 ( \1087 , \1086 );
and \U$841 ( \1088 , RIbe27d78_6, RIbe28c00_37);
nor \U$842 ( \1089 , RIbe27d78_6, RIbe28c00_37);
nor \U$843 ( \1090 , \1088 , \1089 );
not \U$844 ( \1091 , \1090 );
or \U$845 ( \1092 , \1087 , \1091 );
not \U$846 ( \1093 , \314 );
xnor \U$847 ( \1094 , RIbe27d78_6, RIbe28c78_38);
or \U$848 ( \1095 , \1093 , \1094 );
nand \U$849 ( \1096 , \1092 , \1095 );
and \U$850 ( \1097 , \1085 , \1096 );
not \U$851 ( \1098 , \1085 );
not \U$852 ( \1099 , \1096 );
and \U$853 ( \1100 , \1098 , \1099 );
nor \U$854 ( \1101 , \1097 , \1100 );
xor \U$855 ( \1102 , \1081 , \1101 );
not \U$856 ( \1103 , \359 );
not \U$857 ( \1104 , \1103 );
xnor \U$858 ( \1105 , RIbe27c10_3, RIbe29308_52);
or \U$859 ( \1106 , \1104 , \1105 );
not \U$860 ( \1107 , \370 );
not \U$861 ( \1108 , RIbe28c00_37);
not \U$862 ( \1109 , RIbe27c10_3);
or \U$863 ( \1110 , \1108 , \1109 );
or \U$864 ( \1111 , RIbe27c10_3, RIbe28c00_37);
nand \U$865 ( \1112 , \1110 , \1111 );
or \U$866 ( \1113 , \1107 , \1112 );
nand \U$867 ( \1114 , \1106 , \1113 );
buf \U$868 ( \1115 , \1042 );
or \U$869 ( \1116 , \1115 , \1094 );
xor \U$870 ( \1117 , RIbe27d78_6, RIbe28318_18);
not \U$871 ( \1118 , \1117 );
or \U$872 ( \1119 , \1093 , \1118 );
nand \U$873 ( \1120 , \1116 , \1119 );
xor \U$874 ( \1121 , \1114 , \1120 );
xnor \U$875 ( \1122 , RIbe27b98_2, RIbe294e8_56);
or \U$876 ( \1123 , \946 , \1122 );
xor \U$877 ( \1124 , RIbe27b98_2, RIbe288b8_30);
not \U$878 ( \1125 , \1124 );
or \U$879 ( \1126 , \542 , \1125 );
nand \U$880 ( \1127 , \1123 , \1126 );
xor \U$881 ( \1128 , \1121 , \1127 );
not \U$882 ( \1129 , \899 );
buf \U$883 ( \1130 , \1129 );
not \U$884 ( \1131 , \1130 );
not \U$885 ( \1132 , \1131 );
and \U$886 ( \1133 , RIbe286d8_26, RIbe296c8_60);
nor \U$887 ( \1134 , RIbe286d8_26, RIbe296c8_60);
nor \U$888 ( \1135 , \1133 , \1134 );
and \U$889 ( \1136 , \1132 , \1135 );
buf \U$890 ( \1137 , \907 );
and \U$891 ( \1138 , \317 , \901 );
and \U$892 ( \1139 , RIbe27ee0_9, RIbe296c8_60);
nor \U$893 ( \1140 , \1138 , \1139 );
and \U$894 ( \1141 , \1137 , \1140 );
nor \U$895 ( \1142 , \1136 , \1141 );
xor \U$896 ( \1143 , RIbe28a98_34, RIbe28de0_41);
not \U$897 ( \1144 , \1143 );
buf \U$898 ( \1145 , \332 );
not \U$899 ( \1146 , \1145 );
or \U$900 ( \1147 , \1144 , \1146 );
not \U$901 ( \1148 , \346 );
not \U$902 ( \1149 , \1148 );
xor \U$903 ( \1150 , RIbe28de0_41, RIbe293f8_54);
nand \U$904 ( \1151 , \1149 , \1150 );
nand \U$905 ( \1152 , \1147 , \1151 );
not \U$906 ( \1153 , \1152 );
nand \U$907 ( \1154 , RIbe27b98_2, RIbe29470_55);
not \U$908 ( \1155 , \1154 );
and \U$909 ( \1156 , \1153 , \1155 );
and \U$910 ( \1157 , \1152 , \1154 );
nor \U$911 ( \1158 , \1156 , \1157 );
xor \U$912 ( \1159 , \1142 , \1158 );
xor \U$913 ( \1160 , \1128 , \1159 );
xnor \U$914 ( \1161 , \1102 , \1160 );
xnor \U$915 ( \1162 , \1075 , \1161 );
not \U$916 ( \1163 , \1037 );
not \U$917 ( \1164 , \300 );
not \U$918 ( \1165 , \1164 );
or \U$919 ( \1166 , \1163 , \1165 );
nand \U$920 ( \1167 , \315 , \1090 );
nand \U$921 ( \1168 , \1166 , \1167 );
not \U$922 ( \1169 , \942 );
not \U$923 ( \1170 , \361 );
or \U$924 ( \1171 , \1169 , \1170 );
xnor \U$925 ( \1172 , RIbe27d00_5, RIbe27d78_6);
not \U$926 ( \1173 , \1172 );
buf \U$927 ( \1174 , \1173 );
xor \U$928 ( \1175 , RIbe27c10_3, RIbe293f8_54);
nand \U$929 ( \1176 , \1174 , \1175 );
nand \U$930 ( \1177 , \1171 , \1176 );
xor \U$931 ( \1178 , \1168 , \1177 );
or \U$932 ( \1179 , \946 , \955 );
xnor \U$933 ( \1180 , RIbe27b98_2, RIbe29470_55);
or \U$934 ( \1181 , \268 , \1180 );
nand \U$935 ( \1182 , \1179 , \1181 );
and \U$936 ( \1183 , \1178 , \1182 );
and \U$937 ( \1184 , \1168 , \1177 );
or \U$938 ( \1185 , \1183 , \1184 );
xnor \U$939 ( \1186 , \1185 , \1096 );
and \U$940 ( \1187 , \466 , \993 );
and \U$941 ( \1188 , \469 , \1016 );
nor \U$942 ( \1189 , \1187 , \1188 );
not \U$943 ( \1190 , \1189 );
not \U$944 ( \1191 , \1190 );
not \U$945 ( \1192 , \982 );
not \U$946 ( \1193 , \979 );
or \U$947 ( \1194 , \1192 , \1193 );
not \U$948 ( \1195 , \1006 );
nand \U$949 ( \1196 , \1195 , \287 );
nand \U$950 ( \1197 , \1194 , \1196 );
not \U$951 ( \1198 , \1197 );
buf \U$952 ( \1199 , \970 );
not \U$953 ( \1200 , \1199 );
nand \U$954 ( \1201 , \967 , \1200 );
and \U$955 ( \1202 , \1201 , RIbe28930_31);
not \U$956 ( \1203 , \1202 );
or \U$957 ( \1204 , \1198 , \1203 );
or \U$958 ( \1205 , \1202 , \1197 );
nand \U$959 ( \1206 , \1204 , \1205 );
not \U$960 ( \1207 , \1206 );
or \U$961 ( \1208 , \1191 , \1207 );
not \U$962 ( \1209 , \1202 );
nand \U$963 ( \1210 , \1209 , \1197 );
nand \U$964 ( \1211 , \1208 , \1210 );
xor \U$965 ( \1212 , \1186 , \1211 );
xor \U$966 ( \1213 , \1168 , \1177 );
xor \U$967 ( \1214 , \1213 , \1182 );
not \U$968 ( \1215 , \928 );
not \U$969 ( \1216 , \925 );
or \U$970 ( \1217 , \1215 , \1216 );
xor \U$971 ( \1218 , RIbe288b8_30, RIbe28de0_41);
nand \U$972 ( \1219 , \347 , \1218 );
nand \U$973 ( \1220 , \1217 , \1219 );
not \U$974 ( \1221 , \948 );
xor \U$975 ( \1222 , \1220 , \1221 );
not \U$976 ( \1223 , \900 );
not \U$977 ( \1224 , \909 );
or \U$978 ( \1225 , \1223 , \1224 );
not \U$979 ( \1226 , \908 );
xnor \U$980 ( \1227 , RIbe28570_23, RIbe296c8_60);
or \U$981 ( \1228 , \1226 , \1227 );
nand \U$982 ( \1229 , \1225 , \1228 );
xor \U$983 ( \1230 , \1222 , \1229 );
and \U$984 ( \1231 , \1214 , \1230 );
not \U$985 ( \1232 , \1189 );
not \U$986 ( \1233 , \1206 );
or \U$987 ( \1234 , \1232 , \1233 );
or \U$988 ( \1235 , \1206 , \1189 );
nand \U$989 ( \1236 , \1234 , \1235 );
xor \U$990 ( \1237 , \1220 , \1221 );
xor \U$991 ( \1238 , \1237 , \1229 );
and \U$992 ( \1239 , \1236 , \1238 );
and \U$993 ( \1240 , \1214 , \1236 );
or \U$994 ( \1241 , \1231 , \1239 , \1240 );
xor \U$995 ( \1242 , \1212 , \1241 );
xor \U$996 ( \1243 , \1220 , \1221 );
and \U$997 ( \1244 , \1243 , \1229 );
and \U$998 ( \1245 , \1220 , \1221 );
or \U$999 ( \1246 , \1244 , \1245 );
not \U$1000 ( \1247 , \1246 );
not \U$1001 ( \1248 , \1247 );
and \U$1002 ( \1249 , \1061 , \1065 );
and \U$1003 ( \1250 , \885 , RIbe28228_16);
nor \U$1004 ( \1251 , \1249 , \1250 );
not \U$1005 ( \1252 , \1251 );
not \U$1006 ( \1253 , \1252 );
not \U$1007 ( \1254 , \1129 );
not \U$1008 ( \1255 , \1254 );
not \U$1009 ( \1256 , \1227 );
and \U$1010 ( \1257 , \1255 , \1256 );
and \U$1011 ( \1258 , \908 , \1135 );
nor \U$1012 ( \1259 , \1257 , \1258 );
not \U$1013 ( \1260 , \1259 );
xor \U$1014 ( \1261 , RIbe28048_12, RIbe280c0_13);
not \U$1015 ( \1262 , \1261 );
buf \U$1016 ( \1263 , \868 );
not \U$1017 ( \1264 , \1263 );
not \U$1018 ( \1265 , \1264 );
not \U$1019 ( \1266 , \1265 );
or \U$1020 ( \1267 , \1262 , \1266 );
not \U$1021 ( \1268 , \863 );
nand \U$1022 ( \1269 , \1268 , \1057 );
nand \U$1023 ( \1270 , \1267 , \1269 );
not \U$1024 ( \1271 , \1270 );
or \U$1025 ( \1272 , \1260 , \1271 );
or \U$1026 ( \1273 , \1259 , \1270 );
nand \U$1027 ( \1274 , \1272 , \1273 );
not \U$1028 ( \1275 , \1274 );
not \U$1029 ( \1276 , \1275 );
or \U$1030 ( \1277 , \1253 , \1276 );
nand \U$1031 ( \1278 , \1274 , \1251 );
nand \U$1032 ( \1279 , \1277 , \1278 );
not \U$1033 ( \1280 , \1279 );
or \U$1034 ( \1281 , \1248 , \1280 );
or \U$1035 ( \1282 , \1279 , \1247 );
nand \U$1036 ( \1283 , \1281 , \1282 );
buf \U$1037 ( \1284 , \924 );
and \U$1038 ( \1285 , \1284 , \1218 );
and \U$1039 ( \1286 , \514 , \1143 );
nor \U$1040 ( \1287 , \1285 , \1286 );
not \U$1041 ( \1288 , \1287 );
not \U$1042 ( \1289 , \1175 );
not \U$1043 ( \1290 , \361 );
or \U$1044 ( \1291 , \1289 , \1290 );
not \U$1045 ( \1292 , \1105 );
nand \U$1046 ( \1293 , \1292 , \370 );
nand \U$1047 ( \1294 , \1291 , \1293 );
not \U$1048 ( \1295 , \255 );
not \U$1049 ( \1296 , \1295 );
or \U$1050 ( \1297 , \1296 , \1180 );
not \U$1051 ( \1298 , \268 );
not \U$1052 ( \1299 , \1298 );
or \U$1053 ( \1300 , \1299 , \1122 );
nand \U$1054 ( \1301 , \1297 , \1300 );
xor \U$1055 ( \1302 , \1294 , \1301 );
not \U$1056 ( \1303 , \1302 );
or \U$1057 ( \1304 , \1288 , \1303 );
or \U$1058 ( \1305 , \1302 , \1287 );
nand \U$1059 ( \1306 , \1304 , \1305 );
xor \U$1060 ( \1307 , \1283 , \1306 );
and \U$1061 ( \1308 , \1242 , \1307 );
and \U$1062 ( \1309 , \1212 , \1241 );
nor \U$1063 ( \1310 , \1308 , \1309 );
or \U$1064 ( \1311 , \1162 , \1310 );
or \U$1065 ( \1312 , \1075 , \1161 );
nand \U$1066 ( \1313 , \1311 , \1312 );
not \U$1067 ( \1314 , \1313 );
not \U$1068 ( \1315 , \1294 );
not \U$1069 ( \1316 , \1301 );
or \U$1070 ( \1317 , \1315 , \1316 );
or \U$1071 ( \1318 , \1301 , \1294 );
not \U$1072 ( \1319 , \1287 );
nand \U$1073 ( \1320 , \1318 , \1319 );
nand \U$1074 ( \1321 , \1317 , \1320 );
not \U$1075 ( \1322 , \1321 );
not \U$1076 ( \1323 , \1322 );
not \U$1077 ( \1324 , \1261 );
not \U$1078 ( \1325 , \1053 );
not \U$1079 ( \1326 , \1325 );
not \U$1080 ( \1327 , \1326 );
or \U$1081 ( \1328 , \1324 , \1327 );
xnor \U$1082 ( \1329 , RIbe280c0_13, RIbe29380_53);
not \U$1083 ( \1330 , \1329 );
nand \U$1084 ( \1331 , \1330 , \869 );
nand \U$1085 ( \1332 , \1328 , \1331 );
not \U$1086 ( \1333 , \1332 );
not \U$1087 ( \1334 , \1012 );
not \U$1088 ( \1335 , \979 );
or \U$1089 ( \1336 , \1334 , \1335 );
xnor \U$1090 ( \1337 , RIbe28570_23, RIbe29038_46);
not \U$1091 ( \1338 , \1337 );
nand \U$1092 ( \1339 , \1338 , \287 );
nand \U$1093 ( \1340 , \1336 , \1339 );
not \U$1094 ( \1341 , \1340 );
not \U$1095 ( \1342 , \1341 );
or \U$1096 ( \1343 , \1333 , \1342 );
or \U$1097 ( \1344 , \1341 , \1332 );
nand \U$1098 ( \1345 , \1343 , \1344 );
not \U$1099 ( \1346 , \1345 );
and \U$1100 ( \1347 , \466 , \1022 );
and \U$1101 ( \1348 , \902 , \387 );
and \U$1102 ( \1349 , RIbe28750_27, RIbe290b0_47);
nor \U$1103 ( \1350 , \1348 , \1349 );
and \U$1104 ( \1351 , \399 , \1350 );
nor \U$1105 ( \1352 , \1347 , \1351 );
not \U$1106 ( \1353 , \1352 );
and \U$1107 ( \1354 , \1346 , \1353 );
and \U$1108 ( \1355 , \1345 , \1352 );
nor \U$1109 ( \1356 , \1354 , \1355 );
not \U$1110 ( \1357 , \1356 );
or \U$1111 ( \1358 , \1323 , \1357 );
not \U$1112 ( \1359 , \1270 );
not \U$1113 ( \1360 , \1259 );
not \U$1114 ( \1361 , \1360 );
or \U$1115 ( \1362 , \1359 , \1361 );
nand \U$1116 ( \1363 , \1274 , \1252 );
nand \U$1117 ( \1364 , \1362 , \1363 );
nand \U$1118 ( \1365 , \1358 , \1364 );
not \U$1119 ( \1366 , \1356 );
nand \U$1120 ( \1367 , \1366 , \1321 );
nand \U$1121 ( \1368 , \1365 , \1367 );
not \U$1122 ( \1369 , \1368 );
not \U$1123 ( \1370 , \1101 );
not \U$1124 ( \1371 , \1081 );
or \U$1125 ( \1372 , \1370 , \1371 );
nand \U$1126 ( \1373 , \1096 , \1085 );
nand \U$1127 ( \1374 , \1372 , \1373 );
not \U$1128 ( \1375 , \1374 );
not \U$1129 ( \1376 , \1375 );
and \U$1130 ( \1377 , \1369 , \1376 );
and \U$1131 ( \1378 , \1368 , \1375 );
nor \U$1132 ( \1379 , \1377 , \1378 );
xor \U$1133 ( \1380 , \1114 , \1120 );
and \U$1134 ( \1381 , \1380 , \1127 );
and \U$1135 ( \1382 , \1114 , \1120 );
or \U$1136 ( \1383 , \1381 , \1382 );
not \U$1137 ( \1384 , \1158 );
not \U$1138 ( \1385 , \1142 );
and \U$1139 ( \1386 , \1384 , \1385 );
not \U$1140 ( \1387 , \1152 );
nor \U$1141 ( \1388 , \1387 , \1154 );
nor \U$1142 ( \1389 , \1386 , \1388 );
xnor \U$1143 ( \1390 , \1383 , \1389 );
not \U$1144 ( \1391 , \1345 );
or \U$1145 ( \1392 , \1391 , \1352 );
not \U$1146 ( \1393 , \1332 );
or \U$1147 ( \1394 , \1341 , \1393 );
nand \U$1148 ( \1395 , \1392 , \1394 );
xnor \U$1149 ( \1396 , \1390 , \1395 );
xnor \U$1150 ( \1397 , \1379 , \1396 );
not \U$1151 ( \1398 , \1397 );
not \U$1152 ( \1399 , \1306 );
not \U$1153 ( \1400 , \1283 );
or \U$1154 ( \1401 , \1399 , \1400 );
not \U$1155 ( \1402 , \1247 );
nand \U$1156 ( \1403 , \1402 , \1279 );
nand \U$1157 ( \1404 , \1401 , \1403 );
not \U$1158 ( \1405 , \1404 );
not \U$1159 ( \1406 , \1405 );
and \U$1160 ( \1407 , \1211 , \1186 );
and \U$1161 ( \1408 , \1185 , \1099 );
nor \U$1162 ( \1409 , \1407 , \1408 );
not \U$1163 ( \1410 , \1409 );
and \U$1164 ( \1411 , \1406 , \1410 );
and \U$1165 ( \1412 , \1409 , \1404 );
not \U$1166 ( \1413 , \1409 );
and \U$1167 ( \1414 , \1413 , \1405 );
or \U$1168 ( \1415 , \1412 , \1414 );
not \U$1169 ( \1416 , \1356 );
not \U$1170 ( \1417 , \1322 );
not \U$1171 ( \1418 , \1364 );
or \U$1172 ( \1419 , \1417 , \1418 );
or \U$1173 ( \1420 , \1364 , \1322 );
nand \U$1174 ( \1421 , \1419 , \1420 );
not \U$1175 ( \1422 , \1421 );
or \U$1176 ( \1423 , \1416 , \1422 );
or \U$1177 ( \1424 , \1421 , \1356 );
nand \U$1178 ( \1425 , \1423 , \1424 );
and \U$1179 ( \1426 , \1415 , \1425 );
nor \U$1180 ( \1427 , \1411 , \1426 );
not \U$1181 ( \1428 , \1117 );
not \U$1182 ( \1429 , \1086 );
or \U$1183 ( \1430 , \1428 , \1429 );
xnor \U$1184 ( \1431 , RIbe27d78_6, RIbe284f8_22);
not \U$1185 ( \1432 , \1431 );
nand \U$1186 ( \1433 , \1432 , \315 );
nand \U$1187 ( \1434 , \1430 , \1433 );
not \U$1188 ( \1435 , \1434 );
and \U$1189 ( \1436 , RIbe27b98_2, RIbe294e8_56);
and \U$1190 ( \1437 , \1435 , \1436 );
not \U$1191 ( \1438 , \1435 );
not \U$1192 ( \1439 , \1436 );
and \U$1193 ( \1440 , \1438 , \1439 );
nor \U$1194 ( \1441 , \1437 , \1440 );
and \U$1195 ( \1442 , \386 , \1350 );
xor \U$1196 ( \1443 , RIbe28840_29, RIbe290b0_47);
and \U$1197 ( \1444 , \399 , \1443 );
nor \U$1198 ( \1445 , \1442 , \1444 );
and \U$1199 ( \1446 , \1441 , \1445 );
not \U$1200 ( \1447 , \1441 );
not \U$1201 ( \1448 , \1445 );
and \U$1202 ( \1449 , \1447 , \1448 );
nor \U$1203 ( \1450 , \1446 , \1449 );
not \U$1204 ( \1451 , \1450 );
not \U$1205 ( \1452 , \1254 );
and \U$1206 ( \1453 , \1452 , \1140 );
and \U$1207 ( \1454 , \901 , \431 );
and \U$1208 ( \1455 , RIbe28048_12, RIbe296c8_60);
nor \U$1209 ( \1456 , \1454 , \1455 );
and \U$1210 ( \1457 , \908 , \1456 );
nor \U$1211 ( \1458 , \1453 , \1457 );
not \U$1212 ( \1459 , \1458 );
not \U$1213 ( \1460 , \1459 );
not \U$1214 ( \1461 , \979 );
not \U$1215 ( \1462 , \1461 );
not \U$1216 ( \1463 , \1337 );
and \U$1217 ( \1464 , \1462 , \1463 );
not \U$1218 ( \1465 , \287 );
not \U$1219 ( \1466 , RIbe29038_46);
not \U$1220 ( \1467 , RIbe286d8_26);
or \U$1221 ( \1468 , \1466 , \1467 );
or \U$1222 ( \1469 , RIbe286d8_26, RIbe29038_46);
nand \U$1223 ( \1470 , \1468 , \1469 );
nor \U$1224 ( \1471 , \1465 , \1470 );
nor \U$1225 ( \1472 , \1464 , \1471 );
not \U$1226 ( \1473 , \1150 );
not \U$1227 ( \1474 , \925 );
or \U$1228 ( \1475 , \1473 , \1474 );
xor \U$1229 ( \1476 , RIbe28de0_41, RIbe29308_52);
nand \U$1230 ( \1477 , \514 , \1476 );
nand \U$1231 ( \1478 , \1475 , \1477 );
not \U$1232 ( \1479 , \1478 );
and \U$1233 ( \1480 , \1472 , \1479 );
not \U$1234 ( \1481 , \1472 );
and \U$1235 ( \1482 , \1481 , \1478 );
nor \U$1236 ( \1483 , \1480 , \1482 );
not \U$1237 ( \1484 , \1483 );
not \U$1238 ( \1485 , \1484 );
or \U$1239 ( \1486 , \1460 , \1485 );
nand \U$1240 ( \1487 , \1483 , \1458 );
nand \U$1241 ( \1488 , \1486 , \1487 );
not \U$1242 ( \1489 , \1488 );
or \U$1243 ( \1490 , \1451 , \1489 );
or \U$1244 ( \1491 , \1488 , \1450 );
nand \U$1245 ( \1492 , \1490 , \1491 );
not \U$1246 ( \1493 , \359 );
not \U$1247 ( \1494 , \1493 );
not \U$1248 ( \1495 , \1494 );
not \U$1249 ( \1496 , \1112 );
and \U$1250 ( \1497 , \1495 , \1496 );
not \U$1251 ( \1498 , \1172 );
and \U$1252 ( \1499 , RIbe28c78_38, RIbe27c10_3);
not \U$1253 ( \1500 , RIbe28c78_38);
and \U$1254 ( \1501 , \1500 , \363 );
nor \U$1255 ( \1502 , \1499 , \1501 );
and \U$1256 ( \1503 , \1498 , \1502 );
nor \U$1257 ( \1504 , \1497 , \1503 );
not \U$1258 ( \1505 , \1504 );
not \U$1259 ( \1506 , \1124 );
not \U$1260 ( \1507 , \258 );
or \U$1261 ( \1508 , \1506 , \1507 );
or \U$1262 ( \1509 , RIbe27b98_2, RIbe28a98_34);
nand \U$1263 ( \1510 , RIbe27b98_2, RIbe28a98_34);
nand \U$1264 ( \1511 , \1509 , \1510 );
not \U$1265 ( \1512 , \1511 );
nand \U$1266 ( \1513 , \1512 , \269 );
nand \U$1267 ( \1514 , \1508 , \1513 );
or \U$1268 ( \1515 , \863 , \1329 );
not \U$1269 ( \1516 , \869 );
not \U$1270 ( \1517 , RIbe280c0_13);
or \U$1271 ( \1518 , \1516 , \1517 );
nand \U$1272 ( \1519 , \1515 , \1518 );
xor \U$1273 ( \1520 , \1514 , \1519 );
not \U$1274 ( \1521 , \1520 );
or \U$1275 ( \1522 , \1505 , \1521 );
or \U$1276 ( \1523 , \1520 , \1504 );
nand \U$1277 ( \1524 , \1522 , \1523 );
not \U$1278 ( \1525 , \1524 );
and \U$1279 ( \1526 , \1492 , \1525 );
not \U$1280 ( \1527 , \1492 );
and \U$1281 ( \1528 , \1527 , \1524 );
nor \U$1282 ( \1529 , \1526 , \1528 );
and \U$1283 ( \1530 , \1102 , \1160 );
and \U$1284 ( \1531 , \1128 , \1159 );
nor \U$1285 ( \1532 , \1530 , \1531 );
not \U$1286 ( \1533 , \1532 );
xor \U$1287 ( \1534 , \1529 , \1533 );
not \U$1288 ( \1535 , \1534 );
and \U$1289 ( \1536 , \1427 , \1535 );
not \U$1290 ( \1537 , \1427 );
and \U$1291 ( \1538 , \1537 , \1534 );
nor \U$1292 ( \1539 , \1536 , \1538 );
not \U$1293 ( \1540 , \1539 );
not \U$1294 ( \1541 , \1540 );
or \U$1295 ( \1542 , \1398 , \1541 );
not \U$1296 ( \1543 , \1397 );
nand \U$1297 ( \1544 , \1543 , \1539 );
nand \U$1298 ( \1545 , \1542 , \1544 );
not \U$1299 ( \1546 , \1545 );
or \U$1300 ( \1547 , \1314 , \1546 );
not \U$1301 ( \1548 , \1397 );
nand \U$1302 ( \1549 , \1548 , \1540 );
nand \U$1303 ( \1550 , \1547 , \1549 );
not \U$1304 ( \1551 , \1476 );
not \U$1305 ( \1552 , \334 );
or \U$1306 ( \1553 , \1551 , \1552 );
xor \U$1307 ( \1554 , RIbe28c00_37, RIbe28de0_41);
nand \U$1308 ( \1555 , \347 , \1554 );
nand \U$1309 ( \1556 , \1553 , \1555 );
nand \U$1310 ( \1557 , RIbe27b98_2, RIbe288b8_30);
xor \U$1311 ( \1558 , \1556 , \1557 );
not \U$1312 ( \1559 , \1456 );
not \U$1313 ( \1560 , \1132 );
or \U$1314 ( \1561 , \1559 , \1560 );
xor \U$1315 ( \1562 , RIbe29380_53, RIbe296c8_60);
nand \U$1316 ( \1563 , \908 , \1562 );
nand \U$1317 ( \1564 , \1561 , \1563 );
xnor \U$1318 ( \1565 , \1558 , \1564 );
not \U$1319 ( \1566 , \256 );
or \U$1320 ( \1567 , \1566 , \1511 );
or \U$1321 ( \1568 , RIbe27b98_2, RIbe293f8_54);
nand \U$1322 ( \1569 , RIbe27b98_2, RIbe293f8_54);
nand \U$1323 ( \1570 , \1568 , \1569 );
or \U$1324 ( \1571 , \268 , \1570 );
nand \U$1325 ( \1572 , \1567 , \1571 );
not \U$1326 ( \1573 , \869 );
not \U$1327 ( \1574 , \1573 );
not \U$1328 ( \1575 , \862 );
not \U$1329 ( \1576 , \1575 );
or \U$1330 ( \1577 , \1574 , \1576 );
nand \U$1331 ( \1578 , \1577 , RIbe280c0_13);
not \U$1332 ( \1579 , \1578 );
not \U$1333 ( \1580 , \1461 );
not \U$1334 ( \1581 , \1470 );
and \U$1335 ( \1582 , \1580 , \1581 );
buf \U$1336 ( \1583 , \284 );
not \U$1337 ( \1584 , \1583 );
xnor \U$1338 ( \1585 , RIbe27ee0_9, RIbe29038_46);
nor \U$1339 ( \1586 , \1584 , \1585 );
nor \U$1340 ( \1587 , \1582 , \1586 );
not \U$1341 ( \1588 , \1587 );
or \U$1342 ( \1589 , \1579 , \1588 );
or \U$1343 ( \1590 , \1587 , \1578 );
nand \U$1344 ( \1591 , \1589 , \1590 );
xor \U$1345 ( \1592 , \1572 , \1591 );
xor \U$1346 ( \1593 , \1565 , \1592 );
not \U$1347 ( \1594 , \1443 );
not \U$1348 ( \1595 , \466 );
or \U$1349 ( \1596 , \1594 , \1595 );
and \U$1350 ( \1597 , RIbe28570_23, RIbe290b0_47);
nor \U$1351 ( \1598 , RIbe28570_23, RIbe290b0_47);
nor \U$1352 ( \1599 , \1597 , \1598 );
nand \U$1353 ( \1600 , \399 , \1599 );
nand \U$1354 ( \1601 , \1596 , \1600 );
not \U$1355 ( \1602 , \1502 );
not \U$1356 ( \1603 , \936 );
or \U$1357 ( \1604 , \1602 , \1603 );
not \U$1358 ( \1605 , RIbe27c10_3);
not \U$1359 ( \1606 , RIbe28318_18);
and \U$1360 ( \1607 , \1605 , \1606 );
and \U$1361 ( \1608 , RIbe27c10_3, RIbe28318_18);
nor \U$1362 ( \1609 , \1607 , \1608 );
nand \U$1363 ( \1610 , \370 , \1609 );
nand \U$1364 ( \1611 , \1604 , \1610 );
xor \U$1365 ( \1612 , \1601 , \1611 );
not \U$1366 ( \1613 , \300 );
not \U$1367 ( \1614 , \1613 );
or \U$1368 ( \1615 , \1614 , \1431 );
xnor \U$1369 ( \1616 , RIbe27d78_6, RIbe28750_27);
or \U$1370 ( \1617 , \670 , \1616 );
nand \U$1371 ( \1618 , \1615 , \1617 );
xnor \U$1372 ( \1619 , \1612 , \1618 );
xor \U$1373 ( \1620 , \1593 , \1619 );
not \U$1374 ( \1621 , \1524 );
not \U$1375 ( \1622 , \1492 );
or \U$1376 ( \1623 , \1621 , \1622 );
not \U$1377 ( \1624 , \1450 );
nand \U$1378 ( \1625 , \1624 , \1488 );
nand \U$1379 ( \1626 , \1623 , \1625 );
and \U$1380 ( \1627 , \1620 , \1626 );
not \U$1381 ( \1628 , \1620 );
not \U$1382 ( \1629 , \1626 );
and \U$1383 ( \1630 , \1628 , \1629 );
nor \U$1384 ( \1631 , \1627 , \1630 );
not \U$1385 ( \1632 , \1379 );
not \U$1386 ( \1633 , \1396 );
and \U$1387 ( \1634 , \1632 , \1633 );
and \U$1388 ( \1635 , \1368 , \1374 );
nor \U$1389 ( \1636 , \1634 , \1635 );
xor \U$1390 ( \1637 , \1631 , \1636 );
or \U$1391 ( \1638 , \1514 , \1519 );
not \U$1392 ( \1639 , \1504 );
nand \U$1393 ( \1640 , \1638 , \1639 );
nand \U$1394 ( \1641 , \1514 , \1519 );
and \U$1395 ( \1642 , \1640 , \1641 );
xor \U$1396 ( \1643 , \1435 , \1642 );
or \U$1397 ( \1644 , \1484 , \1458 );
or \U$1398 ( \1645 , \1472 , \1479 );
nand \U$1399 ( \1646 , \1644 , \1645 );
xnor \U$1400 ( \1647 , \1643 , \1646 );
not \U$1401 ( \1648 , \1395 );
not \U$1402 ( \1649 , \1390 );
or \U$1403 ( \1650 , \1648 , \1649 );
not \U$1404 ( \1651 , \1389 );
nand \U$1405 ( \1652 , \1651 , \1383 );
nand \U$1406 ( \1653 , \1650 , \1652 );
not \U$1407 ( \1654 , \1653 );
and \U$1408 ( \1655 , \1448 , \1441 );
and \U$1409 ( \1656 , \1435 , \1436 );
nor \U$1410 ( \1657 , \1655 , \1656 );
not \U$1411 ( \1658 , \1657 );
and \U$1412 ( \1659 , \1654 , \1658 );
and \U$1413 ( \1660 , \1653 , \1657 );
nor \U$1414 ( \1661 , \1659 , \1660 );
xor \U$1415 ( \1662 , \1647 , \1661 );
xor \U$1416 ( \1663 , \1637 , \1662 );
or \U$1417 ( \1664 , \1427 , \1534 );
or \U$1418 ( \1665 , \1529 , \1532 );
nand \U$1419 ( \1666 , \1664 , \1665 );
xor \U$1420 ( \1667 , \1663 , \1666 );
nor \U$1421 ( \1668 , \1550 , \1667 );
not \U$1422 ( \1669 , \1668 );
and \U$1423 ( \1670 , \1545 , \1313 );
not \U$1424 ( \1671 , \1545 );
not \U$1425 ( \1672 , \1313 );
and \U$1426 ( \1673 , \1671 , \1672 );
nor \U$1427 ( \1674 , \1670 , \1673 );
not \U$1428 ( \1675 , \1674 );
xor \U$1429 ( \1676 , \1220 , \1221 );
xor \U$1430 ( \1677 , \1676 , \1229 );
xor \U$1431 ( \1678 , \1214 , \1236 );
xor \U$1432 ( \1679 , \1677 , \1678 );
not \U$1433 ( \1680 , \1679 );
xnor \U$1434 ( \1681 , \996 , \975 );
xor \U$1435 ( \1682 , \875 , \893 );
xor \U$1436 ( \1683 , \1682 , \911 );
nand \U$1437 ( \1684 , \1681 , \1683 );
xor \U$1438 ( \1685 , \930 , \944 );
xor \U$1439 ( \1686 , \1685 , \957 );
and \U$1440 ( \1687 , \1684 , \1686 );
nor \U$1441 ( \1688 , \1681 , \1683 );
nor \U$1442 ( \1689 , \1687 , \1688 );
not \U$1443 ( \1690 , \1689 );
xnor \U$1444 ( \1691 , \914 , \1001 );
not \U$1445 ( \1692 , \1691 );
or \U$1446 ( \1693 , \1690 , \1692 );
or \U$1447 ( \1694 , \1691 , \1689 );
nand \U$1448 ( \1695 , \1693 , \1694 );
not \U$1449 ( \1696 , \1695 );
or \U$1450 ( \1697 , \1680 , \1696 );
not \U$1451 ( \1698 , \1689 );
nand \U$1452 ( \1699 , \1698 , \1691 );
nand \U$1453 ( \1700 , \1697 , \1699 );
not \U$1454 ( \1701 , \1700 );
and \U$1455 ( \1702 , \1005 , \1072 );
not \U$1456 ( \1703 , \1005 );
not \U$1457 ( \1704 , \1072 );
and \U$1458 ( \1705 , \1703 , \1704 );
nor \U$1459 ( \1706 , \1702 , \1705 );
not \U$1460 ( \1707 , \1706 );
xnor \U$1461 ( \1708 , \1060 , \1067 );
not \U$1462 ( \1709 , RIbe282a0_17);
not \U$1463 ( \1710 , RIbe28de0_41);
and \U$1464 ( \1711 , \1709 , \1710 );
and \U$1465 ( \1712 , RIbe282a0_17, RIbe28de0_41);
nor \U$1466 ( \1713 , \1711 , \1712 );
and \U$1467 ( \1714 , \1284 , \1713 );
and \U$1468 ( \1715 , \514 , \921 );
nor \U$1469 ( \1716 , \1714 , \1715 );
nand \U$1470 ( \1717 , RIbe27b98_2, RIbe29740_61);
xor \U$1471 ( \1718 , \1716 , \1717 );
and \U$1472 ( \1719 , RIbe284f8_22, RIbe296c8_60);
nor \U$1473 ( \1720 , RIbe284f8_22, RIbe296c8_60);
nor \U$1474 ( \1721 , \1719 , \1720 );
and \U$1475 ( \1722 , \1452 , \1721 );
and \U$1476 ( \1723 , \908 , \905 );
nor \U$1477 ( \1724 , \1722 , \1723 );
and \U$1478 ( \1725 , \1718 , \1724 );
and \U$1479 ( \1726 , \1716 , \1717 );
nor \U$1480 ( \1727 , \1725 , \1726 );
and \U$1481 ( \1728 , RIbe27b98_2, RIbe297b8_62);
xor \U$1482 ( \1729 , \1728 , \1051 );
and \U$1483 ( \1730 , \1727 , \1729 );
and \U$1484 ( \1731 , \1051 , \1728 );
nor \U$1485 ( \1732 , \1730 , \1731 );
xor \U$1486 ( \1733 , \1708 , \1732 );
buf \U$1487 ( \1734 , \267 );
not \U$1488 ( \1735 , \1734 );
not \U$1489 ( \1736 , \1735 );
not \U$1490 ( \1737 , \949 );
and \U$1491 ( \1738 , \1736 , \1737 );
not \U$1492 ( \1739 , RIbe27b98_2);
not \U$1493 ( \1740 , RIbe297b8_62);
and \U$1494 ( \1741 , \1739 , \1740 );
nor \U$1495 ( \1742 , \1741 , \1728 );
and \U$1496 ( \1743 , \546 , \1742 );
nor \U$1497 ( \1744 , \1738 , \1743 );
not \U$1498 ( \1745 , \1093 );
not \U$1499 ( \1746 , \1049 );
not \U$1500 ( \1747 , \1746 );
and \U$1501 ( \1748 , \1745 , \1747 );
not \U$1502 ( \1749 , RIbe27d78_6);
not \U$1503 ( \1750 , RIbe28a98_34);
and \U$1504 ( \1751 , \1749 , \1750 );
and \U$1505 ( \1752 , RIbe27d78_6, RIbe28a98_34);
nor \U$1506 ( \1753 , \1751 , \1752 );
and \U$1507 ( \1754 , \1044 , \1753 );
nor \U$1508 ( \1755 , \1748 , \1754 );
xnor \U$1509 ( \1756 , \1744 , \1755 );
and \U$1510 ( \1757 , RIbe294e8_56, RIbe27c10_3);
not \U$1511 ( \1758 , RIbe294e8_56);
and \U$1512 ( \1759 , \1758 , \363 );
nor \U$1513 ( \1760 , \1757 , \1759 );
and \U$1514 ( \1761 , \361 , \1760 );
and \U$1515 ( \1762 , \370 , \934 );
nor \U$1516 ( \1763 , \1761 , \1762 );
or \U$1517 ( \1764 , \1756 , \1763 );
or \U$1518 ( \1765 , \1744 , \1755 );
nand \U$1519 ( \1766 , \1764 , \1765 );
xor \U$1520 ( \1767 , RIbe28b88_36, RIbe29290_51);
buf \U$1521 ( \1768 , \1767 );
buf \U$1522 ( \1769 , \1768 );
not \U$1523 ( \1770 , \1769 );
not \U$1524 ( \1771 , \1770 );
nor \U$1525 ( \1772 , RIbe28a20_33, RIbe28b88_36);
not \U$1526 ( \1773 , \1772 );
and \U$1527 ( \1774 , RIbe29290_51, RIbe28a20_33);
not \U$1528 ( \1775 , RIbe29290_51);
and \U$1529 ( \1776 , \1775 , RIbe28b88_36);
nor \U$1530 ( \1777 , \1774 , \1776 );
nand \U$1531 ( \1778 , \1773 , \1777 );
not \U$1532 ( \1779 , \1778 );
buf \U$1533 ( \1780 , \1779 );
buf \U$1534 ( \1781 , \1780 );
not \U$1535 ( \1782 , \1781 );
not \U$1536 ( \1783 , \1782 );
or \U$1537 ( \1784 , \1771 , \1783 );
nand \U$1538 ( \1785 , \1784 , RIbe28a20_33);
not \U$1539 ( \1786 , \1785 );
not \U$1540 ( \1787 , RIbe28048_12);
not \U$1541 ( \1788 , RIbe28930_31);
and \U$1542 ( \1789 , \1787 , \1788 );
and \U$1543 ( \1790 , RIbe28048_12, RIbe28930_31);
nor \U$1544 ( \1791 , \1789 , \1790 );
not \U$1545 ( \1792 , \1791 );
buf \U$1546 ( \1793 , \965 );
not \U$1547 ( \1794 , \1793 );
or \U$1548 ( \1795 , \1792 , \1794 );
not \U$1549 ( \1796 , \968 );
buf \U$1550 ( \1797 , \970 );
nand \U$1551 ( \1798 , \1796 , \1797 );
nand \U$1552 ( \1799 , \1795 , \1798 );
not \U$1553 ( \1800 , \1799 );
and \U$1554 ( \1801 , RIbe28c78_38, RIbe29038_46);
nor \U$1555 ( \1802 , RIbe28c78_38, RIbe29038_46);
nor \U$1556 ( \1803 , \1801 , \1802 );
and \U$1557 ( \1804 , \979 , \1803 );
buf \U$1558 ( \1805 , \1583 );
and \U$1559 ( \1806 , \1805 , \977 );
nor \U$1560 ( \1807 , \1804 , \1806 );
not \U$1561 ( \1808 , \1807 );
or \U$1562 ( \1809 , \1800 , \1808 );
or \U$1563 ( \1810 , \1807 , \1799 );
nand \U$1564 ( \1811 , \1809 , \1810 );
not \U$1565 ( \1812 , \1811 );
or \U$1566 ( \1813 , \1786 , \1812 );
not \U$1567 ( \1814 , \1807 );
nand \U$1568 ( \1815 , \1814 , \1799 );
nand \U$1569 ( \1816 , \1813 , \1815 );
not \U$1570 ( \1817 , \1816 );
and \U$1571 ( \1818 , RIbe280c0_13, RIbe28840_29);
not \U$1572 ( \1819 , RIbe280c0_13);
and \U$1573 ( \1820 , \1819 , \364 );
nor \U$1574 ( \1821 , \1818 , \1820 );
not \U$1575 ( \1822 , \1821 );
not \U$1576 ( \1823 , \1054 );
or \U$1577 ( \1824 , \1822 , \1823 );
not \U$1578 ( \1825 , \865 );
nand \U$1579 ( \1826 , \1825 , \869 );
nand \U$1580 ( \1827 , \1824 , \1826 );
xor \U$1581 ( \1828 , RIbe290b0_47, RIbe29308_52);
not \U$1582 ( \1829 , \1828 );
not \U$1583 ( \1830 , \466 );
or \U$1584 ( \1831 , \1829 , \1830 );
nand \U$1585 ( \1832 , \399 , \985 );
nand \U$1586 ( \1833 , \1831 , \1832 );
xor \U$1587 ( \1834 , \1827 , \1833 );
not \U$1588 ( \1835 , \1061 );
and \U$1589 ( \1836 , \304 , RIbe28228_16);
and \U$1590 ( \1837 , \888 , RIbe286d8_26);
nor \U$1591 ( \1838 , \1836 , \1837 );
or \U$1592 ( \1839 , \1835 , \1838 );
or \U$1593 ( \1840 , \886 , \882 );
nand \U$1594 ( \1841 , \1839 , \1840 );
and \U$1595 ( \1842 , \1834 , \1841 );
and \U$1596 ( \1843 , \1827 , \1833 );
nor \U$1597 ( \1844 , \1842 , \1843 );
not \U$1598 ( \1845 , \1844 );
or \U$1599 ( \1846 , \1817 , \1845 );
or \U$1600 ( \1847 , \1816 , \1844 );
nand \U$1601 ( \1848 , \1846 , \1847 );
and \U$1602 ( \1849 , \1766 , \1848 );
not \U$1603 ( \1850 , \1816 );
nor \U$1604 ( \1851 , \1850 , \1844 );
nor \U$1605 ( \1852 , \1849 , \1851 );
and \U$1606 ( \1853 , \1733 , \1852 );
and \U$1607 ( \1854 , \1708 , \1732 );
or \U$1608 ( \1855 , \1853 , \1854 );
not \U$1609 ( \1856 , \1855 );
or \U$1610 ( \1857 , \1707 , \1856 );
or \U$1611 ( \1858 , \1706 , \1855 );
nand \U$1612 ( \1859 , \1857 , \1858 );
not \U$1613 ( \1860 , \1859 );
or \U$1614 ( \1861 , \1701 , \1860 );
not \U$1615 ( \1862 , \1855 );
nand \U$1616 ( \1863 , \1862 , \1706 );
nand \U$1617 ( \1864 , \1861 , \1863 );
xor \U$1618 ( \1865 , \1415 , \1425 );
and \U$1619 ( \1866 , \1864 , \1865 );
xor \U$1620 ( \1867 , \1162 , \1310 );
xor \U$1621 ( \1868 , \1865 , \1864 );
and \U$1622 ( \1869 , \1867 , \1868 );
nor \U$1623 ( \1870 , \1866 , \1869 );
nand \U$1624 ( \1871 , \1675 , \1870 );
and \U$1625 ( \1872 , \1669 , \1871 );
or \U$1626 ( \1873 , \1647 , \1661 );
not \U$1627 ( \1874 , \1653 );
or \U$1628 ( \1875 , \1874 , \1657 );
nand \U$1629 ( \1876 , \1873 , \1875 );
not \U$1630 ( \1877 , \1572 );
not \U$1631 ( \1878 , \1591 );
or \U$1632 ( \1879 , \1877 , \1878 );
not \U$1633 ( \1880 , \1587 );
nand \U$1634 ( \1881 , \1880 , \1578 );
nand \U$1635 ( \1882 , \1879 , \1881 );
not \U$1636 ( \1883 , \1564 );
xnor \U$1637 ( \1884 , \1556 , \1557 );
not \U$1638 ( \1885 , \1884 );
or \U$1639 ( \1886 , \1883 , \1885 );
not \U$1640 ( \1887 , \1557 );
nand \U$1641 ( \1888 , \1887 , \1556 );
nand \U$1642 ( \1889 , \1886 , \1888 );
xor \U$1643 ( \1890 , \1882 , \1889 );
xor \U$1644 ( \1891 , RIbe27b98_2, RIbe29308_52);
not \U$1645 ( \1892 , \1891 );
not \U$1646 ( \1893 , \1298 );
or \U$1647 ( \1894 , \1892 , \1893 );
not \U$1648 ( \1895 , \1570 );
nand \U$1649 ( \1896 , \1895 , \256 );
nand \U$1650 ( \1897 , \1894 , \1896 );
xor \U$1651 ( \1898 , RIbe28c78_38, RIbe28de0_41);
not \U$1652 ( \1899 , \1898 );
not \U$1653 ( \1900 , \514 );
or \U$1654 ( \1901 , \1899 , \1900 );
nand \U$1655 ( \1902 , \1284 , \1554 );
nand \U$1656 ( \1903 , \1901 , \1902 );
xnor \U$1657 ( \1904 , \1897 , \1903 );
and \U$1658 ( \1905 , \466 , \1599 );
xor \U$1659 ( \1906 , RIbe286d8_26, RIbe290b0_47);
and \U$1660 ( \1907 , \469 , \1906 );
nor \U$1661 ( \1908 , \1905 , \1907 );
xor \U$1662 ( \1909 , \1904 , \1908 );
and \U$1663 ( \1910 , \1890 , \1909 );
not \U$1664 ( \1911 , \1890 );
not \U$1665 ( \1912 , \1909 );
and \U$1666 ( \1913 , \1911 , \1912 );
nor \U$1667 ( \1914 , \1910 , \1913 );
and \U$1668 ( \1915 , \1884 , \1564 );
not \U$1669 ( \1916 , \1884 );
not \U$1670 ( \1917 , \1564 );
and \U$1671 ( \1918 , \1916 , \1917 );
or \U$1672 ( \1919 , \1915 , \1918 );
not \U$1673 ( \1920 , \1919 );
not \U$1674 ( \1921 , \1920 );
not \U$1675 ( \1922 , \1592 );
or \U$1676 ( \1923 , \1921 , \1922 );
not \U$1677 ( \1924 , \1619 );
xnor \U$1678 ( \1925 , \1919 , \1592 );
nand \U$1679 ( \1926 , \1924 , \1925 );
nand \U$1680 ( \1927 , \1923 , \1926 );
xor \U$1681 ( \1928 , \1914 , \1927 );
and \U$1682 ( \1929 , \1876 , \1928 );
not \U$1683 ( \1930 , \1876 );
not \U$1684 ( \1931 , \1928 );
and \U$1685 ( \1932 , \1930 , \1931 );
nor \U$1686 ( \1933 , \1929 , \1932 );
not \U$1687 ( \1934 , \1562 );
not \U$1688 ( \1935 , \1132 );
or \U$1689 ( \1936 , \1934 , \1935 );
buf \U$1690 ( \1937 , \895 );
not \U$1691 ( \1938 , \1937 );
not \U$1692 ( \1939 , \1938 );
nand \U$1693 ( \1940 , \1939 , RIbe296c8_60);
nand \U$1694 ( \1941 , \1936 , \1940 );
not \U$1695 ( \1942 , \360 );
not \U$1696 ( \1943 , \1609 );
not \U$1697 ( \1944 , \1943 );
and \U$1698 ( \1945 , \1942 , \1944 );
xor \U$1699 ( \1946 , RIbe27c10_3, RIbe284f8_22);
and \U$1700 ( \1947 , \370 , \1946 );
nor \U$1701 ( \1948 , \1945 , \1947 );
nand \U$1702 ( \1949 , \1941 , \1948 );
not \U$1703 ( \1950 , \1949 );
nor \U$1704 ( \1951 , \1941 , \1948 );
nor \U$1705 ( \1952 , \1950 , \1951 );
not \U$1706 ( \1953 , \1952 );
or \U$1707 ( \1954 , \1611 , \1601 );
nand \U$1708 ( \1955 , \1954 , \1618 );
nand \U$1709 ( \1956 , \1601 , \1611 );
nand \U$1710 ( \1957 , \1955 , \1956 );
not \U$1711 ( \1958 , \1957 );
and \U$1712 ( \1959 , \1953 , \1958 );
and \U$1713 ( \1960 , \1957 , \1952 );
nor \U$1714 ( \1961 , \1959 , \1960 );
not \U$1715 ( \1962 , \1510 );
xor \U$1716 ( \1963 , RIbe27d78_6, RIbe28840_29);
not \U$1717 ( \1964 , \1963 );
not \U$1718 ( \1965 , \314 );
or \U$1719 ( \1966 , \1964 , \1965 );
or \U$1720 ( \1967 , \301 , \1616 );
nand \U$1721 ( \1968 , \1966 , \1967 );
not \U$1722 ( \1969 , \1968 );
not \U$1723 ( \1970 , \1461 );
not \U$1724 ( \1971 , \1585 );
and \U$1725 ( \1972 , \1970 , \1971 );
and \U$1726 ( \1973 , RIbe28048_12, RIbe29038_46);
nor \U$1727 ( \1974 , RIbe28048_12, RIbe29038_46);
nor \U$1728 ( \1975 , \1973 , \1974 );
and \U$1729 ( \1976 , \1583 , \1975 );
nor \U$1730 ( \1977 , \1972 , \1976 );
not \U$1731 ( \1978 , \1977 );
or \U$1732 ( \1979 , \1969 , \1978 );
or \U$1733 ( \1980 , \1977 , \1968 );
nand \U$1734 ( \1981 , \1979 , \1980 );
not \U$1735 ( \1982 , \1981 );
or \U$1736 ( \1983 , \1962 , \1982 );
or \U$1737 ( \1984 , \1981 , \1510 );
nand \U$1738 ( \1985 , \1983 , \1984 );
xor \U$1739 ( \1986 , \1961 , \1985 );
not \U$1740 ( \1987 , \1646 );
not \U$1741 ( \1988 , \1643 );
or \U$1742 ( \1989 , \1987 , \1988 );
or \U$1743 ( \1990 , \1642 , \1435 );
nand \U$1744 ( \1991 , \1989 , \1990 );
xor \U$1745 ( \1992 , \1986 , \1991 );
and \U$1746 ( \1993 , \1933 , \1992 );
not \U$1747 ( \1994 , \1933 );
not \U$1748 ( \1995 , \1992 );
and \U$1749 ( \1996 , \1994 , \1995 );
nor \U$1750 ( \1997 , \1993 , \1996 );
or \U$1751 ( \1998 , \1631 , \1636 );
or \U$1752 ( \1999 , \1629 , \1620 );
nand \U$1753 ( \2000 , \1998 , \1999 );
and \U$1754 ( \2001 , \1997 , \2000 );
and \U$1755 ( \2002 , \1933 , \1992 );
nor \U$1756 ( \2003 , \2001 , \2002 );
not \U$1757 ( \2004 , \1909 );
not \U$1758 ( \2005 , \1890 );
or \U$1759 ( \2006 , \2004 , \2005 );
nand \U$1760 ( \2007 , \1882 , \1889 );
nand \U$1761 ( \2008 , \2006 , \2007 );
not \U$1762 ( \2009 , \2008 );
not \U$1763 ( \2010 , \1510 );
or \U$1764 ( \2011 , \1968 , \2010 );
not \U$1765 ( \2012 , \1977 );
nand \U$1766 ( \2013 , \2011 , \2012 );
nand \U$1767 ( \2014 , \1968 , \2010 );
and \U$1768 ( \2015 , \2013 , \2014 );
not \U$1769 ( \2016 , \2015 );
not \U$1770 ( \2017 , \2016 );
not \U$1771 ( \2018 , \1137 );
not \U$1772 ( \2019 , \2018 );
not \U$1773 ( \2020 , \1132 );
not \U$1774 ( \2021 , \2020 );
or \U$1775 ( \2022 , \2019 , \2021 );
nand \U$1776 ( \2023 , \2022 , RIbe296c8_60);
not \U$1777 ( \2024 , \1898 );
not \U$1778 ( \2025 , \1145 );
or \U$1779 ( \2026 , \2024 , \2025 );
nand \U$1780 ( \2027 , \1149 , \510 );
nand \U$1781 ( \2028 , \2026 , \2027 );
xor \U$1782 ( \2029 , \2023 , \2028 );
not \U$1783 ( \2030 , \1569 );
xor \U$1784 ( \2031 , \2029 , \2030 );
not \U$1785 ( \2032 , \2031 );
not \U$1786 ( \2033 , \2032 );
or \U$1787 ( \2034 , \2017 , \2033 );
nand \U$1788 ( \2035 , \2031 , \2015 );
nand \U$1789 ( \2036 , \2034 , \2035 );
not \U$1790 ( \2037 , \1904 );
not \U$1791 ( \2038 , \1908 );
and \U$1792 ( \2039 , \2037 , \2038 );
and \U$1793 ( \2040 , \1897 , \1903 );
nor \U$1794 ( \2041 , \2039 , \2040 );
xor \U$1795 ( \2042 , \2036 , \2041 );
not \U$1796 ( \2043 , \2042 );
or \U$1797 ( \2044 , \2009 , \2043 );
or \U$1798 ( \2045 , \2042 , \2008 );
nand \U$1799 ( \2046 , \2044 , \2045 );
xor \U$1800 ( \2047 , \1961 , \1985 );
and \U$1801 ( \2048 , \2047 , \1991 );
and \U$1802 ( \2049 , \1961 , \1985 );
or \U$1803 ( \2050 , \2048 , \2049 );
xor \U$1804 ( \2051 , \2046 , \2050 );
not \U$1805 ( \2052 , \1115 );
and \U$1806 ( \2053 , \2052 , \1963 );
and \U$1807 ( \2054 , \314 , \554 );
nor \U$1808 ( \2055 , \2053 , \2054 );
and \U$1809 ( \2056 , \546 , \1891 );
and \U$1810 ( \2057 , \1298 , \549 );
nor \U$1811 ( \2058 , \2056 , \2057 );
xor \U$1812 ( \2059 , \2055 , \2058 );
not \U$1813 ( \2060 , \1941 );
xor \U$1814 ( \2061 , \2059 , \2060 );
not \U$1815 ( \2062 , \1946 );
not \U$1816 ( \2063 , \1494 );
not \U$1817 ( \2064 , \2063 );
or \U$1818 ( \2065 , \2062 , \2064 );
nand \U$1819 ( \2066 , \370 , \563 );
nand \U$1820 ( \2067 , \2065 , \2066 );
not \U$1821 ( \2068 , \1906 );
not \U$1822 ( \2069 , \466 );
or \U$1823 ( \2070 , \2068 , \2069 );
not \U$1824 ( \2071 , \468 );
nand \U$1825 ( \2072 , \2071 , \526 );
nand \U$1826 ( \2073 , \2070 , \2072 );
xor \U$1827 ( \2074 , \2067 , \2073 );
not \U$1828 ( \2075 , \1975 );
not \U$1829 ( \2076 , \979 );
or \U$1830 ( \2077 , \2075 , \2076 );
nand \U$1831 ( \2078 , \1583 , \492 );
nand \U$1832 ( \2079 , \2077 , \2078 );
xnor \U$1833 ( \2080 , \2074 , \2079 );
xnor \U$1834 ( \2081 , \2061 , \2080 );
and \U$1835 ( \2082 , \1957 , \1949 );
nor \U$1836 ( \2083 , \2082 , \1951 );
xor \U$1837 ( \2084 , \2081 , \2083 );
xor \U$1838 ( \2085 , \2051 , \2084 );
and \U$1839 ( \2086 , \1876 , \1928 );
and \U$1840 ( \2087 , \1914 , \1927 );
nor \U$1841 ( \2088 , \2086 , \2087 );
and \U$1842 ( \2089 , \2085 , \2088 );
not \U$1843 ( \2090 , \2085 );
not \U$1844 ( \2091 , \2088 );
and \U$1845 ( \2092 , \2090 , \2091 );
nor \U$1846 ( \2093 , \2089 , \2092 );
nand \U$1847 ( \2094 , \2003 , \2093 );
xnor \U$1848 ( \2095 , \1997 , \2000 );
xor \U$1849 ( \2096 , \1637 , \1662 );
and \U$1850 ( \2097 , \2096 , \1666 );
and \U$1851 ( \2098 , \1637 , \1662 );
nor \U$1852 ( \2099 , \2097 , \2098 );
nand \U$1853 ( \2100 , \2095 , \2099 );
and \U$1854 ( \2101 , \1872 , \2094 , \2100 );
and \U$1855 ( \2102 , \2085 , \2091 );
and \U$1856 ( \2103 , \2051 , \2084 );
nor \U$1857 ( \2104 , \2102 , \2103 );
not \U$1858 ( \2105 , \2050 );
not \U$1859 ( \2106 , \2046 );
or \U$1860 ( \2107 , \2105 , \2106 );
not \U$1861 ( \2108 , \2008 );
or \U$1862 ( \2109 , \2108 , \2042 );
nand \U$1863 ( \2110 , \2107 , \2109 );
or \U$1864 ( \2111 , \2081 , \2083 );
or \U$1865 ( \2112 , \2061 , \2080 );
nand \U$1866 ( \2113 , \2111 , \2112 );
xor \U$1867 ( \2114 , \2110 , \2113 );
not \U$1868 ( \2115 , \2036 );
or \U$1869 ( \2116 , \2115 , \2041 );
or \U$1870 ( \2117 , \2032 , \2015 );
nand \U$1871 ( \2118 , \2116 , \2117 );
not \U$1872 ( \2119 , \2073 );
not \U$1873 ( \2120 , \2079 );
or \U$1874 ( \2121 , \2119 , \2120 );
or \U$1875 ( \2122 , \2079 , \2073 );
nand \U$1876 ( \2123 , \2122 , \2067 );
nand \U$1877 ( \2124 , \2121 , \2123 );
not \U$1878 ( \2125 , \2124 );
and \U$1879 ( \2126 , \2125 , \536 );
and \U$1880 ( \2127 , \2124 , \497 );
nor \U$1881 ( \2128 , \2126 , \2127 );
xor \U$1882 ( \2129 , \2023 , \2028 );
not \U$1883 ( \2130 , \1569 );
and \U$1884 ( \2131 , \2129 , \2130 );
and \U$1885 ( \2132 , \2023 , \2028 );
or \U$1886 ( \2133 , \2131 , \2132 );
not \U$1887 ( \2134 , \2133 );
xor \U$1888 ( \2135 , \2128 , \2134 );
xor \U$1889 ( \2136 , \2118 , \2135 );
xnor \U$1890 ( \2137 , \522 , \529 );
xor \U$1891 ( \2138 , \2055 , \2058 );
and \U$1892 ( \2139 , \2138 , \2060 );
and \U$1893 ( \2140 , \2055 , \2058 );
or \U$1894 ( \2141 , \2139 , \2140 );
xnor \U$1895 ( \2142 , \2137 , \2141 );
xor \U$1896 ( \2143 , \551 , \557 );
xor \U$1897 ( \2144 , \2143 , \566 );
xor \U$1898 ( \2145 , \2142 , \2144 );
xor \U$1899 ( \2146 , \2136 , \2145 );
xnor \U$1900 ( \2147 , \2114 , \2146 );
nand \U$1901 ( \2148 , \2104 , \2147 );
xor \U$1902 ( \2149 , \533 , \508 );
or \U$1903 ( \2150 , \2128 , \2134 );
or \U$1904 ( \2151 , \2125 , \497 );
nand \U$1905 ( \2152 , \2150 , \2151 );
xor \U$1906 ( \2153 , \2149 , \2152 );
or \U$1907 ( \2154 , \2142 , \2144 );
or \U$1908 ( \2155 , \2137 , \2141 );
nand \U$1909 ( \2156 , \2154 , \2155 );
xor \U$1910 ( \2157 , \2153 , \2156 );
xor \U$1911 ( \2158 , \569 , \570 );
xor \U$1912 ( \2159 , \2158 , \572 );
xor \U$1913 ( \2160 , \2157 , \2159 );
and \U$1914 ( \2161 , \2136 , \2145 );
and \U$1915 ( \2162 , \2118 , \2135 );
nor \U$1916 ( \2163 , \2161 , \2162 );
and \U$1917 ( \2164 , \2160 , \2163 );
not \U$1918 ( \2165 , \2160 );
not \U$1919 ( \2166 , \2163 );
and \U$1920 ( \2167 , \2165 , \2166 );
nor \U$1921 ( \2168 , \2164 , \2167 );
and \U$1922 ( \2169 , \2114 , \2146 );
and \U$1923 ( \2170 , \2110 , \2113 );
nor \U$1924 ( \2171 , \2169 , \2170 );
nand \U$1925 ( \2172 , \2168 , \2171 );
and \U$1926 ( \2173 , \2148 , \2172 );
and \U$1927 ( \2174 , \2160 , \2166 );
and \U$1928 ( \2175 , \2157 , \2159 );
nor \U$1929 ( \2176 , \2174 , \2175 );
xor \U$1930 ( \2177 , \380 , \409 );
and \U$1931 ( \2178 , \2153 , \2156 );
and \U$1932 ( \2179 , \2149 , \2152 );
nor \U$1933 ( \2180 , \2178 , \2179 );
not \U$1934 ( \2181 , \2180 );
and \U$1935 ( \2182 , \2177 , \2181 );
not \U$1936 ( \2183 , \2177 );
and \U$1937 ( \2184 , \2183 , \2180 );
nor \U$1938 ( \2185 , \2182 , \2184 );
and \U$1939 ( \2186 , \429 , \436 );
not \U$1940 ( \2187 , \429 );
and \U$1941 ( \2188 , \2187 , \461 );
nor \U$1942 ( \2189 , \2186 , \2188 );
xor \U$1943 ( \2190 , \2189 , \538 );
xor \U$1944 ( \2191 , \2190 , \575 );
xnor \U$1945 ( \2192 , \2185 , \2191 );
nand \U$1946 ( \2193 , \2176 , \2192 );
and \U$1947 ( \2194 , \2173 , \2193 );
and \U$1948 ( \2195 , \2185 , \2191 );
and \U$1949 ( \2196 , \2181 , \2177 );
nor \U$1950 ( \2197 , \2195 , \2196 );
xor \U$1951 ( \2198 , \412 , \488 );
not \U$1952 ( \2199 , \580 );
xor \U$1953 ( \2200 , \2198 , \2199 );
nand \U$1954 ( \2201 , \2197 , \2200 );
and \U$1955 ( \2202 , \2101 , \2194 , \2201 );
not \U$1956 ( \2203 , \2202 );
xnor \U$1957 ( \2204 , \1859 , \1700 );
xnor \U$1958 ( \2205 , \1242 , \1307 );
xor \U$1959 ( \2206 , \2204 , \2205 );
not \U$1960 ( \2207 , RIbe28138_14);
not \U$1961 ( \2208 , RIbe28de0_41);
and \U$1962 ( \2209 , \2207 , \2208 );
and \U$1963 ( \2210 , RIbe28138_14, RIbe28de0_41);
nor \U$1964 ( \2211 , \2209 , \2210 );
and \U$1965 ( \2212 , \1284 , \2211 );
and \U$1966 ( \2213 , \349 , \1713 );
nor \U$1967 ( \2214 , \2212 , \2213 );
and \U$1968 ( \2215 , RIbe290b0_47, RIbe293f8_54);
nor \U$1969 ( \2216 , RIbe290b0_47, RIbe293f8_54);
nor \U$1970 ( \2217 , \2215 , \2216 );
not \U$1971 ( \2218 , \2217 );
nor \U$1972 ( \2219 , \2218 , \524 );
and \U$1973 ( \2220 , \399 , \1828 );
nor \U$1974 ( \2221 , \2219 , \2220 );
xor \U$1975 ( \2222 , \2214 , \2221 );
and \U$1976 ( \2223 , \363 , \919 );
and \U$1977 ( \2224 , RIbe27c10_3, RIbe29470_55);
nor \U$1978 ( \2225 , \2223 , \2224 );
and \U$1979 ( \2226 , \361 , \2225 );
and \U$1980 ( \2227 , \370 , \1760 );
nor \U$1981 ( \2228 , \2226 , \2227 );
and \U$1982 ( \2229 , \2222 , \2228 );
and \U$1983 ( \2230 , \2214 , \2221 );
nor \U$1984 ( \2231 , \2229 , \2230 );
not \U$1985 ( \2232 , \2231 );
not \U$1986 ( \2233 , RIbe28228_16);
not \U$1987 ( \2234 , RIbe28570_23);
and \U$1988 ( \2235 , \2233 , \2234 );
and \U$1989 ( \2236 , RIbe28228_16, RIbe28570_23);
nor \U$1990 ( \2237 , \2235 , \2236 );
not \U$1991 ( \2238 , \2237 );
not \U$1992 ( \2239 , \1061 );
or \U$1993 ( \2240 , \2238 , \2239 );
or \U$1994 ( \2241 , \886 , \1838 );
nand \U$1995 ( \2242 , \2240 , \2241 );
not \U$1996 ( \2243 , \2242 );
not \U$1997 ( \2244 , RIbe28318_18);
and \U$1998 ( \2245 , \901 , \2244 );
and \U$1999 ( \2246 , RIbe28318_18, RIbe296c8_60);
nor \U$2000 ( \2247 , \2245 , \2246 );
not \U$2001 ( \2248 , \2247 );
not \U$2002 ( \2249 , \1452 );
or \U$2003 ( \2250 , \2248 , \2249 );
nand \U$2004 ( \2251 , \1137 , \1721 );
nand \U$2005 ( \2252 , \2250 , \2251 );
not \U$2006 ( \2253 , \283 );
not \U$2007 ( \2254 , RIbe29038_46);
not \U$2008 ( \2255 , RIbe28c00_37);
or \U$2009 ( \2256 , \2254 , \2255 );
or \U$2010 ( \2257 , RIbe28c00_37, RIbe29038_46);
nand \U$2011 ( \2258 , \2256 , \2257 );
not \U$2012 ( \2259 , \2258 );
and \U$2013 ( \2260 , \2253 , \2259 );
and \U$2014 ( \2261 , \287 , \1803 );
nor \U$2015 ( \2262 , \2260 , \2261 );
xnor \U$2016 ( \2263 , \2252 , \2262 );
not \U$2017 ( \2264 , \2263 );
or \U$2018 ( \2265 , \2243 , \2264 );
not \U$2019 ( \2266 , \2262 );
nand \U$2020 ( \2267 , \2266 , \2252 );
nand \U$2021 ( \2268 , \2265 , \2267 );
not \U$2022 ( \2269 , \2268 );
and \U$2023 ( \2270 , RIbe28a20_33, \388 );
not \U$2024 ( \2271 , RIbe28a20_33);
and \U$2025 ( \2272 , \2271 , RIbe29380_53);
nor \U$2026 ( \2273 , \2270 , \2272 );
not \U$2027 ( \2274 , \2273 );
not \U$2028 ( \2275 , \2274 );
buf \U$2029 ( \2276 , \1780 );
not \U$2030 ( \2277 , \2276 );
or \U$2031 ( \2278 , \2275 , \2277 );
nand \U$2032 ( \2279 , \1769 , RIbe28a20_33);
nand \U$2033 ( \2280 , \2278 , \2279 );
not \U$2034 ( \2281 , \2280 );
not \U$2035 ( \2282 , \2281 );
and \U$2036 ( \2283 , \2269 , \2282 );
and \U$2037 ( \2284 , \2268 , \2281 );
nor \U$2038 ( \2285 , \2283 , \2284 );
not \U$2039 ( \2286 , \2285 );
not \U$2040 ( \2287 , \2286 );
or \U$2041 ( \2288 , \2232 , \2287 );
nand \U$2042 ( \2289 , \2268 , \2280 );
nand \U$2043 ( \2290 , \2288 , \2289 );
not \U$2044 ( \2291 , \2290 );
xnor \U$2045 ( \2292 , \1727 , \1729 );
not \U$2046 ( \2293 , \2292 );
and \U$2047 ( \2294 , \2291 , \2293 );
and \U$2048 ( \2295 , \2290 , \2292 );
nor \U$2049 ( \2296 , \2294 , \2295 );
xor \U$2050 ( \2297 , \1827 , \1833 );
xor \U$2051 ( \2298 , \2297 , \1841 );
not \U$2052 ( \2299 , RIbe27ee0_9);
not \U$2053 ( \2300 , RIbe28930_31);
and \U$2054 ( \2301 , \2299 , \2300 );
and \U$2055 ( \2302 , RIbe27ee0_9, RIbe28930_31);
nor \U$2056 ( \2303 , \2301 , \2302 );
and \U$2057 ( \2304 , \966 , \2303 );
and \U$2058 ( \2305 , \971 , \1791 );
nor \U$2059 ( \2306 , \2304 , \2305 );
not \U$2060 ( \2307 , \2306 );
not \U$2061 ( \2308 , \2307 );
not \U$2062 ( \2309 , \259 );
xnor \U$2063 ( \2310 , RIbe27b98_2, RIbe29740_61);
not \U$2064 ( \2311 , \2310 );
and \U$2065 ( \2312 , \2309 , \2311 );
and \U$2066 ( \2313 , \1298 , \1742 );
nor \U$2067 ( \2314 , \2312 , \2313 );
not \U$2068 ( \2315 , \1093 );
not \U$2069 ( \2316 , \1753 );
not \U$2070 ( \2317 , \2316 );
and \U$2071 ( \2318 , \2315 , \2317 );
not \U$2072 ( \2319 , RIbe27d78_6);
not \U$2073 ( \2320 , RIbe288b8_30);
and \U$2074 ( \2321 , \2319 , \2320 );
and \U$2075 ( \2322 , RIbe27d78_6, RIbe288b8_30);
nor \U$2076 ( \2323 , \2321 , \2322 );
and \U$2077 ( \2324 , \1613 , \2323 );
nor \U$2078 ( \2325 , \2318 , \2324 );
and \U$2079 ( \2326 , \2314 , \2325 );
not \U$2080 ( \2327 , \2314 );
not \U$2081 ( \2328 , \2325 );
and \U$2082 ( \2329 , \2327 , \2328 );
nor \U$2083 ( \2330 , \2326 , \2329 );
not \U$2084 ( \2331 , \2330 );
or \U$2085 ( \2332 , \2308 , \2331 );
not \U$2086 ( \2333 , \2314 );
nand \U$2087 ( \2334 , \2333 , \2328 );
nand \U$2088 ( \2335 , \2332 , \2334 );
xor \U$2089 ( \2336 , \2298 , \2335 );
xor \U$2090 ( \2337 , \1811 , \1785 );
and \U$2091 ( \2338 , \2336 , \2337 );
and \U$2092 ( \2339 , \2298 , \2335 );
nor \U$2093 ( \2340 , \2338 , \2339 );
or \U$2094 ( \2341 , \2296 , \2340 );
not \U$2095 ( \2342 , \2290 );
or \U$2096 ( \2343 , \2342 , \2292 );
nand \U$2097 ( \2344 , \2341 , \2343 );
xor \U$2098 ( \2345 , \1708 , \1732 );
xor \U$2099 ( \2346 , \2345 , \1852 );
not \U$2100 ( \2347 , \2346 );
and \U$2101 ( \2348 , \2344 , \2347 );
not \U$2102 ( \2349 , \2344 );
and \U$2103 ( \2350 , \2349 , \2346 );
nor \U$2104 ( \2351 , \2348 , \2350 );
xor \U$2105 ( \2352 , \1695 , \1679 );
and \U$2106 ( \2353 , \2351 , \2352 );
and \U$2107 ( \2354 , \2344 , \2347 );
nor \U$2108 ( \2355 , \2353 , \2354 );
and \U$2109 ( \2356 , \2206 , \2355 );
and \U$2110 ( \2357 , \2204 , \2205 );
or \U$2111 ( \2358 , \2356 , \2357 );
xnor \U$2112 ( \2359 , \1868 , \1867 );
nand \U$2113 ( \2360 , \2358 , \2359 );
not \U$2114 ( \2361 , \2360 );
xor \U$2115 ( \2362 , RIbe28228_16, RIbe294e8_56);
and \U$2116 ( \2363 , \879 , \2362 );
and \U$2117 ( \2364 , RIbe28228_16, RIbe288b8_30);
nor \U$2118 ( \2365 , RIbe28228_16, RIbe288b8_30);
nor \U$2119 ( \2366 , \2364 , \2365 );
and \U$2120 ( \2367 , \887 , \2366 );
nor \U$2121 ( \2368 , \2363 , \2367 );
buf \U$2122 ( \2369 , \1263 );
not \U$2123 ( \2370 , \2369 );
xor \U$2124 ( \2371 , RIbe280c0_13, RIbe29470_55);
not \U$2125 ( \2372 , \2371 );
or \U$2126 ( \2373 , \2370 , \2372 );
and \U$2127 ( \2374 , RIbe280c0_13, \951 );
not \U$2128 ( \2375 , RIbe280c0_13);
and \U$2129 ( \2376 , \2375 , RIbe282a0_17);
nor \U$2130 ( \2377 , \2374 , \2376 );
not \U$2131 ( \2378 , \2377 );
not \U$2132 ( \2379 , \859 );
buf \U$2133 ( \2380 , \2379 );
nand \U$2134 ( \2381 , \2378 , \2380 );
nand \U$2135 ( \2382 , \2373 , \2381 );
and \U$2136 ( \2383 , \2368 , \2382 );
not \U$2137 ( \2384 , \2368 );
not \U$2138 ( \2385 , \2382 );
and \U$2139 ( \2386 , \2384 , \2385 );
or \U$2140 ( \2387 , \2383 , \2386 );
not \U$2141 ( \2388 , \282 );
not \U$2142 ( \2389 , \2388 );
xnor \U$2143 ( \2390 , RIbe29038_46, RIbe295d8_58);
not \U$2144 ( \2391 , \2390 );
and \U$2145 ( \2392 , \2389 , \2391 );
not \U$2146 ( \2393 , RIbe29038_46);
not \U$2147 ( \2394 , RIbe29740_61);
and \U$2148 ( \2395 , \2393 , \2394 );
and \U$2149 ( \2396 , RIbe29038_46, RIbe29740_61);
nor \U$2150 ( \2397 , \2395 , \2396 );
and \U$2151 ( \2398 , \1805 , \2397 );
nor \U$2152 ( \2399 , \2392 , \2398 );
not \U$2153 ( \2400 , \2399 );
and \U$2154 ( \2401 , \2387 , \2400 );
not \U$2155 ( \2402 , \2387 );
and \U$2156 ( \2403 , \2402 , \2399 );
nor \U$2157 ( \2404 , \2401 , \2403 );
not \U$2158 ( \2405 , \2404 );
xor \U$2159 ( \2406 , RIbe296c8_60, RIbe297b8_62);
not \U$2160 ( \2407 , \2406 );
not \U$2161 ( \2408 , \1130 );
or \U$2162 ( \2409 , \2407 , \2408 );
not \U$2163 ( \2410 , RIbe28138_14);
not \U$2164 ( \2411 , RIbe296c8_60);
and \U$2165 ( \2412 , \2410 , \2411 );
and \U$2166 ( \2413 , RIbe28138_14, RIbe296c8_60);
nor \U$2167 ( \2414 , \2412 , \2413 );
nand \U$2168 ( \2415 , \908 , \2414 );
nand \U$2169 ( \2416 , \2409 , \2415 );
not \U$2170 ( \2417 , \2416 );
and \U$2171 ( \2418 , RIbe27d78_6, RIbe29a10_67);
not \U$2172 ( \2419 , RIbe27d78_6);
not \U$2173 ( \2420 , RIbe29a10_67);
and \U$2174 ( \2421 , \2419 , \2420 );
nor \U$2175 ( \2422 , \2418 , \2421 );
not \U$2176 ( \2423 , \2422 );
not \U$2177 ( \2424 , \1086 );
or \U$2178 ( \2425 , \2423 , \2424 );
not \U$2179 ( \2426 , RIbe27d78_6);
not \U$2180 ( \2427 , RIbe29b00_69);
and \U$2181 ( \2428 , \2426 , \2427 );
and \U$2182 ( \2429 , RIbe27d78_6, RIbe29b00_69);
nor \U$2183 ( \2430 , \2428 , \2429 );
nand \U$2184 ( \2431 , \315 , \2430 );
nand \U$2185 ( \2432 , \2425 , \2431 );
xor \U$2186 ( \2433 , \2417 , \2432 );
xor \U$2187 ( \2434 , RIbe27b98_2, RIbe298a8_64);
not \U$2188 ( \2435 , \2434 );
not \U$2189 ( \2436 , \256 );
or \U$2190 ( \2437 , \2435 , \2436 );
xnor \U$2191 ( \2438 , RIbe29998_66, RIbe27b98_2);
not \U$2192 ( \2439 , \2438 );
nand \U$2193 ( \2440 , \2439 , \269 );
nand \U$2194 ( \2441 , \2437 , \2440 );
not \U$2195 ( \2442 , \2441 );
xor \U$2196 ( \2443 , \2433 , \2442 );
not \U$2197 ( \2444 , \2443 );
and \U$2198 ( \2445 , RIbe27e68_8, RIbe28048_12);
not \U$2199 ( \2446 , RIbe27e68_8);
and \U$2200 ( \2447 , \2446 , \431 );
nor \U$2201 ( \2448 , \2445 , \2447 );
not \U$2202 ( \2449 , \2448 );
not \U$2203 ( \2450 , RIbe27e68_8);
nor \U$2204 ( \2451 , RIbe27f58_10, RIbe27fd0_11);
not \U$2205 ( \2452 , \2451 );
or \U$2206 ( \2453 , \2450 , \2452 );
not \U$2207 ( \2454 , RIbe27e68_8);
nand \U$2208 ( \2455 , \2454 , RIbe27fd0_11, RIbe27f58_10);
nand \U$2209 ( \2456 , \2453 , \2455 );
buf \U$2210 ( \2457 , \2456 );
buf \U$2211 ( \2458 , \2457 );
buf \U$2212 ( \2459 , \2458 );
not \U$2213 ( \2460 , \2459 );
or \U$2214 ( \2461 , \2449 , \2460 );
xor \U$2215 ( \2462 , RIbe27f58_10, RIbe27fd0_11);
buf \U$2216 ( \2463 , \2462 );
buf \U$2217 ( \2464 , \2463 );
and \U$2218 ( \2465 , RIbe27e68_8, RIbe29380_53);
not \U$2219 ( \2466 , RIbe27e68_8);
and \U$2220 ( \2467 , \2466 , \388 );
nor \U$2221 ( \2468 , \2465 , \2467 );
nand \U$2222 ( \2469 , \2464 , \2468 );
nand \U$2223 ( \2470 , \2461 , \2469 );
xor \U$2224 ( \2471 , RIbe28a20_33, RIbe29308_52);
not \U$2225 ( \2472 , \2471 );
not \U$2226 ( \2473 , \1781 );
or \U$2227 ( \2474 , \2472 , \2473 );
buf \U$2228 ( \2475 , \1768 );
buf \U$2229 ( \2476 , \2475 );
and \U$2230 ( \2477 , RIbe28a20_33, RIbe28c00_37);
not \U$2231 ( \2478 , RIbe28a20_33);
not \U$2232 ( \2479 , RIbe28c00_37);
and \U$2233 ( \2480 , \2478 , \2479 );
nor \U$2234 ( \2481 , \2477 , \2480 );
nand \U$2235 ( \2482 , \2476 , \2481 );
nand \U$2236 ( \2483 , \2474 , \2482 );
xor \U$2237 ( \2484 , \2470 , \2483 );
and \U$2238 ( \2485 , RIbe28930_31, RIbe28a98_34);
nor \U$2239 ( \2486 , RIbe28930_31, RIbe28a98_34);
nor \U$2240 ( \2487 , \2485 , \2486 );
and \U$2241 ( \2488 , \966 , \2487 );
not \U$2242 ( \2489 , RIbe293f8_54);
and \U$2243 ( \2490 , \973 , \2489 );
and \U$2244 ( \2491 , RIbe28930_31, RIbe293f8_54);
nor \U$2245 ( \2492 , \2490 , \2491 );
and \U$2246 ( \2493 , \1199 , \2492 );
nor \U$2247 ( \2494 , \2488 , \2493 );
and \U$2248 ( \2495 , \2484 , \2494 );
not \U$2249 ( \2496 , \2484 );
not \U$2250 ( \2497 , \2494 );
and \U$2251 ( \2498 , \2496 , \2497 );
or \U$2252 ( \2499 , \2495 , \2498 );
not \U$2253 ( \2500 , \2499 );
or \U$2254 ( \2501 , \2444 , \2500 );
or \U$2255 ( \2502 , \2499 , \2443 );
nand \U$2256 ( \2503 , \2501 , \2502 );
not \U$2257 ( \2504 , \2503 );
or \U$2258 ( \2505 , \2405 , \2504 );
or \U$2259 ( \2506 , \2503 , \2404 );
nand \U$2260 ( \2507 , \2505 , \2506 );
not \U$2261 ( \2508 , \2507 );
xnor \U$2262 ( \2509 , RIbe28480_21, RIbe28750_27);
not \U$2263 ( \2510 , \2509 );
not \U$2264 ( \2511 , \2510 );
xor \U$2265 ( \2512 , RIbe28480_21, RIbe287c8_28);
not \U$2266 ( \2513 , RIbe287c8_28);
nand \U$2267 ( \2514 , \2513 , RIbe285e8_24);
not \U$2268 ( \2515 , RIbe285e8_24);
nand \U$2269 ( \2516 , \2515 , RIbe287c8_28);
and \U$2270 ( \2517 , \2512 , \2514 , \2516 );
buf \U$2271 ( \2518 , \2517 );
buf \U$2272 ( \2519 , \2518 );
buf \U$2273 ( \2520 , \2519 );
not \U$2274 ( \2521 , \2520 );
or \U$2275 ( \2522 , \2511 , \2521 );
xnor \U$2276 ( \2523 , RIbe28480_21, RIbe28840_29);
not \U$2277 ( \2524 , \2523 );
xor \U$2278 ( \2525 , RIbe285e8_24, RIbe287c8_28);
not \U$2279 ( \2526 , \2525 );
not \U$2280 ( \2527 , \2526 );
nand \U$2281 ( \2528 , \2524 , \2527 );
nand \U$2282 ( \2529 , \2522 , \2528 );
not \U$2283 ( \2530 , RIbe288b8_30);
not \U$2284 ( \2531 , RIbe28930_31);
and \U$2285 ( \2532 , \2530 , \2531 );
and \U$2286 ( \2533 , RIbe288b8_30, RIbe28930_31);
nor \U$2287 ( \2534 , \2532 , \2533 );
not \U$2288 ( \2535 , \2534 );
not \U$2289 ( \2536 , \966 );
or \U$2290 ( \2537 , \2535 , \2536 );
nand \U$2291 ( \2538 , \1199 , \2487 );
nand \U$2292 ( \2539 , \2537 , \2538 );
xor \U$2293 ( \2540 , \2529 , \2539 );
and \U$2294 ( \2541 , RIbe28b88_36, RIbe28c00_37);
not \U$2295 ( \2542 , RIbe28b88_36);
and \U$2296 ( \2543 , \2542 , \2479 );
nor \U$2297 ( \2544 , \2541 , \2543 );
not \U$2298 ( \2545 , \2544 );
not \U$2299 ( \2546 , RIbe28b10_35);
nand \U$2300 ( \2547 , \2546 , RIbe28390_19);
nor \U$2301 ( \2548 , RIbe28390_19, RIbe28b88_36);
not \U$2302 ( \2549 , \2548 );
nand \U$2303 ( \2550 , RIbe28b10_35, RIbe28b88_36);
and \U$2304 ( \2551 , \2547 , \2549 , \2550 );
buf \U$2305 ( \2552 , \2551 );
buf \U$2306 ( \2553 , \2552 );
buf \U$2307 ( \2554 , \2553 );
not \U$2308 ( \2555 , \2554 );
or \U$2309 ( \2556 , \2545 , \2555 );
xor \U$2310 ( \2557 , RIbe28390_19, RIbe28b10_35);
buf \U$2311 ( \2558 , \2557 );
buf \U$2312 ( \2559 , \2558 );
buf \U$2313 ( \2560 , \2559 );
buf \U$2314 ( \2561 , \2560 );
not \U$2315 ( \2562 , RIbe28b88_36);
not \U$2316 ( \2563 , RIbe28c78_38);
and \U$2317 ( \2564 , \2562 , \2563 );
and \U$2318 ( \2565 , RIbe28b88_36, RIbe28c78_38);
nor \U$2319 ( \2566 , \2564 , \2565 );
nand \U$2320 ( \2567 , \2561 , \2566 );
nand \U$2321 ( \2568 , \2556 , \2567 );
not \U$2322 ( \2569 , \2568 );
and \U$2323 ( \2570 , \2540 , \2569 );
not \U$2324 ( \2571 , \2540 );
and \U$2325 ( \2572 , \2571 , \2568 );
or \U$2326 ( \2573 , \2570 , \2572 );
not \U$2327 ( \2574 , \2573 );
not \U$2328 ( \2575 , \2574 );
not \U$2329 ( \2576 , RIbe27c10_3);
not \U$2330 ( \2577 , RIbe27c88_4);
and \U$2331 ( \2578 , \2576 , \2577 );
and \U$2332 ( \2579 , RIbe27c10_3, RIbe27c88_4);
nor \U$2333 ( \2580 , \2578 , \2579 );
not \U$2334 ( \2581 , \2580 );
not \U$2335 ( \2582 , \361 );
or \U$2336 ( \2583 , \2581 , \2582 );
xnor \U$2337 ( \2584 , RIbe27df0_7, RIbe27c10_3);
not \U$2338 ( \2585 , \2584 );
nand \U$2339 ( \2586 , \2585 , \369 );
nand \U$2340 ( \2587 , \2583 , \2586 );
not \U$2341 ( \2588 , \2587 );
nand \U$2342 ( \2589 , RIbe27b20_1, RIbe27b98_2);
not \U$2343 ( \2590 , \2589 );
and \U$2344 ( \2591 , \2588 , \2590 );
and \U$2345 ( \2592 , \2587 , \2589 );
nor \U$2346 ( \2593 , \2591 , \2592 );
not \U$2347 ( \2594 , RIbe27e68_8);
or \U$2348 ( \2595 , \2594 , RIbe27ee0_9);
or \U$2349 ( \2596 , \317 , RIbe27e68_8);
nand \U$2350 ( \2597 , \2595 , \2596 );
not \U$2351 ( \2598 , \2597 );
buf \U$2352 ( \2599 , \2457 );
buf \U$2353 ( \2600 , \2599 );
not \U$2354 ( \2601 , \2600 );
or \U$2355 ( \2602 , \2598 , \2601 );
buf \U$2356 ( \2603 , \2463 );
nand \U$2357 ( \2604 , \2603 , \2448 );
nand \U$2358 ( \2605 , \2602 , \2604 );
xor \U$2359 ( \2606 , \2593 , \2605 );
not \U$2360 ( \2607 , \2606 );
xor \U$2361 ( \2608 , RIbe28570_23, RIbe285e8_24);
not \U$2362 ( \2609 , \2608 );
and \U$2363 ( \2610 , RIbe27e68_8, RIbe285e8_24);
not \U$2364 ( \2611 , RIbe27e68_8);
and \U$2365 ( \2612 , \2611 , RIbe28660_25);
nor \U$2366 ( \2613 , \2610 , \2612 );
nor \U$2367 ( \2614 , RIbe285e8_24, RIbe28660_25);
not \U$2368 ( \2615 , \2614 );
nand \U$2369 ( \2616 , \2613 , \2615 );
buf \U$2370 ( \2617 , \2616 );
not \U$2371 ( \2618 , \2617 );
not \U$2372 ( \2619 , \2618 );
or \U$2373 ( \2620 , \2609 , \2619 );
xnor \U$2374 ( \2621 , RIbe286d8_26, RIbe285e8_24);
not \U$2375 ( \2622 , \2621 );
xor \U$2376 ( \2623 , RIbe27e68_8, RIbe28660_25);
buf \U$2377 ( \2624 , \2623 );
buf \U$2378 ( \2625 , \2624 );
buf \U$2379 ( \2626 , \2625 );
nand \U$2380 ( \2627 , \2622 , \2626 );
nand \U$2381 ( \2628 , \2620 , \2627 );
and \U$2382 ( \2629 , RIbe28390_19, RIbe28318_18);
not \U$2383 ( \2630 , RIbe28390_19);
and \U$2384 ( \2631 , \2630 , \2244 );
nor \U$2385 ( \2632 , \2629 , \2631 );
not \U$2386 ( \2633 , \2632 );
xor \U$2387 ( \2634 , RIbe28408_20, RIbe28480_21);
not \U$2388 ( \2635 , \2634 );
xor \U$2389 ( \2636 , RIbe28390_19, RIbe28408_20);
nand \U$2390 ( \2637 , \2635 , \2636 );
buf \U$2391 ( \2638 , \2637 );
not \U$2392 ( \2639 , \2638 );
buf \U$2393 ( \2640 , \2639 );
not \U$2394 ( \2641 , \2640 );
or \U$2395 ( \2642 , \2633 , \2641 );
xnor \U$2396 ( \2643 , RIbe28390_19, RIbe284f8_22);
not \U$2397 ( \2644 , \2643 );
not \U$2398 ( \2645 , \2634 );
buf \U$2399 ( \2646 , \2645 );
not \U$2400 ( \2647 , \2646 );
buf \U$2401 ( \2648 , \2647 );
nand \U$2402 ( \2649 , \2644 , \2648 );
nand \U$2403 ( \2650 , \2642 , \2649 );
xor \U$2404 ( \2651 , \2628 , \2650 );
xnor \U$2405 ( \2652 , RIbe280c0_13, RIbe28138_14);
or \U$2406 ( \2653 , \1575 , \2652 );
or \U$2407 ( \2654 , \1573 , \2377 );
nand \U$2408 ( \2655 , \2653 , \2654 );
xor \U$2409 ( \2656 , \2651 , \2655 );
not \U$2410 ( \2657 , \2656 );
or \U$2411 ( \2658 , \2607 , \2657 );
or \U$2412 ( \2659 , \2656 , \2606 );
nand \U$2413 ( \2660 , \2658 , \2659 );
not \U$2414 ( \2661 , \2660 );
or \U$2415 ( \2662 , \2575 , \2661 );
not \U$2416 ( \2663 , \2606 );
nand \U$2417 ( \2664 , \2663 , \2656 );
nand \U$2418 ( \2665 , \2662 , \2664 );
not \U$2419 ( \2666 , \2665 );
not \U$2420 ( \2667 , \2519 );
or \U$2421 ( \2668 , \2667 , \2523 );
xnor \U$2422 ( \2669 , RIbe28480_21, RIbe28570_23);
xnor \U$2423 ( \2670 , RIbe285e8_24, RIbe287c8_28);
not \U$2424 ( \2671 , \2670 );
not \U$2425 ( \2672 , \2671 );
or \U$2426 ( \2673 , \2669 , \2672 );
nand \U$2427 ( \2674 , \2668 , \2673 );
and \U$2428 ( \2675 , RIbe28cf0_39, RIbe27b98_2);
xor \U$2429 ( \2676 , RIbe28d68_40, RIbe28de0_41);
not \U$2430 ( \2677 , \2676 );
not \U$2431 ( \2678 , \332 );
or \U$2432 ( \2679 , \2677 , \2678 );
xor \U$2433 ( \2680 , RIbe27c88_4, RIbe28de0_41);
nand \U$2434 ( \2681 , \514 , \2680 );
nand \U$2435 ( \2682 , \2679 , \2681 );
xor \U$2436 ( \2683 , \2675 , \2682 );
not \U$2437 ( \2684 , \2683 );
and \U$2438 ( \2685 , \2674 , \2684 );
not \U$2439 ( \2686 , \2674 );
and \U$2440 ( \2687 , \2686 , \2683 );
nor \U$2441 ( \2688 , \2685 , \2687 );
not \U$2442 ( \2689 , \2688 );
not \U$2443 ( \2690 , \2689 );
buf \U$2444 ( \2691 , \2559 );
not \U$2445 ( \2692 , \2691 );
not \U$2446 ( \2693 , \2692 );
and \U$2447 ( \2694 , RIbe28b88_36, \2244 );
not \U$2448 ( \2695 , RIbe28b88_36);
and \U$2449 ( \2696 , \2695 , RIbe28318_18);
nor \U$2450 ( \2697 , \2694 , \2696 );
not \U$2451 ( \2698 , \2697 );
and \U$2452 ( \2699 , \2693 , \2698 );
not \U$2453 ( \2700 , \2552 );
not \U$2454 ( \2701 , \2700 );
buf \U$2455 ( \2702 , \2701 );
and \U$2456 ( \2703 , \2702 , \2566 );
nor \U$2457 ( \2704 , \2699 , \2703 );
not \U$2458 ( \2705 , \2704 );
xor \U$2459 ( \2706 , RIbe28ed0_43, RIbe28f48_44);
buf \U$2460 ( \2707 , \2706 );
not \U$2461 ( \2708 , \2707 );
not \U$2462 ( \2709 , \2708 );
and \U$2463 ( \2710 , RIbe28ed0_43, RIbe27fd0_11);
not \U$2464 ( \2711 , RIbe28ed0_43);
and \U$2465 ( \2712 , \2711 , RIbe28f48_44);
nor \U$2466 ( \2713 , \2710 , \2712 );
nor \U$2467 ( \2714 , RIbe27fd0_11, RIbe28f48_44);
not \U$2468 ( \2715 , \2714 );
nand \U$2469 ( \2716 , \2713 , \2715 );
buf \U$2470 ( \2717 , \2716 );
buf \U$2471 ( \2718 , \2717 );
not \U$2472 ( \2719 , \2718 );
or \U$2473 ( \2720 , \2709 , \2719 );
nand \U$2474 ( \2721 , \2720 , RIbe27fd0_11);
not \U$2475 ( \2722 , \2721 );
not \U$2476 ( \2723 , RIbe290b0_47);
not \U$2477 ( \2724 , RIbe29128_48);
and \U$2478 ( \2725 , \2723 , \2724 );
and \U$2479 ( \2726 , RIbe290b0_47, RIbe29128_48);
nor \U$2480 ( \2727 , \2725 , \2726 );
not \U$2481 ( \2728 , \2727 );
not \U$2482 ( \2729 , \383 );
buf \U$2483 ( \2730 , \2729 );
buf \U$2484 ( \2731 , \2730 );
not \U$2485 ( \2732 , \2731 );
or \U$2486 ( \2733 , \2728 , \2732 );
not \U$2487 ( \2734 , RIbe290b0_47);
not \U$2488 ( \2735 , RIbe291a0_49);
and \U$2489 ( \2736 , \2734 , \2735 );
and \U$2490 ( \2737 , RIbe290b0_47, RIbe291a0_49);
nor \U$2491 ( \2738 , \2736 , \2737 );
nand \U$2492 ( \2739 , \2071 , \2738 );
nand \U$2493 ( \2740 , \2733 , \2739 );
not \U$2494 ( \2741 , \2740 );
not \U$2495 ( \2742 , \2741 );
or \U$2496 ( \2743 , \2722 , \2742 );
not \U$2497 ( \2744 , \2721 );
nand \U$2498 ( \2745 , \2744 , \2740 );
nand \U$2499 ( \2746 , \2743 , \2745 );
not \U$2500 ( \2747 , \2746 );
or \U$2501 ( \2748 , \2705 , \2747 );
or \U$2502 ( \2749 , \2746 , \2704 );
nand \U$2503 ( \2750 , \2748 , \2749 );
not \U$2504 ( \2751 , \2750 );
not \U$2505 ( \2752 , \2751 );
or \U$2506 ( \2753 , \2690 , \2752 );
nand \U$2507 ( \2754 , \2688 , \2750 );
nand \U$2508 ( \2755 , \2753 , \2754 );
xor \U$2509 ( \2756 , RIbe27ee0_9, RIbe285e8_24);
not \U$2510 ( \2757 , \2756 );
buf \U$2511 ( \2758 , \2623 );
not \U$2512 ( \2759 , \2758 );
or \U$2513 ( \2760 , \2757 , \2759 );
not \U$2514 ( \2761 , \2617 );
not \U$2515 ( \2762 , \2761 );
or \U$2516 ( \2763 , \2762 , \2621 );
nand \U$2517 ( \2764 , \2760 , \2763 );
or \U$2518 ( \2765 , \360 , \2584 );
not \U$2519 ( \2766 , RIbe29218_50);
not \U$2520 ( \2767 , RIbe27c10_3);
or \U$2521 ( \2768 , \2766 , \2767 );
or \U$2522 ( \2769 , RIbe27c10_3, RIbe29218_50);
nand \U$2523 ( \2770 , \2768 , \2769 );
or \U$2524 ( \2771 , \1107 , \2770 );
nand \U$2525 ( \2772 , \2765 , \2771 );
xor \U$2526 ( \2773 , \2764 , \2772 );
not \U$2527 ( \2774 , \2640 );
or \U$2528 ( \2775 , \2774 , \2643 );
buf \U$2529 ( \2776 , \2634 );
buf \U$2530 ( \2777 , \2776 );
not \U$2531 ( \2778 , \2777 );
not \U$2532 ( \2779 , RIbe28390_19);
and \U$2533 ( \2780 , RIbe28750_27, \2779 );
not \U$2534 ( \2781 , RIbe28750_27);
and \U$2535 ( \2782 , \2781 , RIbe28390_19);
nor \U$2536 ( \2783 , \2780 , \2782 );
or \U$2537 ( \2784 , \2778 , \2783 );
nand \U$2538 ( \2785 , \2775 , \2784 );
xor \U$2539 ( \2786 , \2773 , \2785 );
not \U$2540 ( \2787 , \2786 );
and \U$2541 ( \2788 , \2755 , \2787 );
not \U$2542 ( \2789 , \2755 );
and \U$2543 ( \2790 , \2789 , \2786 );
nor \U$2544 ( \2791 , \2788 , \2790 );
not \U$2545 ( \2792 , \2791 );
or \U$2546 ( \2793 , \2666 , \2792 );
or \U$2547 ( \2794 , \2665 , \2791 );
nand \U$2548 ( \2795 , \2793 , \2794 );
not \U$2549 ( \2796 , \2795 );
or \U$2550 ( \2797 , \2508 , \2796 );
not \U$2551 ( \2798 , \2665 );
or \U$2552 ( \2799 , \2798 , \2791 );
nand \U$2553 ( \2800 , \2797 , \2799 );
not \U$2554 ( \2801 , \2746 );
or \U$2555 ( \2802 , \2801 , \2704 );
not \U$2556 ( \2803 , \2740 );
or \U$2557 ( \2804 , \2803 , \2744 );
nand \U$2558 ( \2805 , \2802 , \2804 );
and \U$2559 ( \2806 , \2683 , \2674 );
and \U$2560 ( \2807 , \2675 , \2682 );
nor \U$2561 ( \2808 , \2806 , \2807 );
not \U$2562 ( \2809 , \2808 );
xor \U$2563 ( \2810 , \2764 , \2772 );
and \U$2564 ( \2811 , \2810 , \2785 );
and \U$2565 ( \2812 , \2764 , \2772 );
or \U$2566 ( \2813 , \2811 , \2812 );
not \U$2567 ( \2814 , \2813 );
or \U$2568 ( \2815 , \2809 , \2814 );
or \U$2569 ( \2816 , \2813 , \2808 );
nand \U$2570 ( \2817 , \2815 , \2816 );
xor \U$2571 ( \2818 , \2805 , \2817 );
not \U$2572 ( \2819 , \2786 );
not \U$2573 ( \2820 , \2755 );
or \U$2574 ( \2821 , \2819 , \2820 );
nand \U$2575 ( \2822 , \2750 , \2689 );
nand \U$2576 ( \2823 , \2821 , \2822 );
and \U$2577 ( \2824 , \2818 , \2823 );
not \U$2578 ( \2825 , \2818 );
not \U$2579 ( \2826 , \2823 );
and \U$2580 ( \2827 , \2825 , \2826 );
nor \U$2581 ( \2828 , \2824 , \2827 );
nand \U$2582 ( \2829 , RIbe27b98_2, RIbe298a8_64);
not \U$2583 ( \2830 , \2829 );
not \U$2584 ( \2831 , \2371 );
not \U$2585 ( \2832 , \2380 );
or \U$2586 ( \2833 , \2831 , \2832 );
xnor \U$2587 ( \2834 , RIbe294e8_56, RIbe280c0_13);
not \U$2588 ( \2835 , \2834 );
nand \U$2589 ( \2836 , \2835 , \869 );
nand \U$2590 ( \2837 , \2833 , \2836 );
not \U$2591 ( \2838 , \2837 );
or \U$2592 ( \2839 , \2830 , \2838 );
or \U$2593 ( \2840 , \2837 , \2829 );
nand \U$2594 ( \2841 , \2839 , \2840 );
and \U$2595 ( \2842 , \979 , \2397 );
not \U$2596 ( \2843 , RIbe29038_46);
not \U$2597 ( \2844 , RIbe297b8_62);
and \U$2598 ( \2845 , \2843 , \2844 );
and \U$2599 ( \2846 , RIbe29038_46, RIbe297b8_62);
nor \U$2600 ( \2847 , \2845 , \2846 );
and \U$2601 ( \2848 , \287 , \2847 );
nor \U$2602 ( \2849 , \2842 , \2848 );
not \U$2603 ( \2850 , \2849 );
and \U$2604 ( \2851 , \2841 , \2850 );
not \U$2605 ( \2852 , \2841 );
and \U$2606 ( \2853 , \2852 , \2849 );
nor \U$2607 ( \2854 , \2851 , \2853 );
not \U$2608 ( \2855 , \2854 );
not \U$2609 ( \2856 , \2680 );
not \U$2610 ( \2857 , \333 );
not \U$2611 ( \2858 , \2857 );
or \U$2612 ( \2859 , \2856 , \2858 );
xor \U$2613 ( \2860 , RIbe27df0_7, RIbe28de0_41);
nand \U$2614 ( \2861 , \514 , \2860 );
nand \U$2615 ( \2862 , \2859 , \2861 );
not \U$2616 ( \2863 , \2481 );
not \U$2617 ( \2864 , \1781 );
or \U$2618 ( \2865 , \2863 , \2864 );
not \U$2619 ( \2866 , RIbe28a20_33);
not \U$2620 ( \2867 , RIbe28c78_38);
and \U$2621 ( \2868 , \2866 , \2867 );
and \U$2622 ( \2869 , RIbe28a20_33, RIbe28c78_38);
nor \U$2623 ( \2870 , \2868 , \2869 );
nand \U$2624 ( \2871 , \1769 , \2870 );
nand \U$2625 ( \2872 , \2865 , \2871 );
xor \U$2626 ( \2873 , \2862 , \2872 );
not \U$2627 ( \2874 , \2414 );
not \U$2628 ( \2875 , \899 );
not \U$2629 ( \2876 , \2875 );
not \U$2630 ( \2877 , \2876 );
not \U$2631 ( \2878 , \2877 );
or \U$2632 ( \2879 , \2874 , \2878 );
and \U$2633 ( \2880 , \901 , \951 );
and \U$2634 ( \2881 , RIbe282a0_17, RIbe296c8_60);
nor \U$2635 ( \2882 , \2880 , \2881 );
nand \U$2636 ( \2883 , \1939 , \2882 );
nand \U$2637 ( \2884 , \2879 , \2883 );
xnor \U$2638 ( \2885 , \2873 , \2884 );
not \U$2639 ( \2886 , \2885 );
or \U$2640 ( \2887 , \2855 , \2886 );
or \U$2641 ( \2888 , \2885 , \2854 );
nand \U$2642 ( \2889 , \2887 , \2888 );
not \U$2643 ( \2890 , \2617 );
not \U$2644 ( \2891 , \2890 );
not \U$2645 ( \2892 , \2756 );
or \U$2646 ( \2893 , \2891 , \2892 );
not \U$2647 ( \2894 , \2626 );
xnor \U$2648 ( \2895 , RIbe28048_12, RIbe285e8_24);
or \U$2649 ( \2896 , \2894 , \2895 );
nand \U$2650 ( \2897 , \2893 , \2896 );
or \U$2651 ( \2898 , \360 , \2770 );
xnor \U$2652 ( \2899 , RIbe27c10_3, RIbe29a10_67);
or \U$2653 ( \2900 , \1107 , \2899 );
nand \U$2654 ( \2901 , \2898 , \2900 );
xor \U$2655 ( \2902 , \2897 , \2901 );
or \U$2656 ( \2903 , \2774 , \2783 );
and \U$2657 ( \2904 , RIbe28390_19, RIbe28840_29);
not \U$2658 ( \2905 , RIbe28390_19);
and \U$2659 ( \2906 , \2905 , \364 );
nor \U$2660 ( \2907 , \2904 , \2906 );
not \U$2661 ( \2908 , \2907 );
or \U$2662 ( \2909 , \2778 , \2908 );
nand \U$2663 ( \2910 , \2903 , \2909 );
xor \U$2664 ( \2911 , \2902 , \2910 );
xor \U$2665 ( \2912 , \2889 , \2911 );
and \U$2666 ( \2913 , \2828 , \2912 );
not \U$2667 ( \2914 , \2828 );
not \U$2668 ( \2915 , \2912 );
and \U$2669 ( \2916 , \2914 , \2915 );
nor \U$2670 ( \2917 , \2913 , \2916 );
xor \U$2671 ( \2918 , \2800 , \2917 );
or \U$2672 ( \2919 , \2499 , \2404 );
nand \U$2673 ( \2920 , \2919 , \2443 );
nand \U$2674 ( \2921 , \2499 , \2404 );
and \U$2675 ( \2922 , \2920 , \2921 );
not \U$2676 ( \2923 , \2922 );
not \U$2677 ( \2924 , \2593 );
and \U$2678 ( \2925 , \2924 , \2605 );
not \U$2679 ( \2926 , \2587 );
nor \U$2680 ( \2927 , \2926 , \2589 );
nor \U$2681 ( \2928 , \2925 , \2927 );
not \U$2682 ( \2929 , \2928 );
xor \U$2683 ( \2930 , \2628 , \2650 );
and \U$2684 ( \2931 , \2930 , \2655 );
and \U$2685 ( \2932 , \2628 , \2650 );
or \U$2686 ( \2933 , \2931 , \2932 );
not \U$2687 ( \2934 , \2933 );
and \U$2688 ( \2935 , \2929 , \2934 );
and \U$2689 ( \2936 , \2928 , \2933 );
nor \U$2690 ( \2937 , \2935 , \2936 );
xnor \U$2691 ( \2938 , RIbe296c8_60, RIbe29740_61);
not \U$2692 ( \2939 , \2938 );
not \U$2693 ( \2940 , \2939 );
not \U$2694 ( \2941 , \900 );
or \U$2695 ( \2942 , \2940 , \2941 );
nand \U$2696 ( \2943 , \1137 , \2406 );
nand \U$2697 ( \2944 , \2942 , \2943 );
xor \U$2698 ( \2945 , RIbe29038_46, RIbe291a0_49);
not \U$2699 ( \2946 , \2945 );
not \U$2700 ( \2947 , \979 );
or \U$2701 ( \2948 , \2946 , \2947 );
not \U$2702 ( \2949 , \2390 );
nand \U$2703 ( \2950 , \2949 , \287 );
nand \U$2704 ( \2951 , \2948 , \2950 );
xor \U$2705 ( \2952 , \2944 , \2951 );
not \U$2706 ( \2953 , \2952 );
not \U$2707 ( \2954 , \2953 );
and \U$2708 ( \2955 , RIbe28228_16, RIbe29470_55);
nor \U$2709 ( \2956 , RIbe28228_16, RIbe29470_55);
nor \U$2710 ( \2957 , \2955 , \2956 );
and \U$2711 ( \2958 , \1061 , \2957 );
and \U$2712 ( \2959 , \885 , \2362 );
nor \U$2713 ( \2960 , \2958 , \2959 );
not \U$2714 ( \2961 , \2960 );
and \U$2715 ( \2962 , \2954 , \2961 );
and \U$2716 ( \2963 , \2951 , \2944 );
nor \U$2717 ( \2964 , \2962 , \2963 );
or \U$2718 ( \2965 , \2937 , \2964 );
not \U$2719 ( \2966 , \2928 );
nand \U$2720 ( \2967 , \2966 , \2933 );
nand \U$2721 ( \2968 , \2965 , \2967 );
not \U$2722 ( \2969 , \2968 );
and \U$2723 ( \2970 , \2923 , \2969 );
and \U$2724 ( \2971 , \2968 , \2922 );
nor \U$2725 ( \2972 , \2970 , \2971 );
not \U$2726 ( \2973 , \2368 );
not \U$2727 ( \2974 , \2385 );
and \U$2728 ( \2975 , \2973 , \2974 );
and \U$2729 ( \2976 , \2385 , \2368 );
nor \U$2730 ( \2977 , \2976 , \2399 );
nor \U$2731 ( \2978 , \2975 , \2977 );
not \U$2732 ( \2979 , \2978 );
not \U$2733 ( \2980 , \2497 );
not \U$2734 ( \2981 , \2484 );
or \U$2735 ( \2982 , \2980 , \2981 );
nand \U$2736 ( \2983 , \2483 , \2470 );
nand \U$2737 ( \2984 , \2982 , \2983 );
not \U$2738 ( \2985 , \2984 );
or \U$2739 ( \2986 , \2979 , \2985 );
or \U$2740 ( \2987 , \2984 , \2978 );
nand \U$2741 ( \2988 , \2986 , \2987 );
not \U$2742 ( \2989 , \2468 );
not \U$2743 ( \2990 , \2600 );
or \U$2744 ( \2991 , \2989 , \2990 );
nand \U$2745 ( \2992 , \2464 , RIbe27e68_8);
nand \U$2746 ( \2993 , \2991 , \2992 );
or \U$2747 ( \2994 , \387 , RIbe295d8_58);
not \U$2748 ( \2995 , RIbe295d8_58);
or \U$2749 ( \2996 , \2995 , RIbe290b0_47);
nand \U$2750 ( \2997 , \2994 , \2996 );
not \U$2751 ( \2998 , \2997 );
not \U$2752 ( \2999 , \399 );
or \U$2753 ( \3000 , \2998 , \2999 );
xor \U$2754 ( \3001 , RIbe290b0_47, RIbe291a0_49);
nand \U$2755 ( \3002 , \3001 , \466 );
nand \U$2756 ( \3003 , \3000 , \3002 );
not \U$2757 ( \3004 , \1296 );
not \U$2758 ( \3005 , \2438 );
and \U$2759 ( \3006 , \3004 , \3005 );
xor \U$2760 ( \3007 , RIbe28d68_40, RIbe27b98_2);
and \U$2761 ( \3008 , \269 , \3007 );
nor \U$2762 ( \3009 , \3006 , \3008 );
not \U$2763 ( \3010 , \3009 );
xor \U$2764 ( \3011 , \3003 , \3010 );
xor \U$2765 ( \3012 , \2993 , \3011 );
xnor \U$2766 ( \3013 , \2988 , \3012 );
xor \U$2767 ( \3014 , \2972 , \3013 );
and \U$2768 ( \3015 , \2918 , \3014 );
and \U$2769 ( \3016 , \2800 , \2917 );
nor \U$2770 ( \3017 , \3015 , \3016 );
not \U$2771 ( \3018 , \3017 );
not \U$2772 ( \3019 , \3018 );
not \U$2773 ( \3020 , \2554 );
not \U$2774 ( \3021 , \3020 );
not \U$2775 ( \3022 , \2697 );
and \U$2776 ( \3023 , \3021 , \3022 );
not \U$2777 ( \3024 , RIbe284f8_22);
not \U$2778 ( \3025 , RIbe28b88_36);
and \U$2779 ( \3026 , \3024 , \3025 );
and \U$2780 ( \3027 , RIbe284f8_22, RIbe28b88_36);
nor \U$2781 ( \3028 , \3026 , \3027 );
and \U$2782 ( \3029 , \2561 , \3028 );
nor \U$2783 ( \3030 , \3023 , \3029 );
not \U$2784 ( \3031 , \3030 );
and \U$2785 ( \3032 , \1044 , \2430 );
not \U$2786 ( \3033 , RIbe27d78_6);
not \U$2787 ( \3034 , RIbe29128_48);
and \U$2788 ( \3035 , \3033 , \3034 );
and \U$2789 ( \3036 , RIbe27d78_6, RIbe29128_48);
nor \U$2790 ( \3037 , \3035 , \3036 );
and \U$2791 ( \3038 , \314 , \3037 );
nor \U$2792 ( \3039 , \3032 , \3038 );
not \U$2793 ( \3040 , \3039 );
and \U$2794 ( \3041 , \3031 , \3040 );
and \U$2795 ( \3042 , \3030 , \3039 );
nor \U$2796 ( \3043 , \3041 , \3042 );
not \U$2797 ( \3044 , \3043 );
not \U$2798 ( \3045 , \2417 );
not \U$2799 ( \3046 , \2442 );
or \U$2800 ( \3047 , \3045 , \3046 );
nand \U$2801 ( \3048 , \3047 , \2432 );
nand \U$2802 ( \3049 , \2441 , \2416 );
nand \U$2803 ( \3050 , \3048 , \3049 );
not \U$2804 ( \3051 , \3050 );
or \U$2805 ( \3052 , \3044 , \3051 );
or \U$2806 ( \3053 , \3050 , \3043 );
nand \U$2807 ( \3054 , \3052 , \3053 );
not \U$2808 ( \3055 , \3054 );
buf \U$2809 ( \3056 , \878 );
and \U$2810 ( \3057 , \3056 , \2366 );
and \U$2811 ( \3058 , \888 , \940 );
and \U$2812 ( \3059 , RIbe28228_16, RIbe28a98_34);
nor \U$2813 ( \3060 , \3058 , \3059 );
and \U$2814 ( \3061 , \885 , \3060 );
nor \U$2815 ( \3062 , \3057 , \3061 );
not \U$2816 ( \3063 , \2492 );
buf \U$2817 ( \3064 , \1793 );
not \U$2818 ( \3065 , \3064 );
or \U$2819 ( \3066 , \3063 , \3065 );
xnor \U$2820 ( \3067 , RIbe28930_31, RIbe29308_52);
not \U$2821 ( \3068 , \3067 );
nand \U$2822 ( \3069 , \3068 , \971 );
nand \U$2823 ( \3070 , \3066 , \3069 );
not \U$2824 ( \3071 , \2667 );
not \U$2825 ( \3072 , \2669 );
and \U$2826 ( \3073 , \3071 , \3072 );
buf \U$2827 ( \3074 , \2525 );
buf \U$2828 ( \3075 , \3074 );
and \U$2829 ( \3076 , RIbe28480_21, RIbe286d8_26);
nor \U$2830 ( \3077 , RIbe28480_21, RIbe286d8_26);
nor \U$2831 ( \3078 , \3076 , \3077 );
and \U$2832 ( \3079 , \3075 , \3078 );
nor \U$2833 ( \3080 , \3073 , \3079 );
xnor \U$2834 ( \3081 , \3070 , \3080 );
xor \U$2835 ( \3082 , \3062 , \3081 );
not \U$2836 ( \3083 , \3082 );
and \U$2837 ( \3084 , \3055 , \3083 );
and \U$2838 ( \3085 , \3054 , \3082 );
nor \U$2839 ( \3086 , \3084 , \3085 );
not \U$2840 ( \3087 , \3086 );
xor \U$2841 ( \3088 , RIbe290b0_47, RIbe29b00_69);
not \U$2842 ( \3089 , \3088 );
not \U$2843 ( \3090 , \2731 );
or \U$2844 ( \3091 , \3089 , \3090 );
nand \U$2845 ( \3092 , \2071 , \2727 );
nand \U$2846 ( \3093 , \3091 , \3092 );
xor \U$2847 ( \3094 , RIbe28cf0_39, RIbe27b98_2);
not \U$2848 ( \3095 , \3094 );
not \U$2849 ( \3096 , \546 );
or \U$2850 ( \3097 , \3095 , \3096 );
nand \U$2851 ( \3098 , \1734 , \2434 );
nand \U$2852 ( \3099 , \3097 , \3098 );
or \U$2853 ( \3100 , \3093 , \3099 );
xor \U$2854 ( \3101 , RIbe28de0_41, RIbe29998_66);
not \U$2855 ( \3102 , \3101 );
buf \U$2856 ( \3103 , \924 );
not \U$2857 ( \3104 , \3103 );
or \U$2858 ( \3105 , \3102 , \3104 );
nand \U$2859 ( \3106 , \514 , \2676 );
nand \U$2860 ( \3107 , \3105 , \3106 );
nand \U$2861 ( \3108 , \3100 , \3107 );
nand \U$2862 ( \3109 , \3099 , \3093 );
nand \U$2863 ( \3110 , \3108 , \3109 );
xor \U$2864 ( \3111 , \3110 , \2568 );
not \U$2865 ( \3112 , \1782 );
not \U$2866 ( \3113 , RIbe28a20_33);
not \U$2867 ( \3114 , RIbe293f8_54);
and \U$2868 ( \3115 , \3113 , \3114 );
and \U$2869 ( \3116 , RIbe28a20_33, RIbe293f8_54);
nor \U$2870 ( \3117 , \3115 , \3116 );
not \U$2871 ( \3118 , \3117 );
not \U$2872 ( \3119 , \3118 );
and \U$2873 ( \3120 , \3112 , \3119 );
not \U$2874 ( \3121 , RIbe28a20_33);
not \U$2875 ( \3122 , RIbe29308_52);
and \U$2876 ( \3123 , \3121 , \3122 );
and \U$2877 ( \3124 , RIbe28a20_33, RIbe29308_52);
nor \U$2878 ( \3125 , \3123 , \3124 );
and \U$2879 ( \3126 , \1769 , \3125 );
nor \U$2880 ( \3127 , \3120 , \3126 );
not \U$2881 ( \3128 , \3127 );
not \U$2882 ( \3129 , \3128 );
not \U$2883 ( \3130 , \2422 );
not \U$2884 ( \3131 , \314 );
or \U$2885 ( \3132 , \3130 , \3131 );
xor \U$2886 ( \3133 , RIbe27d78_6, RIbe29218_50);
nand \U$2887 ( \3134 , \1613 , \3133 );
nand \U$2888 ( \3135 , \3132 , \3134 );
not \U$2889 ( \3136 , \3135 );
not \U$2890 ( \3137 , \2718 );
xnor \U$2891 ( \3138 , RIbe29380_53, RIbe27fd0_11);
not \U$2892 ( \3139 , \3138 );
and \U$2893 ( \3140 , \3137 , \3139 );
and \U$2894 ( \3141 , \2707 , RIbe27fd0_11);
nor \U$2895 ( \3142 , \3140 , \3141 );
not \U$2896 ( \3143 , \3142 );
or \U$2897 ( \3144 , \3136 , \3143 );
or \U$2898 ( \3145 , \3135 , \3142 );
nand \U$2899 ( \3146 , \3144 , \3145 );
not \U$2900 ( \3147 , \3146 );
or \U$2901 ( \3148 , \3129 , \3147 );
not \U$2902 ( \3149 , \3142 );
nand \U$2903 ( \3150 , \3149 , \3135 );
nand \U$2904 ( \3151 , \3148 , \3150 );
and \U$2905 ( \3152 , \3111 , \3151 );
and \U$2906 ( \3153 , \3110 , \2568 );
nor \U$2907 ( \3154 , \3152 , \3153 );
not \U$2908 ( \3155 , \3154 );
and \U$2909 ( \3156 , \3087 , \3155 );
not \U$2910 ( \3157 , \3082 );
and \U$2911 ( \3158 , \3054 , \3157 );
nor \U$2912 ( \3159 , \3156 , \3158 );
and \U$2913 ( \3160 , \282 , \2847 );
xor \U$2914 ( \3161 , RIbe28138_14, RIbe29038_46);
and \U$2915 ( \3162 , \287 , \3161 );
nor \U$2916 ( \3163 , \3160 , \3162 );
not \U$2917 ( \3164 , \259 );
not \U$2918 ( \3165 , \3007 );
not \U$2919 ( \3166 , \3165 );
and \U$2920 ( \3167 , \3164 , \3166 );
xor \U$2921 ( \3168 , RIbe27c88_4, RIbe27b98_2);
and \U$2922 ( \3169 , \1298 , \3168 );
nor \U$2923 ( \3170 , \3167 , \3169 );
xor \U$2924 ( \3171 , \3163 , \3170 );
and \U$2925 ( \3172 , \1452 , \2882 );
and \U$2926 ( \3173 , RIbe296c8_60, RIbe29470_55);
not \U$2927 ( \3174 , RIbe296c8_60);
and \U$2928 ( \3175 , \3174 , \919 );
nor \U$2929 ( \3176 , \3173 , \3175 );
and \U$2930 ( \3177 , \908 , \3176 );
nor \U$2931 ( \3178 , \3172 , \3177 );
xor \U$2932 ( \3179 , \3171 , \3178 );
not \U$2933 ( \3180 , \2997 );
not \U$2934 ( \3181 , \466 );
or \U$2935 ( \3182 , \3180 , \3181 );
and \U$2936 ( \3183 , RIbe290b0_47, RIbe29740_61);
not \U$2937 ( \3184 , RIbe290b0_47);
not \U$2938 ( \3185 , RIbe29740_61);
and \U$2939 ( \3186 , \3184 , \3185 );
nor \U$2940 ( \3187 , \3183 , \3186 );
nand \U$2941 ( \3188 , \2071 , \3187 );
nand \U$2942 ( \3189 , \3182 , \3188 );
not \U$2943 ( \3190 , \2870 );
not \U$2944 ( \3191 , \2276 );
or \U$2945 ( \3192 , \3190 , \3191 );
xnor \U$2946 ( \3193 , RIbe28318_18, RIbe28a20_33);
not \U$2947 ( \3194 , \3193 );
nand \U$2948 ( \3195 , \3194 , \2476 );
nand \U$2949 ( \3196 , \3192 , \3195 );
not \U$2950 ( \3197 , \3196 );
and \U$2951 ( \3198 , \3189 , \3197 );
not \U$2952 ( \3199 , \3189 );
and \U$2953 ( \3200 , \3199 , \3196 );
or \U$2954 ( \3201 , \3198 , \3200 );
and \U$2955 ( \3202 , \3201 , \3030 );
not \U$2956 ( \3203 , \3201 );
not \U$2957 ( \3204 , \3030 );
and \U$2958 ( \3205 , \3203 , \3204 );
nor \U$2959 ( \3206 , \3202 , \3205 );
xor \U$2960 ( \3207 , \3179 , \3206 );
not \U$2961 ( \3208 , \3207 );
not \U$2962 ( \3209 , \2817 );
not \U$2963 ( \3210 , \2805 );
or \U$2964 ( \3211 , \3209 , \3210 );
not \U$2965 ( \3212 , \2808 );
nand \U$2966 ( \3213 , \3212 , \2813 );
nand \U$2967 ( \3214 , \3211 , \3213 );
not \U$2968 ( \3215 , \3214 );
not \U$2969 ( \3216 , \3215 );
or \U$2970 ( \3217 , \3208 , \3216 );
or \U$2971 ( \3218 , \3215 , \3207 );
nand \U$2972 ( \3219 , \3217 , \3218 );
xnor \U$2973 ( \3220 , \3159 , \3219 );
or \U$2974 ( \3221 , \2972 , \3013 );
not \U$2975 ( \3222 , \2968 );
or \U$2976 ( \3223 , \3222 , \2922 );
nand \U$2977 ( \3224 , \3221 , \3223 );
xnor \U$2978 ( \3225 , \3220 , \3224 );
not \U$2979 ( \3226 , \3225 );
not \U$2980 ( \3227 , \3226 );
not \U$2981 ( \3228 , \3154 );
and \U$2982 ( \3229 , \3086 , \3228 );
not \U$2983 ( \3230 , \3086 );
and \U$2984 ( \3231 , \3230 , \3154 );
nor \U$2985 ( \3232 , \3229 , \3231 );
not \U$2986 ( \3233 , \3232 );
not \U$2987 ( \3234 , \3233 );
not \U$2988 ( \3235 , RIbe280c0_13);
not \U$2989 ( \3236 , RIbe297b8_62);
and \U$2990 ( \3237 , \3235 , \3236 );
and \U$2991 ( \3238 , RIbe280c0_13, RIbe297b8_62);
nor \U$2992 ( \3239 , \3237 , \3238 );
not \U$2993 ( \3240 , \3239 );
not \U$2994 ( \3241 , \862 );
or \U$2995 ( \3242 , \3240 , \3241 );
not \U$2996 ( \3243 , \2652 );
nand \U$2997 ( \3244 , \3243 , \869 );
nand \U$2998 ( \3245 , \3242 , \3244 );
not \U$2999 ( \3246 , \3245 );
xor \U$3000 ( \3247 , RIbe29bf0_71, RIbe29c68_72);
buf \U$3001 ( \3248 , \3247 );
buf \U$3002 ( \3249 , \3248 );
not \U$3003 ( \3250 , \3249 );
not \U$3004 ( \3251 , \3250 );
not \U$3005 ( \3252 , \3247 );
xor \U$3006 ( \3253 , RIbe28f48_44, RIbe29bf0_71);
nand \U$3007 ( \3254 , \3252 , \3253 );
buf \U$3008 ( \3255 , \3254 );
not \U$3009 ( \3256 , \3255 );
not \U$3010 ( \3257 , \3256 );
not \U$3011 ( \3258 , \3257 );
or \U$3012 ( \3259 , \3251 , \3258 );
nand \U$3013 ( \3260 , \3259 , RIbe28f48_44);
xor \U$3014 ( \3261 , RIbe285e8_24, RIbe28840_29);
not \U$3015 ( \3262 , \3261 );
not \U$3016 ( \3263 , \2618 );
or \U$3017 ( \3264 , \3262 , \3263 );
nand \U$3018 ( \3265 , \2626 , \2608 );
nand \U$3019 ( \3266 , \3264 , \3265 );
nor \U$3020 ( \3267 , \3260 , \3266 );
or \U$3021 ( \3268 , \3246 , \3267 );
nand \U$3022 ( \3269 , \3260 , \3266 );
nand \U$3023 ( \3270 , \3268 , \3269 );
not \U$3024 ( \3271 , \3270 );
xor \U$3025 ( \3272 , RIbe28228_16, RIbe282a0_17);
not \U$3026 ( \3273 , \3272 );
not \U$3027 ( \3274 , \1061 );
or \U$3028 ( \3275 , \3273 , \3274 );
nand \U$3029 ( \3276 , \885 , \2957 );
nand \U$3030 ( \3277 , \3275 , \3276 );
xor \U$3031 ( \3278 , RIbe29038_46, RIbe29128_48);
not \U$3032 ( \3279 , \3278 );
not \U$3033 ( \3280 , \979 );
or \U$3034 ( \3281 , \3279 , \3280 );
nand \U$3035 ( \3282 , \1805 , \2945 );
nand \U$3036 ( \3283 , \3281 , \3282 );
xor \U$3037 ( \3284 , \3277 , \3283 );
xnor \U$3038 ( \3285 , RIbe295d8_58, RIbe296c8_60);
or \U$3039 ( \3286 , \2020 , \3285 );
or \U$3040 ( \3287 , \1226 , \2938 );
nand \U$3041 ( \3288 , \3286 , \3287 );
and \U$3042 ( \3289 , \3284 , \3288 );
and \U$3043 ( \3290 , \3277 , \3283 );
or \U$3044 ( \3291 , \3289 , \3290 );
not \U$3045 ( \3292 , \3291 );
or \U$3046 ( \3293 , \3271 , \3292 );
xor \U$3047 ( \3294 , RIbe27d78_6, RIbe27df0_7);
not \U$3048 ( \3295 , \3294 );
not \U$3049 ( \3296 , \2052 );
or \U$3050 ( \3297 , \3295 , \3296 );
nand \U$3051 ( \3298 , \315 , \3133 );
nand \U$3052 ( \3299 , \3297 , \3298 );
not \U$3053 ( \3300 , \3094 );
not \U$3054 ( \3301 , \1298 );
or \U$3055 ( \3302 , \3300 , \3301 );
or \U$3056 ( \3303 , RIbe27b20_1, RIbe27b98_2);
and \U$3057 ( \3304 , \3303 , \2589 );
nand \U$3058 ( \3305 , \546 , \3304 );
nand \U$3059 ( \3306 , \3302 , \3305 );
xor \U$3060 ( \3307 , \3299 , \3306 );
not \U$3061 ( \3308 , \2597 );
not \U$3062 ( \3309 , \2464 );
or \U$3063 ( \3310 , \3308 , \3309 );
not \U$3064 ( \3311 , \2600 );
xnor \U$3065 ( \3312 , RIbe27e68_8, RIbe286d8_26);
or \U$3066 ( \3313 , \3311 , \3312 );
nand \U$3067 ( \3314 , \3310 , \3313 );
and \U$3068 ( \3315 , \3307 , \3314 );
and \U$3069 ( \3316 , \3299 , \3306 );
nor \U$3070 ( \3317 , \3315 , \3316 );
not \U$3071 ( \3318 , \3317 );
xor \U$3072 ( \3319 , \3270 , \3291 );
nand \U$3073 ( \3320 , \3318 , \3319 );
nand \U$3074 ( \3321 , \3293 , \3320 );
not \U$3075 ( \3322 , \3321 );
and \U$3076 ( \3323 , \2540 , \2569 );
and \U$3077 ( \3324 , \2539 , \2529 );
nor \U$3078 ( \3325 , \3323 , \3324 );
not \U$3079 ( \3326 , \3325 );
nand \U$3080 ( \3327 , RIbe27b98_2, RIbe29b78_70);
not \U$3081 ( \3328 , \3327 );
not \U$3082 ( \3329 , RIbe28de0_41);
not \U$3083 ( \3330 , RIbe298a8_64);
and \U$3084 ( \3331 , \3329 , \3330 );
and \U$3085 ( \3332 , RIbe28de0_41, RIbe298a8_64);
nor \U$3086 ( \3333 , \3331 , \3332 );
not \U$3087 ( \3334 , \3333 );
not \U$3088 ( \3335 , \332 );
or \U$3089 ( \3336 , \3334 , \3335 );
nand \U$3090 ( \3337 , \514 , \3101 );
nand \U$3091 ( \3338 , \3336 , \3337 );
not \U$3092 ( \3339 , \3338 );
or \U$3093 ( \3340 , \3328 , \3339 );
or \U$3094 ( \3341 , \3338 , \3327 );
nand \U$3095 ( \3342 , \3340 , \3341 );
not \U$3096 ( \3343 , \3342 );
buf \U$3097 ( \3344 , \2518 );
not \U$3098 ( \3345 , \3344 );
xnor \U$3099 ( \3346 , RIbe28480_21, RIbe284f8_22);
or \U$3100 ( \3347 , \3345 , \3346 );
or \U$3101 ( \3348 , \2672 , \2509 );
nand \U$3102 ( \3349 , \3347 , \3348 );
not \U$3103 ( \3350 , \3349 );
or \U$3104 ( \3351 , \3343 , \3350 );
not \U$3105 ( \3352 , \3327 );
nand \U$3106 ( \3353 , \3352 , \3338 );
nand \U$3107 ( \3354 , \3351 , \3353 );
not \U$3108 ( \3355 , \3354 );
not \U$3109 ( \3356 , \524 );
not \U$3110 ( \3357 , RIbe29a10_67);
not \U$3111 ( \3358 , RIbe290b0_47);
or \U$3112 ( \3359 , \3357 , \3358 );
or \U$3113 ( \3360 , RIbe290b0_47, RIbe29a10_67);
nand \U$3114 ( \3361 , \3359 , \3360 );
not \U$3115 ( \3362 , \3361 );
and \U$3116 ( \3363 , \3356 , \3362 );
and \U$3117 ( \3364 , \469 , \3088 );
nor \U$3118 ( \3365 , \3363 , \3364 );
and \U$3119 ( \3366 , RIbe28a20_33, RIbe28a98_34);
not \U$3120 ( \3367 , RIbe28a20_33);
and \U$3121 ( \3368 , \3367 , \940 );
nor \U$3122 ( \3369 , \3366 , \3368 );
not \U$3123 ( \3370 , \3369 );
not \U$3124 ( \3371 , \2276 );
or \U$3125 ( \3372 , \3370 , \3371 );
nand \U$3126 ( \3373 , \2475 , \3117 );
nand \U$3127 ( \3374 , \3372 , \3373 );
xor \U$3128 ( \3375 , RIbe27fd0_11, RIbe28048_12);
not \U$3129 ( \3376 , \3375 );
not \U$3130 ( \3377 , \2717 );
buf \U$3131 ( \3378 , \3377 );
not \U$3132 ( \3379 , \3378 );
or \U$3133 ( \3380 , \3376 , \3379 );
not \U$3134 ( \3381 , \3138 );
nand \U$3135 ( \3382 , \3381 , \2707 );
nand \U$3136 ( \3383 , \3380 , \3382 );
nor \U$3137 ( \3384 , \3374 , \3383 );
or \U$3138 ( \3385 , \3365 , \3384 );
nand \U$3139 ( \3386 , \3374 , \3383 );
nand \U$3140 ( \3387 , \3385 , \3386 );
not \U$3141 ( \3388 , \3387 );
or \U$3142 ( \3389 , \3355 , \3388 );
or \U$3143 ( \3390 , \3354 , \3387 );
and \U$3144 ( \3391 , RIbe27c10_3, RIbe28d68_40);
nor \U$3145 ( \3392 , RIbe27c10_3, RIbe28d68_40);
nor \U$3146 ( \3393 , \3391 , \3392 );
not \U$3147 ( \3394 , \3393 );
not \U$3148 ( \3395 , \361 );
or \U$3149 ( \3396 , \3394 , \3395 );
nand \U$3150 ( \3397 , \370 , \2580 );
nand \U$3151 ( \3398 , \3396 , \3397 );
xor \U$3152 ( \3399 , RIbe28b88_36, RIbe29308_52);
not \U$3153 ( \3400 , \3399 );
buf \U$3154 ( \3401 , \2552 );
buf \U$3155 ( \3402 , \3401 );
not \U$3156 ( \3403 , \3402 );
or \U$3157 ( \3404 , \3400 , \3403 );
nand \U$3158 ( \3405 , \2561 , \2544 );
nand \U$3159 ( \3406 , \3404 , \3405 );
xor \U$3160 ( \3407 , \3398 , \3406 );
not \U$3161 ( \3408 , \2638 );
not \U$3162 ( \3409 , \3408 );
xnor \U$3163 ( \3410 , RIbe28390_19, RIbe28c78_38);
or \U$3164 ( \3411 , \3409 , \3410 );
not \U$3165 ( \3412 , \2648 );
not \U$3166 ( \3413 , \2632 );
or \U$3167 ( \3414 , \3412 , \3413 );
nand \U$3168 ( \3415 , \3411 , \3414 );
and \U$3169 ( \3416 , \3407 , \3415 );
and \U$3170 ( \3417 , \3398 , \3406 );
or \U$3171 ( \3418 , \3416 , \3417 );
nand \U$3172 ( \3419 , \3390 , \3418 );
nand \U$3173 ( \3420 , \3389 , \3419 );
not \U$3174 ( \3421 , \3420 );
or \U$3175 ( \3422 , \3326 , \3421 );
or \U$3176 ( \3423 , \3325 , \3420 );
nand \U$3177 ( \3424 , \3422 , \3423 );
not \U$3178 ( \3425 , \3424 );
or \U$3179 ( \3426 , \3322 , \3425 );
not \U$3180 ( \3427 , \3325 );
nand \U$3181 ( \3428 , \3427 , \3420 );
nand \U$3182 ( \3429 , \3426 , \3428 );
not \U$3183 ( \3430 , \3429 );
or \U$3184 ( \3431 , \3234 , \3430 );
xor \U$3185 ( \3432 , \3099 , \3107 );
xor \U$3186 ( \3433 , \3093 , \3432 );
and \U$3187 ( \3434 , \3146 , \3127 );
not \U$3188 ( \3435 , \3146 );
and \U$3189 ( \3436 , \3435 , \3128 );
or \U$3190 ( \3437 , \3434 , \3436 );
xor \U$3191 ( \3438 , \3433 , \3437 );
not \U$3192 ( \3439 , \2960 );
not \U$3193 ( \3440 , \2952 );
or \U$3194 ( \3441 , \3439 , \3440 );
or \U$3195 ( \3442 , \2952 , \2960 );
nand \U$3196 ( \3443 , \3441 , \3442 );
and \U$3197 ( \3444 , \3438 , \3443 );
and \U$3198 ( \3445 , \3433 , \3437 );
or \U$3199 ( \3446 , \3444 , \3445 );
and \U$3200 ( \3447 , \3110 , \2569 );
not \U$3201 ( \3448 , \3110 );
and \U$3202 ( \3449 , \3448 , \2568 );
nor \U$3203 ( \3450 , \3447 , \3449 );
xor \U$3204 ( \3451 , \3450 , \3151 );
xnor \U$3205 ( \3452 , \3446 , \3451 );
xor \U$3206 ( \3453 , \2964 , \2937 );
and \U$3207 ( \3454 , \3452 , \3453 );
not \U$3208 ( \3455 , \3446 );
nor \U$3209 ( \3456 , \3455 , \3451 );
nor \U$3210 ( \3457 , \3454 , \3456 );
not \U$3211 ( \3458 , \3457 );
xnor \U$3212 ( \3459 , \3429 , \3232 );
nand \U$3213 ( \3460 , \3458 , \3459 );
nand \U$3214 ( \3461 , \3431 , \3460 );
not \U$3215 ( \3462 , \3461 );
not \U$3216 ( \3463 , \3462 );
or \U$3217 ( \3464 , \3227 , \3463 );
nand \U$3218 ( \3465 , \3461 , \3225 );
nand \U$3219 ( \3466 , \3464 , \3465 );
not \U$3220 ( \3467 , \3466 );
or \U$3221 ( \3468 , \3019 , \3467 );
nand \U$3222 ( \3469 , \3461 , \3226 );
nand \U$3223 ( \3470 , \3468 , \3469 );
nand \U$3224 ( \3471 , RIbe27b98_2, RIbe29998_66);
not \U$3225 ( \3472 , \3471 );
not \U$3226 ( \3473 , \2860 );
not \U$3227 ( \3474 , \3103 );
or \U$3228 ( \3475 , \3473 , \3474 );
xor \U$3229 ( \3476 , RIbe28de0_41, RIbe29218_50);
nand \U$3230 ( \3477 , \347 , \3476 );
nand \U$3231 ( \3478 , \3475 , \3477 );
not \U$3232 ( \3479 , \3478 );
or \U$3233 ( \3480 , \3472 , \3479 );
or \U$3234 ( \3481 , \3471 , \3478 );
nand \U$3235 ( \3482 , \3480 , \3481 );
buf \U$3236 ( \3483 , \2518 );
not \U$3237 ( \3484 , \3483 );
not \U$3238 ( \3485 , \3484 );
and \U$3239 ( \3486 , \3485 , \3078 );
and \U$3240 ( \3487 , RIbe27ee0_9, RIbe28480_21);
nor \U$3241 ( \3488 , RIbe27ee0_9, RIbe28480_21);
nor \U$3242 ( \3489 , \3487 , \3488 );
and \U$3243 ( \3490 , \2527 , \3489 );
nor \U$3244 ( \3491 , \3486 , \3490 );
and \U$3245 ( \3492 , \3482 , \3491 );
not \U$3246 ( \3493 , \3482 );
not \U$3247 ( \3494 , \3491 );
and \U$3248 ( \3495 , \3493 , \3494 );
nor \U$3249 ( \3496 , \3492 , \3495 );
not \U$3250 ( \3497 , \3496 );
not \U$3251 ( \3498 , \2618 );
not \U$3252 ( \3499 , \3498 );
not \U$3253 ( \3500 , \2895 );
and \U$3254 ( \3501 , \3499 , \3500 );
not \U$3255 ( \3502 , \2625 );
and \U$3256 ( \3503 , RIbe285e8_24, \388 );
not \U$3257 ( \3504 , RIbe285e8_24);
and \U$3258 ( \3505 , \3504 , RIbe29380_53);
nor \U$3259 ( \3506 , \3503 , \3505 );
nor \U$3260 ( \3507 , \3502 , \3506 );
nor \U$3261 ( \3508 , \3501 , \3507 );
not \U$3262 ( \3509 , \1325 );
not \U$3263 ( \3510 , \2834 );
and \U$3264 ( \3511 , \3509 , \3510 );
xnor \U$3265 ( \3512 , RIbe280c0_13, RIbe288b8_30);
nor \U$3266 ( \3513 , \1264 , \3512 );
nor \U$3267 ( \3514 , \3511 , \3513 );
xor \U$3268 ( \3515 , \3508 , \3514 );
and \U$3269 ( \3516 , \1061 , \3060 );
or \U$3270 ( \3517 , \888 , RIbe293f8_54);
or \U$3271 ( \3518 , \2489 , RIbe28228_16);
nand \U$3272 ( \3519 , \3517 , \3518 );
and \U$3273 ( \3520 , \885 , \3519 );
nor \U$3274 ( \3521 , \3516 , \3520 );
xor \U$3275 ( \3522 , \3515 , \3521 );
not \U$3276 ( \3523 , \3522 );
not \U$3277 ( \3524 , \3523 );
not \U$3278 ( \3525 , \1093 );
xnor \U$3279 ( \3526 , RIbe27d78_6, RIbe291a0_49);
not \U$3280 ( \3527 , \3526 );
and \U$3281 ( \3528 , \3525 , \3527 );
and \U$3282 ( \3529 , \1613 , \3037 );
nor \U$3283 ( \3530 , \3528 , \3529 );
not \U$3284 ( \3531 , \967 );
not \U$3285 ( \3532 , \3067 );
and \U$3286 ( \3533 , \3531 , \3532 );
and \U$3287 ( \3534 , RIbe28930_31, RIbe28c00_37);
nor \U$3288 ( \3535 , RIbe28930_31, RIbe28c00_37);
nor \U$3289 ( \3536 , \3534 , \3535 );
and \U$3290 ( \3537 , \971 , \3536 );
nor \U$3291 ( \3538 , \3533 , \3537 );
xor \U$3292 ( \3539 , \3530 , \3538 );
not \U$3293 ( \3540 , \2603 );
and \U$3294 ( \3541 , \3311 , \3540 );
nor \U$3295 ( \3542 , \3541 , \2594 );
xor \U$3296 ( \3543 , \3539 , \3542 );
not \U$3297 ( \3544 , \3543 );
or \U$3298 ( \3545 , \3524 , \3544 );
or \U$3299 ( \3546 , \3543 , \3523 );
nand \U$3300 ( \3547 , \3545 , \3546 );
not \U$3301 ( \3548 , \3547 );
or \U$3302 ( \3549 , \3497 , \3548 );
or \U$3303 ( \3550 , \3496 , \3547 );
nand \U$3304 ( \3551 , \3549 , \3550 );
not \U$3305 ( \3552 , \3551 );
not \U$3306 ( \3553 , \2911 );
not \U$3307 ( \3554 , \2889 );
or \U$3308 ( \3555 , \3553 , \3554 );
not \U$3309 ( \3556 , \2885 );
nand \U$3310 ( \3557 , \3556 , \2854 );
nand \U$3311 ( \3558 , \3555 , \3557 );
not \U$3312 ( \3559 , \3012 );
not \U$3313 ( \3560 , \2988 );
or \U$3314 ( \3561 , \3559 , \3560 );
not \U$3315 ( \3562 , \2978 );
nand \U$3316 ( \3563 , \3562 , \2984 );
nand \U$3317 ( \3564 , \3561 , \3563 );
xor \U$3318 ( \3565 , \3558 , \3564 );
not \U$3319 ( \3566 , \3565 );
or \U$3320 ( \3567 , \3552 , \3566 );
nand \U$3321 ( \3568 , \3564 , \3558 );
nand \U$3322 ( \3569 , \3567 , \3568 );
not \U$3323 ( \3570 , \2907 );
not \U$3324 ( \3571 , \2640 );
or \U$3325 ( \3572 , \3570 , \3571 );
not \U$3326 ( \3573 , RIbe28390_19);
not \U$3327 ( \3574 , RIbe28570_23);
and \U$3328 ( \3575 , \3573 , \3574 );
and \U$3329 ( \3576 , RIbe28390_19, RIbe28570_23);
nor \U$3330 ( \3577 , \3575 , \3576 );
nand \U$3331 ( \3578 , \2648 , \3577 );
nand \U$3332 ( \3579 , \3572 , \3578 );
not \U$3333 ( \3580 , \3579 );
not \U$3334 ( \3581 , \2899 );
not \U$3335 ( \3582 , \3581 );
not \U$3336 ( \3583 , \1493 );
or \U$3337 ( \3584 , \3582 , \3583 );
and \U$3338 ( \3585 , RIbe29b00_69, RIbe27c10_3);
not \U$3339 ( \3586 , RIbe29b00_69);
and \U$3340 ( \3587 , \3586 , \363 );
nor \U$3341 ( \3588 , \3585 , \3587 );
nand \U$3342 ( \3589 , \370 , \3588 );
nand \U$3343 ( \3590 , \3584 , \3589 );
not \U$3344 ( \3591 , \3590 );
or \U$3345 ( \3592 , \3580 , \3591 );
and \U$3346 ( \3593 , \2702 , \3028 );
not \U$3347 ( \3594 , \2692 );
xor \U$3348 ( \3595 , RIbe28750_27, RIbe28b88_36);
and \U$3349 ( \3596 , \3594 , \3595 );
nor \U$3350 ( \3597 , \3593 , \3596 );
not \U$3351 ( \3598 , \3597 );
not \U$3352 ( \3599 , \3579 );
not \U$3353 ( \3600 , \3591 );
or \U$3354 ( \3601 , \3599 , \3600 );
nand \U$3355 ( \3602 , \3580 , \3590 );
nand \U$3356 ( \3603 , \3601 , \3602 );
nand \U$3357 ( \3604 , \3598 , \3603 );
nand \U$3358 ( \3605 , \3592 , \3604 );
not \U$3359 ( \3606 , \3482 );
not \U$3360 ( \3607 , \3494 );
or \U$3361 ( \3608 , \3606 , \3607 );
not \U$3362 ( \3609 , \3471 );
nand \U$3363 ( \3610 , \3609 , \3478 );
nand \U$3364 ( \3611 , \3608 , \3610 );
not \U$3365 ( \3612 , \3595 );
not \U$3366 ( \3613 , \2554 );
or \U$3367 ( \3614 , \3612 , \3613 );
xnor \U$3368 ( \3615 , RIbe28b88_36, RIbe28840_29);
not \U$3369 ( \3616 , \3615 );
nand \U$3370 ( \3617 , \3616 , \2691 );
nand \U$3371 ( \3618 , \3614 , \3617 );
and \U$3372 ( \3619 , \3611 , \3618 );
not \U$3373 ( \3620 , \3611 );
not \U$3374 ( \3621 , \3618 );
and \U$3375 ( \3622 , \3620 , \3621 );
or \U$3376 ( \3623 , \3619 , \3622 );
xor \U$3377 ( \3624 , \3605 , \3623 );
not \U$3378 ( \3625 , \3062 );
not \U$3379 ( \3626 , \3625 );
not \U$3380 ( \3627 , \3081 );
or \U$3381 ( \3628 , \3626 , \3627 );
not \U$3382 ( \3629 , \3080 );
nand \U$3383 ( \3630 , \3629 , \3070 );
nand \U$3384 ( \3631 , \3628 , \3630 );
not \U$3385 ( \3632 , \3631 );
not \U$3386 ( \3633 , \3009 );
not \U$3387 ( \3634 , \2993 );
not \U$3388 ( \3635 , \3634 );
or \U$3389 ( \3636 , \3633 , \3635 );
nand \U$3390 ( \3637 , \3636 , \3003 );
nand \U$3391 ( \3638 , \3010 , \2993 );
nand \U$3392 ( \3639 , \3637 , \3638 );
not \U$3393 ( \3640 , \2862 );
not \U$3394 ( \3641 , \2872 );
or \U$3395 ( \3642 , \3640 , \3641 );
or \U$3396 ( \3643 , \2872 , \2862 );
nand \U$3397 ( \3644 , \3643 , \2884 );
nand \U$3398 ( \3645 , \3642 , \3644 );
xor \U$3399 ( \3646 , \3639 , \3645 );
not \U$3400 ( \3647 , \3646 );
or \U$3401 ( \3648 , \3632 , \3647 );
nand \U$3402 ( \3649 , \3645 , \3639 );
nand \U$3403 ( \3650 , \3648 , \3649 );
and \U$3404 ( \3651 , \3624 , \3650 );
not \U$3405 ( \3652 , \3624 );
not \U$3406 ( \3653 , \3650 );
and \U$3407 ( \3654 , \3652 , \3653 );
nor \U$3408 ( \3655 , \3651 , \3654 );
xor \U$3409 ( \3656 , \3508 , \3514 );
and \U$3410 ( \3657 , \3656 , \3521 );
and \U$3411 ( \3658 , \3508 , \3514 );
or \U$3412 ( \3659 , \3657 , \3658 );
xor \U$3413 ( \3660 , \3530 , \3538 );
and \U$3414 ( \3661 , \3660 , \3542 );
and \U$3415 ( \3662 , \3530 , \3538 );
or \U$3416 ( \3663 , \3661 , \3662 );
xor \U$3417 ( \3664 , \3659 , \3663 );
xor \U$3418 ( \3665 , \3163 , \3170 );
and \U$3419 ( \3666 , \3665 , \3178 );
and \U$3420 ( \3667 , \3163 , \3170 );
or \U$3421 ( \3668 , \3666 , \3667 );
xor \U$3422 ( \3669 , \3664 , \3668 );
not \U$3423 ( \3670 , \3669 );
and \U$3424 ( \3671 , \3655 , \3670 );
not \U$3425 ( \3672 , \3655 );
and \U$3426 ( \3673 , \3672 , \3669 );
nor \U$3427 ( \3674 , \3671 , \3673 );
xnor \U$3428 ( \3675 , \3569 , \3674 );
not \U$3429 ( \3676 , \3543 );
nand \U$3430 ( \3677 , \3522 , \3496 );
nand \U$3431 ( \3678 , \3676 , \3677 );
not \U$3432 ( \3679 , \3496 );
nand \U$3433 ( \3680 , \3679 , \3523 );
and \U$3434 ( \3681 , \3678 , \3680 );
not \U$3435 ( \3682 , \3681 );
not \U$3436 ( \3683 , \3597 );
not \U$3437 ( \3684 , \3603 );
or \U$3438 ( \3685 , \3683 , \3684 );
or \U$3439 ( \3686 , \3603 , \3597 );
nand \U$3440 ( \3687 , \3685 , \3686 );
not \U$3441 ( \3688 , \3687 );
xor \U$3442 ( \3689 , \2897 , \2901 );
and \U$3443 ( \3690 , \3689 , \2910 );
and \U$3444 ( \3691 , \2897 , \2901 );
or \U$3445 ( \3692 , \3690 , \3691 );
not \U$3446 ( \3693 , \2850 );
not \U$3447 ( \3694 , \2841 );
or \U$3448 ( \3695 , \3693 , \3694 );
not \U$3449 ( \3696 , \2829 );
nand \U$3450 ( \3697 , \3696 , \2837 );
nand \U$3451 ( \3698 , \3695 , \3697 );
and \U$3452 ( \3699 , \3692 , \3698 );
not \U$3453 ( \3700 , \3692 );
not \U$3454 ( \3701 , \3698 );
and \U$3455 ( \3702 , \3700 , \3701 );
nor \U$3456 ( \3703 , \3699 , \3702 );
not \U$3457 ( \3704 , \3703 );
or \U$3458 ( \3705 , \3688 , \3704 );
nand \U$3459 ( \3706 , \3698 , \3692 );
nand \U$3460 ( \3707 , \3705 , \3706 );
not \U$3461 ( \3708 , \3707 );
or \U$3462 ( \3709 , \3682 , \3708 );
or \U$3463 ( \3710 , \3707 , \3681 );
nand \U$3464 ( \3711 , \3709 , \3710 );
not \U$3465 ( \3712 , \2638 );
and \U$3466 ( \3713 , \3712 , \3577 );
buf \U$3467 ( \3714 , \2776 );
and \U$3468 ( \3715 , RIbe28390_19, RIbe286d8_26);
nor \U$3469 ( \3716 , RIbe28390_19, RIbe286d8_26);
nor \U$3470 ( \3717 , \3715 , \3716 );
and \U$3471 ( \3718 , \3714 , \3717 );
nor \U$3472 ( \3719 , \3713 , \3718 );
not \U$3473 ( \3720 , \3161 );
not \U$3474 ( \3721 , \979 );
or \U$3475 ( \3722 , \3720 , \3721 );
xnor \U$3476 ( \3723 , RIbe29038_46, RIbe282a0_17);
not \U$3477 ( \3724 , \3723 );
nand \U$3478 ( \3725 , \3724 , \287 );
nand \U$3479 ( \3726 , \3722 , \3725 );
not \U$3480 ( \3727 , \3176 );
not \U$3481 ( \3728 , \1130 );
or \U$3482 ( \3729 , \3727 , \3728 );
and \U$3483 ( \3730 , RIbe294e8_56, RIbe296c8_60);
nor \U$3484 ( \3731 , RIbe294e8_56, RIbe296c8_60);
nor \U$3485 ( \3732 , \3730 , \3731 );
nand \U$3486 ( \3733 , \908 , \3732 );
nand \U$3487 ( \3734 , \3729 , \3733 );
xor \U$3488 ( \3735 , \3726 , \3734 );
xnor \U$3489 ( \3736 , \3719 , \3735 );
not \U$3490 ( \3737 , \3476 );
not \U$3491 ( \3738 , \332 );
or \U$3492 ( \3739 , \3737 , \3738 );
xor \U$3493 ( \3740 , RIbe28de0_41, RIbe29a10_67);
nand \U$3494 ( \3741 , \1149 , \3740 );
nand \U$3495 ( \3742 , \3739 , \3741 );
not \U$3496 ( \3743 , \314 );
xor \U$3497 ( \3744 , RIbe27d78_6, RIbe295d8_58);
not \U$3498 ( \3745 , \3744 );
or \U$3499 ( \3746 , \3743 , \3745 );
or \U$3500 ( \3747 , \300 , \3526 );
nand \U$3501 ( \3748 , \3746 , \3747 );
xor \U$3502 ( \3749 , \3742 , \3748 );
not \U$3503 ( \3750 , \2276 );
or \U$3504 ( \3751 , \3750 , \3193 );
not \U$3505 ( \3752 , RIbe284f8_22);
and \U$3506 ( \3753 , RIbe28a20_33, \3752 );
not \U$3507 ( \3754 , RIbe28a20_33);
and \U$3508 ( \3755 , \3754 , RIbe284f8_22);
nor \U$3509 ( \3756 , \3753 , \3755 );
or \U$3510 ( \3757 , \1770 , \3756 );
nand \U$3511 ( \3758 , \3751 , \3757 );
xor \U$3512 ( \3759 , \3749 , \3758 );
xor \U$3513 ( \3760 , \3736 , \3759 );
not \U$3514 ( \3761 , \3489 );
not \U$3515 ( \3762 , \2520 );
or \U$3516 ( \3763 , \3761 , \3762 );
and \U$3517 ( \3764 , RIbe28480_21, \431 );
not \U$3518 ( \3765 , RIbe28480_21);
and \U$3519 ( \3766 , \3765 , RIbe28048_12);
nor \U$3520 ( \3767 , \3764 , \3766 );
or \U$3521 ( \3768 , \2672 , \3767 );
nand \U$3522 ( \3769 , \3763 , \3768 );
not \U$3523 ( \3770 , \3168 );
not \U$3524 ( \3771 , \258 );
or \U$3525 ( \3772 , \3770 , \3771 );
and \U$3526 ( \3773 , RIbe27df0_7, \713 );
not \U$3527 ( \3774 , RIbe27df0_7);
and \U$3528 ( \3775 , \3774 , RIbe27b98_2);
nor \U$3529 ( \3776 , \3773 , \3775 );
not \U$3530 ( \3777 , \3776 );
nand \U$3531 ( \3778 , \3777 , \1298 );
nand \U$3532 ( \3779 , \3772 , \3778 );
not \U$3533 ( \3780 , \3187 );
not \U$3534 ( \3781 , \466 );
or \U$3535 ( \3782 , \3780 , \3781 );
xnor \U$3536 ( \3783 , RIbe297b8_62, RIbe290b0_47);
not \U$3537 ( \3784 , \3783 );
nand \U$3538 ( \3785 , \3784 , \469 );
nand \U$3539 ( \3786 , \3782 , \3785 );
xor \U$3540 ( \3787 , \3779 , \3786 );
xor \U$3541 ( \3788 , \3769 , \3787 );
xor \U$3542 ( \3789 , \3760 , \3788 );
xnor \U$3543 ( \3790 , \3711 , \3789 );
xnor \U$3544 ( \3791 , \3675 , \3790 );
not \U$3545 ( \3792 , \3791 );
xor \U$3546 ( \3793 , \3565 , \3551 );
not \U$3547 ( \3794 , \3793 );
not \U$3548 ( \3795 , \3050 );
not \U$3549 ( \3796 , \3043 );
not \U$3550 ( \3797 , \3796 );
or \U$3551 ( \3798 , \3795 , \3797 );
or \U$3552 ( \3799 , \3204 , \3039 );
nand \U$3553 ( \3800 , \3798 , \3799 );
not \U$3554 ( \3801 , \3800 );
xor \U$3555 ( \3802 , \3631 , \3646 );
not \U$3556 ( \3803 , \3802 );
not \U$3557 ( \3804 , \3803 );
or \U$3558 ( \3805 , \3801 , \3804 );
not \U$3559 ( \3806 , \3800 );
nand \U$3560 ( \3807 , \3806 , \3802 );
nand \U$3561 ( \3808 , \3805 , \3807 );
not \U$3562 ( \3809 , \3808 );
xnor \U$3563 ( \3810 , \3687 , \3703 );
not \U$3564 ( \3811 , \3810 );
and \U$3565 ( \3812 , \3809 , \3811 );
and \U$3566 ( \3813 , \3808 , \3810 );
nor \U$3567 ( \3814 , \3812 , \3813 );
not \U$3568 ( \3815 , \3814 );
not \U$3569 ( \3816 , \2912 );
not \U$3570 ( \3817 , \2828 );
or \U$3571 ( \3818 , \3816 , \3817 );
nand \U$3572 ( \3819 , \2818 , \2823 );
nand \U$3573 ( \3820 , \3818 , \3819 );
not \U$3574 ( \3821 , \3820 );
or \U$3575 ( \3822 , \3815 , \3821 );
or \U$3576 ( \3823 , \3820 , \3814 );
nand \U$3577 ( \3824 , \3822 , \3823 );
not \U$3578 ( \3825 , \3824 );
or \U$3579 ( \3826 , \3794 , \3825 );
not \U$3580 ( \3827 , \3814 );
nand \U$3581 ( \3828 , \3827 , \3820 );
nand \U$3582 ( \3829 , \3826 , \3828 );
not \U$3583 ( \3830 , \3829 );
not \U$3584 ( \3831 , \3830 );
not \U$3585 ( \3832 , \3224 );
not \U$3586 ( \3833 , \3220 );
or \U$3587 ( \3834 , \3832 , \3833 );
not \U$3588 ( \3835 , \3159 );
nand \U$3589 ( \3836 , \3835 , \3219 );
nand \U$3590 ( \3837 , \3834 , \3836 );
not \U$3591 ( \3838 , \3837 );
and \U$3592 ( \3839 , \3056 , \3519 );
not \U$3593 ( \3840 , RIbe29308_52);
and \U$3594 ( \3841 , \888 , \3840 );
and \U$3595 ( \3842 , RIbe28228_16, RIbe29308_52);
nor \U$3596 ( \3843 , \3841 , \3842 );
and \U$3597 ( \3844 , \885 , \3843 );
nor \U$3598 ( \3845 , \3839 , \3844 );
not \U$3599 ( \3846 , \1054 );
not \U$3600 ( \3847 , \3846 );
not \U$3601 ( \3848 , \3512 );
and \U$3602 ( \3849 , \3847 , \3848 );
and \U$3603 ( \3850 , RIbe280c0_13, RIbe28a98_34);
not \U$3604 ( \3851 , RIbe280c0_13);
and \U$3605 ( \3852 , \3851 , \940 );
nor \U$3606 ( \3853 , \3850 , \3852 );
and \U$3607 ( \3854 , \1265 , \3853 );
nor \U$3608 ( \3855 , \3849 , \3854 );
xor \U$3609 ( \3856 , \3845 , \3855 );
and \U$3610 ( \3857 , \1793 , \3536 );
not \U$3611 ( \3858 , RIbe28c78_38);
not \U$3612 ( \3859 , RIbe28930_31);
or \U$3613 ( \3860 , \3858 , \3859 );
or \U$3614 ( \3861 , RIbe28930_31, RIbe28c78_38);
nand \U$3615 ( \3862 , \3860 , \3861 );
not \U$3616 ( \3863 , \3862 );
and \U$3617 ( \3864 , \971 , \3863 );
nor \U$3618 ( \3865 , \3857 , \3864 );
xor \U$3619 ( \3866 , \3856 , \3865 );
not \U$3620 ( \3867 , \3866 );
not \U$3621 ( \3868 , \3196 );
not \U$3622 ( \3869 , \3204 );
or \U$3623 ( \3870 , \3868 , \3869 );
not \U$3624 ( \3871 , \3197 );
not \U$3625 ( \3872 , \3030 );
or \U$3626 ( \3873 , \3871 , \3872 );
nand \U$3627 ( \3874 , \3873 , \3189 );
nand \U$3628 ( \3875 , \3870 , \3874 );
not \U$3629 ( \3876 , \3875 );
not \U$3630 ( \3877 , \3588 );
not \U$3631 ( \3878 , \361 );
or \U$3632 ( \3879 , \3877 , \3878 );
xor \U$3633 ( \3880 , RIbe27c10_3, RIbe29128_48);
nand \U$3634 ( \3881 , \1173 , \3880 );
nand \U$3635 ( \3882 , \3879 , \3881 );
and \U$3636 ( \3883 , RIbe28d68_40, RIbe27b98_2);
nor \U$3637 ( \3884 , \3882 , \3883 );
not \U$3638 ( \3885 , \3884 );
nand \U$3639 ( \3886 , \3882 , \3883 );
nand \U$3640 ( \3887 , \3885 , \3886 );
not \U$3641 ( \3888 , \2891 );
not \U$3642 ( \3889 , \3506 );
and \U$3643 ( \3890 , \3888 , \3889 );
and \U$3644 ( \3891 , \2758 , RIbe285e8_24);
nor \U$3645 ( \3892 , \3890 , \3891 );
xnor \U$3646 ( \3893 , \3887 , \3892 );
not \U$3647 ( \3894 , \3893 );
or \U$3648 ( \3895 , \3876 , \3894 );
or \U$3649 ( \3896 , \3893 , \3875 );
nand \U$3650 ( \3897 , \3895 , \3896 );
not \U$3651 ( \3898 , \3897 );
or \U$3652 ( \3899 , \3867 , \3898 );
or \U$3653 ( \3900 , \3897 , \3866 );
nand \U$3654 ( \3901 , \3899 , \3900 );
not \U$3655 ( \3902 , \3901 );
not \U$3656 ( \3903 , \3207 );
not \U$3657 ( \3904 , \3214 );
or \U$3658 ( \3905 , \3903 , \3904 );
or \U$3659 ( \3906 , \3206 , \3179 );
nand \U$3660 ( \3907 , \3905 , \3906 );
not \U$3661 ( \3908 , \3907 );
not \U$3662 ( \3909 , \3908 );
or \U$3663 ( \3910 , \3902 , \3909 );
not \U$3664 ( \3911 , \3901 );
nand \U$3665 ( \3912 , \3911 , \3907 );
nand \U$3666 ( \3913 , \3910 , \3912 );
not \U$3667 ( \3914 , \3810 );
not \U$3668 ( \3915 , \3914 );
not \U$3669 ( \3916 , \3808 );
or \U$3670 ( \3917 , \3915 , \3916 );
nand \U$3671 ( \3918 , \3802 , \3800 );
nand \U$3672 ( \3919 , \3917 , \3918 );
and \U$3673 ( \3920 , \3913 , \3919 );
not \U$3674 ( \3921 , \3913 );
not \U$3675 ( \3922 , \3919 );
and \U$3676 ( \3923 , \3921 , \3922 );
nor \U$3677 ( \3924 , \3920 , \3923 );
not \U$3678 ( \3925 , \3924 );
not \U$3679 ( \3926 , \3925 );
or \U$3680 ( \3927 , \3838 , \3926 );
not \U$3681 ( \3928 , \3837 );
nand \U$3682 ( \3929 , \3928 , \3924 );
nand \U$3683 ( \3930 , \3927 , \3929 );
not \U$3684 ( \3931 , \3930 );
or \U$3685 ( \3932 , \3831 , \3931 );
or \U$3686 ( \3933 , \3930 , \3830 );
nand \U$3687 ( \3934 , \3932 , \3933 );
not \U$3688 ( \3935 , \3934 );
or \U$3689 ( \3936 , \3792 , \3935 );
or \U$3690 ( \3937 , \3791 , \3934 );
nand \U$3691 ( \3938 , \3936 , \3937 );
xor \U$3692 ( \3939 , \3470 , \3938 );
not \U$3693 ( \3940 , \3466 );
not \U$3694 ( \3941 , \3017 );
and \U$3695 ( \3942 , \3940 , \3941 );
and \U$3696 ( \3943 , \3466 , \3017 );
nor \U$3697 ( \3944 , \3942 , \3943 );
not \U$3698 ( \3945 , \3944 );
not \U$3699 ( \3946 , \3945 );
xor \U$3700 ( \3947 , \3424 , \3321 );
not \U$3701 ( \3948 , \3947 );
not \U$3702 ( \3949 , \1793 );
not \U$3703 ( \3950 , \3949 );
not \U$3704 ( \3951 , RIbe294e8_56);
not \U$3705 ( \3952 , RIbe28930_31);
or \U$3706 ( \3953 , \3951 , \3952 );
or \U$3707 ( \3954 , RIbe28930_31, RIbe294e8_56);
nand \U$3708 ( \3955 , \3953 , \3954 );
not \U$3709 ( \3956 , \3955 );
and \U$3710 ( \3957 , \3950 , \3956 );
and \U$3711 ( \3958 , \971 , \2534 );
nor \U$3712 ( \3959 , \3957 , \3958 );
not \U$3713 ( \3960 , \3402 );
not \U$3714 ( \3961 , \3960 );
not \U$3715 ( \3962 , RIbe28b88_36);
not \U$3716 ( \3963 , RIbe293f8_54);
and \U$3717 ( \3964 , \3962 , \3963 );
and \U$3718 ( \3965 , RIbe28b88_36, RIbe293f8_54);
nor \U$3719 ( \3966 , \3964 , \3965 );
not \U$3720 ( \3967 , \3966 );
not \U$3721 ( \3968 , \3967 );
and \U$3722 ( \3969 , \3961 , \3968 );
not \U$3723 ( \3970 , RIbe28b88_36);
or \U$3724 ( \3971 , \3970 , RIbe29308_52);
or \U$3725 ( \3972 , \3840 , RIbe28b88_36);
nand \U$3726 ( \3973 , \3971 , \3972 );
and \U$3727 ( \3974 , \2560 , \3973 );
nor \U$3728 ( \3975 , \3969 , \3974 );
xor \U$3729 ( \3976 , \3959 , \3975 );
not \U$3730 ( \3977 , \3976 );
xnor \U$3731 ( \3978 , RIbe290b0_47, RIbe29218_50);
or \U$3732 ( \3979 , \467 , \3978 );
not \U$3733 ( \3980 , \399 );
or \U$3734 ( \3981 , \3980 , \3361 );
nand \U$3735 ( \3982 , \3979 , \3981 );
not \U$3736 ( \3983 , \3982 );
xor \U$3737 ( \3984 , RIbe27b98_2, RIbe29b78_70);
not \U$3738 ( \3985 , \3984 );
not \U$3739 ( \3986 , \1295 );
or \U$3740 ( \3987 , \3985 , \3986 );
nand \U$3741 ( \3988 , \1734 , \3304 );
nand \U$3742 ( \3989 , \3987 , \3988 );
xor \U$3743 ( \3990 , RIbe28de0_41, RIbe28cf0_39);
and \U$3744 ( \3991 , \1284 , \3990 );
and \U$3745 ( \3992 , \514 , \3333 );
nor \U$3746 ( \3993 , \3991 , \3992 );
not \U$3747 ( \3994 , \3993 );
and \U$3748 ( \3995 , \3989 , \3994 );
not \U$3749 ( \3996 , \3989 );
and \U$3750 ( \3997 , \3996 , \3993 );
nor \U$3751 ( \3998 , \3995 , \3997 );
not \U$3752 ( \3999 , \3998 );
or \U$3753 ( \4000 , \3983 , \3999 );
nand \U$3754 ( \4001 , \3989 , \3994 );
nand \U$3755 ( \4002 , \4000 , \4001 );
not \U$3756 ( \4003 , \4002 );
or \U$3757 ( \4004 , \3977 , \4003 );
not \U$3758 ( \4005 , \3959 );
not \U$3759 ( \4006 , \3975 );
nand \U$3760 ( \4007 , \4005 , \4006 );
nand \U$3761 ( \4008 , \4004 , \4007 );
not \U$3762 ( \4009 , RIbe28930_31);
not \U$3763 ( \4010 , RIbe29470_55);
and \U$3764 ( \4011 , \4009 , \4010 );
and \U$3765 ( \4012 , RIbe28930_31, RIbe29470_55);
nor \U$3766 ( \4013 , \4011 , \4012 );
not \U$3767 ( \4014 , \4013 );
or \U$3768 ( \4015 , \967 , \4014 );
not \U$3769 ( \4016 , \1797 );
or \U$3770 ( \4017 , \4016 , \3955 );
nand \U$3771 ( \4018 , \4015 , \4017 );
not \U$3772 ( \4019 , \4018 );
and \U$3773 ( \4020 , RIbe28390_19, RIbe28c00_37);
not \U$3774 ( \4021 , RIbe28390_19);
and \U$3775 ( \4022 , \4021 , \2479 );
nor \U$3776 ( \4023 , \4020 , \4022 );
not \U$3777 ( \4024 , \4023 );
not \U$3778 ( \4025 , \2640 );
or \U$3779 ( \4026 , \4024 , \4025 );
not \U$3780 ( \4027 , \3410 );
nand \U$3781 ( \4028 , \4027 , \2777 );
nand \U$3782 ( \4029 , \4026 , \4028 );
not \U$3783 ( \4030 , \4029 );
not \U$3784 ( \4031 , \2718 );
and \U$3785 ( \4032 , RIbe27fd0_11, \317 );
not \U$3786 ( \4033 , RIbe27fd0_11);
and \U$3787 ( \4034 , \4033 , RIbe27ee0_9);
nor \U$3788 ( \4035 , \4032 , \4034 );
not \U$3789 ( \4036 , \4035 );
and \U$3790 ( \4037 , \4031 , \4036 );
and \U$3791 ( \4038 , \2707 , \3375 );
nor \U$3792 ( \4039 , \4037 , \4038 );
not \U$3793 ( \4040 , \4039 );
or \U$3794 ( \4041 , \4030 , \4040 );
or \U$3795 ( \4042 , \4029 , \4039 );
nand \U$3796 ( \4043 , \4041 , \4042 );
not \U$3797 ( \4044 , \4043 );
or \U$3798 ( \4045 , \4019 , \4044 );
not \U$3799 ( \4046 , \4039 );
nand \U$3800 ( \4047 , \4046 , \4029 );
nand \U$3801 ( \4048 , \4045 , \4047 );
xor \U$3802 ( \4049 , RIbe285e8_24, RIbe28750_27);
not \U$3803 ( \4050 , \4049 );
not \U$3804 ( \4051 , \2618 );
or \U$3805 ( \4052 , \4050 , \4051 );
nand \U$3806 ( \4053 , \2758 , \3261 );
nand \U$3807 ( \4054 , \4052 , \4053 );
not \U$3808 ( \4055 , \4054 );
not \U$3809 ( \4056 , RIbe27c88_4);
not \U$3810 ( \4057 , RIbe27d78_6);
and \U$3811 ( \4058 , \4056 , \4057 );
and \U$3812 ( \4059 , RIbe27c88_4, RIbe27d78_6);
nor \U$3813 ( \4060 , \4058 , \4059 );
not \U$3814 ( \4061 , \4060 );
not \U$3815 ( \4062 , \1164 );
or \U$3816 ( \4063 , \4061 , \4062 );
nand \U$3817 ( \4064 , \315 , \3294 );
nand \U$3818 ( \4065 , \4063 , \4064 );
not \U$3819 ( \4066 , \4065 );
or \U$3820 ( \4067 , \4055 , \4066 );
or \U$3821 ( \4068 , \4065 , \4054 );
xor \U$3822 ( \4069 , RIbe28318_18, RIbe28480_21);
not \U$3823 ( \4070 , \4069 );
not \U$3824 ( \4071 , \2519 );
or \U$3825 ( \4072 , \4070 , \4071 );
not \U$3826 ( \4073 , \3346 );
nand \U$3827 ( \4074 , \4073 , \2527 );
nand \U$3828 ( \4075 , \4072 , \4074 );
nand \U$3829 ( \4076 , \4068 , \4075 );
nand \U$3830 ( \4077 , \4067 , \4076 );
or \U$3831 ( \4078 , \4048 , \4077 );
not \U$3832 ( \4079 , \360 );
not \U$3833 ( \4080 , RIbe29998_66);
not \U$3834 ( \4081 , RIbe27c10_3);
or \U$3835 ( \4082 , \4080 , \4081 );
or \U$3836 ( \4083 , RIbe27c10_3, RIbe29998_66);
nand \U$3837 ( \4084 , \4082 , \4083 );
not \U$3838 ( \4085 , \4084 );
and \U$3839 ( \4086 , \4079 , \4085 );
and \U$3840 ( \4087 , \1174 , \3393 );
nor \U$3841 ( \4088 , \4086 , \4087 );
xor \U$3842 ( \4089 , RIbe27e68_8, RIbe28570_23);
not \U$3843 ( \4090 , \4089 );
not \U$3844 ( \4091 , \2459 );
or \U$3845 ( \4092 , \4090 , \4091 );
not \U$3846 ( \4093 , \3312 );
nand \U$3847 ( \4094 , \4093 , \2464 );
nand \U$3848 ( \4095 , \4092 , \4094 );
and \U$3849 ( \4096 , RIbe28138_14, RIbe28228_16);
nor \U$3850 ( \4097 , RIbe28138_14, RIbe28228_16);
nor \U$3851 ( \4098 , \4096 , \4097 );
not \U$3852 ( \4099 , \4098 );
not \U$3853 ( \4100 , \3056 );
or \U$3854 ( \4101 , \4099 , \4100 );
nand \U$3855 ( \4102 , \885 , \3272 );
nand \U$3856 ( \4103 , \4101 , \4102 );
nor \U$3857 ( \4104 , \4095 , \4103 );
or \U$3858 ( \4105 , \4088 , \4104 );
nand \U$3859 ( \4106 , \4095 , \4103 );
nand \U$3860 ( \4107 , \4105 , \4106 );
nand \U$3861 ( \4108 , \4078 , \4107 );
nand \U$3862 ( \4109 , \4048 , \4077 );
nand \U$3863 ( \4110 , \4108 , \4109 );
xor \U$3864 ( \4111 , \4008 , \4110 );
not \U$3865 ( \4112 , \4111 );
not \U$3866 ( \4113 , \3317 );
not \U$3867 ( \4114 , \3319 );
or \U$3868 ( \4115 , \4113 , \4114 );
or \U$3869 ( \4116 , \3319 , \3317 );
nand \U$3870 ( \4117 , \4115 , \4116 );
not \U$3871 ( \4118 , \4117 );
or \U$3872 ( \4119 , \4112 , \4118 );
nand \U$3873 ( \4120 , \4110 , \4008 );
nand \U$3874 ( \4121 , \4119 , \4120 );
not \U$3875 ( \4122 , \4121 );
xor \U$3876 ( \4123 , \3387 , \3354 );
xnor \U$3877 ( \4124 , \4123 , \3418 );
not \U$3878 ( \4125 , \3384 );
nand \U$3879 ( \4126 , \4125 , \3386 );
not \U$3880 ( \4127 , \4126 );
not \U$3881 ( \4128 , \3365 );
and \U$3882 ( \4129 , \4127 , \4128 );
and \U$3883 ( \4130 , \4126 , \3365 );
nor \U$3884 ( \4131 , \4129 , \4130 );
xor \U$3885 ( \4132 , RIbe291a0_49, RIbe296c8_60);
not \U$3886 ( \4133 , \4132 );
not \U$3887 ( \4134 , \1130 );
or \U$3888 ( \4135 , \4133 , \4134 );
not \U$3889 ( \4136 , \3285 );
nand \U$3890 ( \4137 , \4136 , \908 );
nand \U$3891 ( \4138 , \4135 , \4137 );
not \U$3892 ( \4139 , \3278 );
not \U$3893 ( \4140 , \287 );
or \U$3894 ( \4141 , \4139 , \4140 );
not \U$3895 ( \4142 , RIbe29038_46);
not \U$3896 ( \4143 , RIbe29b00_69);
and \U$3897 ( \4144 , \4142 , \4143 );
and \U$3898 ( \4145 , RIbe29038_46, RIbe29b00_69);
nor \U$3899 ( \4146 , \4144 , \4145 );
nand \U$3900 ( \4147 , \979 , \4146 );
nand \U$3901 ( \4148 , \4141 , \4147 );
xor \U$3902 ( \4149 , \4138 , \4148 );
and \U$3903 ( \4150 , RIbe28a20_33, RIbe288b8_30);
not \U$3904 ( \4151 , RIbe28a20_33);
and \U$3905 ( \4152 , \4151 , \931 );
nor \U$3906 ( \4153 , \4150 , \4152 );
not \U$3907 ( \4154 , \4153 );
not \U$3908 ( \4155 , \1781 );
or \U$3909 ( \4156 , \4154 , \4155 );
not \U$3910 ( \4157 , \3369 );
or \U$3911 ( \4158 , \1770 , \4157 );
nand \U$3912 ( \4159 , \4156 , \4158 );
and \U$3913 ( \4160 , \4149 , \4159 );
and \U$3914 ( \4161 , \4138 , \4148 );
or \U$3915 ( \4162 , \4160 , \4161 );
or \U$3916 ( \4163 , \4131 , \4162 );
not \U$3917 ( \4164 , \1325 );
not \U$3918 ( \4165 , RIbe29740_61);
not \U$3919 ( \4166 , RIbe280c0_13);
or \U$3920 ( \4167 , \4165 , \4166 );
or \U$3921 ( \4168 , RIbe280c0_13, RIbe29740_61);
nand \U$3922 ( \4169 , \4167 , \4168 );
not \U$3923 ( \4170 , \4169 );
and \U$3924 ( \4171 , \4164 , \4170 );
and \U$3925 ( \4172 , \869 , \3239 );
nor \U$3926 ( \4173 , \4171 , \4172 );
not \U$3927 ( \4174 , \4173 );
not \U$3928 ( \4175 , \4174 );
not \U$3929 ( \4176 , \3255 );
xnor \U$3930 ( \4177 , RIbe29380_53, RIbe28f48_44);
not \U$3931 ( \4178 , \4177 );
and \U$3932 ( \4179 , \4176 , \4178 );
buf \U$3933 ( \4180 , \3248 );
buf \U$3934 ( \4181 , \4180 );
and \U$3935 ( \4182 , \4181 , RIbe28f48_44);
nor \U$3936 ( \4183 , \4179 , \4182 );
nand \U$3937 ( \4184 , RIbe27b98_2, RIbe29ce0_73);
and \U$3938 ( \4185 , \4183 , \4184 );
not \U$3939 ( \4186 , \4183 );
not \U$3940 ( \4187 , \4184 );
and \U$3941 ( \4188 , \4186 , \4187 );
nor \U$3942 ( \4189 , \4185 , \4188 );
not \U$3943 ( \4190 , \4189 );
or \U$3944 ( \4191 , \4175 , \4190 );
not \U$3945 ( \4192 , \4183 );
nand \U$3946 ( \4193 , \4192 , \4187 );
nand \U$3947 ( \4194 , \4191 , \4193 );
not \U$3948 ( \4195 , \4194 );
nand \U$3949 ( \4196 , \4131 , \4162 );
nand \U$3950 ( \4197 , \4195 , \4196 );
nand \U$3951 ( \4198 , \4163 , \4197 );
nand \U$3952 ( \4199 , \4124 , \4198 );
xor \U$3953 ( \4200 , \3299 , \3306 );
xor \U$3954 ( \4201 , \4200 , \3314 );
not \U$3955 ( \4202 , \4201 );
not \U$3956 ( \4203 , \3349 );
and \U$3957 ( \4204 , \3342 , \4203 );
not \U$3958 ( \4205 , \3342 );
and \U$3959 ( \4206 , \4205 , \3349 );
nor \U$3960 ( \4207 , \4204 , \4206 );
xor \U$3961 ( \4208 , \3398 , \3406 );
xor \U$3962 ( \4209 , \4208 , \3415 );
xnor \U$3963 ( \4210 , \4207 , \4209 );
not \U$3964 ( \4211 , \4210 );
or \U$3965 ( \4212 , \4202 , \4211 );
not \U$3966 ( \4213 , \4207 );
nand \U$3967 ( \4214 , \4213 , \4209 );
nand \U$3968 ( \4215 , \4212 , \4214 );
and \U$3969 ( \4216 , \4199 , \4215 );
nor \U$3970 ( \4217 , \4124 , \4198 );
nor \U$3971 ( \4218 , \4216 , \4217 );
not \U$3972 ( \4219 , \4218 );
or \U$3973 ( \4220 , \4122 , \4219 );
or \U$3974 ( \4221 , \4218 , \4121 );
nand \U$3975 ( \4222 , \4220 , \4221 );
not \U$3976 ( \4223 , \4222 );
or \U$3977 ( \4224 , \3948 , \4223 );
not \U$3978 ( \4225 , \4218 );
nand \U$3979 ( \4226 , \4225 , \4121 );
nand \U$3980 ( \4227 , \4224 , \4226 );
not \U$3981 ( \4228 , \4227 );
not \U$3982 ( \4229 , \3459 );
not \U$3983 ( \4230 , \3457 );
and \U$3984 ( \4231 , \4229 , \4230 );
and \U$3985 ( \4232 , \3459 , \3457 );
nor \U$3986 ( \4233 , \4231 , \4232 );
not \U$3987 ( \4234 , \4233 );
or \U$3988 ( \4235 , \4228 , \4234 );
or \U$3989 ( \4236 , \4233 , \4227 );
nand \U$3990 ( \4237 , \4235 , \4236 );
xor \U$3991 ( \4238 , \2795 , \2507 );
not \U$3992 ( \4239 , \4238 );
and \U$3993 ( \4240 , \3959 , \3975 );
not \U$3994 ( \4241 , \3959 );
and \U$3995 ( \4242 , \4241 , \4006 );
nor \U$3996 ( \4243 , \4240 , \4242 );
xor \U$3997 ( \4244 , \4002 , \4243 );
xor \U$3998 ( \4245 , \3277 , \3283 );
xor \U$3999 ( \4246 , \4245 , \3288 );
not \U$4000 ( \4247 , \3267 );
nand \U$4001 ( \4248 , \4247 , \3269 );
not \U$4002 ( \4249 , \4248 );
not \U$4003 ( \4250 , \3245 );
and \U$4004 ( \4251 , \4249 , \4250 );
and \U$4005 ( \4252 , \4248 , \3245 );
nor \U$4006 ( \4253 , \4251 , \4252 );
not \U$4007 ( \4254 , \4253 );
and \U$4008 ( \4255 , \4246 , \4254 );
not \U$4009 ( \4256 , \4246 );
and \U$4010 ( \4257 , \4256 , \4253 );
nor \U$4011 ( \4258 , \4255 , \4257 );
and \U$4012 ( \4259 , \4244 , \4258 );
and \U$4013 ( \4260 , \4246 , \4254 );
nor \U$4014 ( \4261 , \4259 , \4260 );
not \U$4015 ( \4262 , \4261 );
not \U$4016 ( \4263 , \2573 );
not \U$4017 ( \4264 , \2660 );
or \U$4018 ( \4265 , \4263 , \4264 );
or \U$4019 ( \4266 , \2660 , \2573 );
nand \U$4020 ( \4267 , \4265 , \4266 );
xor \U$4021 ( \4268 , \3433 , \3437 );
xor \U$4022 ( \4269 , \4268 , \3443 );
nor \U$4023 ( \4270 , \4267 , \4269 );
not \U$4024 ( \4271 , \4270 );
and \U$4025 ( \4272 , \4262 , \4271 );
buf \U$4026 ( \4273 , \4269 );
and \U$4027 ( \4274 , \4267 , \4273 );
nor \U$4028 ( \4275 , \4272 , \4274 );
not \U$4029 ( \4276 , \4275 );
not \U$4030 ( \4277 , \3453 );
xor \U$4031 ( \4278 , \3446 , \3451 );
not \U$4032 ( \4279 , \4278 );
or \U$4033 ( \4280 , \4277 , \4279 );
or \U$4034 ( \4281 , \4278 , \3453 );
nand \U$4035 ( \4282 , \4280 , \4281 );
not \U$4036 ( \4283 , \4282 );
or \U$4037 ( \4284 , \4276 , \4283 );
or \U$4038 ( \4285 , \4275 , \4282 );
nand \U$4039 ( \4286 , \4284 , \4285 );
not \U$4040 ( \4287 , \4286 );
or \U$4041 ( \4288 , \4239 , \4287 );
not \U$4042 ( \4289 , \4275 );
nand \U$4043 ( \4290 , \4289 , \4282 );
nand \U$4044 ( \4291 , \4288 , \4290 );
nand \U$4045 ( \4292 , \4237 , \4291 );
not \U$4046 ( \4293 , \4233 );
nand \U$4047 ( \4294 , \4293 , \4227 );
and \U$4048 ( \4295 , \4292 , \4294 );
xor \U$4049 ( \4296 , \3824 , \3793 );
not \U$4050 ( \4297 , \4296 );
and \U$4051 ( \4298 , \4295 , \4297 );
not \U$4052 ( \4299 , \4295 );
and \U$4053 ( \4300 , \4299 , \4296 );
nor \U$4054 ( \4301 , \4298 , \4300 );
not \U$4055 ( \4302 , \4301 );
or \U$4056 ( \4303 , \3946 , \4302 );
not \U$4057 ( \4304 , \4295 );
nand \U$4058 ( \4305 , \4304 , \4296 );
nand \U$4059 ( \4306 , \4303 , \4305 );
nor \U$4060 ( \4307 , \3939 , \4306 );
not \U$4061 ( \4308 , \4307 );
not \U$4062 ( \4309 , \3944 );
not \U$4063 ( \4310 , \4301 );
or \U$4064 ( \4311 , \4309 , \4310 );
or \U$4065 ( \4312 , \4301 , \3944 );
nand \U$4066 ( \4313 , \4311 , \4312 );
not \U$4067 ( \4314 , \4313 );
not \U$4068 ( \4315 , \4261 );
xor \U$4069 ( \4316 , \4273 , \4267 );
not \U$4070 ( \4317 , \4316 );
or \U$4071 ( \4318 , \4315 , \4317 );
or \U$4072 ( \4319 , \4316 , \4261 );
nand \U$4073 ( \4320 , \4318 , \4319 );
not \U$4074 ( \4321 , \4320 );
xor \U$4075 ( \4322 , \4258 , \4244 );
not \U$4076 ( \4323 , \4322 );
not \U$4077 ( \4324 , \4201 );
and \U$4078 ( \4325 , \4210 , \4324 );
not \U$4079 ( \4326 , \4210 );
and \U$4080 ( \4327 , \4326 , \4201 );
nor \U$4081 ( \4328 , \4325 , \4327 );
not \U$4082 ( \4329 , \4328 );
xor \U$4083 ( \4330 , RIbe288b8_30, RIbe28b88_36);
not \U$4084 ( \4331 , \4330 );
not \U$4085 ( \4332 , \2702 );
or \U$4086 ( \4333 , \4331 , \4332 );
and \U$4087 ( \4334 , RIbe28a98_34, RIbe28b88_36);
nor \U$4088 ( \4335 , RIbe28a98_34, RIbe28b88_36);
nor \U$4089 ( \4336 , \4334 , \4335 );
nand \U$4090 ( \4337 , \2560 , \4336 );
nand \U$4091 ( \4338 , \4333 , \4337 );
not \U$4092 ( \4339 , \4338 );
not \U$4093 ( \4340 , \1614 );
xor \U$4094 ( \4341 , RIbe27d78_6, RIbe28d68_40);
not \U$4095 ( \4342 , \4341 );
not \U$4096 ( \4343 , \4342 );
and \U$4097 ( \4344 , \4340 , \4343 );
and \U$4098 ( \4345 , \315 , \4060 );
nor \U$4099 ( \4346 , \4344 , \4345 );
xor \U$4100 ( \4347 , \4339 , \4346 );
not \U$4101 ( \4348 , \1566 );
xor \U$4102 ( \4349 , RIbe27b98_2, RIbe29ce0_73);
and \U$4103 ( \4350 , \4348 , \4349 );
and \U$4104 ( \4351 , \1298 , \3984 );
nor \U$4105 ( \4352 , \4350 , \4351 );
and \U$4106 ( \4353 , \4347 , \4352 );
and \U$4107 ( \4354 , \4339 , \4346 );
or \U$4108 ( \4355 , \4353 , \4354 );
not \U$4109 ( \4356 , \4355 );
not \U$4110 ( \4357 , \4173 );
not \U$4111 ( \4358 , \4189 );
or \U$4112 ( \4359 , \4357 , \4358 );
or \U$4113 ( \4360 , \4189 , \4173 );
nand \U$4114 ( \4361 , \4359 , \4360 );
not \U$4115 ( \4362 , \4361 );
or \U$4116 ( \4363 , \4356 , \4362 );
or \U$4117 ( \4364 , \4361 , \4355 );
nand \U$4118 ( \4365 , \4363 , \4364 );
not \U$4119 ( \4366 , \4365 );
not \U$4120 ( \4367 , \2718 );
not \U$4121 ( \4368 , RIbe27fd0_11);
not \U$4122 ( \4369 , RIbe28570_23);
and \U$4123 ( \4370 , \4368 , \4369 );
and \U$4124 ( \4371 , RIbe27fd0_11, RIbe28570_23);
nor \U$4125 ( \4372 , \4370 , \4371 );
not \U$4126 ( \4373 , \4372 );
not \U$4127 ( \4374 , \4373 );
and \U$4128 ( \4375 , \4367 , \4374 );
xnor \U$4129 ( \4376 , RIbe27fd0_11, RIbe286d8_26);
not \U$4130 ( \4377 , \4376 );
and \U$4131 ( \4378 , \2707 , \4377 );
nor \U$4132 ( \4379 , \4375 , \4378 );
not \U$4133 ( \4380 , RIbe27ee0_9);
not \U$4134 ( \4381 , RIbe28f48_44);
and \U$4135 ( \4382 , \4380 , \4381 );
and \U$4136 ( \4383 , RIbe27ee0_9, RIbe28f48_44);
nor \U$4137 ( \4384 , \4382 , \4383 );
and \U$4138 ( \4385 , \3256 , \4384 );
and \U$4139 ( \4386 , RIbe28f48_44, RIbe28048_12);
not \U$4140 ( \4387 , RIbe28f48_44);
and \U$4141 ( \4388 , \4387 , \431 );
nor \U$4142 ( \4389 , \4386 , \4388 );
and \U$4143 ( \4390 , \4181 , \4389 );
nor \U$4144 ( \4391 , \4385 , \4390 );
xor \U$4145 ( \4392 , \4379 , \4391 );
xor \U$4146 ( \4393 , RIbe29038_46, RIbe29218_50);
and \U$4147 ( \4394 , \282 , \4393 );
not \U$4148 ( \4395 , RIbe29038_46);
not \U$4149 ( \4396 , RIbe29a10_67);
and \U$4150 ( \4397 , \4395 , \4396 );
and \U$4151 ( \4398 , RIbe29038_46, RIbe29a10_67);
nor \U$4152 ( \4399 , \4397 , \4398 );
and \U$4153 ( \4400 , \1805 , \4399 );
nor \U$4154 ( \4401 , \4394 , \4400 );
and \U$4155 ( \4402 , \4392 , \4401 );
and \U$4156 ( \4403 , \4379 , \4391 );
or \U$4157 ( \4404 , \4402 , \4403 );
not \U$4158 ( \4405 , \4404 );
not \U$4159 ( \4406 , \4405 );
xor \U$4160 ( \4407 , RIbe28de0_41, RIbe29b78_70);
and \U$4161 ( \4408 , \332 , \4407 );
xor \U$4162 ( \4409 , RIbe28de0_41, RIbe27b20_1);
and \U$4163 ( \4410 , \514 , \4409 );
nor \U$4164 ( \4411 , \4408 , \4410 );
not \U$4165 ( \4412 , \4411 );
not \U$4166 ( \4413 , \4412 );
xor \U$4167 ( \4414 , RIbe29d58_74, RIbe27b98_2);
not \U$4168 ( \4415 , \4414 );
not \U$4169 ( \4416 , \258 );
or \U$4170 ( \4417 , \4415 , \4416 );
nand \U$4171 ( \4418 , \269 , \4349 );
nand \U$4172 ( \4419 , \4417 , \4418 );
xnor \U$4173 ( \4420 , RIbe28c00_37, RIbe28480_21);
or \U$4174 ( \4421 , \3484 , \4420 );
xnor \U$4175 ( \4422 , RIbe28c78_38, RIbe28480_21);
or \U$4176 ( \4423 , \2672 , \4422 );
nand \U$4177 ( \4424 , \4421 , \4423 );
xor \U$4178 ( \4425 , \4419 , \4424 );
not \U$4179 ( \4426 , \4425 );
or \U$4180 ( \4427 , \4413 , \4426 );
nand \U$4181 ( \4428 , \4419 , \4424 );
nand \U$4182 ( \4429 , \4427 , \4428 );
xor \U$4183 ( \4430 , RIbe28228_16, RIbe29740_61);
not \U$4184 ( \4431 , \4430 );
not \U$4185 ( \4432 , \1061 );
or \U$4186 ( \4433 , \4431 , \4432 );
and \U$4187 ( \4434 , RIbe28228_16, RIbe297b8_62);
nor \U$4188 ( \4435 , RIbe28228_16, RIbe297b8_62);
nor \U$4189 ( \4436 , \4434 , \4435 );
nand \U$4190 ( \4437 , \885 , \4436 );
nand \U$4191 ( \4438 , \4433 , \4437 );
not \U$4192 ( \4439 , \4438 );
xor \U$4193 ( \4440 , RIbe28750_27, RIbe27e68_8);
not \U$4194 ( \4441 , \4440 );
not \U$4195 ( \4442 , \2457 );
not \U$4196 ( \4443 , \4442 );
not \U$4197 ( \4444 , \4443 );
or \U$4198 ( \4445 , \4441 , \4444 );
not \U$4199 ( \4446 , \2464 );
not \U$4200 ( \4447 , \4446 );
xor \U$4201 ( \4448 , RIbe28840_29, RIbe27e68_8);
nand \U$4202 ( \4449 , \4447 , \4448 );
nand \U$4203 ( \4450 , \4445 , \4449 );
not \U$4204 ( \4451 , \4450 );
or \U$4205 ( \4452 , \4439 , \4451 );
or \U$4206 ( \4453 , \4450 , \4438 );
xor \U$4207 ( \4454 , RIbe29b00_69, RIbe296c8_60);
not \U$4208 ( \4455 , \4454 );
not \U$4209 ( \4456 , \1452 );
or \U$4210 ( \4457 , \4455 , \4456 );
xor \U$4211 ( \4458 , RIbe29128_48, RIbe296c8_60);
nand \U$4212 ( \4459 , \1137 , \4458 );
nand \U$4213 ( \4460 , \4457 , \4459 );
nand \U$4214 ( \4461 , \4453 , \4460 );
nand \U$4215 ( \4462 , \4452 , \4461 );
xor \U$4216 ( \4463 , \4429 , \4462 );
not \U$4217 ( \4464 , \4463 );
or \U$4218 ( \4465 , \4406 , \4464 );
nand \U$4219 ( \4466 , \4429 , \4462 );
nand \U$4220 ( \4467 , \4465 , \4466 );
not \U$4221 ( \4468 , \4467 );
or \U$4222 ( \4469 , \4366 , \4468 );
not \U$4223 ( \4470 , \4355 );
nand \U$4224 ( \4471 , \4470 , \4361 );
nand \U$4225 ( \4472 , \4469 , \4471 );
not \U$4226 ( \4473 , \4472 );
or \U$4227 ( \4474 , \4329 , \4473 );
or \U$4228 ( \4475 , \4472 , \4328 );
nand \U$4229 ( \4476 , \4474 , \4475 );
not \U$4230 ( \4477 , \4476 );
or \U$4231 ( \4478 , \4323 , \4477 );
not \U$4232 ( \4479 , \4328 );
nand \U$4233 ( \4480 , \4479 , \4472 );
nand \U$4234 ( \4481 , \4478 , \4480 );
not \U$4235 ( \4482 , \4124 );
not \U$4236 ( \4483 , \4215 );
or \U$4237 ( \4484 , \4482 , \4483 );
or \U$4238 ( \4485 , \4215 , \4124 );
nand \U$4239 ( \4486 , \4484 , \4485 );
not \U$4240 ( \4487 , \4486 );
not \U$4241 ( \4488 , \4198 );
and \U$4242 ( \4489 , \4487 , \4488 );
and \U$4243 ( \4490 , \4486 , \4198 );
nor \U$4244 ( \4491 , \4489 , \4490 );
not \U$4245 ( \4492 , \4491 );
and \U$4246 ( \4493 , \4481 , \4492 );
not \U$4247 ( \4494 , \4481 );
and \U$4248 ( \4495 , \4494 , \4491 );
nor \U$4249 ( \4496 , \4493 , \4495 );
not \U$4250 ( \4497 , \4496 );
or \U$4251 ( \4498 , \4321 , \4497 );
nand \U$4252 ( \4499 , \4481 , \4492 );
nand \U$4253 ( \4500 , \4498 , \4499 );
not \U$4254 ( \4501 , \4500 );
xnor \U$4255 ( \4502 , \4222 , \3947 );
xnor \U$4256 ( \4503 , \4111 , \4117 );
not \U$4257 ( \4504 , \4503 );
not \U$4258 ( \4505 , \4504 );
xor \U$4259 ( \4506 , \4077 , \4107 );
xnor \U$4260 ( \4507 , \4506 , \4048 );
not \U$4261 ( \4508 , \4018 );
and \U$4262 ( \4509 , \4043 , \4508 );
not \U$4263 ( \4510 , \4043 );
and \U$4264 ( \4511 , \4510 , \4018 );
nor \U$4265 ( \4512 , \4509 , \4511 );
not \U$4266 ( \4513 , \4106 );
nor \U$4267 ( \4514 , \4513 , \4104 );
xor \U$4268 ( \4515 , \4514 , \4088 );
xor \U$4269 ( \4516 , \4512 , \4515 );
xnor \U$4270 ( \4517 , \3998 , \3982 );
and \U$4271 ( \4518 , \4516 , \4517 );
and \U$4272 ( \4519 , \4512 , \4515 );
or \U$4273 ( \4520 , \4518 , \4519 );
xor \U$4274 ( \4521 , \4507 , \4520 );
xor \U$4275 ( \4522 , \4138 , \4148 );
xor \U$4276 ( \4523 , \4522 , \4159 );
xor \U$4277 ( \4524 , \4065 , \4054 );
xor \U$4278 ( \4525 , \4524 , \4075 );
xor \U$4279 ( \4526 , \4523 , \4525 );
not \U$4280 ( \4527 , \1494 );
xnor \U$4281 ( \4528 , RIbe298a8_64, RIbe27c10_3);
not \U$4282 ( \4529 , \4528 );
and \U$4283 ( \4530 , \4527 , \4529 );
not \U$4284 ( \4531 , \1498 );
nor \U$4285 ( \4532 , \4531 , \4084 );
nor \U$4286 ( \4533 , \4530 , \4532 );
not \U$4287 ( \4534 , \524 );
xnor \U$4288 ( \4535 , RIbe27df0_7, RIbe290b0_47);
not \U$4289 ( \4536 , \4535 );
and \U$4290 ( \4537 , \4534 , \4536 );
nor \U$4291 ( \4538 , \468 , \3978 );
nor \U$4292 ( \4539 , \4537 , \4538 );
xor \U$4293 ( \4540 , \4533 , \4539 );
not \U$4294 ( \4541 , \3402 );
not \U$4295 ( \4542 , \4541 );
not \U$4296 ( \4543 , \4336 );
not \U$4297 ( \4544 , \4543 );
and \U$4298 ( \4545 , \4542 , \4544 );
and \U$4299 ( \4546 , \3594 , \3966 );
nor \U$4300 ( \4547 , \4545 , \4546 );
and \U$4301 ( \4548 , \4540 , \4547 );
and \U$4302 ( \4549 , \4533 , \4539 );
or \U$4303 ( \4550 , \4548 , \4549 );
not \U$4304 ( \4551 , \4550 );
and \U$4305 ( \4552 , \4526 , \4551 );
and \U$4306 ( \4553 , \4523 , \4525 );
or \U$4307 ( \4554 , \4552 , \4553 );
not \U$4308 ( \4555 , \4554 );
and \U$4309 ( \4556 , \4521 , \4555 );
and \U$4310 ( \4557 , \4507 , \4520 );
or \U$4311 ( \4558 , \4556 , \4557 );
not \U$4312 ( \4559 , \4558 );
not \U$4313 ( \4560 , \4559 );
and \U$4314 ( \4561 , \1061 , \4436 );
and \U$4315 ( \4562 , \885 , \4098 );
nor \U$4316 ( \4563 , \4561 , \4562 );
not \U$4317 ( \4564 , \4563 );
not \U$4318 ( \4565 , \4564 );
not \U$4319 ( \4566 , \4448 );
not \U$4320 ( \4567 , \2600 );
or \U$4321 ( \4568 , \4566 , \4567 );
nand \U$4322 ( \4569 , \2603 , \4089 );
nand \U$4323 ( \4570 , \4568 , \4569 );
not \U$4324 ( \4571 , \4570 );
xor \U$4325 ( \4572 , RIbe29dd0_75, RIbe29e48_76);
not \U$4326 ( \4573 , \4572 );
xor \U$4327 ( \4574 , RIbe29c68_72, RIbe29dd0_75);
nand \U$4328 ( \4575 , \4573 , \4574 );
buf \U$4329 ( \4576 , \4575 );
buf \U$4330 ( \4577 , \4576 );
not \U$4331 ( \4578 , \4577 );
not \U$4332 ( \4579 , \4578 );
buf \U$4333 ( \4580 , \4572 );
not \U$4334 ( \4581 , \4580 );
nand \U$4335 ( \4582 , \4579 , \4581 );
and \U$4336 ( \4583 , \4582 , RIbe29c68_72);
not \U$4337 ( \4584 , \4583 );
or \U$4338 ( \4585 , \4571 , \4584 );
or \U$4339 ( \4586 , \4583 , \4570 );
nand \U$4340 ( \4587 , \4585 , \4586 );
not \U$4341 ( \4588 , \4587 );
or \U$4342 ( \4589 , \4565 , \4588 );
not \U$4343 ( \4590 , \4583 );
nand \U$4344 ( \4591 , \4590 , \4570 );
nand \U$4345 ( \4592 , \4589 , \4591 );
not \U$4346 ( \4593 , RIbe28390_19);
not \U$4347 ( \4594 , RIbe29308_52);
and \U$4348 ( \4595 , \4593 , \4594 );
and \U$4349 ( \4596 , RIbe28390_19, RIbe29308_52);
nor \U$4350 ( \4597 , \4595 , \4596 );
not \U$4351 ( \4598 , \4597 );
not \U$4352 ( \4599 , \2640 );
or \U$4353 ( \4600 , \4598 , \4599 );
nand \U$4354 ( \4601 , \2777 , \4023 );
nand \U$4355 ( \4602 , \4600 , \4601 );
not \U$4356 ( \4603 , \2626 );
not \U$4357 ( \4604 , \4049 );
or \U$4358 ( \4605 , \4603 , \4604 );
xnor \U$4359 ( \4606 , RIbe285e8_24, RIbe284f8_22);
or \U$4360 ( \4607 , \3498 , \4606 );
nand \U$4361 ( \4608 , \4605 , \4607 );
nor \U$4362 ( \4609 , \4602 , \4608 );
not \U$4363 ( \4610 , \1325 );
xnor \U$4364 ( \4611 , RIbe280c0_13, RIbe295d8_58);
not \U$4365 ( \4612 , \4611 );
and \U$4366 ( \4613 , \4610 , \4612 );
nor \U$4367 ( \4614 , \1573 , \4169 );
nor \U$4368 ( \4615 , \4613 , \4614 );
or \U$4369 ( \4616 , \4609 , \4615 );
nand \U$4370 ( \4617 , \4602 , \4608 );
nand \U$4371 ( \4618 , \4616 , \4617 );
not \U$4372 ( \4619 , \4618 );
not \U$4373 ( \4620 , \4389 );
not \U$4374 ( \4621 , \3256 );
or \U$4375 ( \4622 , \4620 , \4621 );
not \U$4376 ( \4623 , \4177 );
nand \U$4377 ( \4624 , \4623 , \3249 );
nand \U$4378 ( \4625 , \4622 , \4624 );
not \U$4379 ( \4626 , \4458 );
not \U$4380 ( \4627 , \2877 );
or \U$4381 ( \4628 , \4626 , \4627 );
nand \U$4382 ( \4629 , \1137 , \4132 );
nand \U$4383 ( \4630 , \4628 , \4629 );
or \U$4384 ( \4631 , \4625 , \4630 );
not \U$4385 ( \4632 , \4399 );
not \U$4386 ( \4633 , \282 );
or \U$4387 ( \4634 , \4632 , \4633 );
nand \U$4388 ( \4635 , \287 , \4146 );
nand \U$4389 ( \4636 , \4634 , \4635 );
nand \U$4390 ( \4637 , \4631 , \4636 );
nand \U$4391 ( \4638 , \4625 , \4630 );
and \U$4392 ( \4639 , \4637 , \4638 );
not \U$4393 ( \4640 , \4639 );
or \U$4394 ( \4641 , \4619 , \4640 );
or \U$4395 ( \4642 , \4618 , \4639 );
nand \U$4396 ( \4643 , \4641 , \4642 );
and \U$4397 ( \4644 , \4592 , \4643 );
not \U$4398 ( \4645 , \4618 );
nor \U$4399 ( \4646 , \4645 , \4639 );
nor \U$4400 ( \4647 , \4644 , \4646 );
not \U$4401 ( \4648 , \4647 );
nand \U$4402 ( \4649 , RIbe27b98_2, RIbe29d58_74);
not \U$4403 ( \4650 , \4409 );
not \U$4404 ( \4651 , \332 );
or \U$4405 ( \4652 , \4650 , \4651 );
nand \U$4406 ( \4653 , \347 , \3990 );
nand \U$4407 ( \4654 , \4652 , \4653 );
xnor \U$4408 ( \4655 , \4649 , \4654 );
not \U$4409 ( \4656 , \4655 );
not \U$4410 ( \4657 , \4069 );
not \U$4411 ( \4658 , \2527 );
or \U$4412 ( \4659 , \4657 , \4658 );
not \U$4413 ( \4660 , \4422 );
nand \U$4414 ( \4661 , \4660 , \2520 );
nand \U$4415 ( \4662 , \4659 , \4661 );
not \U$4416 ( \4663 , \4662 );
or \U$4417 ( \4664 , \4656 , \4663 );
not \U$4418 ( \4665 , \4649 );
nand \U$4419 ( \4666 , \4665 , \4654 );
nand \U$4420 ( \4667 , \4664 , \4666 );
and \U$4421 ( \4668 , \4667 , \4006 );
not \U$4422 ( \4669 , \4667 );
and \U$4423 ( \4670 , \4669 , \3975 );
or \U$4424 ( \4671 , \4668 , \4670 );
not \U$4425 ( \4672 , \4671 );
not \U$4426 ( \4673 , \2708 );
not \U$4427 ( \4674 , \4035 );
and \U$4428 ( \4675 , \4673 , \4674 );
not \U$4429 ( \4676 , \3378 );
nor \U$4430 ( \4677 , \4676 , \4376 );
nor \U$4431 ( \4678 , \4675 , \4677 );
not \U$4432 ( \4679 , \3750 );
xor \U$4433 ( \4680 , RIbe28a20_33, RIbe294e8_56);
not \U$4434 ( \4681 , \4680 );
not \U$4435 ( \4682 , \4681 );
and \U$4436 ( \4683 , \4679 , \4682 );
and \U$4437 ( \4684 , \1769 , \4153 );
nor \U$4438 ( \4685 , \4683 , \4684 );
xor \U$4439 ( \4686 , \4678 , \4685 );
and \U$4440 ( \4687 , RIbe28930_31, RIbe282a0_17);
not \U$4441 ( \4688 , RIbe28930_31);
and \U$4442 ( \4689 , \4688 , \951 );
nor \U$4443 ( \4690 , \4687 , \4689 );
and \U$4444 ( \4691 , \966 , \4690 );
and \U$4445 ( \4692 , \1199 , \4013 );
nor \U$4446 ( \4693 , \4691 , \4692 );
and \U$4447 ( \4694 , \4686 , \4693 );
and \U$4448 ( \4695 , \4678 , \4685 );
or \U$4449 ( \4696 , \4694 , \4695 );
not \U$4450 ( \4697 , \4696 );
not \U$4451 ( \4698 , \4697 );
or \U$4452 ( \4699 , \4672 , \4698 );
nand \U$4453 ( \4700 , \4667 , \3975 );
nand \U$4454 ( \4701 , \4699 , \4700 );
not \U$4455 ( \4702 , \4701 );
or \U$4456 ( \4703 , \4648 , \4702 );
or \U$4457 ( \4704 , \4701 , \4647 );
nand \U$4458 ( \4705 , \4703 , \4704 );
not \U$4459 ( \4706 , \4705 );
or \U$4460 ( \4707 , \4131 , \4162 );
nand \U$4461 ( \4708 , \4707 , \4196 );
xnor \U$4462 ( \4709 , \4708 , \4194 );
not \U$4463 ( \4710 , \4709 );
or \U$4464 ( \4711 , \4706 , \4710 );
not \U$4465 ( \4712 , \4647 );
nand \U$4466 ( \4713 , \4712 , \4701 );
nand \U$4467 ( \4714 , \4711 , \4713 );
not \U$4468 ( \4715 , \4714 );
not \U$4469 ( \4716 , \4715 );
or \U$4470 ( \4717 , \4560 , \4716 );
nand \U$4471 ( \4718 , \4558 , \4714 );
nand \U$4472 ( \4719 , \4717 , \4718 );
not \U$4473 ( \4720 , \4719 );
or \U$4474 ( \4721 , \4505 , \4720 );
nand \U$4475 ( \4722 , \4714 , \4559 );
nand \U$4476 ( \4723 , \4721 , \4722 );
xnor \U$4477 ( \4724 , \4502 , \4723 );
not \U$4478 ( \4725 , \4724 );
or \U$4479 ( \4726 , \4501 , \4725 );
not \U$4480 ( \4727 , \4502 );
nand \U$4481 ( \4728 , \4727 , \4723 );
nand \U$4482 ( \4729 , \4726 , \4728 );
not \U$4483 ( \4730 , \4729 );
not \U$4484 ( \4731 , \4291 );
not \U$4485 ( \4732 , \4731 );
not \U$4486 ( \4733 , \4237 );
or \U$4487 ( \4734 , \4732 , \4733 );
not \U$4488 ( \4735 , \4237 );
nand \U$4489 ( \4736 , \4735 , \4291 );
nand \U$4490 ( \4737 , \4734 , \4736 );
and \U$4491 ( \4738 , \2918 , \3014 );
not \U$4492 ( \4739 , \2918 );
not \U$4493 ( \4740 , \3014 );
and \U$4494 ( \4741 , \4739 , \4740 );
nor \U$4495 ( \4742 , \4738 , \4741 );
and \U$4496 ( \4743 , \4737 , \4742 );
not \U$4497 ( \4744 , \4737 );
not \U$4498 ( \4745 , \4742 );
and \U$4499 ( \4746 , \4744 , \4745 );
nor \U$4500 ( \4747 , \4743 , \4746 );
not \U$4501 ( \4748 , \4747 );
or \U$4502 ( \4749 , \4730 , \4748 );
nand \U$4503 ( \4750 , \4737 , \4742 );
nand \U$4504 ( \4751 , \4749 , \4750 );
not \U$4505 ( \4752 , \4751 );
nand \U$4506 ( \4753 , \4314 , \4752 );
nand \U$4507 ( \4754 , \4308 , \4753 );
xor \U$4508 ( \4755 , \4500 , \4724 );
not \U$4509 ( \4756 , \4755 );
xor \U$4510 ( \4757 , \4286 , \4238 );
xor \U$4511 ( \4758 , \4476 , \4322 );
not \U$4512 ( \4759 , \4758 );
xor \U$4513 ( \4760 , \4678 , \4685 );
xor \U$4514 ( \4761 , \4760 , \4693 );
xor \U$4515 ( \4762 , \4625 , \4636 );
xnor \U$4516 ( \4763 , \4762 , \4630 );
xor \U$4517 ( \4764 , \4761 , \4763 );
and \U$4518 ( \4765 , \4587 , \4563 );
not \U$4519 ( \4766 , \4587 );
and \U$4520 ( \4767 , \4766 , \4564 );
nor \U$4521 ( \4768 , \4765 , \4767 );
and \U$4522 ( \4769 , \4764 , \4768 );
and \U$4523 ( \4770 , \4761 , \4763 );
or \U$4524 ( \4771 , \4769 , \4770 );
xor \U$4525 ( \4772 , \4655 , \4662 );
not \U$4526 ( \4773 , \4772 );
xor \U$4527 ( \4774 , \4533 , \4539 );
xor \U$4528 ( \4775 , \4774 , \4547 );
nand \U$4529 ( \4776 , \4773 , \4775 );
not \U$4530 ( \4777 , \4609 );
nand \U$4531 ( \4778 , \4777 , \4617 );
xor \U$4532 ( \4779 , \4778 , \4615 );
and \U$4533 ( \4780 , \4776 , \4779 );
not \U$4534 ( \4781 , \4772 );
nor \U$4535 ( \4782 , \4781 , \4775 );
nor \U$4536 ( \4783 , \4780 , \4782 );
xor \U$4537 ( \4784 , \4771 , \4783 );
xor \U$4538 ( \4785 , \4512 , \4515 );
xor \U$4539 ( \4786 , \4785 , \4517 );
and \U$4540 ( \4787 , \4784 , \4786 );
and \U$4541 ( \4788 , \4771 , \4783 );
nor \U$4542 ( \4789 , \4787 , \4788 );
xor \U$4543 ( \4790 , RIbe294e8_56, RIbe28b88_36);
not \U$4544 ( \4791 , \4790 );
not \U$4545 ( \4792 , \2554 );
or \U$4546 ( \4793 , \4791 , \4792 );
nand \U$4547 ( \4794 , \2560 , \4330 );
nand \U$4548 ( \4795 , \4793 , \4794 );
not \U$4549 ( \4796 , \2758 );
xor \U$4550 ( \4797 , RIbe28318_18, RIbe285e8_24);
not \U$4551 ( \4798 , \4797 );
or \U$4552 ( \4799 , \4796 , \4798 );
xor \U$4553 ( \4800 , RIbe28c78_38, RIbe285e8_24);
not \U$4554 ( \4801 , \4800 );
or \U$4555 ( \4802 , \2762 , \4801 );
nand \U$4556 ( \4803 , \4799 , \4802 );
or \U$4557 ( \4804 , \4795 , \4803 );
not \U$4558 ( \4805 , RIbe29128_48);
not \U$4559 ( \4806 , RIbe280c0_13);
or \U$4560 ( \4807 , \4805 , \4806 );
or \U$4561 ( \4808 , RIbe280c0_13, RIbe29128_48);
nand \U$4562 ( \4809 , \4807 , \4808 );
or \U$4563 ( \4810 , \863 , \4809 );
xnor \U$4564 ( \4811 , RIbe280c0_13, RIbe291a0_49);
or \U$4565 ( \4812 , \1516 , \4811 );
nand \U$4566 ( \4813 , \4810 , \4812 );
nand \U$4567 ( \4814 , \4804 , \4813 );
nand \U$4568 ( \4815 , \4795 , \4803 );
and \U$4569 ( \4816 , \4814 , \4815 );
not \U$4570 ( \4817 , \4816 );
not \U$4571 ( \4818 , \4817 );
xor \U$4572 ( \4819 , RIbe27e68_8, RIbe284f8_22);
not \U$4573 ( \4820 , \4819 );
not \U$4574 ( \4821 , \4443 );
or \U$4575 ( \4822 , \4820 , \4821 );
nand \U$4576 ( \4823 , \4447 , \4440 );
nand \U$4577 ( \4824 , \4822 , \4823 );
xor \U$4578 ( \4825 , RIbe27b98_2, RIbe29ec0_77);
not \U$4579 ( \4826 , \4825 );
not \U$4580 ( \4827 , \255 );
buf \U$4581 ( \4828 , \4827 );
not \U$4582 ( \4829 , \4828 );
or \U$4583 ( \4830 , \4826 , \4829 );
nand \U$4584 ( \4831 , \269 , \4414 );
nand \U$4585 ( \4832 , \4830 , \4831 );
nor \U$4586 ( \4833 , \4824 , \4832 );
and \U$4587 ( \4834 , RIbe2a028_80, RIbe29fb0_79);
not \U$4588 ( \4835 , RIbe2a028_80);
and \U$4589 ( \4836 , \4835 , RIbe29e48_76);
nor \U$4590 ( \4837 , \4834 , \4836 );
not \U$4591 ( \4838 , \4837 );
nand \U$4592 ( \4839 , RIbe29e48_76, RIbe29fb0_79);
nand \U$4593 ( \4840 , \4838 , \4839 );
buf \U$4594 ( \4841 , \4840 );
not \U$4595 ( \4842 , \4841 );
buf \U$4596 ( \4843 , \4842 );
not \U$4597 ( \4844 , RIbe29fb0_79);
not \U$4598 ( \4845 , RIbe2a028_80);
and \U$4599 ( \4846 , \4844 , \4845 );
and \U$4600 ( \4847 , RIbe29fb0_79, RIbe2a028_80);
nor \U$4601 ( \4848 , \4846 , \4847 );
buf \U$4602 ( \4849 , \4848 );
buf \U$4603 ( \4850 , \4849 );
buf \U$4604 ( \4851 , \4850 );
or \U$4605 ( \4852 , \4843 , \4851 );
nand \U$4606 ( \4853 , \4852 , RIbe29e48_76);
not \U$4607 ( \4854 , \4853 );
or \U$4608 ( \4855 , \4833 , \4854 );
nand \U$4609 ( \4856 , \4824 , \4832 );
nand \U$4610 ( \4857 , \4855 , \4856 );
and \U$4611 ( \4858 , RIbe28480_21, RIbe29308_52);
nor \U$4612 ( \4859 , RIbe28480_21, RIbe29308_52);
nor \U$4613 ( \4860 , \4858 , \4859 );
not \U$4614 ( \4861 , \4860 );
not \U$4615 ( \4862 , \2519 );
or \U$4616 ( \4863 , \4861 , \4862 );
not \U$4617 ( \4864 , \4420 );
nand \U$4618 ( \4865 , \4864 , \3075 );
nand \U$4619 ( \4866 , \4863 , \4865 );
not \U$4620 ( \4867 , \4866 );
and \U$4621 ( \4868 , RIbe29f38_78, RIbe27b98_2);
xor \U$4622 ( \4869 , RIbe28de0_41, RIbe29ce0_73);
not \U$4623 ( \4870 , \4869 );
not \U$4624 ( \4871 , \331 );
or \U$4625 ( \4872 , \4870 , \4871 );
nand \U$4626 ( \4873 , \347 , \4407 );
nand \U$4627 ( \4874 , \4872 , \4873 );
xor \U$4628 ( \4875 , \4868 , \4874 );
not \U$4629 ( \4876 , \4875 );
or \U$4630 ( \4877 , \4867 , \4876 );
nand \U$4631 ( \4878 , \4874 , \4868 );
nand \U$4632 ( \4879 , \4877 , \4878 );
not \U$4633 ( \4880 , \4879 );
and \U$4634 ( \4881 , \4857 , \4880 );
not \U$4635 ( \4882 , \4857 );
and \U$4636 ( \4883 , \4882 , \4879 );
or \U$4637 ( \4884 , \4881 , \4883 );
not \U$4638 ( \4885 , \4884 );
or \U$4639 ( \4886 , \4818 , \4885 );
not \U$4640 ( \4887 , \4880 );
nand \U$4641 ( \4888 , \4887 , \4857 );
nand \U$4642 ( \4889 , \4886 , \4888 );
not \U$4643 ( \4890 , \4889 );
xor \U$4644 ( \4891 , RIbe28840_29, RIbe27fd0_11);
not \U$4645 ( \4892 , \4891 );
not \U$4646 ( \4893 , \2717 );
not \U$4647 ( \4894 , \4893 );
or \U$4648 ( \4895 , \4892 , \4894 );
not \U$4649 ( \4896 , \2706 );
not \U$4650 ( \4897 , \4896 );
nand \U$4651 ( \4898 , \4897 , \4372 );
nand \U$4652 ( \4899 , \4895 , \4898 );
not \U$4653 ( \4900 , \4899 );
not \U$4654 ( \4901 , RIbe28930_31);
not \U$4655 ( \4902 , RIbe297b8_62);
and \U$4656 ( \4903 , \4901 , \4902 );
and \U$4657 ( \4904 , RIbe28930_31, RIbe297b8_62);
nor \U$4658 ( \4905 , \4903 , \4904 );
not \U$4659 ( \4906 , \4905 );
not \U$4660 ( \4907 , \966 );
or \U$4661 ( \4908 , \4906 , \4907 );
not \U$4662 ( \4909 , RIbe28138_14);
not \U$4663 ( \4910 , RIbe28930_31);
and \U$4664 ( \4911 , \4909 , \4910 );
and \U$4665 ( \4912 , RIbe28138_14, RIbe28930_31);
nor \U$4666 ( \4913 , \4911 , \4912 );
nand \U$4667 ( \4914 , \1797 , \4913 );
nand \U$4668 ( \4915 , \4908 , \4914 );
not \U$4669 ( \4916 , \4915 );
or \U$4670 ( \4917 , \4900 , \4916 );
or \U$4671 ( \4918 , \4915 , \4899 );
xor \U$4672 ( \4919 , RIbe298a8_64, RIbe27d78_6);
not \U$4673 ( \4920 , \4919 );
not \U$4674 ( \4921 , \1164 );
or \U$4675 ( \4922 , \4920 , \4921 );
xor \U$4676 ( \4923 , RIbe27d78_6, RIbe29998_66);
nand \U$4677 ( \4924 , \315 , \4923 );
nand \U$4678 ( \4925 , \4922 , \4924 );
nand \U$4679 ( \4926 , \4918 , \4925 );
nand \U$4680 ( \4927 , \4917 , \4926 );
not \U$4681 ( \4928 , \4927 );
xor \U$4682 ( \4929 , RIbe27c10_3, RIbe28cf0_39);
not \U$4683 ( \4930 , \4929 );
not \U$4684 ( \4931 , \1103 );
or \U$4685 ( \4932 , \4930 , \4931 );
not \U$4686 ( \4933 , \4528 );
nand \U$4687 ( \4934 , \4933 , \370 );
nand \U$4688 ( \4935 , \4932 , \4934 );
xnor \U$4689 ( \4936 , \4935 , \4338 );
not \U$4690 ( \4937 , \4936 );
or \U$4691 ( \4938 , \4928 , \4937 );
nand \U$4692 ( \4939 , \4339 , \4935 );
nand \U$4693 ( \4940 , \4938 , \4939 );
xor \U$4694 ( \4941 , \4339 , \4346 );
xor \U$4695 ( \4942 , \4941 , \4352 );
xor \U$4696 ( \4943 , \4940 , \4942 );
or \U$4697 ( \4944 , \4890 , \4943 );
not \U$4698 ( \4945 , \4940 );
or \U$4699 ( \4946 , \4945 , \4942 );
nand \U$4700 ( \4947 , \4944 , \4946 );
not \U$4701 ( \4948 , \4947 );
xor \U$4702 ( \4949 , \4523 , \4525 );
not \U$4703 ( \4950 , \4550 );
xor \U$4704 ( \4951 , \4949 , \4950 );
xor \U$4705 ( \4952 , \4365 , \4467 );
not \U$4706 ( \4953 , \4952 );
and \U$4707 ( \4954 , \4951 , \4953 );
not \U$4708 ( \4955 , \4951 );
and \U$4709 ( \4956 , \4955 , \4952 );
or \U$4710 ( \4957 , \4954 , \4956 );
not \U$4711 ( \4958 , \4957 );
or \U$4712 ( \4959 , \4948 , \4958 );
not \U$4713 ( \4960 , \4953 );
nand \U$4714 ( \4961 , \4960 , \4951 );
nand \U$4715 ( \4962 , \4959 , \4961 );
xor \U$4716 ( \4963 , \4789 , \4962 );
not \U$4717 ( \4964 , \4963 );
or \U$4718 ( \4965 , \4759 , \4964 );
nand \U$4719 ( \4966 , \4962 , \4789 );
nand \U$4720 ( \4967 , \4965 , \4966 );
not \U$4721 ( \4968 , \4967 );
not \U$4722 ( \4969 , \4503 );
not \U$4723 ( \4970 , \4719 );
or \U$4724 ( \4971 , \4969 , \4970 );
or \U$4725 ( \4972 , \4719 , \4503 );
nand \U$4726 ( \4973 , \4971 , \4972 );
xor \U$4727 ( \4974 , \4507 , \4520 );
xor \U$4728 ( \4975 , \4974 , \4555 );
not \U$4729 ( \4976 , \4975 );
not \U$4730 ( \4977 , \4976 );
xnor \U$4731 ( \4978 , \4705 , \4709 );
not \U$4732 ( \4979 , \4978 );
and \U$4733 ( \4980 , \4643 , \4592 );
not \U$4734 ( \4981 , \4643 );
not \U$4735 ( \4982 , \4592 );
and \U$4736 ( \4983 , \4981 , \4982 );
nor \U$4737 ( \4984 , \4980 , \4983 );
not \U$4738 ( \4985 , \4984 );
not \U$4739 ( \4986 , \4696 );
not \U$4740 ( \4987 , \4671 );
or \U$4741 ( \4988 , \4986 , \4987 );
or \U$4742 ( \4989 , \4671 , \4696 );
nand \U$4743 ( \4990 , \4988 , \4989 );
not \U$4744 ( \4991 , \4990 );
not \U$4745 ( \4992 , \4797 );
not \U$4746 ( \4993 , \2890 );
or \U$4747 ( \4994 , \4992 , \4993 );
not \U$4748 ( \4995 , \4606 );
nand \U$4749 ( \4996 , \4995 , \2758 );
nand \U$4750 ( \4997 , \4994 , \4996 );
not \U$4751 ( \4998 , \4997 );
or \U$4752 ( \4999 , \1325 , \4811 );
or \U$4753 ( \5000 , \1516 , \4611 );
nand \U$4754 ( \5001 , \4999 , \5000 );
not \U$4755 ( \5002 , \5001 );
or \U$4756 ( \5003 , \4998 , \5002 );
or \U$4757 ( \5004 , \4997 , \5001 );
xor \U$4758 ( \5005 , RIbe293f8_54, RIbe28390_19);
not \U$4759 ( \5006 , \5005 );
not \U$4760 ( \5007 , \2640 );
or \U$4761 ( \5008 , \5006 , \5007 );
nand \U$4762 ( \5009 , \3714 , \4597 );
nand \U$4763 ( \5010 , \5008 , \5009 );
nand \U$4764 ( \5011 , \5004 , \5010 );
nand \U$4765 ( \5012 , \5003 , \5011 );
not \U$4766 ( \5013 , \5012 );
not \U$4767 ( \5014 , \4913 );
not \U$4768 ( \5015 , \966 );
or \U$4769 ( \5016 , \5014 , \5015 );
nand \U$4770 ( \5017 , \971 , \4690 );
nand \U$4771 ( \5018 , \5016 , \5017 );
not \U$4772 ( \5019 , \5018 );
nand \U$4773 ( \5020 , RIbe27b98_2, RIbe29ec0_77);
not \U$4774 ( \5021 , \5020 );
xor \U$4775 ( \5022 , RIbe29c68_72, RIbe29380_53);
not \U$4776 ( \5023 , \5022 );
not \U$4777 ( \5024 , \4576 );
not \U$4778 ( \5025 , \5024 );
or \U$4779 ( \5026 , \5023 , \5025 );
nand \U$4780 ( \5027 , \4580 , RIbe29c68_72);
nand \U$4781 ( \5028 , \5026 , \5027 );
not \U$4782 ( \5029 , \5028 );
or \U$4783 ( \5030 , \5021 , \5029 );
or \U$4784 ( \5031 , \5028 , \5020 );
nand \U$4785 ( \5032 , \5030 , \5031 );
not \U$4786 ( \5033 , \5032 );
or \U$4787 ( \5034 , \5019 , \5033 );
not \U$4788 ( \5035 , \5020 );
nand \U$4789 ( \5036 , \5035 , \5028 );
nand \U$4790 ( \5037 , \5034 , \5036 );
not \U$4791 ( \5038 , \5037 );
not \U$4792 ( \5039 , \5038 );
or \U$4793 ( \5040 , \5013 , \5039 );
or \U$4794 ( \5041 , \5038 , \5012 );
nand \U$4795 ( \5042 , \5040 , \5041 );
not \U$4796 ( \5043 , \5042 );
not \U$4797 ( \5044 , \4923 );
not \U$4798 ( \5045 , \1044 );
or \U$4799 ( \5046 , \5044 , \5045 );
nand \U$4800 ( \5047 , \314 , \4341 );
nand \U$4801 ( \5048 , \5046 , \5047 );
not \U$4802 ( \5049 , \5048 );
xor \U$4803 ( \5050 , RIbe29470_55, RIbe28a20_33);
not \U$4804 ( \5051 , \5050 );
not \U$4805 ( \5052 , \1781 );
or \U$4806 ( \5053 , \5051 , \5052 );
xor \U$4807 ( \5054 , RIbe28b88_36, RIbe29290_51);
buf \U$4808 ( \5055 , \5054 );
nand \U$4809 ( \5056 , \5055 , \4680 );
nand \U$4810 ( \5057 , \5053 , \5056 );
not \U$4811 ( \5058 , \5057 );
or \U$4812 ( \5059 , \5049 , \5058 );
or \U$4813 ( \5060 , \5057 , \5048 );
not \U$4814 ( \5061 , RIbe27c88_4);
not \U$4815 ( \5062 , RIbe290b0_47);
and \U$4816 ( \5063 , \5061 , \5062 );
and \U$4817 ( \5064 , RIbe27c88_4, RIbe290b0_47);
nor \U$4818 ( \5065 , \5063 , \5064 );
not \U$4819 ( \5066 , \5065 );
not \U$4820 ( \5067 , \525 );
or \U$4821 ( \5068 , \5066 , \5067 );
not \U$4822 ( \5069 , \4535 );
nand \U$4823 ( \5070 , \5069 , \399 );
nand \U$4824 ( \5071 , \5068 , \5070 );
nand \U$4825 ( \5072 , \5060 , \5071 );
nand \U$4826 ( \5073 , \5059 , \5072 );
not \U$4827 ( \5074 , \5073 );
or \U$4828 ( \5075 , \5043 , \5074 );
nand \U$4829 ( \5076 , \5037 , \5012 );
nand \U$4830 ( \5077 , \5075 , \5076 );
not \U$4831 ( \5078 , \5077 );
not \U$4832 ( \5079 , \5078 );
and \U$4833 ( \5080 , \4991 , \5079 );
and \U$4834 ( \5081 , \4990 , \5078 );
nor \U$4835 ( \5082 , \5080 , \5081 );
not \U$4836 ( \5083 , \5082 );
not \U$4837 ( \5084 , \5083 );
or \U$4838 ( \5085 , \4985 , \5084 );
not \U$4839 ( \5086 , \5078 );
nand \U$4840 ( \5087 , \5086 , \4990 );
nand \U$4841 ( \5088 , \5085 , \5087 );
not \U$4842 ( \5089 , \5088 );
or \U$4843 ( \5090 , \4979 , \5089 );
or \U$4844 ( \5091 , \5088 , \4978 );
nand \U$4845 ( \5092 , \5090 , \5091 );
not \U$4846 ( \5093 , \5092 );
or \U$4847 ( \5094 , \4977 , \5093 );
not \U$4848 ( \5095 , \4978 );
nand \U$4849 ( \5096 , \5095 , \5088 );
nand \U$4850 ( \5097 , \5094 , \5096 );
nor \U$4851 ( \5098 , \4973 , \5097 );
not \U$4852 ( \5099 , \5098 );
not \U$4853 ( \5100 , \5099 );
or \U$4854 ( \5101 , \4968 , \5100 );
nand \U$4855 ( \5102 , \5097 , \4973 );
nand \U$4856 ( \5103 , \5101 , \5102 );
xor \U$4857 ( \5104 , \4757 , \5103 );
not \U$4858 ( \5105 , \5104 );
or \U$4859 ( \5106 , \4756 , \5105 );
nand \U$4860 ( \5107 , \5103 , \4757 );
nand \U$4861 ( \5108 , \5106 , \5107 );
xor \U$4862 ( \5109 , \4747 , \4729 );
nand \U$4863 ( \5110 , \5108 , \5109 );
or \U$4864 ( \5111 , \4754 , \5110 );
not \U$4865 ( \5112 , \4307 );
nand \U$4866 ( \5113 , \4313 , \4751 );
not \U$4867 ( \5114 , \5113 );
and \U$4868 ( \5115 , \5112 , \5114 );
nand \U$4869 ( \5116 , \3939 , \4306 );
or \U$4870 ( \5117 , \3675 , \3790 );
nand \U$4871 ( \5118 , \3569 , \3674 );
nand \U$4872 ( \5119 , \5117 , \5118 );
not \U$4873 ( \5120 , \3670 );
not \U$4874 ( \5121 , \3655 );
or \U$4875 ( \5122 , \5120 , \5121 );
nand \U$4876 ( \5123 , \3624 , \3650 );
nand \U$4877 ( \5124 , \5122 , \5123 );
or \U$4878 ( \5125 , \524 , \3783 );
xnor \U$4879 ( \5126 , RIbe28138_14, RIbe290b0_47);
or \U$4880 ( \5127 , \468 , \5126 );
nand \U$4881 ( \5128 , \5125 , \5127 );
not \U$4882 ( \5129 , \3756 );
not \U$4883 ( \5130 , \5129 );
not \U$4884 ( \5131 , \2276 );
or \U$4885 ( \5132 , \5130 , \5131 );
xor \U$4886 ( \5133 , RIbe28a20_33, RIbe28750_27);
nand \U$4887 ( \5134 , \1769 , \5133 );
nand \U$4888 ( \5135 , \5132 , \5134 );
xor \U$4889 ( \5136 , \5128 , \5135 );
not \U$4890 ( \5137 , \3880 );
not \U$4891 ( \5138 , \936 );
or \U$4892 ( \5139 , \5137 , \5138 );
not \U$4893 ( \5140 , RIbe27c10_3);
not \U$4894 ( \5141 , RIbe291a0_49);
and \U$4895 ( \5142 , \5140 , \5141 );
and \U$4896 ( \5143 , RIbe27c10_3, RIbe291a0_49);
nor \U$4897 ( \5144 , \5142 , \5143 );
nand \U$4898 ( \5145 , \370 , \5144 );
nand \U$4899 ( \5146 , \5139 , \5145 );
xor \U$4900 ( \5147 , \5136 , \5146 );
not \U$4901 ( \5148 , \2758 );
not \U$4902 ( \5149 , \5148 );
not \U$4903 ( \5150 , \2617 );
or \U$4904 ( \5151 , \5149 , \5150 );
nand \U$4905 ( \5152 , \5151 , RIbe285e8_24);
and \U$4906 ( \5153 , RIbe27d78_6, RIbe29740_61);
not \U$4907 ( \5154 , RIbe27d78_6);
and \U$4908 ( \5155 , \5154 , \3185 );
nor \U$4909 ( \5156 , \5153 , \5155 );
not \U$4910 ( \5157 , \5156 );
not \U$4911 ( \5158 , \315 );
or \U$4912 ( \5159 , \5157 , \5158 );
nand \U$4913 ( \5160 , \1164 , \3744 );
nand \U$4914 ( \5161 , \5159 , \5160 );
xor \U$4915 ( \5162 , \5152 , \5161 );
or \U$4916 ( \5163 , \946 , \3776 );
xnor \U$4917 ( \5164 , RIbe29218_50, RIbe27b98_2);
or \U$4918 ( \5165 , \1735 , \5164 );
nand \U$4919 ( \5166 , \5163 , \5165 );
xor \U$4920 ( \5167 , \5162 , \5166 );
not \U$4921 ( \5168 , \5167 );
or \U$4922 ( \5169 , \283 , \3723 );
xnor \U$4923 ( \5170 , RIbe29470_55, RIbe29038_46);
or \U$4924 ( \5171 , \1465 , \5170 );
nand \U$4925 ( \5172 , \5169 , \5171 );
not \U$4926 ( \5173 , \5172 );
not \U$4927 ( \5174 , \3949 );
not \U$4928 ( \5175 , \3862 );
and \U$4929 ( \5176 , \5174 , \5175 );
not \U$4930 ( \5177 , \1199 );
not \U$4931 ( \5178 , RIbe28930_31);
not \U$4932 ( \5179 , RIbe28318_18);
or \U$4933 ( \5180 , \5178 , \5179 );
or \U$4934 ( \5181 , RIbe28318_18, RIbe28930_31);
nand \U$4935 ( \5182 , \5180 , \5181 );
nor \U$4936 ( \5183 , \5177 , \5182 );
nor \U$4937 ( \5184 , \5176 , \5183 );
not \U$4938 ( \5185 , \5184 );
or \U$4939 ( \5186 , \5173 , \5185 );
or \U$4940 ( \5187 , \5172 , \5184 );
nand \U$4941 ( \5188 , \5186 , \5187 );
not \U$4942 ( \5189 , \5188 );
nand \U$4943 ( \5190 , \900 , \3732 );
not \U$4944 ( \5191 , RIbe296c8_60);
not \U$4945 ( \5192 , RIbe288b8_30);
or \U$4946 ( \5193 , \5191 , \5192 );
or \U$4947 ( \5194 , RIbe288b8_30, RIbe296c8_60);
nand \U$4948 ( \5195 , \5193 , \5194 );
not \U$4949 ( \5196 , \5195 );
nand \U$4950 ( \5197 , \5196 , \1137 );
and \U$4951 ( \5198 , \5190 , \5197 );
not \U$4952 ( \5199 , \5198 );
and \U$4953 ( \5200 , \5189 , \5199 );
and \U$4954 ( \5201 , \5188 , \5198 );
nor \U$4955 ( \5202 , \5200 , \5201 );
not \U$4956 ( \5203 , \5202 );
or \U$4957 ( \5204 , \5168 , \5203 );
or \U$4958 ( \5205 , \5202 , \5167 );
nand \U$4959 ( \5206 , \5204 , \5205 );
xor \U$4960 ( \5207 , \5147 , \5206 );
not \U$4961 ( \5208 , \886 );
and \U$4962 ( \5209 , RIbe28228_16, \2479 );
not \U$4963 ( \5210 , RIbe28228_16);
and \U$4964 ( \5211 , \5210 , RIbe28c00_37);
nor \U$4965 ( \5212 , \5209 , \5211 );
not \U$4966 ( \5213 , \5212 );
and \U$4967 ( \5214 , \5208 , \5213 );
and \U$4968 ( \5215 , \1061 , \3843 );
nor \U$4969 ( \5216 , \5214 , \5215 );
not \U$4970 ( \5217 , \3412 );
and \U$4971 ( \5218 , RIbe28390_19, RIbe27ee0_9);
not \U$4972 ( \5219 , RIbe28390_19);
and \U$4973 ( \5220 , \5219 , \317 );
nor \U$4974 ( \5221 , \5218 , \5220 );
not \U$4975 ( \5222 , \5221 );
not \U$4976 ( \5223 , \5222 );
and \U$4977 ( \5224 , \5217 , \5223 );
and \U$4978 ( \5225 , \3712 , \3717 );
nor \U$4979 ( \5226 , \5224 , \5225 );
xor \U$4980 ( \5227 , \5216 , \5226 );
and \U$4981 ( \5228 , \862 , \3853 );
xnor \U$4982 ( \5229 , RIbe280c0_13, RIbe293f8_54);
not \U$4983 ( \5230 , \5229 );
and \U$4984 ( \5231 , \1265 , \5230 );
nor \U$4985 ( \5232 , \5228 , \5231 );
xor \U$4986 ( \5233 , \5227 , \5232 );
not \U$4987 ( \5234 , \5233 );
not \U$4988 ( \5235 , \3758 );
not \U$4989 ( \5236 , \3749 );
or \U$4990 ( \5237 , \5235 , \5236 );
nand \U$4991 ( \5238 , \3742 , \3748 );
nand \U$4992 ( \5239 , \5237 , \5238 );
not \U$4993 ( \5240 , \5239 );
or \U$4994 ( \5241 , \2667 , \3767 );
and \U$4995 ( \5242 , RIbe28480_21, \388 );
not \U$4996 ( \5243 , RIbe28480_21);
and \U$4997 ( \5244 , \5243 , RIbe29380_53);
nor \U$4998 ( \5245 , \5242 , \5244 );
or \U$4999 ( \5246 , \5245 , \2672 );
nand \U$5000 ( \5247 , \5241 , \5246 );
not \U$5001 ( \5248 , \5247 );
and \U$5002 ( \5249 , RIbe27c88_4, RIbe27b98_2);
not \U$5003 ( \5250 , \3740 );
not \U$5004 ( \5251 , \3103 );
or \U$5005 ( \5252 , \5250 , \5251 );
xor \U$5006 ( \5253 , RIbe28de0_41, RIbe29b00_69);
nand \U$5007 ( \5254 , \514 , \5253 );
nand \U$5008 ( \5255 , \5252 , \5254 );
xor \U$5009 ( \5256 , \5249 , \5255 );
not \U$5010 ( \5257 , \5256 );
not \U$5011 ( \5258 , \5257 );
or \U$5012 ( \5259 , \5248 , \5258 );
or \U$5013 ( \5260 , \5257 , \5247 );
nand \U$5014 ( \5261 , \5259 , \5260 );
not \U$5015 ( \5262 , \5261 );
not \U$5016 ( \5263 , \5262 );
or \U$5017 ( \5264 , \5240 , \5263 );
not \U$5018 ( \5265 , \5239 );
nand \U$5019 ( \5266 , \5265 , \5261 );
nand \U$5020 ( \5267 , \5264 , \5266 );
not \U$5021 ( \5268 , \5267 );
or \U$5022 ( \5269 , \5234 , \5268 );
or \U$5023 ( \5270 , \5267 , \5233 );
nand \U$5024 ( \5271 , \5269 , \5270 );
xor \U$5025 ( \5272 , \5207 , \5271 );
xnor \U$5026 ( \5273 , \5124 , \5272 );
not \U$5027 ( \5274 , \5273 );
not \U$5028 ( \5275 , \3913 );
or \U$5029 ( \5276 , \5275 , \3922 );
nand \U$5030 ( \5277 , \3907 , \3901 );
nand \U$5031 ( \5278 , \5276 , \5277 );
not \U$5032 ( \5279 , \5278 );
or \U$5033 ( \5280 , \5274 , \5279 );
or \U$5034 ( \5281 , \5278 , \5273 );
nand \U$5035 ( \5282 , \5280 , \5281 );
xor \U$5036 ( \5283 , \5119 , \5282 );
not \U$5037 ( \5284 , \3789 );
not \U$5038 ( \5285 , \3711 );
or \U$5039 ( \5286 , \5284 , \5285 );
not \U$5040 ( \5287 , \3681 );
nand \U$5041 ( \5288 , \5287 , \3707 );
nand \U$5042 ( \5289 , \5286 , \5288 );
not \U$5043 ( \5290 , \2560 );
and \U$5044 ( \5291 , RIbe28570_23, RIbe28b88_36);
nor \U$5045 ( \5292 , RIbe28570_23, RIbe28b88_36);
nor \U$5046 ( \5293 , \5291 , \5292 );
not \U$5047 ( \5294 , \5293 );
or \U$5048 ( \5295 , \5290 , \5294 );
or \U$5049 ( \5296 , \3960 , \3615 );
nand \U$5050 ( \5297 , \5295 , \5296 );
and \U$5051 ( \5298 , \3618 , \5297 );
not \U$5052 ( \5299 , \5298 );
not \U$5053 ( \5300 , \5297 );
nand \U$5054 ( \5301 , \5300 , \3621 );
nand \U$5055 ( \5302 , \5299 , \5301 );
not \U$5056 ( \5303 , \3786 );
not \U$5057 ( \5304 , \3779 );
or \U$5058 ( \5305 , \5303 , \5304 );
or \U$5059 ( \5306 , \3786 , \3779 );
nand \U$5060 ( \5307 , \5306 , \3769 );
nand \U$5061 ( \5308 , \5305 , \5307 );
xnor \U$5062 ( \5309 , \5302 , \5308 );
xor \U$5063 ( \5310 , \3659 , \3663 );
and \U$5064 ( \5311 , \5310 , \3668 );
and \U$5065 ( \5312 , \3659 , \3663 );
or \U$5066 ( \5313 , \5311 , \5312 );
xor \U$5067 ( \5314 , \5309 , \5313 );
not \U$5068 ( \5315 , \3605 );
not \U$5069 ( \5316 , \3623 );
or \U$5070 ( \5317 , \5315 , \5316 );
nand \U$5071 ( \5318 , \3611 , \3621 );
nand \U$5072 ( \5319 , \5317 , \5318 );
xor \U$5073 ( \5320 , \5314 , \5319 );
not \U$5074 ( \5321 , \5320 );
and \U$5075 ( \5322 , \5289 , \5321 );
not \U$5076 ( \5323 , \5289 );
and \U$5077 ( \5324 , \5323 , \5320 );
nor \U$5078 ( \5325 , \5322 , \5324 );
xor \U$5079 ( \5326 , \3736 , \3759 );
and \U$5080 ( \5327 , \5326 , \3788 );
and \U$5081 ( \5328 , \3736 , \3759 );
nor \U$5082 ( \5329 , \5327 , \5328 );
not \U$5083 ( \5330 , \3875 );
not \U$5084 ( \5331 , \3893 );
not \U$5085 ( \5332 , \5331 );
or \U$5086 ( \5333 , \5330 , \5332 );
not \U$5087 ( \5334 , \3866 );
nand \U$5088 ( \5335 , \5334 , \3897 );
nand \U$5089 ( \5336 , \5333 , \5335 );
not \U$5090 ( \5337 , \5336 );
or \U$5091 ( \5338 , \3884 , \3892 );
nand \U$5092 ( \5339 , \5338 , \3886 );
not \U$5093 ( \5340 , \3734 );
not \U$5094 ( \5341 , \3726 );
or \U$5095 ( \5342 , \5340 , \5341 );
not \U$5096 ( \5343 , \3719 );
nand \U$5097 ( \5344 , \5343 , \3735 );
nand \U$5098 ( \5345 , \5342 , \5344 );
xor \U$5099 ( \5346 , \5339 , \5345 );
not \U$5100 ( \5347 , \5346 );
xor \U$5101 ( \5348 , \3845 , \3855 );
and \U$5102 ( \5349 , \5348 , \3865 );
and \U$5103 ( \5350 , \3845 , \3855 );
or \U$5104 ( \5351 , \5349 , \5350 );
not \U$5105 ( \5352 , \5351 );
and \U$5106 ( \5353 , \5347 , \5352 );
and \U$5107 ( \5354 , \5346 , \5351 );
nor \U$5108 ( \5355 , \5353 , \5354 );
not \U$5109 ( \5356 , \5355 );
or \U$5110 ( \5357 , \5337 , \5356 );
or \U$5111 ( \5358 , \5355 , \5336 );
nand \U$5112 ( \5359 , \5357 , \5358 );
not \U$5113 ( \5360 , \5359 );
xor \U$5114 ( \5361 , \5329 , \5360 );
xor \U$5115 ( \5362 , \5325 , \5361 );
not \U$5116 ( \5363 , \3829 );
not \U$5117 ( \5364 , \3930 );
or \U$5118 ( \5365 , \5363 , \5364 );
nand \U$5119 ( \5366 , \3924 , \3837 );
nand \U$5120 ( \5367 , \5365 , \5366 );
xor \U$5121 ( \5368 , \5362 , \5367 );
xor \U$5122 ( \5369 , \5283 , \5368 );
not \U$5123 ( \5370 , \3470 );
not \U$5124 ( \5371 , \3938 );
or \U$5125 ( \5372 , \5370 , \5371 );
not \U$5126 ( \5373 , \3791 );
nand \U$5127 ( \5374 , \5373 , \3934 );
nand \U$5128 ( \5375 , \5372 , \5374 );
nand \U$5129 ( \5376 , \5369 , \5375 );
nand \U$5130 ( \5377 , \5116 , \5376 );
nor \U$5131 ( \5378 , \5115 , \5377 );
nand \U$5132 ( \5379 , \5111 , \5378 );
and \U$5133 ( \5380 , \5368 , \5283 );
and \U$5134 ( \5381 , \5362 , \5367 );
nor \U$5135 ( \5382 , \5380 , \5381 );
not \U$5136 ( \5383 , \5351 );
and \U$5137 ( \5384 , \5346 , \5383 );
and \U$5138 ( \5385 , \5339 , \5345 );
nor \U$5139 ( \5386 , \5384 , \5385 );
and \U$5140 ( \5387 , \5308 , \5301 );
nor \U$5141 ( \5388 , \5387 , \5298 );
or \U$5142 ( \5389 , RIbe28a98_34, RIbe296c8_60);
nand \U$5143 ( \5390 , RIbe28a98_34, RIbe296c8_60);
nand \U$5144 ( \5391 , \5389 , \5390 );
nor \U$5145 ( \5392 , \1938 , \5391 );
nor \U$5146 ( \5393 , \1131 , \5195 );
nor \U$5147 ( \5394 , \5392 , \5393 );
not \U$5148 ( \5395 , \5394 );
not \U$5149 ( \5396 , \5133 );
not \U$5150 ( \5397 , \2276 );
or \U$5151 ( \5398 , \5396 , \5397 );
and \U$5152 ( \5399 , RIbe28a20_33, RIbe28840_29);
not \U$5153 ( \5400 , RIbe28a20_33);
and \U$5154 ( \5401 , \5400 , \364 );
nor \U$5155 ( \5402 , \5399 , \5401 );
nand \U$5156 ( \5403 , \1769 , \5402 );
nand \U$5157 ( \5404 , \5398 , \5403 );
not \U$5158 ( \5405 , \5404 );
or \U$5159 ( \5406 , \5395 , \5405 );
or \U$5160 ( \5407 , \5404 , \5394 );
nand \U$5161 ( \5408 , \5406 , \5407 );
or \U$5162 ( \5409 , \3345 , \5245 );
not \U$5163 ( \5410 , RIbe28480_21);
or \U$5164 ( \5411 , \5410 , \2672 );
nand \U$5165 ( \5412 , \5409 , \5411 );
and \U$5166 ( \5413 , \5408 , \5412 );
not \U$5167 ( \5414 , \5408 );
not \U$5168 ( \5415 , \5412 );
and \U$5169 ( \5416 , \5414 , \5415 );
nor \U$5170 ( \5417 , \5413 , \5416 );
xnor \U$5171 ( \5418 , \5388 , \5417 );
xnor \U$5172 ( \5419 , \5386 , \5418 );
not \U$5173 ( \5420 , \5419 );
not \U$5174 ( \5421 , \5336 );
not \U$5175 ( \5422 , \5355 );
not \U$5176 ( \5423 , \5422 );
or \U$5177 ( \5424 , \5421 , \5423 );
not \U$5178 ( \5425 , \5329 );
nand \U$5179 ( \5426 , \5425 , \5359 );
nand \U$5180 ( \5427 , \5424 , \5426 );
not \U$5181 ( \5428 , \5427 );
or \U$5182 ( \5429 , \5420 , \5428 );
or \U$5183 ( \5430 , \5427 , \5419 );
nand \U$5184 ( \5431 , \5429 , \5430 );
not \U$5185 ( \5432 , \5233 );
not \U$5186 ( \5433 , \5432 );
not \U$5187 ( \5434 , \5267 );
or \U$5188 ( \5435 , \5433 , \5434 );
not \U$5189 ( \5436 , \5262 );
nand \U$5190 ( \5437 , \5436 , \5239 );
nand \U$5191 ( \5438 , \5435 , \5437 );
xor \U$5192 ( \5439 , \5216 , \5226 );
and \U$5193 ( \5440 , \5439 , \5232 );
and \U$5194 ( \5441 , \5216 , \5226 );
or \U$5195 ( \5442 , \5440 , \5441 );
not \U$5196 ( \5443 , \5442 );
xor \U$5197 ( \5444 , \5152 , \5161 );
and \U$5198 ( \5445 , \5444 , \5166 );
and \U$5199 ( \5446 , \5152 , \5161 );
or \U$5200 ( \5447 , \5445 , \5446 );
and \U$5201 ( \5448 , \5247 , \5256 );
and \U$5202 ( \5449 , \5249 , \5255 );
nor \U$5203 ( \5450 , \5448 , \5449 );
xnor \U$5204 ( \5451 , \5447 , \5450 );
not \U$5205 ( \5452 , \5451 );
or \U$5206 ( \5453 , \5443 , \5452 );
or \U$5207 ( \5454 , \5451 , \5442 );
nand \U$5208 ( \5455 , \5453 , \5454 );
xor \U$5209 ( \5456 , \5438 , \5455 );
not \U$5210 ( \5457 , \5128 );
not \U$5211 ( \5458 , \5135 );
or \U$5212 ( \5459 , \5457 , \5458 );
or \U$5213 ( \5460 , \5135 , \5128 );
nand \U$5214 ( \5461 , \5460 , \5146 );
nand \U$5215 ( \5462 , \5459 , \5461 );
not \U$5216 ( \5463 , \5198 );
nand \U$5217 ( \5464 , \5463 , \5188 );
not \U$5218 ( \5465 , \5184 );
nand \U$5219 ( \5466 , \5465 , \5172 );
nand \U$5220 ( \5467 , \5464 , \5466 );
xor \U$5221 ( \5468 , \5462 , \5467 );
or \U$5222 ( \5469 , \385 , \5126 );
not \U$5223 ( \5470 , \2071 );
and \U$5224 ( \5471 , \387 , RIbe282a0_17);
and \U$5225 ( \5472 , \951 , RIbe290b0_47);
nor \U$5226 ( \5473 , \5471 , \5472 );
or \U$5227 ( \5474 , \5470 , \5473 );
nand \U$5228 ( \5475 , \5469 , \5474 );
or \U$5229 ( \5476 , \1575 , \5229 );
xnor \U$5230 ( \5477 , RIbe280c0_13, RIbe29308_52);
or \U$5231 ( \5478 , \1573 , \5477 );
nand \U$5232 ( \5479 , \5476 , \5478 );
xor \U$5233 ( \5480 , \5475 , \5479 );
not \U$5234 ( \5481 , \5293 );
not \U$5235 ( \5482 , \3402 );
or \U$5236 ( \5483 , \5481 , \5482 );
and \U$5237 ( \5484 , \3970 , \304 );
and \U$5238 ( \5485 , RIbe286d8_26, RIbe28b88_36);
nor \U$5239 ( \5486 , \5484 , \5485 );
nand \U$5240 ( \5487 , \2691 , \5486 );
nand \U$5241 ( \5488 , \5483 , \5487 );
xor \U$5242 ( \5489 , \5480 , \5488 );
xor \U$5243 ( \5490 , \5468 , \5489 );
xor \U$5244 ( \5491 , \5456 , \5490 );
xnor \U$5245 ( \5492 , \5431 , \5491 );
not \U$5246 ( \5493 , \5361 );
not \U$5247 ( \5494 , \5325 );
or \U$5248 ( \5495 , \5493 , \5494 );
nand \U$5249 ( \5496 , \5321 , \5289 );
nand \U$5250 ( \5497 , \5495 , \5496 );
not \U$5251 ( \5498 , \5497 );
not \U$5252 ( \5499 , \5498 );
not \U$5253 ( \5500 , \5272 );
not \U$5254 ( \5501 , \5124 );
or \U$5255 ( \5502 , \5500 , \5501 );
nand \U$5256 ( \5503 , \5207 , \5271 );
nand \U$5257 ( \5504 , \5502 , \5503 );
not \U$5258 ( \5505 , \5313 );
not \U$5259 ( \5506 , \5505 );
not \U$5260 ( \5507 , \5309 );
not \U$5261 ( \5508 , \5507 );
not \U$5262 ( \5509 , \5319 );
or \U$5263 ( \5510 , \5508 , \5509 );
or \U$5264 ( \5511 , \5319 , \5507 );
nand \U$5265 ( \5512 , \5510 , \5511 );
not \U$5266 ( \5513 , \5512 );
or \U$5267 ( \5514 , \5506 , \5513 );
nand \U$5268 ( \5515 , \5319 , \5309 );
nand \U$5269 ( \5516 , \5514 , \5515 );
not \U$5270 ( \5517 , \5516 );
not \U$5271 ( \5518 , \5147 );
not \U$5272 ( \5519 , \5206 );
or \U$5273 ( \5520 , \5518 , \5519 );
not \U$5274 ( \5521 , \5202 );
nand \U$5275 ( \5522 , \5521 , \5167 );
nand \U$5276 ( \5523 , \5520 , \5522 );
not \U$5277 ( \5524 , \5523 );
and \U$5278 ( \5525 , RIbe27b98_2, RIbe27df0_7);
not \U$5279 ( \5526 , \5525 );
not \U$5280 ( \5527 , \5170 );
not \U$5281 ( \5528 , \5527 );
not \U$5282 ( \5529 , \282 );
or \U$5283 ( \5530 , \5528 , \5529 );
not \U$5284 ( \5531 , RIbe29038_46);
not \U$5285 ( \5532 , RIbe294e8_56);
and \U$5286 ( \5533 , \5531 , \5532 );
and \U$5287 ( \5534 , RIbe29038_46, RIbe294e8_56);
nor \U$5288 ( \5535 , \5533 , \5534 );
nand \U$5289 ( \5536 , \287 , \5535 );
nand \U$5290 ( \5537 , \5530 , \5536 );
not \U$5291 ( \5538 , \5537 );
not \U$5292 ( \5539 , \5538 );
or \U$5293 ( \5540 , \5526 , \5539 );
not \U$5294 ( \5541 , \5525 );
nand \U$5295 ( \5542 , \5541 , \5537 );
nand \U$5296 ( \5543 , \5540 , \5542 );
nand \U$5297 ( \5544 , \361 , \5144 );
or \U$5298 ( \5545 , \363 , RIbe295d8_58);
or \U$5299 ( \5546 , \2995 , RIbe27c10_3);
nand \U$5300 ( \5547 , \5545 , \5546 );
nand \U$5301 ( \5548 , \1174 , \5547 );
and \U$5302 ( \5549 , \5544 , \5548 );
xor \U$5303 ( \5550 , \5543 , \5549 );
not \U$5304 ( \5551 , \5550 );
not \U$5305 ( \5552 , \5551 );
not \U$5306 ( \5553 , \5221 );
not \U$5307 ( \5554 , \2639 );
or \U$5308 ( \5555 , \5553 , \5554 );
not \U$5309 ( \5556 , RIbe28048_12);
not \U$5310 ( \5557 , RIbe28390_19);
and \U$5311 ( \5558 , \5556 , \5557 );
and \U$5312 ( \5559 , RIbe28048_12, RIbe28390_19);
nor \U$5313 ( \5560 , \5558 , \5559 );
nand \U$5314 ( \5561 , \3714 , \5560 );
nand \U$5315 ( \5562 , \5555 , \5561 );
not \U$5316 ( \5563 , \5156 );
not \U$5317 ( \5564 , \1164 );
or \U$5318 ( \5565 , \5563 , \5564 );
xor \U$5319 ( \5566 , RIbe27d78_6, RIbe297b8_62);
nand \U$5320 ( \5567 , \315 , \5566 );
nand \U$5321 ( \5568 , \5565 , \5567 );
xor \U$5322 ( \5569 , \5562 , \5568 );
and \U$5323 ( \5570 , RIbe284f8_22, RIbe28930_31);
nor \U$5324 ( \5571 , RIbe284f8_22, RIbe28930_31);
nor \U$5325 ( \5572 , \5570 , \5571 );
and \U$5326 ( \5573 , \971 , \5572 );
not \U$5327 ( \5574 , \1793 );
nor \U$5328 ( \5575 , \5574 , \5182 );
nor \U$5329 ( \5576 , \5573 , \5575 );
not \U$5330 ( \5577 , \5576 );
and \U$5331 ( \5578 , \5569 , \5577 );
not \U$5332 ( \5579 , \5569 );
and \U$5333 ( \5580 , \5579 , \5576 );
nor \U$5334 ( \5581 , \5578 , \5580 );
not \U$5335 ( \5582 , \5581 );
not \U$5336 ( \5583 , \5582 );
or \U$5337 ( \5584 , \5552 , \5583 );
nand \U$5338 ( \5585 , \5550 , \5581 );
nand \U$5339 ( \5586 , \5584 , \5585 );
not \U$5340 ( \5587 , \5253 );
not \U$5341 ( \5588 , \925 );
or \U$5342 ( \5589 , \5587 , \5588 );
and \U$5343 ( \5590 , RIbe28de0_41, RIbe29128_48);
not \U$5344 ( \5591 , RIbe28de0_41);
not \U$5345 ( \5592 , RIbe29128_48);
and \U$5346 ( \5593 , \5591 , \5592 );
nor \U$5347 ( \5594 , \5590 , \5593 );
nand \U$5348 ( \5595 , \514 , \5594 );
nand \U$5349 ( \5596 , \5589 , \5595 );
not \U$5350 ( \5597 , \3056 );
or \U$5351 ( \5598 , \5597 , \5212 );
xnor \U$5352 ( \5599 , RIbe28228_16, RIbe28c78_38);
or \U$5353 ( \5600 , \886 , \5599 );
nand \U$5354 ( \5601 , \5598 , \5600 );
xor \U$5355 ( \5602 , \5596 , \5601 );
or \U$5356 ( \5603 , \1566 , \5164 );
and \U$5357 ( \5604 , RIbe27b98_2, RIbe29a10_67);
not \U$5358 ( \5605 , RIbe27b98_2);
and \U$5359 ( \5606 , \5605 , \2420 );
nor \U$5360 ( \5607 , \5604 , \5606 );
not \U$5361 ( \5608 , \5607 );
or \U$5362 ( \5609 , \542 , \5608 );
nand \U$5363 ( \5610 , \5603 , \5609 );
xor \U$5364 ( \5611 , \5602 , \5610 );
xnor \U$5365 ( \5612 , \5586 , \5611 );
not \U$5366 ( \5613 , \5612 );
and \U$5367 ( \5614 , \5524 , \5613 );
and \U$5368 ( \5615 , \5612 , \5523 );
nor \U$5369 ( \5616 , \5614 , \5615 );
not \U$5370 ( \5617 , \5616 );
and \U$5371 ( \5618 , \5517 , \5617 );
and \U$5372 ( \5619 , \5516 , \5616 );
nor \U$5373 ( \5620 , \5618 , \5619 );
xnor \U$5374 ( \5621 , \5504 , \5620 );
not \U$5375 ( \5622 , \5621 );
and \U$5376 ( \5623 , \5499 , \5622 );
and \U$5377 ( \5624 , \5621 , \5498 );
nor \U$5378 ( \5625 , \5623 , \5624 );
xor \U$5379 ( \5626 , \5492 , \5625 );
not \U$5380 ( \5627 , \5278 );
not \U$5381 ( \5628 , \5627 );
not \U$5382 ( \5629 , \5273 );
and \U$5383 ( \5630 , \5628 , \5629 );
and \U$5384 ( \5631 , \5282 , \5119 );
nor \U$5385 ( \5632 , \5630 , \5631 );
xor \U$5386 ( \5633 , \5626 , \5632 );
nand \U$5387 ( \5634 , \5382 , \5633 );
or \U$5388 ( \5635 , \5488 , \5479 );
nand \U$5389 ( \5636 , \5635 , \5475 );
nand \U$5390 ( \5637 , \5488 , \5479 );
and \U$5391 ( \5638 , \5636 , \5637 );
not \U$5392 ( \5639 , \5537 );
not \U$5393 ( \5640 , \5525 );
or \U$5394 ( \5641 , \5639 , \5640 );
not \U$5395 ( \5642 , \5544 );
not \U$5396 ( \5643 , \5548 );
or \U$5397 ( \5644 , \5642 , \5643 );
nand \U$5398 ( \5645 , \5644 , \5543 );
nand \U$5399 ( \5646 , \5641 , \5645 );
and \U$5400 ( \5647 , \5646 , \5415 );
not \U$5401 ( \5648 , \5646 );
and \U$5402 ( \5649 , \5648 , \5412 );
or \U$5403 ( \5650 , \5647 , \5649 );
xnor \U$5404 ( \5651 , \5638 , \5650 );
not \U$5405 ( \5652 , \5611 );
not \U$5406 ( \5653 , \5586 );
or \U$5407 ( \5654 , \5652 , \5653 );
not \U$5408 ( \5655 , \5582 );
nand \U$5409 ( \5656 , \5655 , \5551 );
nand \U$5410 ( \5657 , \5654 , \5656 );
xor \U$5411 ( \5658 , \5651 , \5657 );
xor \U$5412 ( \5659 , \5596 , \5601 );
and \U$5413 ( \5660 , \5659 , \5610 );
and \U$5414 ( \5661 , \5596 , \5601 );
or \U$5415 ( \5662 , \5660 , \5661 );
not \U$5416 ( \5663 , \5568 );
not \U$5417 ( \5664 , \5562 );
or \U$5418 ( \5665 , \5663 , \5664 );
nand \U$5419 ( \5666 , \5569 , \5577 );
nand \U$5420 ( \5667 , \5665 , \5666 );
xor \U$5421 ( \5668 , \5662 , \5667 );
not \U$5422 ( \5669 , \5599 );
not \U$5423 ( \5670 , \5669 );
not \U$5424 ( \5671 , \3056 );
or \U$5425 ( \5672 , \5670 , \5671 );
and \U$5426 ( \5673 , RIbe28228_16, RIbe28318_18);
not \U$5427 ( \5674 , RIbe28228_16);
and \U$5428 ( \5675 , \5674 , \2244 );
nor \U$5429 ( \5676 , \5673 , \5675 );
nand \U$5430 ( \5677 , \885 , \5676 );
nand \U$5431 ( \5678 , \5672 , \5677 );
not \U$5432 ( \5679 , \5607 );
not \U$5433 ( \5680 , \256 );
or \U$5434 ( \5681 , \5679 , \5680 );
xnor \U$5435 ( \5682 , RIbe29b00_69, RIbe27b98_2);
not \U$5436 ( \5683 , \5682 );
nand \U$5437 ( \5684 , \5683 , \1734 );
nand \U$5438 ( \5685 , \5681 , \5684 );
xor \U$5439 ( \5686 , \5678 , \5685 );
not \U$5440 ( \5687 , \1131 );
not \U$5441 ( \5688 , \5391 );
and \U$5442 ( \5689 , \5687 , \5688 );
and \U$5443 ( \5690 , RIbe293f8_54, RIbe296c8_60);
nor \U$5444 ( \5691 , RIbe293f8_54, RIbe296c8_60);
nor \U$5445 ( \5692 , \5690 , \5691 );
and \U$5446 ( \5693 , \1137 , \5692 );
nor \U$5447 ( \5694 , \5689 , \5693 );
not \U$5448 ( \5695 , \5694 );
and \U$5449 ( \5696 , \5686 , \5695 );
not \U$5450 ( \5697 , \5686 );
and \U$5451 ( \5698 , \5697 , \5694 );
nor \U$5452 ( \5699 , \5696 , \5698 );
xor \U$5453 ( \5700 , \5668 , \5699 );
xor \U$5454 ( \5701 , \5658 , \5700 );
or \U$5455 ( \5702 , \5386 , \5418 );
or \U$5456 ( \5703 , \5388 , \5417 );
nand \U$5457 ( \5704 , \5702 , \5703 );
and \U$5458 ( \5705 , \5456 , \5490 );
and \U$5459 ( \5706 , \5438 , \5455 );
nor \U$5460 ( \5707 , \5705 , \5706 );
xnor \U$5461 ( \5708 , \5704 , \5707 );
xnor \U$5462 ( \5709 , \5701 , \5708 );
not \U$5463 ( \5710 , \5709 );
not \U$5464 ( \5711 , \5621 );
not \U$5465 ( \5712 , \5497 );
or \U$5466 ( \5713 , \5711 , \5712 );
not \U$5467 ( \5714 , \5620 );
nand \U$5468 ( \5715 , \5714 , \5504 );
nand \U$5469 ( \5716 , \5713 , \5715 );
not \U$5470 ( \5717 , \5716 );
or \U$5471 ( \5718 , \5710 , \5717 );
or \U$5472 ( \5719 , \5709 , \5716 );
nand \U$5473 ( \5720 , \5718 , \5719 );
xor \U$5474 ( \5721 , \5462 , \5467 );
and \U$5475 ( \5722 , \5721 , \5489 );
and \U$5476 ( \5723 , \5462 , \5467 );
nor \U$5477 ( \5724 , \5722 , \5723 );
not \U$5478 ( \5725 , \5724 );
not \U$5479 ( \5726 , \5442 );
not \U$5480 ( \5727 , \5726 );
not \U$5481 ( \5728 , \5451 );
or \U$5482 ( \5729 , \5727 , \5728 );
not \U$5483 ( \5730 , \5450 );
nand \U$5484 ( \5731 , \5730 , \5447 );
nand \U$5485 ( \5732 , \5729 , \5731 );
not \U$5486 ( \5733 , \5732 );
nand \U$5487 ( \5734 , \5408 , \5415 );
not \U$5488 ( \5735 , \5394 );
nand \U$5489 ( \5736 , \5735 , \5404 );
and \U$5490 ( \5737 , \5734 , \5736 );
not \U$5491 ( \5738 , \5566 );
not \U$5492 ( \5739 , \1042 );
not \U$5493 ( \5740 , \5739 );
or \U$5494 ( \5741 , \5738 , \5740 );
xor \U$5495 ( \5742 , RIbe27d78_6, RIbe28138_14);
nand \U$5496 ( \5743 , \314 , \5742 );
nand \U$5497 ( \5744 , \5741 , \5743 );
not \U$5498 ( \5745 , \5535 );
not \U$5499 ( \5746 , \282 );
or \U$5500 ( \5747 , \5745 , \5746 );
not \U$5501 ( \5748 , RIbe288b8_30);
not \U$5502 ( \5749 , RIbe29038_46);
and \U$5503 ( \5750 , \5748 , \5749 );
and \U$5504 ( \5751 , RIbe288b8_30, RIbe29038_46);
nor \U$5505 ( \5752 , \5750 , \5751 );
nand \U$5506 ( \5753 , \1583 , \5752 );
nand \U$5507 ( \5754 , \5747 , \5753 );
xor \U$5508 ( \5755 , \5744 , \5754 );
and \U$5509 ( \5756 , \1793 , \5572 );
and \U$5510 ( \5757 , RIbe28750_27, RIbe28930_31);
not \U$5511 ( \5758 , RIbe28750_27);
and \U$5512 ( \5759 , \5758 , \973 );
nor \U$5513 ( \5760 , \5757 , \5759 );
and \U$5514 ( \5761 , \971 , \5760 );
nor \U$5515 ( \5762 , \5756 , \5761 );
and \U$5516 ( \5763 , \5755 , \5762 );
not \U$5517 ( \5764 , \5755 );
not \U$5518 ( \5765 , \5762 );
and \U$5519 ( \5766 , \5764 , \5765 );
nor \U$5520 ( \5767 , \5763 , \5766 );
and \U$5521 ( \5768 , \5737 , \5767 );
not \U$5522 ( \5769 , \5737 );
not \U$5523 ( \5770 , \5767 );
and \U$5524 ( \5771 , \5769 , \5770 );
nor \U$5525 ( \5772 , \5768 , \5771 );
not \U$5526 ( \5773 , \5772 );
and \U$5527 ( \5774 , \5733 , \5773 );
not \U$5528 ( \5775 , \5733 );
and \U$5529 ( \5776 , \5775 , \5772 );
nor \U$5530 ( \5777 , \5774 , \5776 );
not \U$5531 ( \5778 , \5777 );
or \U$5532 ( \5779 , \5725 , \5778 );
or \U$5533 ( \5780 , \5724 , \5777 );
nand \U$5534 ( \5781 , \5779 , \5780 );
not \U$5535 ( \5782 , \5402 );
not \U$5536 ( \5783 , \2276 );
or \U$5537 ( \5784 , \5782 , \5783 );
xnor \U$5538 ( \5785 , RIbe28a20_33, RIbe28570_23);
not \U$5539 ( \5786 , \5785 );
nand \U$5540 ( \5787 , \5786 , \2476 );
nand \U$5541 ( \5788 , \5784 , \5787 );
not \U$5542 ( \5789 , \5547 );
not \U$5543 ( \5790 , \361 );
or \U$5544 ( \5791 , \5789 , \5790 );
not \U$5545 ( \5792 , RIbe27c10_3);
not \U$5546 ( \5793 , RIbe29740_61);
and \U$5547 ( \5794 , \5792 , \5793 );
and \U$5548 ( \5795 , RIbe27c10_3, RIbe29740_61);
nor \U$5549 ( \5796 , \5794 , \5795 );
nand \U$5550 ( \5797 , \1174 , \5796 );
nand \U$5551 ( \5798 , \5791 , \5797 );
xor \U$5552 ( \5799 , \5788 , \5798 );
or \U$5553 ( \5800 , \524 , \5473 );
and \U$5554 ( \5801 , RIbe290b0_47, \919 );
not \U$5555 ( \5802 , RIbe290b0_47);
and \U$5556 ( \5803 , \5802 , RIbe29470_55);
nor \U$5557 ( \5804 , \5801 , \5803 );
or \U$5558 ( \5805 , \5470 , \5804 );
nand \U$5559 ( \5806 , \5800 , \5805 );
xor \U$5560 ( \5807 , \5799 , \5806 );
not \U$5561 ( \5808 , \5807 );
not \U$5562 ( \5809 , \5486 );
not \U$5563 ( \5810 , \2702 );
or \U$5564 ( \5811 , \5809 , \5810 );
and \U$5565 ( \5812 , RIbe28b88_36, RIbe27ee0_9);
not \U$5566 ( \5813 , RIbe28b88_36);
and \U$5567 ( \5814 , \5813 , \317 );
nor \U$5568 ( \5815 , \5812 , \5814 );
nand \U$5569 ( \5816 , \2560 , \5815 );
nand \U$5570 ( \5817 , \5811 , \5816 );
not \U$5571 ( \5818 , \1265 );
not \U$5572 ( \5819 , RIbe280c0_13);
not \U$5573 ( \5820 , RIbe28c00_37);
and \U$5574 ( \5821 , \5819 , \5820 );
and \U$5575 ( \5822 , RIbe280c0_13, RIbe28c00_37);
nor \U$5576 ( \5823 , \5821 , \5822 );
not \U$5577 ( \5824 , \5823 );
or \U$5578 ( \5825 , \5818 , \5824 );
not \U$5579 ( \5826 , \5477 );
nand \U$5580 ( \5827 , \5826 , \862 );
nand \U$5581 ( \5828 , \5825 , \5827 );
xor \U$5582 ( \5829 , \5817 , \5828 );
and \U$5583 ( \5830 , \2640 , \5560 );
buf \U$5584 ( \5831 , \3714 );
and \U$5585 ( \5832 , RIbe28390_19, RIbe29380_53);
nor \U$5586 ( \5833 , RIbe28390_19, RIbe29380_53);
nor \U$5587 ( \5834 , \5832 , \5833 );
and \U$5588 ( \5835 , \5831 , \5834 );
nor \U$5589 ( \5836 , \5830 , \5835 );
not \U$5590 ( \5837 , \5836 );
and \U$5591 ( \5838 , \5829 , \5837 );
not \U$5592 ( \5839 , \5829 );
and \U$5593 ( \5840 , \5839 , \5836 );
nor \U$5594 ( \5841 , \5838 , \5840 );
nand \U$5595 ( \5842 , RIbe27b98_2, RIbe29218_50);
not \U$5596 ( \5843 , \5594 );
not \U$5597 ( \5844 , \925 );
or \U$5598 ( \5845 , \5843 , \5844 );
xor \U$5599 ( \5846 , RIbe291a0_49, RIbe28de0_41);
nand \U$5600 ( \5847 , \514 , \5846 );
nand \U$5601 ( \5848 , \5845 , \5847 );
xor \U$5602 ( \5849 , \5842 , \5848 );
not \U$5603 ( \5850 , \2672 );
not \U$5604 ( \5851 , \3484 );
or \U$5605 ( \5852 , \5850 , \5851 );
nand \U$5606 ( \5853 , \5852 , RIbe28480_21);
xnor \U$5607 ( \5854 , \5849 , \5853 );
and \U$5608 ( \5855 , \5841 , \5854 );
not \U$5609 ( \5856 , \5841 );
not \U$5610 ( \5857 , \5854 );
and \U$5611 ( \5858 , \5856 , \5857 );
or \U$5612 ( \5859 , \5855 , \5858 );
not \U$5613 ( \5860 , \5859 );
or \U$5614 ( \5861 , \5808 , \5860 );
or \U$5615 ( \5862 , \5859 , \5807 );
nand \U$5616 ( \5863 , \5861 , \5862 );
not \U$5617 ( \5864 , \5863 );
and \U$5618 ( \5865 , \5781 , \5864 );
not \U$5619 ( \5866 , \5781 );
and \U$5620 ( \5867 , \5866 , \5863 );
nor \U$5621 ( \5868 , \5865 , \5867 );
not \U$5622 ( \5869 , \5868 );
not \U$5623 ( \5870 , \5869 );
not \U$5624 ( \5871 , \5616 );
not \U$5625 ( \5872 , \5871 );
not \U$5626 ( \5873 , \5516 );
or \U$5627 ( \5874 , \5872 , \5873 );
not \U$5628 ( \5875 , \5612 );
nand \U$5629 ( \5876 , \5875 , \5523 );
nand \U$5630 ( \5877 , \5874 , \5876 );
not \U$5631 ( \5878 , \5877 );
not \U$5632 ( \5879 , \5878 );
or \U$5633 ( \5880 , \5870 , \5879 );
nand \U$5634 ( \5881 , \5877 , \5868 );
nand \U$5635 ( \5882 , \5880 , \5881 );
not \U$5636 ( \5883 , \5491 );
not \U$5637 ( \5884 , \5431 );
or \U$5638 ( \5885 , \5883 , \5884 );
not \U$5639 ( \5886 , \5419 );
nand \U$5640 ( \5887 , \5886 , \5427 );
nand \U$5641 ( \5888 , \5885 , \5887 );
xor \U$5642 ( \5889 , \5882 , \5888 );
not \U$5643 ( \5890 , \5889 );
and \U$5644 ( \5891 , \5720 , \5890 );
not \U$5645 ( \5892 , \5720 );
and \U$5646 ( \5893 , \5892 , \5889 );
nor \U$5647 ( \5894 , \5891 , \5893 );
xor \U$5648 ( \5895 , \5492 , \5625 );
and \U$5649 ( \5896 , \5895 , \5632 );
and \U$5650 ( \5897 , \5492 , \5625 );
or \U$5651 ( \5898 , \5896 , \5897 );
nand \U$5652 ( \5899 , \5894 , \5898 );
and \U$5653 ( \5900 , \5634 , \5899 );
and \U$5654 ( \5901 , \5668 , \5699 );
and \U$5655 ( \5902 , \5662 , \5667 );
nor \U$5656 ( \5903 , \5901 , \5902 );
not \U$5657 ( \5904 , \5903 );
and \U$5658 ( \5905 , \282 , \5752 );
and \U$5659 ( \5906 , \290 , \940 );
and \U$5660 ( \5907 , RIbe28a98_34, RIbe29038_46);
nor \U$5661 ( \5908 , \5906 , \5907 );
and \U$5662 ( \5909 , \287 , \5908 );
nor \U$5663 ( \5910 , \5905 , \5909 );
nand \U$5664 ( \5911 , RIbe27b98_2, RIbe29a10_67);
not \U$5665 ( \5912 , \5911 );
not \U$5666 ( \5913 , \5804 );
not \U$5667 ( \5914 , \5913 );
not \U$5668 ( \5915 , \466 );
or \U$5669 ( \5916 , \5914 , \5915 );
xor \U$5670 ( \5917 , RIbe290b0_47, RIbe294e8_56);
nand \U$5671 ( \5918 , \2071 , \5917 );
nand \U$5672 ( \5919 , \5916 , \5918 );
not \U$5673 ( \5920 , \5919 );
or \U$5674 ( \5921 , \5912 , \5920 );
or \U$5675 ( \5922 , \5919 , \5911 );
nand \U$5676 ( \5923 , \5921 , \5922 );
xnor \U$5677 ( \5924 , \5910 , \5923 );
and \U$5678 ( \5925 , \2640 , \5834 );
and \U$5679 ( \5926 , \2777 , RIbe28390_19);
nor \U$5680 ( \5927 , \5925 , \5926 );
not \U$5681 ( \5928 , \5927 );
not \U$5682 ( \5929 , \5742 );
not \U$5683 ( \5930 , \1164 );
or \U$5684 ( \5931 , \5929 , \5930 );
xor \U$5685 ( \5932 , RIbe27d78_6, RIbe282a0_17);
nand \U$5686 ( \5933 , \315 , \5932 );
nand \U$5687 ( \5934 , \5931 , \5933 );
not \U$5688 ( \5935 , \5692 );
not \U$5689 ( \5936 , \1452 );
or \U$5690 ( \5937 , \5935 , \5936 );
xnor \U$5691 ( \5938 , RIbe29308_52, RIbe296c8_60);
not \U$5692 ( \5939 , \5938 );
nand \U$5693 ( \5940 , \5939 , \1137 );
nand \U$5694 ( \5941 , \5937 , \5940 );
xor \U$5695 ( \5942 , \5934 , \5941 );
not \U$5696 ( \5943 , \5942 );
or \U$5697 ( \5944 , \5928 , \5943 );
or \U$5698 ( \5945 , \5942 , \5927 );
nand \U$5699 ( \5946 , \5944 , \5945 );
not \U$5700 ( \5947 , \5946 );
not \U$5701 ( \5948 , \5842 );
or \U$5702 ( \5949 , \5848 , \5948 );
nand \U$5703 ( \5950 , \5949 , \5853 );
nand \U$5704 ( \5951 , \5848 , \5948 );
and \U$5705 ( \5952 , \5950 , \5951 );
not \U$5706 ( \5953 , \5952 );
and \U$5707 ( \5954 , \5947 , \5953 );
and \U$5708 ( \5955 , \5946 , \5952 );
nor \U$5709 ( \5956 , \5954 , \5955 );
and \U$5710 ( \5957 , \5924 , \5956 );
not \U$5711 ( \5958 , \5924 );
not \U$5712 ( \5959 , \5956 );
and \U$5713 ( \5960 , \5958 , \5959 );
or \U$5714 ( \5961 , \5957 , \5960 );
not \U$5715 ( \5962 , \5961 );
or \U$5716 ( \5963 , \5904 , \5962 );
or \U$5717 ( \5964 , \5961 , \5903 );
nand \U$5718 ( \5965 , \5963 , \5964 );
not \U$5719 ( \5966 , \5965 );
not \U$5720 ( \5967 , \5638 );
not \U$5721 ( \5968 , \5967 );
not \U$5722 ( \5969 , \5650 );
or \U$5723 ( \5970 , \5968 , \5969 );
nand \U$5724 ( \5971 , \5646 , \5412 );
nand \U$5725 ( \5972 , \5970 , \5971 );
or \U$5726 ( \5973 , \1566 , \5682 );
or \U$5727 ( \5974 , RIbe27b98_2, RIbe29128_48);
nand \U$5728 ( \5975 , RIbe27b98_2, RIbe29128_48);
nand \U$5729 ( \5976 , \5974 , \5975 );
not \U$5730 ( \5977 , \5976 );
nand \U$5731 ( \5978 , \5977 , \1734 );
nand \U$5732 ( \5979 , \5973 , \5978 );
not \U$5733 ( \5980 , \5979 );
not \U$5734 ( \5981 , \1770 );
xnor \U$5735 ( \5982 , RIbe286d8_26, RIbe28a20_33);
not \U$5736 ( \5983 , \5982 );
and \U$5737 ( \5984 , \5981 , \5983 );
not \U$5738 ( \5985 , \2276 );
nor \U$5739 ( \5986 , \5985 , \5785 );
nor \U$5740 ( \5987 , \5984 , \5986 );
not \U$5741 ( \5988 , \5987 );
or \U$5742 ( \5989 , \5980 , \5988 );
or \U$5743 ( \5990 , \5987 , \5979 );
nand \U$5744 ( \5991 , \5989 , \5990 );
not \U$5745 ( \5992 , \5991 );
nand \U$5746 ( \5993 , \1793 , \5760 );
and \U$5747 ( \5994 , RIbe28930_31, \364 );
not \U$5748 ( \5995 , RIbe28930_31);
and \U$5749 ( \5996 , \5995 , RIbe28840_29);
nor \U$5750 ( \5997 , \5994 , \5996 );
not \U$5751 ( \5998 , \5997 );
nand \U$5752 ( \5999 , \5998 , \1797 );
and \U$5753 ( \6000 , \5993 , \5999 );
not \U$5754 ( \6001 , \6000 );
and \U$5755 ( \6002 , \5992 , \6001 );
and \U$5756 ( \6003 , \5991 , \6000 );
nor \U$5757 ( \6004 , \6002 , \6003 );
not \U$5758 ( \6005 , \5676 );
not \U$5759 ( \6006 , \1061 );
or \U$5760 ( \6007 , \6005 , \6006 );
xnor \U$5761 ( \6008 , RIbe284f8_22, RIbe28228_16);
not \U$5762 ( \6009 , \6008 );
nand \U$5763 ( \6010 , \6009 , \885 );
nand \U$5764 ( \6011 , \6007 , \6010 );
not \U$5765 ( \6012 , \1148 );
xnor \U$5766 ( \6013 , RIbe28de0_41, RIbe295d8_58);
not \U$5767 ( \6014 , \6013 );
and \U$5768 ( \6015 , \6012 , \6014 );
and \U$5769 ( \6016 , \1145 , \5846 );
nor \U$5770 ( \6017 , \6015 , \6016 );
xnor \U$5771 ( \6018 , \6011 , \6017 );
and \U$5772 ( \6019 , \936 , \5796 );
not \U$5773 ( \6020 , RIbe27c10_3);
not \U$5774 ( \6021 , RIbe297b8_62);
and \U$5775 ( \6022 , \6020 , \6021 );
and \U$5776 ( \6023 , RIbe27c10_3, RIbe297b8_62);
nor \U$5777 ( \6024 , \6022 , \6023 );
and \U$5778 ( \6025 , \1498 , \6024 );
nor \U$5779 ( \6026 , \6019 , \6025 );
not \U$5780 ( \6027 , \6026 );
and \U$5781 ( \6028 , \6018 , \6027 );
not \U$5782 ( \6029 , \6018 );
and \U$5783 ( \6030 , \6029 , \6026 );
nor \U$5784 ( \6031 , \6028 , \6030 );
and \U$5785 ( \6032 , \6004 , \6031 );
not \U$5786 ( \6033 , \6004 );
not \U$5787 ( \6034 , \6031 );
and \U$5788 ( \6035 , \6033 , \6034 );
nor \U$5789 ( \6036 , \6032 , \6035 );
xor \U$5790 ( \6037 , \5972 , \6036 );
not \U$5791 ( \6038 , \6037 );
and \U$5792 ( \6039 , \5966 , \6038 );
and \U$5793 ( \6040 , \5965 , \6037 );
nor \U$5794 ( \6041 , \6039 , \6040 );
not \U$5795 ( \6042 , \5863 );
not \U$5796 ( \6043 , \5781 );
or \U$5797 ( \6044 , \6042 , \6043 );
not \U$5798 ( \6045 , \5724 );
nand \U$5799 ( \6046 , \6045 , \5777 );
nand \U$5800 ( \6047 , \6044 , \6046 );
xnor \U$5801 ( \6048 , \6041 , \6047 );
not \U$5802 ( \6049 , \5701 );
not \U$5803 ( \6050 , \5708 );
or \U$5804 ( \6051 , \6049 , \6050 );
not \U$5805 ( \6052 , \5707 );
nand \U$5806 ( \6053 , \6052 , \5704 );
nand \U$5807 ( \6054 , \6051 , \6053 );
not \U$5808 ( \6055 , \6054 );
and \U$5809 ( \6056 , \6048 , \6055 );
not \U$5810 ( \6057 , \6048 );
and \U$5811 ( \6058 , \6057 , \6054 );
nor \U$5812 ( \6059 , \6056 , \6058 );
not \U$5813 ( \6060 , \6059 );
not \U$5814 ( \6061 , \5700 );
not \U$5815 ( \6062 , \5658 );
or \U$5816 ( \6063 , \6061 , \6062 );
nand \U$5817 ( \6064 , \5651 , \5657 );
nand \U$5818 ( \6065 , \6063 , \6064 );
not \U$5819 ( \6066 , \6065 );
not \U$5820 ( \6067 , \5737 );
not \U$5821 ( \6068 , \5767 );
and \U$5822 ( \6069 , \6067 , \6068 );
not \U$5823 ( \6070 , \5733 );
and \U$5824 ( \6071 , \6070 , \5772 );
nor \U$5825 ( \6072 , \6069 , \6071 );
not \U$5826 ( \6073 , \6072 );
and \U$5827 ( \6074 , \6066 , \6073 );
and \U$5828 ( \6075 , \6065 , \6072 );
nor \U$5829 ( \6076 , \6074 , \6075 );
not \U$5830 ( \6077 , \5854 );
not \U$5831 ( \6078 , \5807 );
or \U$5832 ( \6079 , \6077 , \6078 );
not \U$5833 ( \6080 , \5857 );
not \U$5834 ( \6081 , \5807 );
not \U$5835 ( \6082 , \6081 );
or \U$5836 ( \6083 , \6080 , \6082 );
nand \U$5837 ( \6084 , \6083 , \5841 );
nand \U$5838 ( \6085 , \6079 , \6084 );
not \U$5839 ( \6086 , \6085 );
not \U$5840 ( \6087 , \5837 );
not \U$5841 ( \6088 , \5829 );
or \U$5842 ( \6089 , \6087 , \6088 );
nand \U$5843 ( \6090 , \5817 , \5828 );
nand \U$5844 ( \6091 , \6089 , \6090 );
not \U$5845 ( \6092 , \6091 );
and \U$5846 ( \6093 , \1326 , \5823 );
not \U$5847 ( \6094 , RIbe280c0_13);
not \U$5848 ( \6095 , RIbe28c78_38);
and \U$5849 ( \6096 , \6094 , \6095 );
and \U$5850 ( \6097 , RIbe280c0_13, RIbe28c78_38);
nor \U$5851 ( \6098 , \6096 , \6097 );
and \U$5852 ( \6099 , \869 , \6098 );
nor \U$5853 ( \6100 , \6093 , \6099 );
not \U$5854 ( \6101 , \5815 );
not \U$5855 ( \6102 , \2702 );
or \U$5856 ( \6103 , \6101 , \6102 );
xor \U$5857 ( \6104 , RIbe28048_12, RIbe28b88_36);
nand \U$5858 ( \6105 , \6104 , \2561 );
nand \U$5859 ( \6106 , \6103 , \6105 );
and \U$5860 ( \6107 , \6100 , \6106 );
not \U$5861 ( \6108 , \6100 );
not \U$5862 ( \6109 , \6106 );
and \U$5863 ( \6110 , \6108 , \6109 );
or \U$5864 ( \6111 , \6107 , \6110 );
not \U$5865 ( \6112 , \6111 );
and \U$5866 ( \6113 , \6092 , \6112 );
and \U$5867 ( \6114 , \6091 , \6111 );
nor \U$5868 ( \6115 , \6113 , \6114 );
not \U$5869 ( \6116 , \6115 );
or \U$5870 ( \6117 , \6086 , \6116 );
or \U$5871 ( \6118 , \6085 , \6115 );
nand \U$5872 ( \6119 , \6117 , \6118 );
not \U$5873 ( \6120 , \6119 );
not \U$5874 ( \6121 , \6120 );
xor \U$5875 ( \6122 , \5788 , \5798 );
and \U$5876 ( \6123 , \6122 , \5806 );
and \U$5877 ( \6124 , \5788 , \5798 );
or \U$5878 ( \6125 , \6123 , \6124 );
not \U$5879 ( \6126 , \5678 );
not \U$5880 ( \6127 , \5685 );
or \U$5881 ( \6128 , \6126 , \6127 );
or \U$5882 ( \6129 , \5678 , \5685 );
nand \U$5883 ( \6130 , \6129 , \5695 );
nand \U$5884 ( \6131 , \6128 , \6130 );
xor \U$5885 ( \6132 , \6125 , \6131 );
not \U$5886 ( \6133 , \5765 );
not \U$5887 ( \6134 , \5755 );
or \U$5888 ( \6135 , \6133 , \6134 );
nand \U$5889 ( \6136 , \5754 , \5744 );
nand \U$5890 ( \6137 , \6135 , \6136 );
xor \U$5891 ( \6138 , \6132 , \6137 );
not \U$5892 ( \6139 , \6138 );
and \U$5893 ( \6140 , \6121 , \6139 );
and \U$5894 ( \6141 , \6120 , \6138 );
nor \U$5895 ( \6142 , \6140 , \6141 );
and \U$5896 ( \6143 , \6076 , \6142 );
not \U$5897 ( \6144 , \6076 );
not \U$5898 ( \6145 , \6142 );
and \U$5899 ( \6146 , \6144 , \6145 );
nor \U$5900 ( \6147 , \6143 , \6146 );
not \U$5901 ( \6148 , \5888 );
not \U$5902 ( \6149 , \5882 );
or \U$5903 ( \6150 , \6148 , \6149 );
nand \U$5904 ( \6151 , \5877 , \5869 );
nand \U$5905 ( \6152 , \6150 , \6151 );
xor \U$5906 ( \6153 , \6147 , \6152 );
not \U$5907 ( \6154 , \6153 );
or \U$5908 ( \6155 , \6060 , \6154 );
or \U$5909 ( \6156 , \6153 , \6059 );
nand \U$5910 ( \6157 , \6155 , \6156 );
not \U$5911 ( \6158 , \5889 );
not \U$5912 ( \6159 , \5720 );
or \U$5913 ( \6160 , \6158 , \6159 );
not \U$5914 ( \6161 , \5709 );
nand \U$5915 ( \6162 , \6161 , \5716 );
nand \U$5916 ( \6163 , \6160 , \6162 );
or \U$5917 ( \6164 , \6157 , \6163 );
not \U$5918 ( \6165 , \6059 );
not \U$5919 ( \6166 , \6165 );
not \U$5920 ( \6167 , \6153 );
or \U$5921 ( \6168 , \6166 , \6167 );
nand \U$5922 ( \6169 , \6152 , \6147 );
nand \U$5923 ( \6170 , \6168 , \6169 );
or \U$5924 ( \6171 , \6076 , \6142 );
not \U$5925 ( \6172 , \6065 );
or \U$5926 ( \6173 , \6172 , \6072 );
nand \U$5927 ( \6174 , \6171 , \6173 );
not \U$5928 ( \6175 , \6174 );
not \U$5929 ( \6176 , \6048 );
not \U$5930 ( \6177 , \6054 );
or \U$5931 ( \6178 , \6176 , \6177 );
not \U$5932 ( \6179 , \6041 );
nand \U$5933 ( \6180 , \6179 , \6047 );
nand \U$5934 ( \6181 , \6178 , \6180 );
not \U$5935 ( \6182 , \6181 );
not \U$5936 ( \6183 , \6182 );
or \U$5937 ( \6184 , \6175 , \6183 );
not \U$5938 ( \6185 , \6174 );
nand \U$5939 ( \6186 , \6185 , \6181 );
nand \U$5940 ( \6187 , \6184 , \6186 );
not \U$5941 ( \6188 , \6037 );
nand \U$5942 ( \6189 , \6188 , \5965 );
not \U$5943 ( \6190 , \5903 );
nand \U$5944 ( \6191 , \6190 , \5961 );
and \U$5945 ( \6192 , \6189 , \6191 );
not \U$5946 ( \6193 , \6192 );
or \U$5947 ( \6194 , \967 , \5997 );
xnor \U$5948 ( \6195 , RIbe28570_23, RIbe28930_31);
or \U$5949 ( \6196 , \1200 , \6195 );
nand \U$5950 ( \6197 , \6194 , \6196 );
or \U$5951 ( \6198 , \3750 , \5982 );
xnor \U$5952 ( \6199 , RIbe27ee0_9, RIbe28a20_33);
or \U$5953 ( \6200 , \1770 , \6199 );
nand \U$5954 ( \6201 , \6198 , \6200 );
xor \U$5955 ( \6202 , \6197 , \6201 );
and \U$5956 ( \6203 , RIbe29038_46, RIbe293f8_54);
not \U$5957 ( \6204 , RIbe29038_46);
and \U$5958 ( \6205 , \6204 , \2489 );
nor \U$5959 ( \6206 , \6203 , \6205 );
not \U$5960 ( \6207 , \6206 );
not \U$5961 ( \6208 , \287 );
or \U$5962 ( \6209 , \6207 , \6208 );
nand \U$5963 ( \6210 , \979 , \5908 );
nand \U$5964 ( \6211 , \6209 , \6210 );
xor \U$5965 ( \6212 , \6202 , \6211 );
or \U$5966 ( \6213 , \1835 , \6008 );
xor \U$5967 ( \6214 , RIbe28228_16, RIbe28750_27);
not \U$5968 ( \6215 , \6214 );
or \U$5969 ( \6216 , \886 , \6215 );
nand \U$5970 ( \6217 , \6213 , \6216 );
not \U$5971 ( \6218 , \6217 );
not \U$5972 ( \6219 , \2640 );
not \U$5973 ( \6220 , \5831 );
and \U$5974 ( \6221 , \6219 , \6220 );
nor \U$5975 ( \6222 , \6221 , \2779 );
not \U$5976 ( \6223 , \6222 );
or \U$5977 ( \6224 , \6218 , \6223 );
or \U$5978 ( \6225 , \6217 , \6222 );
nand \U$5979 ( \6226 , \6224 , \6225 );
not \U$5980 ( \6227 , \6226 );
not \U$5981 ( \6228 , \6109 );
and \U$5982 ( \6229 , \6227 , \6228 );
and \U$5983 ( \6230 , \6226 , \6109 );
nor \U$5984 ( \6231 , \6229 , \6230 );
not \U$5985 ( \6232 , \6231 );
not \U$5986 ( \6233 , RIbe28048_12);
not \U$5987 ( \6234 , RIbe28b88_36);
and \U$5988 ( \6235 , \6233 , \6234 );
and \U$5989 ( \6236 , RIbe28048_12, RIbe28b88_36);
nor \U$5990 ( \6237 , \6235 , \6236 );
and \U$5991 ( \6238 , \3402 , \6237 );
and \U$5992 ( \6239 , \3970 , \388 );
and \U$5993 ( \6240 , RIbe28b88_36, RIbe29380_53);
nor \U$5994 ( \6241 , \6239 , \6240 );
and \U$5995 ( \6242 , \2561 , \6241 );
nor \U$5996 ( \6243 , \6238 , \6242 );
not \U$5997 ( \6244 , \5917 );
not \U$5998 ( \6245 , \466 );
or \U$5999 ( \6246 , \6244 , \6245 );
xor \U$6000 ( \6247 , RIbe288b8_30, RIbe290b0_47);
nand \U$6001 ( \6248 , \399 , \6247 );
nand \U$6002 ( \6249 , \6246 , \6248 );
not \U$6003 ( \6250 , \6249 );
not \U$6004 ( \6251 , \6098 );
nor \U$6005 ( \6252 , \6251 , \863 );
and \U$6006 ( \6253 , RIbe280c0_13, RIbe28318_18);
nor \U$6007 ( \6254 , RIbe280c0_13, RIbe28318_18);
nor \U$6008 ( \6255 , \6253 , \6254 );
and \U$6009 ( \6256 , \869 , \6255 );
nor \U$6010 ( \6257 , \6252 , \6256 );
not \U$6011 ( \6258 , \6257 );
or \U$6012 ( \6259 , \6250 , \6258 );
or \U$6013 ( \6260 , \6257 , \6249 );
nand \U$6014 ( \6261 , \6259 , \6260 );
and \U$6015 ( \6262 , \6243 , \6261 );
not \U$6016 ( \6263 , \6243 );
not \U$6017 ( \6264 , \6261 );
and \U$6018 ( \6265 , \6263 , \6264 );
or \U$6019 ( \6266 , \6262 , \6265 );
not \U$6020 ( \6267 , \6266 );
or \U$6021 ( \6268 , \6232 , \6267 );
or \U$6022 ( \6269 , \6266 , \6231 );
nand \U$6023 ( \6270 , \6268 , \6269 );
xor \U$6024 ( \6271 , \6212 , \6270 );
not \U$6025 ( \6272 , \5924 );
not \U$6026 ( \6273 , \5959 );
or \U$6027 ( \6274 , \6272 , \6273 );
not \U$6028 ( \6275 , \5952 );
nand \U$6029 ( \6276 , \6275 , \5946 );
nand \U$6030 ( \6277 , \6274 , \6276 );
not \U$6031 ( \6278 , \6277 );
or \U$6032 ( \6279 , \2876 , \5938 );
and \U$6033 ( \6280 , RIbe296c8_60, \2479 );
not \U$6034 ( \6281 , RIbe296c8_60);
and \U$6035 ( \6282 , \6281 , RIbe28c00_37);
nor \U$6036 ( \6283 , \6280 , \6282 );
or \U$6037 ( \6284 , \1938 , \6283 );
nand \U$6038 ( \6285 , \6279 , \6284 );
nand \U$6039 ( \6286 , RIbe27b98_2, RIbe29b00_69);
not \U$6040 ( \6287 , \6286 );
not \U$6041 ( \6288 , \6013 );
not \U$6042 ( \6289 , \6288 );
not \U$6043 ( \6290 , \2857 );
or \U$6044 ( \6291 , \6289 , \6290 );
not \U$6045 ( \6292 , RIbe28de0_41);
not \U$6046 ( \6293 , RIbe29740_61);
and \U$6047 ( \6294 , \6292 , \6293 );
and \U$6048 ( \6295 , RIbe28de0_41, RIbe29740_61);
nor \U$6049 ( \6296 , \6294 , \6295 );
nand \U$6050 ( \6297 , \347 , \6296 );
nand \U$6051 ( \6298 , \6291 , \6297 );
not \U$6052 ( \6299 , \6298 );
or \U$6053 ( \6300 , \6287 , \6299 );
or \U$6054 ( \6301 , \6298 , \6286 );
nand \U$6055 ( \6302 , \6300 , \6301 );
xor \U$6056 ( \6303 , \6285 , \6302 );
not \U$6057 ( \6304 , \6303 );
not \U$6058 ( \6305 , \5987 );
not \U$6059 ( \6306 , \6305 );
not \U$6060 ( \6307 , \5979 );
or \U$6061 ( \6308 , \6306 , \6307 );
not \U$6062 ( \6309 , \6000 );
nand \U$6063 ( \6310 , \6309 , \5991 );
nand \U$6064 ( \6311 , \6308 , \6310 );
not \U$6065 ( \6312 , \6311 );
not \U$6066 ( \6313 , \6312 );
or \U$6067 ( \6314 , \6304 , \6313 );
not \U$6068 ( \6315 , \6303 );
nand \U$6069 ( \6316 , \6315 , \6311 );
nand \U$6070 ( \6317 , \6314 , \6316 );
not \U$6071 ( \6318 , \6317 );
not \U$6072 ( \6319 , \6024 );
not \U$6073 ( \6320 , \1493 );
or \U$6074 ( \6321 , \6319 , \6320 );
not \U$6075 ( \6322 , RIbe27c10_3);
not \U$6076 ( \6323 , RIbe28138_14);
and \U$6077 ( \6324 , \6322 , \6323 );
and \U$6078 ( \6325 , RIbe27c10_3, RIbe28138_14);
nor \U$6079 ( \6326 , \6324 , \6325 );
nand \U$6080 ( \6327 , \370 , \6326 );
nand \U$6081 ( \6328 , \6321 , \6327 );
not \U$6082 ( \6329 , \5932 );
not \U$6083 ( \6330 , \1086 );
or \U$6084 ( \6331 , \6329 , \6330 );
xnor \U$6085 ( \6332 , RIbe29470_55, RIbe27d78_6);
not \U$6086 ( \6333 , \6332 );
nand \U$6087 ( \6334 , \6333 , \315 );
nand \U$6088 ( \6335 , \6331 , \6334 );
xor \U$6089 ( \6336 , \6328 , \6335 );
or \U$6090 ( \6337 , \946 , \5976 );
or \U$6091 ( \6338 , RIbe27b98_2, RIbe291a0_49);
nand \U$6092 ( \6339 , RIbe27b98_2, RIbe291a0_49);
nand \U$6093 ( \6340 , \6338 , \6339 );
or \U$6094 ( \6341 , \1299 , \6340 );
nand \U$6095 ( \6342 , \6337 , \6341 );
xnor \U$6096 ( \6343 , \6336 , \6342 );
not \U$6097 ( \6344 , \6343 );
and \U$6098 ( \6345 , \6318 , \6344 );
and \U$6099 ( \6346 , \6317 , \6343 );
nor \U$6100 ( \6347 , \6345 , \6346 );
not \U$6101 ( \6348 , \6347 );
or \U$6102 ( \6349 , \6278 , \6348 );
or \U$6103 ( \6350 , \6277 , \6347 );
nand \U$6104 ( \6351 , \6349 , \6350 );
xor \U$6105 ( \6352 , \6271 , \6351 );
not \U$6106 ( \6353 , \6352 );
or \U$6107 ( \6354 , \6193 , \6353 );
or \U$6108 ( \6355 , \6352 , \6192 );
nand \U$6109 ( \6356 , \6354 , \6355 );
not \U$6110 ( \6357 , \5927 );
not \U$6111 ( \6358 , \6357 );
not \U$6112 ( \6359 , \5942 );
or \U$6113 ( \6360 , \6358 , \6359 );
nand \U$6114 ( \6361 , \5941 , \5934 );
nand \U$6115 ( \6362 , \6360 , \6361 );
not \U$6116 ( \6363 , \6027 );
not \U$6117 ( \6364 , \6018 );
or \U$6118 ( \6365 , \6363 , \6364 );
not \U$6119 ( \6366 , \6017 );
nand \U$6120 ( \6367 , \6366 , \6011 );
nand \U$6121 ( \6368 , \6365 , \6367 );
not \U$6122 ( \6369 , \6368 );
xnor \U$6123 ( \6370 , \6362 , \6369 );
not \U$6124 ( \6371 , \5911 );
not \U$6125 ( \6372 , \6371 );
not \U$6126 ( \6373 , \5919 );
or \U$6127 ( \6374 , \6372 , \6373 );
not \U$6128 ( \6375 , \5910 );
nand \U$6129 ( \6376 , \6375 , \5923 );
nand \U$6130 ( \6377 , \6374 , \6376 );
and \U$6131 ( \6378 , \6370 , \6377 );
not \U$6132 ( \6379 , \6370 );
not \U$6133 ( \6380 , \6377 );
and \U$6134 ( \6381 , \6379 , \6380 );
nor \U$6135 ( \6382 , \6378 , \6381 );
not \U$6136 ( \6383 , \6125 );
not \U$6137 ( \6384 , \6131 );
or \U$6138 ( \6385 , \6383 , \6384 );
or \U$6139 ( \6386 , \6125 , \6131 );
nand \U$6140 ( \6387 , \6386 , \6137 );
nand \U$6141 ( \6388 , \6385 , \6387 );
not \U$6142 ( \6389 , \6111 );
not \U$6143 ( \6390 , \6389 );
not \U$6144 ( \6391 , \6091 );
or \U$6145 ( \6392 , \6390 , \6391 );
not \U$6146 ( \6393 , \6100 );
nand \U$6147 ( \6394 , \6393 , \6109 );
nand \U$6148 ( \6395 , \6392 , \6394 );
xor \U$6149 ( \6396 , \6388 , \6395 );
xnor \U$6150 ( \6397 , \6382 , \6396 );
not \U$6151 ( \6398 , \5972 );
or \U$6152 ( \6399 , \6398 , \6036 );
or \U$6153 ( \6400 , \6004 , \6034 );
nand \U$6154 ( \6401 , \6399 , \6400 );
not \U$6155 ( \6402 , \6085 );
not \U$6156 ( \6403 , \6115 );
not \U$6157 ( \6404 , \6403 );
or \U$6158 ( \6405 , \6402 , \6404 );
nand \U$6159 ( \6406 , \6119 , \6138 );
nand \U$6160 ( \6407 , \6405 , \6406 );
xor \U$6161 ( \6408 , \6401 , \6407 );
xnor \U$6162 ( \6409 , \6397 , \6408 );
xor \U$6163 ( \6410 , \6356 , \6409 );
xor \U$6164 ( \6411 , \6187 , \6410 );
or \U$6165 ( \6412 , \6170 , \6411 );
nand \U$6166 ( \6413 , \5900 , \6164 , \6412 );
nor \U$6167 ( \6414 , \5369 , \5375 );
nor \U$6168 ( \6415 , \6413 , \6414 );
nand \U$6169 ( \6416 , \5379 , \6415 );
nand \U$6170 ( \6417 , \6163 , \6157 );
not \U$6171 ( \6418 , \6417 );
not \U$6172 ( \6419 , \5899 );
not \U$6173 ( \6420 , \5633 );
not \U$6174 ( \6421 , \5382 );
nand \U$6175 ( \6422 , \6420 , \6421 );
or \U$6176 ( \6423 , \6419 , \6422 );
or \U$6177 ( \6424 , \5894 , \5898 );
nand \U$6178 ( \6425 , \6423 , \6424 );
nand \U$6179 ( \6426 , \6425 , \6164 );
not \U$6180 ( \6427 , \6426 );
or \U$6181 ( \6428 , \6418 , \6427 );
nand \U$6182 ( \6429 , \6428 , \6412 );
nand \U$6183 ( \6430 , \6170 , \6411 );
nand \U$6184 ( \6431 , \6416 , \6429 , \6430 );
not \U$6185 ( \6432 , \6271 );
not \U$6186 ( \6433 , \6351 );
or \U$6187 ( \6434 , \6432 , \6433 );
not \U$6188 ( \6435 , \6277 );
or \U$6189 ( \6436 , \6435 , \6347 );
nand \U$6190 ( \6437 , \6434 , \6436 );
not \U$6191 ( \6438 , \6437 );
not \U$6192 ( \6439 , \6438 );
not \U$6193 ( \6440 , \6343 );
not \U$6194 ( \6441 , \6440 );
not \U$6195 ( \6442 , \6317 );
or \U$6196 ( \6443 , \6441 , \6442 );
not \U$6197 ( \6444 , \6312 );
nand \U$6198 ( \6445 , \6444 , \6303 );
nand \U$6199 ( \6446 , \6443 , \6445 );
not \U$6200 ( \6447 , \6212 );
not \U$6201 ( \6448 , \6270 );
or \U$6202 ( \6449 , \6447 , \6448 );
not \U$6203 ( \6450 , \6231 );
nand \U$6204 ( \6451 , \6450 , \6266 );
nand \U$6205 ( \6452 , \6449 , \6451 );
xor \U$6206 ( \6453 , \6446 , \6452 );
not \U$6207 ( \6454 , \6328 );
not \U$6208 ( \6455 , \6335 );
or \U$6209 ( \6456 , \6454 , \6455 );
nand \U$6210 ( \6457 , \6336 , \6342 );
nand \U$6211 ( \6458 , \6456 , \6457 );
not \U$6212 ( \6459 , \6285 );
not \U$6213 ( \6460 , \6302 );
or \U$6214 ( \6461 , \6459 , \6460 );
not \U$6215 ( \6462 , \6286 );
nand \U$6216 ( \6463 , \6462 , \6298 );
nand \U$6217 ( \6464 , \6461 , \6463 );
xor \U$6218 ( \6465 , \6458 , \6464 );
not \U$6219 ( \6466 , \5975 );
not \U$6220 ( \6467 , \6283 );
not \U$6221 ( \6468 , \6467 );
not \U$6222 ( \6469 , \1452 );
or \U$6223 ( \6470 , \6468 , \6469 );
not \U$6224 ( \6471 , RIbe28c78_38);
not \U$6225 ( \6472 , RIbe296c8_60);
and \U$6226 ( \6473 , \6471 , \6472 );
and \U$6227 ( \6474 , RIbe28c78_38, RIbe296c8_60);
nor \U$6228 ( \6475 , \6473 , \6474 );
nand \U$6229 ( \6476 , \1137 , \6475 );
nand \U$6230 ( \6477 , \6470 , \6476 );
not \U$6231 ( \6478 , \6477 );
or \U$6232 ( \6479 , \6466 , \6478 );
or \U$6233 ( \6480 , \6477 , \5975 );
nand \U$6234 ( \6481 , \6479 , \6480 );
and \U$6235 ( \6482 , \862 , \6255 );
and \U$6236 ( \6483 , \1517 , \3752 );
and \U$6237 ( \6484 , RIbe280c0_13, RIbe284f8_22);
nor \U$6238 ( \6485 , \6483 , \6484 );
and \U$6239 ( \6486 , \869 , \6485 );
nor \U$6240 ( \6487 , \6482 , \6486 );
not \U$6241 ( \6488 , \6487 );
and \U$6242 ( \6489 , \6481 , \6488 );
not \U$6243 ( \6490 , \6481 );
and \U$6244 ( \6491 , \6490 , \6487 );
nor \U$6245 ( \6492 , \6489 , \6491 );
xor \U$6246 ( \6493 , \6465 , \6492 );
not \U$6247 ( \6494 , \6493 );
and \U$6248 ( \6495 , \6453 , \6494 );
not \U$6249 ( \6496 , \6453 );
and \U$6250 ( \6497 , \6496 , \6493 );
nor \U$6251 ( \6498 , \6495 , \6497 );
not \U$6252 ( \6499 , \6498 );
and \U$6253 ( \6500 , \6439 , \6499 );
xnor \U$6254 ( \6501 , \6437 , \6498 );
not \U$6255 ( \6502 , \6397 );
and \U$6256 ( \6503 , \6408 , \6502 );
and \U$6257 ( \6504 , \6401 , \6407 );
nor \U$6258 ( \6505 , \6503 , \6504 );
not \U$6259 ( \6506 , \6505 );
and \U$6260 ( \6507 , \6501 , \6506 );
nor \U$6261 ( \6508 , \6500 , \6507 );
not \U$6262 ( \6509 , \6508 );
not \U$6263 ( \6510 , \6509 );
not \U$6264 ( \6511 , \6241 );
not \U$6265 ( \6512 , \2702 );
or \U$6266 ( \6513 , \6511 , \6512 );
nand \U$6267 ( \6514 , \2561 , RIbe28b88_36);
nand \U$6268 ( \6515 , \6513 , \6514 );
not \U$6269 ( \6516 , \6515 );
xor \U$6270 ( \6517 , \6197 , \6201 );
and \U$6271 ( \6518 , \6517 , \6211 );
and \U$6272 ( \6519 , \6197 , \6201 );
or \U$6273 ( \6520 , \6518 , \6519 );
xor \U$6274 ( \6521 , \6516 , \6520 );
or \U$6275 ( \6522 , \6264 , \6243 );
not \U$6276 ( \6523 , \6249 );
or \U$6277 ( \6524 , \6523 , \6257 );
nand \U$6278 ( \6525 , \6522 , \6524 );
and \U$6279 ( \6526 , \6521 , \6525 );
not \U$6280 ( \6527 , \6521 );
not \U$6281 ( \6528 , \6525 );
and \U$6282 ( \6529 , \6527 , \6528 );
nor \U$6283 ( \6530 , \6526 , \6529 );
not \U$6284 ( \6531 , \6530 );
not \U$6285 ( \6532 , \6377 );
not \U$6286 ( \6533 , \6370 );
or \U$6287 ( \6534 , \6532 , \6533 );
not \U$6288 ( \6535 , \6369 );
nand \U$6289 ( \6536 , \6535 , \6362 );
nand \U$6290 ( \6537 , \6534 , \6536 );
not \U$6291 ( \6538 , \6537 );
not \U$6292 ( \6539 , \6226 );
not \U$6293 ( \6540 , \6539 );
not \U$6294 ( \6541 , \6109 );
and \U$6295 ( \6542 , \6540 , \6541 );
not \U$6296 ( \6543 , \6222 );
and \U$6297 ( \6544 , \6217 , \6543 );
nor \U$6298 ( \6545 , \6542 , \6544 );
not \U$6299 ( \6546 , \6545 );
and \U$6300 ( \6547 , \6538 , \6546 );
and \U$6301 ( \6548 , \6537 , \6545 );
nor \U$6302 ( \6549 , \6547 , \6548 );
not \U$6303 ( \6550 , \6549 );
not \U$6304 ( \6551 , \6550 );
or \U$6305 ( \6552 , \6531 , \6551 );
not \U$6306 ( \6553 , \6537 );
or \U$6307 ( \6554 , \6553 , \6545 );
nand \U$6308 ( \6555 , \6552 , \6554 );
and \U$6309 ( \6556 , \363 , \951 );
and \U$6310 ( \6557 , RIbe27c10_3, RIbe282a0_17);
nor \U$6311 ( \6558 , \6556 , \6557 );
and \U$6312 ( \6559 , \2063 , \6558 );
and \U$6313 ( \6560 , \1174 , \2225 );
nor \U$6314 ( \6561 , \6559 , \6560 );
not \U$6315 ( \6562 , \6561 );
not \U$6316 ( \6563 , \6562 );
and \U$6317 ( \6564 , \314 , \2323 );
and \U$6318 ( \6565 , RIbe27d78_6, RIbe294e8_56);
nor \U$6319 ( \6566 , RIbe27d78_6, RIbe294e8_56);
nor \U$6320 ( \6567 , \6565 , \6566 );
and \U$6321 ( \6568 , \1044 , \6567 );
nor \U$6322 ( \6569 , \6564 , \6568 );
not \U$6323 ( \6570 , \6569 );
xor \U$6324 ( \6571 , RIbe295d8_58, RIbe27b98_2);
not \U$6325 ( \6572 , \6571 );
not \U$6326 ( \6573 , \546 );
or \U$6327 ( \6574 , \6572 , \6573 );
not \U$6328 ( \6575 , \2310 );
nand \U$6329 ( \6576 , \6575 , \1298 );
nand \U$6330 ( \6577 , \6574 , \6576 );
not \U$6331 ( \6578 , \6577 );
or \U$6332 ( \6579 , \6570 , \6578 );
or \U$6333 ( \6580 , \6577 , \6569 );
nand \U$6334 ( \6581 , \6579 , \6580 );
not \U$6335 ( \6582 , \6581 );
not \U$6336 ( \6583 , \6582 );
or \U$6337 ( \6584 , \6563 , \6583 );
nand \U$6338 ( \6585 , \6581 , \6561 );
nand \U$6339 ( \6586 , \6584 , \6585 );
xor \U$6340 ( \6587 , RIbe28de0_41, RIbe297b8_62);
not \U$6341 ( \6588 , \6587 );
not \U$6342 ( \6589 , \1284 );
or \U$6343 ( \6590 , \6588 , \6589 );
nand \U$6344 ( \6591 , \514 , \2211 );
nand \U$6345 ( \6592 , \6590 , \6591 );
not \U$6346 ( \6593 , \6592 );
not \U$6347 ( \6594 , \6339 );
and \U$6348 ( \6595 , \6593 , \6594 );
and \U$6349 ( \6596 , \6592 , \6339 );
nor \U$6350 ( \6597 , \6595 , \6596 );
and \U$6351 ( \6598 , \2877 , \6475 );
and \U$6352 ( \6599 , \908 , \2247 );
nor \U$6353 ( \6600 , \6598 , \6599 );
xnor \U$6354 ( \6601 , \6597 , \6600 );
not \U$6355 ( \6602 , \6601 );
and \U$6356 ( \6603 , \6586 , \6602 );
not \U$6357 ( \6604 , \6586 );
and \U$6358 ( \6605 , \6604 , \6601 );
nor \U$6359 ( \6606 , \6603 , \6605 );
not \U$6360 ( \6607 , \283 );
and \U$6361 ( \6608 , RIbe29038_46, RIbe29308_52);
nor \U$6362 ( \6609 , RIbe29038_46, RIbe29308_52);
nor \U$6363 ( \6610 , \6608 , \6609 );
not \U$6364 ( \6611 , \6610 );
not \U$6365 ( \6612 , \6611 );
and \U$6366 ( \6613 , \6607 , \6612 );
nor \U$6367 ( \6614 , \1465 , \2258 );
nor \U$6368 ( \6615 , \6613 , \6614 );
not \U$6369 ( \6616 , \6615 );
xnor \U$6370 ( \6617 , RIbe28048_12, RIbe28a20_33);
or \U$6371 ( \6618 , \3750 , \6617 );
not \U$6372 ( \6619 , \2476 );
or \U$6373 ( \6620 , \6619 , \2273 );
nand \U$6374 ( \6621 , \6618 , \6620 );
xnor \U$6375 ( \6622 , RIbe286d8_26, RIbe28930_31);
or \U$6376 ( \6623 , \967 , \6622 );
not \U$6377 ( \6624 , \2303 );
or \U$6378 ( \6625 , \972 , \6624 );
nand \U$6379 ( \6626 , \6623 , \6625 );
or \U$6380 ( \6627 , \6621 , \6626 );
not \U$6381 ( \6628 , \6627 );
and \U$6382 ( \6629 , \6621 , \6626 );
nor \U$6383 ( \6630 , \6628 , \6629 );
not \U$6384 ( \6631 , \6630 );
or \U$6385 ( \6632 , \6616 , \6631 );
or \U$6386 ( \6633 , \6630 , \6615 );
nand \U$6387 ( \6634 , \6632 , \6633 );
xnor \U$6388 ( \6635 , \6606 , \6634 );
not \U$6389 ( \6636 , \6635 );
and \U$6390 ( \6637 , \6521 , \6525 );
and \U$6391 ( \6638 , \6516 , \6520 );
nor \U$6392 ( \6639 , \6637 , \6638 );
not \U$6393 ( \6640 , \6639 );
and \U$6394 ( \6641 , \1054 , \6485 );
and \U$6395 ( \6642 , \1517 , \902 );
and \U$6396 ( \6643 , RIbe280c0_13, RIbe28750_27);
nor \U$6397 ( \6644 , \6642 , \6643 );
and \U$6398 ( \6645 , \869 , \6644 );
nor \U$6399 ( \6646 , \6641 , \6645 );
nand \U$6400 ( \6647 , \4541 , \2692 );
and \U$6401 ( \6648 , \6647 , RIbe28b88_36);
xor \U$6402 ( \6649 , \6646 , \6648 );
xor \U$6403 ( \6650 , RIbe28a98_34, RIbe290b0_47);
and \U$6404 ( \6651 , \466 , \6650 );
and \U$6405 ( \6652 , \469 , \2217 );
nor \U$6406 ( \6653 , \6651 , \6652 );
xor \U$6407 ( \6654 , \6649 , \6653 );
not \U$6408 ( \6655 , \6654 );
not \U$6409 ( \6656 , RIbe28228_16);
not \U$6410 ( \6657 , RIbe28840_29);
and \U$6411 ( \6658 , \6656 , \6657 );
and \U$6412 ( \6659 , RIbe28228_16, RIbe28840_29);
nor \U$6413 ( \6660 , \6658 , \6659 );
and \U$6414 ( \6661 , \1061 , \6660 );
and \U$6415 ( \6662 , \885 , \2237 );
nor \U$6416 ( \6663 , \6661 , \6662 );
not \U$6417 ( \6664 , \6663 );
not \U$6418 ( \6665 , \6515 );
or \U$6419 ( \6666 , \6664 , \6665 );
or \U$6420 ( \6667 , \6515 , \6663 );
nand \U$6421 ( \6668 , \6666 , \6667 );
not \U$6422 ( \6669 , \6214 );
not \U$6423 ( \6670 , \1061 );
or \U$6424 ( \6671 , \6669 , \6670 );
nand \U$6425 ( \6672 , \885 , \6660 );
nand \U$6426 ( \6673 , \6671 , \6672 );
or \U$6427 ( \6674 , \1782 , \6199 );
or \U$6428 ( \6675 , \1770 , \6617 );
nand \U$6429 ( \6676 , \6674 , \6675 );
xor \U$6430 ( \6677 , \6673 , \6676 );
or \U$6431 ( \6678 , \967 , \6195 );
or \U$6432 ( \6679 , \1200 , \6622 );
nand \U$6433 ( \6680 , \6678 , \6679 );
and \U$6434 ( \6681 , \6677 , \6680 );
and \U$6435 ( \6682 , \6673 , \6676 );
or \U$6436 ( \6683 , \6681 , \6682 );
xor \U$6437 ( \6684 , \6668 , \6683 );
not \U$6438 ( \6685 , \6684 );
or \U$6439 ( \6686 , \6655 , \6685 );
or \U$6440 ( \6687 , \6684 , \6654 );
nand \U$6441 ( \6688 , \6686 , \6687 );
not \U$6442 ( \6689 , \6688 );
or \U$6443 ( \6690 , \6640 , \6689 );
or \U$6444 ( \6691 , \6639 , \6688 );
nand \U$6445 ( \6692 , \6690 , \6691 );
not \U$6446 ( \6693 , \6692 );
or \U$6447 ( \6694 , \6636 , \6693 );
or \U$6448 ( \6695 , \6692 , \6635 );
nand \U$6449 ( \6696 , \6694 , \6695 );
xnor \U$6450 ( \6697 , \6555 , \6696 );
not \U$6451 ( \6698 , \6697 );
and \U$6452 ( \6699 , \332 , \6296 );
and \U$6453 ( \6700 , \347 , \6587 );
nor \U$6454 ( \6701 , \6699 , \6700 );
and \U$6455 ( \6702 , \2063 , \6326 );
and \U$6456 ( \6703 , \370 , \6558 );
nor \U$6457 ( \6704 , \6702 , \6703 );
xor \U$6458 ( \6705 , \6701 , \6704 );
not \U$6459 ( \6706 , \6247 );
not \U$6460 ( \6707 , \466 );
or \U$6461 ( \6708 , \6706 , \6707 );
nand \U$6462 ( \6709 , \399 , \6650 );
nand \U$6463 ( \6710 , \6708 , \6709 );
not \U$6464 ( \6711 , \6710 );
xor \U$6465 ( \6712 , \6705 , \6711 );
not \U$6466 ( \6713 , \6712 );
not \U$6467 ( \6714 , \6713 );
not \U$6468 ( \6715 , \6206 );
not \U$6469 ( \6716 , \979 );
or \U$6470 ( \6717 , \6715 , \6716 );
nand \U$6471 ( \6718 , \287 , \6610 );
nand \U$6472 ( \6719 , \6717 , \6718 );
not \U$6473 ( \6720 , \6719 );
and \U$6474 ( \6721 , \315 , \6567 );
not \U$6475 ( \6722 , \5739 );
nor \U$6476 ( \6723 , \6722 , \6332 );
nor \U$6477 ( \6724 , \6721 , \6723 );
not \U$6478 ( \6725 , \6724 );
or \U$6479 ( \6726 , \6720 , \6725 );
or \U$6480 ( \6727 , \6719 , \6724 );
nand \U$6481 ( \6728 , \6726 , \6727 );
not \U$6482 ( \6729 , \6728 );
not \U$6483 ( \6730 , \946 );
not \U$6484 ( \6731 , \6340 );
and \U$6485 ( \6732 , \6730 , \6731 );
and \U$6486 ( \6733 , \1298 , \6571 );
nor \U$6487 ( \6734 , \6732 , \6733 );
not \U$6488 ( \6735 , \6734 );
and \U$6489 ( \6736 , \6729 , \6735 );
and \U$6490 ( \6737 , \6728 , \6734 );
nor \U$6491 ( \6738 , \6736 , \6737 );
nand \U$6492 ( \6739 , \6714 , \6738 );
xor \U$6493 ( \6740 , \6673 , \6676 );
xor \U$6494 ( \6741 , \6740 , \6680 );
and \U$6495 ( \6742 , \6739 , \6741 );
not \U$6496 ( \6743 , \6738 );
nand \U$6497 ( \6744 , \6743 , \6713 );
not \U$6498 ( \6745 , \6744 );
nor \U$6499 ( \6746 , \6742 , \6745 );
not \U$6500 ( \6747 , \6746 );
not \U$6501 ( \6748 , \6747 );
not \U$6502 ( \6749 , \6492 );
not \U$6503 ( \6750 , \6465 );
or \U$6504 ( \6751 , \6749 , \6750 );
nand \U$6505 ( \6752 , \6464 , \6458 );
nand \U$6506 ( \6753 , \6751 , \6752 );
not \U$6507 ( \6754 , \6753 );
not \U$6508 ( \6755 , \6754 );
or \U$6509 ( \6756 , \6748 , \6755 );
nand \U$6510 ( \6757 , \6753 , \6746 );
nand \U$6511 ( \6758 , \6756 , \6757 );
not \U$6512 ( \6759 , \6734 );
not \U$6513 ( \6760 , \6759 );
not \U$6514 ( \6761 , \6728 );
or \U$6515 ( \6762 , \6760 , \6761 );
not \U$6516 ( \6763 , \6724 );
nand \U$6517 ( \6764 , \6763 , \6719 );
nand \U$6518 ( \6765 , \6762 , \6764 );
not \U$6519 ( \6766 , \6488 );
not \U$6520 ( \6767 , \6481 );
or \U$6521 ( \6768 , \6766 , \6767 );
not \U$6522 ( \6769 , \5975 );
nand \U$6523 ( \6770 , \6769 , \6477 );
nand \U$6524 ( \6771 , \6768 , \6770 );
xor \U$6525 ( \6772 , \6765 , \6771 );
xor \U$6526 ( \6773 , \6701 , \6704 );
not \U$6527 ( \6774 , \6710 );
and \U$6528 ( \6775 , \6773 , \6774 );
and \U$6529 ( \6776 , \6701 , \6704 );
or \U$6530 ( \6777 , \6775 , \6776 );
not \U$6531 ( \6778 , \6777 );
xor \U$6532 ( \6779 , \6772 , \6778 );
xnor \U$6533 ( \6780 , \6758 , \6779 );
not \U$6534 ( \6781 , \6780 );
not \U$6535 ( \6782 , \6493 );
not \U$6536 ( \6783 , \6453 );
or \U$6537 ( \6784 , \6782 , \6783 );
nand \U$6538 ( \6785 , \6452 , \6446 );
nand \U$6539 ( \6786 , \6784 , \6785 );
not \U$6540 ( \6787 , \6786 );
or \U$6541 ( \6788 , \6781 , \6787 );
or \U$6542 ( \6789 , \6786 , \6780 );
nand \U$6543 ( \6790 , \6788 , \6789 );
not \U$6544 ( \6791 , \6790 );
not \U$6545 ( \6792 , \6530 );
not \U$6546 ( \6793 , \6549 );
or \U$6547 ( \6794 , \6792 , \6793 );
or \U$6548 ( \6795 , \6549 , \6530 );
nand \U$6549 ( \6796 , \6794 , \6795 );
not \U$6550 ( \6797 , \6796 );
nand \U$6551 ( \6798 , \6739 , \6744 );
not \U$6552 ( \6799 , \6741 );
and \U$6553 ( \6800 , \6798 , \6799 );
not \U$6554 ( \6801 , \6798 );
and \U$6555 ( \6802 , \6801 , \6741 );
nor \U$6556 ( \6803 , \6800 , \6802 );
not \U$6557 ( \6804 , \6396 );
not \U$6558 ( \6805 , \6382 );
or \U$6559 ( \6806 , \6804 , \6805 );
nand \U$6560 ( \6807 , \6395 , \6388 );
nand \U$6561 ( \6808 , \6806 , \6807 );
xor \U$6562 ( \6809 , \6803 , \6808 );
not \U$6563 ( \6810 , \6809 );
or \U$6564 ( \6811 , \6797 , \6810 );
nand \U$6565 ( \6812 , \6808 , \6803 );
nand \U$6566 ( \6813 , \6811 , \6812 );
not \U$6567 ( \6814 , \6813 );
not \U$6568 ( \6815 , \6814 );
or \U$6569 ( \6816 , \6791 , \6815 );
or \U$6570 ( \6817 , \6790 , \6814 );
nand \U$6571 ( \6818 , \6816 , \6817 );
not \U$6572 ( \6819 , \6818 );
or \U$6573 ( \6820 , \6698 , \6819 );
or \U$6574 ( \6821 , \6697 , \6818 );
nand \U$6575 ( \6822 , \6820 , \6821 );
not \U$6576 ( \6823 , \6822 );
or \U$6577 ( \6824 , \6510 , \6823 );
not \U$6578 ( \6825 , \6697 );
nand \U$6579 ( \6826 , \6825 , \6818 );
nand \U$6580 ( \6827 , \6824 , \6826 );
not \U$6581 ( \6828 , \6827 );
not \U$6582 ( \6829 , \6639 );
not \U$6583 ( \6830 , \6829 );
not \U$6584 ( \6831 , \6688 );
or \U$6585 ( \6832 , \6830 , \6831 );
not \U$6586 ( \6833 , \6654 );
nand \U$6587 ( \6834 , \6833 , \6684 );
nand \U$6588 ( \6835 , \6832 , \6834 );
xor \U$6589 ( \6836 , \2214 , \2221 );
xor \U$6590 ( \6837 , \6836 , \2228 );
xor \U$6591 ( \6838 , \6646 , \6648 );
and \U$6592 ( \6839 , \6838 , \6653 );
and \U$6593 ( \6840 , \6646 , \6648 );
or \U$6594 ( \6841 , \6839 , \6840 );
xor \U$6595 ( \6842 , \6837 , \6841 );
not \U$6596 ( \6843 , \2306 );
not \U$6597 ( \6844 , \2330 );
or \U$6598 ( \6845 , \6843 , \6844 );
or \U$6599 ( \6846 , \2330 , \2306 );
nand \U$6600 ( \6847 , \6845 , \6846 );
not \U$6601 ( \6848 , \6847 );
xor \U$6602 ( \6849 , \6842 , \6848 );
not \U$6603 ( \6850 , \6849 );
xor \U$6604 ( \6851 , \6835 , \6850 );
xor \U$6605 ( \6852 , \2263 , \2242 );
and \U$6606 ( \6853 , \1326 , \6644 );
and \U$6607 ( \6854 , \869 , \1821 );
nor \U$6608 ( \6855 , \6853 , \6854 );
not \U$6609 ( \6856 , \6855 );
and \U$6610 ( \6857 , RIbe295d8_58, RIbe27b98_2);
not \U$6611 ( \6858 , \6857 );
not \U$6612 ( \6859 , \2280 );
or \U$6613 ( \6860 , \6858 , \6859 );
or \U$6614 ( \6861 , \2280 , \6857 );
nand \U$6615 ( \6862 , \6860 , \6861 );
not \U$6616 ( \6863 , \6862 );
or \U$6617 ( \6864 , \6856 , \6863 );
or \U$6618 ( \6865 , \6862 , \6855 );
nand \U$6619 ( \6866 , \6864 , \6865 );
xnor \U$6620 ( \6867 , \6852 , \6866 );
xor \U$6621 ( \6868 , \6765 , \6771 );
and \U$6622 ( \6869 , \6868 , \6778 );
and \U$6623 ( \6870 , \6765 , \6771 );
nor \U$6624 ( \6871 , \6869 , \6870 );
xor \U$6625 ( \6872 , \6867 , \6871 );
xor \U$6626 ( \6873 , \6851 , \6872 );
or \U$6627 ( \6874 , \6582 , \6561 );
not \U$6628 ( \6875 , \6577 );
or \U$6629 ( \6876 , \6875 , \6569 );
nand \U$6630 ( \6877 , \6874 , \6876 );
not \U$6631 ( \6878 , \6877 );
not \U$6632 ( \6879 , \6878 );
or \U$6633 ( \6880 , \6597 , \6600 );
not \U$6634 ( \6881 , \6592 );
or \U$6635 ( \6882 , \6881 , \6339 );
nand \U$6636 ( \6883 , \6880 , \6882 );
not \U$6637 ( \6884 , \6883 );
not \U$6638 ( \6885 , \6615 );
and \U$6639 ( \6886 , \6627 , \6885 );
nor \U$6640 ( \6887 , \6886 , \6629 );
not \U$6641 ( \6888 , \6887 );
and \U$6642 ( \6889 , \6884 , \6888 );
and \U$6643 ( \6890 , \6883 , \6887 );
nor \U$6644 ( \6891 , \6889 , \6890 );
not \U$6645 ( \6892 , \6891 );
not \U$6646 ( \6893 , \6892 );
or \U$6647 ( \6894 , \6879 , \6893 );
nand \U$6648 ( \6895 , \6877 , \6891 );
nand \U$6649 ( \6896 , \6894 , \6895 );
not \U$6650 ( \6897 , \6668 );
not \U$6651 ( \6898 , \6683 );
or \U$6652 ( \6899 , \6897 , \6898 );
or \U$6653 ( \6900 , \6516 , \6663 );
nand \U$6654 ( \6901 , \6899 , \6900 );
xor \U$6655 ( \6902 , \6896 , \6901 );
not \U$6656 ( \6903 , \6634 );
not \U$6657 ( \6904 , \6606 );
or \U$6658 ( \6905 , \6903 , \6904 );
not \U$6659 ( \6906 , \6586 );
or \U$6660 ( \6907 , \6906 , \6601 );
nand \U$6661 ( \6908 , \6905 , \6907 );
xor \U$6662 ( \6909 , \6902 , \6908 );
not \U$6663 ( \6910 , \6779 );
not \U$6664 ( \6911 , \6758 );
or \U$6665 ( \6912 , \6910 , \6911 );
or \U$6666 ( \6913 , \6754 , \6746 );
nand \U$6667 ( \6914 , \6912 , \6913 );
and \U$6668 ( \6915 , \6909 , \6914 );
not \U$6669 ( \6916 , \6909 );
not \U$6670 ( \6917 , \6914 );
and \U$6671 ( \6918 , \6916 , \6917 );
nor \U$6672 ( \6919 , \6915 , \6918 );
not \U$6673 ( \6920 , \6696 );
not \U$6674 ( \6921 , \6555 );
or \U$6675 ( \6922 , \6920 , \6921 );
not \U$6676 ( \6923 , \6635 );
nand \U$6677 ( \6924 , \6923 , \6692 );
nand \U$6678 ( \6925 , \6922 , \6924 );
and \U$6679 ( \6926 , \6919 , \6925 );
not \U$6680 ( \6927 , \6919 );
not \U$6681 ( \6928 , \6925 );
and \U$6682 ( \6929 , \6927 , \6928 );
nor \U$6683 ( \6930 , \6926 , \6929 );
xor \U$6684 ( \6931 , \6873 , \6930 );
not \U$6685 ( \6932 , \6931 );
and \U$6686 ( \6933 , \6790 , \6813 );
not \U$6687 ( \6934 , \6780 );
and \U$6688 ( \6935 , \6786 , \6934 );
nor \U$6689 ( \6936 , \6933 , \6935 );
not \U$6690 ( \6937 , \6936 );
and \U$6691 ( \6938 , \6932 , \6937 );
and \U$6692 ( \6939 , \6931 , \6936 );
nor \U$6693 ( \6940 , \6938 , \6939 );
nand \U$6694 ( \6941 , \6828 , \6940 );
not \U$6695 ( \6942 , \6822 );
not \U$6696 ( \6943 , \6508 );
and \U$6697 ( \6944 , \6942 , \6943 );
and \U$6698 ( \6945 , \6822 , \6508 );
nor \U$6699 ( \6946 , \6944 , \6945 );
not \U$6700 ( \6947 , \6501 );
not \U$6701 ( \6948 , \6505 );
and \U$6702 ( \6949 , \6947 , \6948 );
and \U$6703 ( \6950 , \6501 , \6505 );
nor \U$6704 ( \6951 , \6949 , \6950 );
not \U$6705 ( \6952 , \6951 );
xor \U$6706 ( \6953 , \6809 , \6796 );
not \U$6707 ( \6954 , \6356 );
not \U$6708 ( \6955 , \6409 );
or \U$6709 ( \6956 , \6954 , \6955 );
not \U$6710 ( \6957 , \6192 );
nand \U$6711 ( \6958 , \6957 , \6352 );
nand \U$6712 ( \6959 , \6956 , \6958 );
xor \U$6713 ( \6960 , \6953 , \6959 );
and \U$6714 ( \6961 , \6952 , \6960 );
and \U$6715 ( \6962 , \6953 , \6959 );
nor \U$6716 ( \6963 , \6961 , \6962 );
nand \U$6717 ( \6964 , \6946 , \6963 );
buf \U$6718 ( \6965 , \6964 );
nand \U$6719 ( \6966 , \6941 , \6965 );
not \U$6720 ( \6967 , \6410 );
not \U$6721 ( \6968 , \6187 );
or \U$6722 ( \6969 , \6967 , \6968 );
nand \U$6723 ( \6970 , \6181 , \6174 );
nand \U$6724 ( \6971 , \6969 , \6970 );
xnor \U$6725 ( \6972 , \6951 , \6960 );
or \U$6726 ( \6973 , \6971 , \6972 );
not \U$6727 ( \6974 , \6931 );
nor \U$6728 ( \6975 , \6974 , \6936 );
and \U$6729 ( \6976 , \6873 , \6930 );
nor \U$6730 ( \6977 , \6975 , \6976 );
xor \U$6731 ( \6978 , \2298 , \2335 );
xor \U$6732 ( \6979 , \6978 , \2337 );
not \U$6733 ( \6980 , \6979 );
not \U$6734 ( \6981 , \6857 );
not \U$6735 ( \6982 , \2281 );
or \U$6736 ( \6983 , \6981 , \6982 );
not \U$6737 ( \6984 , \6855 );
nand \U$6738 ( \6985 , \6984 , \6862 );
nand \U$6739 ( \6986 , \6983 , \6985 );
not \U$6740 ( \6987 , \6986 );
xor \U$6741 ( \6988 , \1716 , \1717 );
xor \U$6742 ( \6989 , \6988 , \1724 );
not \U$6743 ( \6990 , \6989 );
or \U$6744 ( \6991 , \6987 , \6990 );
or \U$6745 ( \6992 , \6989 , \6986 );
nand \U$6746 ( \6993 , \6991 , \6992 );
xor \U$6747 ( \6994 , \1756 , \1763 );
xnor \U$6748 ( \6995 , \6993 , \6994 );
xor \U$6749 ( \6996 , \6980 , \6995 );
not \U$6750 ( \6997 , \6866 );
not \U$6751 ( \6998 , \6852 );
or \U$6752 ( \6999 , \6997 , \6998 );
or \U$6753 ( \7000 , \6871 , \6867 );
nand \U$6754 ( \7001 , \6999 , \7000 );
xnor \U$6755 ( \7002 , \6996 , \7001 );
not \U$6756 ( \7003 , \7002 );
not \U$6757 ( \7004 , \6925 );
not \U$6758 ( \7005 , \6919 );
or \U$6759 ( \7006 , \7004 , \7005 );
nand \U$6760 ( \7007 , \6914 , \6909 );
nand \U$6761 ( \7008 , \7006 , \7007 );
not \U$6762 ( \7009 , \7008 );
or \U$6763 ( \7010 , \7003 , \7009 );
or \U$6764 ( \7011 , \7008 , \7002 );
nand \U$6765 ( \7012 , \7010 , \7011 );
not \U$6766 ( \7013 , \7012 );
xor \U$6767 ( \7014 , \6896 , \6901 );
and \U$6768 ( \7015 , \7014 , \6908 );
and \U$6769 ( \7016 , \6896 , \6901 );
nor \U$6770 ( \7017 , \7015 , \7016 );
not \U$6771 ( \7018 , \6877 );
not \U$6772 ( \7019 , \6892 );
or \U$6773 ( \7020 , \7018 , \7019 );
not \U$6774 ( \7021 , \6887 );
nand \U$6775 ( \7022 , \7021 , \6883 );
nand \U$6776 ( \7023 , \7020 , \7022 );
and \U$6777 ( \7024 , \2231 , \2285 );
not \U$6778 ( \7025 , \2231 );
and \U$6779 ( \7026 , \7025 , \2286 );
or \U$6780 ( \7027 , \7024 , \7026 );
xor \U$6781 ( \7028 , \7023 , \7027 );
xor \U$6782 ( \7029 , \6837 , \6841 );
not \U$6783 ( \7030 , \6847 );
and \U$6784 ( \7031 , \7029 , \7030 );
and \U$6785 ( \7032 , \6837 , \6841 );
or \U$6786 ( \7033 , \7031 , \7032 );
not \U$6787 ( \7034 , \7033 );
xor \U$6788 ( \7035 , \7028 , \7034 );
and \U$6789 ( \7036 , \7017 , \7035 );
not \U$6790 ( \7037 , \7017 );
not \U$6791 ( \7038 , \7035 );
and \U$6792 ( \7039 , \7037 , \7038 );
nor \U$6793 ( \7040 , \7036 , \7039 );
xor \U$6794 ( \7041 , \6835 , \6850 );
and \U$6795 ( \7042 , \7041 , \6872 );
and \U$6796 ( \7043 , \6835 , \6850 );
nor \U$6797 ( \7044 , \7042 , \7043 );
not \U$6798 ( \7045 , \7044 );
xor \U$6799 ( \7046 , \7040 , \7045 );
not \U$6800 ( \7047 , \7046 );
and \U$6801 ( \7048 , \7013 , \7047 );
and \U$6802 ( \7049 , \7046 , \7012 );
nor \U$6803 ( \7050 , \7048 , \7049 );
nand \U$6804 ( \7051 , \6977 , \7050 );
nand \U$6805 ( \7052 , \6973 , \7051 );
nor \U$6806 ( \7053 , \6966 , \7052 );
xnor \U$6807 ( \7054 , \2296 , \2340 );
xor \U$6808 ( \7055 , \7023 , \7027 );
and \U$6809 ( \7056 , \7055 , \7034 );
and \U$6810 ( \7057 , \7023 , \7027 );
nor \U$6811 ( \7058 , \7056 , \7057 );
xor \U$6812 ( \7059 , \7054 , \7058 );
xor \U$6813 ( \7060 , \1848 , \1766 );
not \U$6814 ( \7061 , \6994 );
not \U$6815 ( \7062 , \6993 );
or \U$6816 ( \7063 , \7061 , \7062 );
not \U$6817 ( \7064 , \6989 );
nand \U$6818 ( \7065 , \7064 , \6986 );
nand \U$6819 ( \7066 , \7063 , \7065 );
xor \U$6820 ( \7067 , \7060 , \7066 );
not \U$6821 ( \7068 , \1688 );
nand \U$6822 ( \7069 , \7068 , \1684 );
xnor \U$6823 ( \7070 , \1686 , \7069 );
xor \U$6824 ( \7071 , \7067 , \7070 );
not \U$6825 ( \7072 , \7071 );
and \U$6826 ( \7073 , \7059 , \7072 );
and \U$6827 ( \7074 , \7054 , \7058 );
or \U$6828 ( \7075 , \7073 , \7074 );
xor \U$6829 ( \7076 , \7060 , \7066 );
and \U$6830 ( \7077 , \7076 , \7070 );
and \U$6831 ( \7078 , \7060 , \7066 );
nor \U$6832 ( \7079 , \7077 , \7078 );
xor \U$6833 ( \7080 , \7075 , \7079 );
xnor \U$6834 ( \7081 , \2351 , \2352 );
xor \U$6835 ( \7082 , \7080 , \7081 );
xor \U$6836 ( \7083 , \7054 , \7058 );
xor \U$6837 ( \7084 , \7083 , \7072 );
not \U$6838 ( \7085 , \7084 );
or \U$6839 ( \7086 , \6980 , \6995 );
not \U$6840 ( \7087 , \6995 );
not \U$6841 ( \7088 , \6980 );
or \U$6842 ( \7089 , \7087 , \7088 );
nand \U$6843 ( \7090 , \7089 , \7001 );
nand \U$6844 ( \7091 , \7086 , \7090 );
or \U$6845 ( \7092 , \7044 , \7040 );
or \U$6846 ( \7093 , \7038 , \7017 );
nand \U$6847 ( \7094 , \7092 , \7093 );
xor \U$6848 ( \7095 , \7091 , \7094 );
and \U$6849 ( \7096 , \7085 , \7095 );
and \U$6850 ( \7097 , \7091 , \7094 );
nor \U$6851 ( \7098 , \7096 , \7097 );
nand \U$6852 ( \7099 , \7082 , \7098 );
not \U$6853 ( \7100 , \7012 );
not \U$6854 ( \7101 , \7100 );
not \U$6855 ( \7102 , \7046 );
and \U$6856 ( \7103 , \7101 , \7102 );
not \U$6857 ( \7104 , \7002 );
and \U$6858 ( \7105 , \7008 , \7104 );
nor \U$6859 ( \7106 , \7103 , \7105 );
not \U$6860 ( \7107 , \7095 );
not \U$6861 ( \7108 , \7084 );
and \U$6862 ( \7109 , \7107 , \7108 );
and \U$6863 ( \7110 , \7095 , \7084 );
nor \U$6864 ( \7111 , \7109 , \7110 );
nand \U$6865 ( \7112 , \7106 , \7111 );
nand \U$6866 ( \7113 , \7099 , \7112 );
xor \U$6867 ( \7114 , \7075 , \7079 );
and \U$6868 ( \7115 , \7114 , \7081 );
and \U$6869 ( \7116 , \7075 , \7079 );
or \U$6870 ( \7117 , \7115 , \7116 );
xor \U$6871 ( \7118 , \2204 , \2205 );
xor \U$6872 ( \7119 , \7118 , \2355 );
and \U$6873 ( \7120 , \7117 , \7119 );
nor \U$6874 ( \7121 , \7113 , \7120 );
and \U$6875 ( \7122 , \7053 , \7121 );
nand \U$6876 ( \7123 , \6431 , \7122 );
not \U$6877 ( \7124 , \7113 );
not \U$6878 ( \7125 , \7124 );
not \U$6879 ( \7126 , \6941 );
not \U$6880 ( \7127 , \6964 );
and \U$6881 ( \7128 , \6971 , \6972 );
not \U$6882 ( \7129 , \7128 );
or \U$6883 ( \7130 , \7127 , \7129 );
not \U$6884 ( \7131 , \6946 );
not \U$6885 ( \7132 , \6963 );
nand \U$6886 ( \7133 , \7131 , \7132 );
nand \U$6887 ( \7134 , \7130 , \7133 );
not \U$6888 ( \7135 , \7134 );
or \U$6889 ( \7136 , \7126 , \7135 );
not \U$6890 ( \7137 , \6940 );
nand \U$6891 ( \7138 , \6827 , \7137 );
nand \U$6892 ( \7139 , \7136 , \7138 );
nand \U$6893 ( \7140 , \7139 , \7051 );
or \U$6894 ( \7141 , \6977 , \7050 );
nand \U$6895 ( \7142 , \7140 , \7141 );
not \U$6896 ( \7143 , \7142 );
or \U$6897 ( \7144 , \7125 , \7143 );
nor \U$6898 ( \7145 , \7106 , \7111 );
and \U$6899 ( \7146 , \7099 , \7145 );
nor \U$6900 ( \7147 , \7082 , \7098 );
nor \U$6901 ( \7148 , \7146 , \7147 );
nand \U$6902 ( \7149 , \7144 , \7148 );
not \U$6903 ( \7150 , \7120 );
nand \U$6904 ( \7151 , \7149 , \7150 );
or \U$6905 ( \7152 , \7117 , \7119 );
nand \U$6906 ( \7153 , \7123 , \7151 , \7152 );
not \U$6907 ( \7154 , \7153 );
or \U$6908 ( \7155 , \2361 , \7154 );
or \U$6909 ( \7156 , \2358 , \2359 );
nand \U$6910 ( \7157 , \7155 , \7156 );
not \U$6911 ( \7158 , \7157 );
or \U$6912 ( \7159 , \2203 , \7158 );
not \U$6913 ( \7160 , \1870 );
nand \U$6914 ( \7161 , \7160 , \1674 );
or \U$6915 ( \7162 , \7161 , \1668 );
nand \U$6916 ( \7163 , \1550 , \1667 );
nand \U$6917 ( \7164 , \7162 , \7163 );
nand \U$6918 ( \7165 , \7164 , \2100 );
or \U$6919 ( \7166 , \2099 , \2095 );
nand \U$6920 ( \7167 , \7165 , \7166 );
not \U$6921 ( \7168 , \7167 );
not \U$6922 ( \7169 , \2094 );
or \U$6923 ( \7170 , \7168 , \7169 );
or \U$6924 ( \7171 , \2003 , \2093 );
nand \U$6925 ( \7172 , \7170 , \7171 );
not \U$6926 ( \7173 , \7172 );
not \U$6927 ( \7174 , \2194 );
or \U$6928 ( \7175 , \7173 , \7174 );
nor \U$6929 ( \7176 , \2147 , \2104 );
and \U$6930 ( \7177 , \7176 , \2172 );
nor \U$6931 ( \7178 , \2171 , \2168 );
nor \U$6932 ( \7179 , \7177 , \7178 );
not \U$6933 ( \7180 , \7179 );
and \U$6934 ( \7181 , \7180 , \2193 );
nor \U$6935 ( \7182 , \2176 , \2192 );
nor \U$6936 ( \7183 , \7181 , \7182 );
nand \U$6937 ( \7184 , \7175 , \7183 );
not \U$6938 ( \7185 , \7184 );
not \U$6939 ( \7186 , \2201 );
or \U$6940 ( \7187 , \7185 , \7186 );
or \U$6941 ( \7188 , \2197 , \2200 );
nand \U$6942 ( \7189 , \7187 , \7188 );
not \U$6943 ( \7190 , \7189 );
nand \U$6944 ( \7191 , \7159 , \7190 );
not \U$6945 ( \7192 , \7191 );
not \U$6946 ( \7193 , \6413 );
or \U$6947 ( \7194 , \5108 , \5109 );
not \U$6948 ( \7195 , \6414 );
nand \U$6949 ( \7196 , \7194 , \7195 );
buf \U$6950 ( \7197 , \4754 );
nor \U$6951 ( \7198 , \7196 , \7197 );
nand \U$6952 ( \7199 , \7193 , \7198 );
nand \U$6953 ( \7200 , \7122 , \2360 );
nor \U$6954 ( \7201 , \7199 , \7200 );
and \U$6955 ( \7202 , \7201 , \2202 );
xor \U$6956 ( \7203 , \4963 , \4758 );
xnor \U$6957 ( \7204 , \5018 , \5032 );
not \U$6958 ( \7205 , \7204 );
xor \U$6959 ( \7206 , \4460 , \4438 );
xor \U$6960 ( \7207 , \7206 , \4450 );
not \U$6961 ( \7208 , \7207 );
or \U$6962 ( \7209 , \7205 , \7208 );
or \U$6963 ( \7210 , \7207 , \7204 );
nand \U$6964 ( \7211 , \7209 , \7210 );
xor \U$6965 ( \7212 , \5010 , \4997 );
xor \U$6966 ( \7213 , \7212 , \5001 );
not \U$6967 ( \7214 , \7213 );
and \U$6968 ( \7215 , \7211 , \7214 );
not \U$6969 ( \7216 , \7211 );
and \U$6970 ( \7217 , \7216 , \7213 );
nor \U$6971 ( \7218 , \7215 , \7217 );
not \U$6972 ( \7219 , \7218 );
not \U$6973 ( \7220 , \7219 );
not \U$6974 ( \7221 , \4832 );
not \U$6975 ( \7222 , \4854 );
or \U$6976 ( \7223 , \7221 , \7222 );
or \U$6977 ( \7224 , \4854 , \4832 );
nand \U$6978 ( \7225 , \7223 , \7224 );
and \U$6979 ( \7226 , \7225 , \4824 );
not \U$6980 ( \7227 , \7225 );
not \U$6981 ( \7228 , \4824 );
and \U$6982 ( \7229 , \7227 , \7228 );
nor \U$6983 ( \7230 , \7226 , \7229 );
not \U$6984 ( \7231 , \7230 );
xor \U$6985 ( \7232 , RIbe29c68_72, RIbe28048_12);
not \U$6986 ( \7233 , \7232 );
not \U$6987 ( \7234 , \5024 );
or \U$6988 ( \7235 , \7233 , \7234 );
not \U$6989 ( \7236 , \4580 );
not \U$6990 ( \7237 , \7236 );
nand \U$6991 ( \7238 , \7237 , \5022 );
nand \U$6992 ( \7239 , \7235 , \7238 );
xor \U$6993 ( \7240 , RIbe29a10_67, RIbe296c8_60);
not \U$6994 ( \7241 , \7240 );
not \U$6995 ( \7242 , \2875 );
or \U$6996 ( \7243 , \7241 , \7242 );
nand \U$6997 ( \7244 , \1939 , \4454 );
nand \U$6998 ( \7245 , \7243 , \7244 );
nor \U$6999 ( \7246 , \7239 , \7245 );
not \U$7000 ( \7247 , \7246 );
nand \U$7001 ( \7248 , \7239 , \7245 );
nand \U$7002 ( \7249 , \7247 , \7248 );
not \U$7003 ( \7250 , \7249 );
not \U$7004 ( \7251 , RIbe28228_16);
not \U$7005 ( \7252 , RIbe295d8_58);
and \U$7006 ( \7253 , \7251 , \7252 );
and \U$7007 ( \7254 , RIbe28228_16, RIbe295d8_58);
nor \U$7008 ( \7255 , \7253 , \7254 );
not \U$7009 ( \7256 , \7255 );
not \U$7010 ( \7257 , \1061 );
or \U$7011 ( \7258 , \7256 , \7257 );
nand \U$7012 ( \7259 , \885 , \4430 );
nand \U$7013 ( \7260 , \7258 , \7259 );
not \U$7014 ( \7261 , \7260 );
and \U$7015 ( \7262 , \7250 , \7261 );
and \U$7016 ( \7263 , \7249 , \7260 );
nor \U$7017 ( \7264 , \7262 , \7263 );
not \U$7018 ( \7265 , \7264 );
and \U$7019 ( \7266 , RIbe28138_14, RIbe28a20_33);
nor \U$7020 ( \7267 , RIbe28138_14, RIbe28a20_33);
nor \U$7021 ( \7268 , \7266 , \7267 );
not \U$7022 ( \7269 , \7268 );
not \U$7023 ( \7270 , \2276 );
or \U$7024 ( \7271 , \7269 , \7270 );
xor \U$7025 ( \7272 , RIbe28a20_33, RIbe282a0_17);
nand \U$7026 ( \7273 , \1769 , \7272 );
nand \U$7027 ( \7274 , \7271 , \7273 );
not \U$7028 ( \7275 , \7274 );
nand \U$7029 ( \7276 , RIbe27b98_2, RIbe2b6a8_128);
and \U$7030 ( \7277 , RIbe28b88_36, RIbe29470_55);
nor \U$7031 ( \7278 , RIbe28b88_36, RIbe29470_55);
nor \U$7032 ( \7279 , \7277 , \7278 );
not \U$7033 ( \7280 , \7279 );
not \U$7034 ( \7281 , \3401 );
or \U$7035 ( \7282 , \7280 , \7281 );
nand \U$7036 ( \7283 , \2691 , \4790 );
nand \U$7037 ( \7284 , \7282 , \7283 );
not \U$7038 ( \7285 , \7284 );
xnor \U$7039 ( \7286 , \7276 , \7285 );
not \U$7040 ( \7287 , \7286 );
or \U$7041 ( \7288 , \7275 , \7287 );
not \U$7042 ( \7289 , \7276 );
nand \U$7043 ( \7290 , \7289 , \7285 );
nand \U$7044 ( \7291 , \7288 , \7290 );
not \U$7045 ( \7292 , \7291 );
or \U$7046 ( \7293 , \7265 , \7292 );
or \U$7047 ( \7294 , \7291 , \7264 );
nand \U$7048 ( \7295 , \7293 , \7294 );
not \U$7049 ( \7296 , \7295 );
or \U$7050 ( \7297 , \7231 , \7296 );
not \U$7051 ( \7298 , \7264 );
nand \U$7052 ( \7299 , \7291 , \7298 );
nand \U$7053 ( \7300 , \7297 , \7299 );
xor \U$7054 ( \7301 , \4875 , \4866 );
xor \U$7055 ( \7302 , RIbe29218_50, RIbe296c8_60);
not \U$7056 ( \7303 , \7302 );
not \U$7057 ( \7304 , \1132 );
or \U$7058 ( \7305 , \7303 , \7304 );
nand \U$7059 ( \7306 , \1137 , \7240 );
nand \U$7060 ( \7307 , \7305 , \7306 );
not \U$7061 ( \7308 , \7307 );
xor \U$7062 ( \7309 , RIbe29b78_70, RIbe27c10_3);
not \U$7063 ( \7310 , \7309 );
not \U$7064 ( \7311 , \1493 );
or \U$7065 ( \7312 , \7310 , \7311 );
xor \U$7066 ( \7313 , RIbe27c10_3, RIbe27b20_1);
nand \U$7067 ( \7314 , \370 , \7313 );
nand \U$7068 ( \7315 , \7312 , \7314 );
and \U$7069 ( \7316 , RIbe28228_16, RIbe291a0_49);
nor \U$7070 ( \7317 , RIbe28228_16, RIbe291a0_49);
nor \U$7071 ( \7318 , \7316 , \7317 );
not \U$7072 ( \7319 , \7318 );
not \U$7073 ( \7320 , \1061 );
or \U$7074 ( \7321 , \7319 , \7320 );
nand \U$7075 ( \7322 , \885 , \7255 );
nand \U$7076 ( \7323 , \7321 , \7322 );
xor \U$7077 ( \7324 , \7315 , \7323 );
not \U$7078 ( \7325 , \7324 );
or \U$7079 ( \7326 , \7308 , \7325 );
nand \U$7080 ( \7327 , \7323 , \7315 );
nand \U$7081 ( \7328 , \7326 , \7327 );
xor \U$7082 ( \7329 , \7301 , \7328 );
not \U$7083 ( \7330 , \4813 );
not \U$7084 ( \7331 , \7330 );
xor \U$7085 ( \7332 , \4803 , \4795 );
not \U$7086 ( \7333 , \7332 );
or \U$7087 ( \7334 , \7331 , \7333 );
or \U$7088 ( \7335 , \7332 , \7330 );
nand \U$7089 ( \7336 , \7334 , \7335 );
and \U$7090 ( \7337 , \7329 , \7336 );
and \U$7091 ( \7338 , \7301 , \7328 );
nor \U$7092 ( \7339 , \7337 , \7338 );
xnor \U$7093 ( \7340 , \7300 , \7339 );
not \U$7094 ( \7341 , \7340 );
or \U$7095 ( \7342 , \7220 , \7341 );
not \U$7096 ( \7343 , \7339 );
nand \U$7097 ( \7344 , \7343 , \7300 );
nand \U$7098 ( \7345 , \7342 , \7344 );
not \U$7099 ( \7346 , RIbe27e68_8);
not \U$7100 ( \7347 , RIbe28c78_38);
and \U$7101 ( \7348 , \7346 , \7347 );
and \U$7102 ( \7349 , RIbe27e68_8, RIbe28c78_38);
nor \U$7103 ( \7350 , \7348 , \7349 );
and \U$7104 ( \7351 , \2600 , \7350 );
and \U$7105 ( \7352 , RIbe27e68_8, RIbe28318_18);
nor \U$7106 ( \7353 , RIbe27e68_8, RIbe28318_18);
nor \U$7107 ( \7354 , \7352 , \7353 );
and \U$7108 ( \7355 , \2464 , \7354 );
nor \U$7109 ( \7356 , \7351 , \7355 );
not \U$7110 ( \7357 , \7356 );
not \U$7111 ( \7358 , \7357 );
and \U$7112 ( \7359 , RIbe28228_16, RIbe29128_48);
nor \U$7113 ( \7360 , RIbe28228_16, RIbe29128_48);
nor \U$7114 ( \7361 , \7359 , \7360 );
not \U$7115 ( \7362 , \7361 );
not \U$7116 ( \7363 , \879 );
or \U$7117 ( \7364 , \7362 , \7363 );
nand \U$7118 ( \7365 , \885 , \7318 );
nand \U$7119 ( \7366 , \7364 , \7365 );
not \U$7120 ( \7367 , \7366 );
buf \U$7121 ( \7368 , \4849 );
xor \U$7122 ( \7369 , RIbe29e48_76, RIbe29380_53);
and \U$7123 ( \7370 , \7368 , \7369 );
buf \U$7124 ( \7371 , \4841 );
not \U$7125 ( \7372 , \7371 );
and \U$7126 ( \7373 , RIbe29e48_76, RIbe28048_12);
not \U$7127 ( \7374 , RIbe29e48_76);
and \U$7128 ( \7375 , \7374 , \431 );
nor \U$7129 ( \7376 , \7373 , \7375 );
and \U$7130 ( \7377 , \7372 , \7376 );
nor \U$7131 ( \7378 , \7370 , \7377 );
not \U$7132 ( \7379 , \7378 );
or \U$7133 ( \7380 , \7367 , \7379 );
or \U$7134 ( \7381 , \7366 , \7378 );
nand \U$7135 ( \7382 , \7380 , \7381 );
not \U$7136 ( \7383 , \7382 );
or \U$7137 ( \7384 , \7358 , \7383 );
not \U$7138 ( \7385 , \7378 );
nand \U$7139 ( \7386 , \7385 , \7366 );
nand \U$7140 ( \7387 , \7384 , \7386 );
not \U$7141 ( \7388 , \7387 );
and \U$7142 ( \7389 , RIbe285e8_24, \3840 );
not \U$7143 ( \7390 , RIbe285e8_24);
and \U$7144 ( \7391 , \7390 , RIbe29308_52);
or \U$7145 ( \7392 , \7389 , \7391 );
not \U$7146 ( \7393 , \7392 );
not \U$7147 ( \7394 , \2618 );
or \U$7148 ( \7395 , \7393 , \7394 );
xor \U$7149 ( \7396 , RIbe28c00_37, RIbe285e8_24);
nand \U$7150 ( \7397 , \2758 , \7396 );
nand \U$7151 ( \7398 , \7395 , \7397 );
not \U$7152 ( \7399 , \7398 );
xor \U$7153 ( \7400 , RIbe298a8_64, RIbe290b0_47);
not \U$7154 ( \7401 , \7400 );
not \U$7155 ( \7402 , \2730 );
or \U$7156 ( \7403 , \7401 , \7402 );
xor \U$7157 ( \7404 , RIbe29998_66, RIbe290b0_47);
nand \U$7158 ( \7405 , \398 , \7404 );
nand \U$7159 ( \7406 , \7403 , \7405 );
xor \U$7160 ( \7407 , RIbe29a10_67, RIbe280c0_13);
not \U$7161 ( \7408 , \7407 );
not \U$7162 ( \7409 , \2379 );
or \U$7163 ( \7410 , \7408 , \7409 );
and \U$7164 ( \7411 , RIbe280c0_13, RIbe29b00_69);
nor \U$7165 ( \7412 , RIbe280c0_13, RIbe29b00_69);
nor \U$7166 ( \7413 , \7411 , \7412 );
nand \U$7167 ( \7414 , \1263 , \7413 );
nand \U$7168 ( \7415 , \7410 , \7414 );
xor \U$7169 ( \7416 , \7406 , \7415 );
not \U$7170 ( \7417 , \7416 );
or \U$7171 ( \7418 , \7399 , \7417 );
nand \U$7172 ( \7419 , \7415 , \7406 );
nand \U$7173 ( \7420 , \7418 , \7419 );
not \U$7174 ( \7421 , \7420 );
not \U$7175 ( \7422 , RIbe28930_31);
not \U$7176 ( \7423 , RIbe295d8_58);
and \U$7177 ( \7424 , \7422 , \7423 );
and \U$7178 ( \7425 , RIbe28930_31, RIbe295d8_58);
nor \U$7179 ( \7426 , \7424 , \7425 );
not \U$7180 ( \7427 , \7426 );
not \U$7181 ( \7428 , \3064 );
or \U$7182 ( \7429 , \7427 , \7428 );
not \U$7183 ( \7430 , RIbe28930_31);
not \U$7184 ( \7431 , RIbe29740_61);
and \U$7185 ( \7432 , \7430 , \7431 );
and \U$7186 ( \7433 , RIbe28930_31, RIbe29740_61);
nor \U$7187 ( \7434 , \7432 , \7433 );
nand \U$7188 ( \7435 , \1797 , \7434 );
nand \U$7189 ( \7436 , \7429 , \7435 );
not \U$7190 ( \7437 , \7436 );
xor \U$7191 ( \7438 , RIbe29ce0_73, RIbe27c10_3);
not \U$7192 ( \7439 , \7438 );
not \U$7193 ( \7440 , \359 );
not \U$7194 ( \7441 , \7440 );
or \U$7195 ( \7442 , \7439 , \7441 );
nand \U$7196 ( \7443 , \369 , \7309 );
nand \U$7197 ( \7444 , \7442 , \7443 );
xor \U$7198 ( \7445 , RIbe297b8_62, RIbe28a20_33);
not \U$7199 ( \7446 , \7445 );
not \U$7200 ( \7447 , \1780 );
or \U$7201 ( \7448 , \7446 , \7447 );
nand \U$7202 ( \7449 , \2475 , \7268 );
nand \U$7203 ( \7450 , \7448 , \7449 );
xor \U$7204 ( \7451 , \7444 , \7450 );
not \U$7205 ( \7452 , \7451 );
or \U$7206 ( \7453 , \7437 , \7452 );
nand \U$7207 ( \7454 , \7450 , \7444 );
nand \U$7208 ( \7455 , \7453 , \7454 );
not \U$7209 ( \7456 , \7455 );
not \U$7210 ( \7457 , \7456 );
or \U$7211 ( \7458 , \7421 , \7457 );
not \U$7212 ( \7459 , \7420 );
nand \U$7213 ( \7460 , \7459 , \7455 );
nand \U$7214 ( \7461 , \7458 , \7460 );
not \U$7215 ( \7462 , \7461 );
or \U$7216 ( \7463 , \7388 , \7462 );
nand \U$7217 ( \7464 , \7455 , \7420 );
nand \U$7218 ( \7465 , \7463 , \7464 );
and \U$7219 ( \7466 , RIbe2aa78_102, RIbe27b98_2);
not \U$7220 ( \7467 , \7466 );
xor \U$7221 ( \7468 , RIbe29ec0_77, RIbe28de0_41);
not \U$7222 ( \7469 , \7468 );
not \U$7223 ( \7470 , \923 );
or \U$7224 ( \7471 , \7469 , \7470 );
xor \U$7225 ( \7472 , RIbe27c10_3, RIbe28e58_42);
xor \U$7226 ( \7473 , RIbe29d58_74, RIbe28de0_41);
nand \U$7227 ( \7474 , \7472 , \7473 );
nand \U$7228 ( \7475 , \7471 , \7474 );
not \U$7229 ( \7476 , \7475 );
or \U$7230 ( \7477 , \7467 , \7476 );
or \U$7231 ( \7478 , \7475 , \7466 );
xor \U$7232 ( \7479 , RIbe28480_21, RIbe28a98_34);
not \U$7233 ( \7480 , \7479 );
not \U$7234 ( \7481 , \2518 );
or \U$7235 ( \7482 , \7480 , \7481 );
not \U$7236 ( \7483 , \2526 );
not \U$7237 ( \7484 , RIbe28480_21);
not \U$7238 ( \7485 , RIbe293f8_54);
and \U$7239 ( \7486 , \7484 , \7485 );
and \U$7240 ( \7487 , RIbe28480_21, RIbe293f8_54);
nor \U$7241 ( \7488 , \7486 , \7487 );
nand \U$7242 ( \7489 , \7483 , \7488 );
nand \U$7243 ( \7490 , \7482 , \7489 );
nand \U$7244 ( \7491 , \7478 , \7490 );
nand \U$7245 ( \7492 , \7477 , \7491 );
not \U$7246 ( \7493 , \7492 );
xor \U$7247 ( \7494 , RIbe27df0_7, RIbe296c8_60);
nand \U$7248 ( \7495 , \897 , \7494 );
not \U$7249 ( \7496 , \7495 );
not \U$7250 ( \7497 , \1937 );
and \U$7251 ( \7498 , \7496 , \7497 );
and \U$7252 ( \7499 , \907 , \7302 );
nor \U$7253 ( \7500 , \7498 , \7499 );
not \U$7254 ( \7501 , \7500 );
xor \U$7255 ( \7502 , RIbe28d68_40, RIbe29038_46);
nand \U$7256 ( \7503 , \276 , \7502 );
or \U$7257 ( \7504 , \7503 , \286 );
xor \U$7258 ( \7505 , RIbe27c88_4, RIbe29038_46);
nand \U$7259 ( \7506 , \284 , \7505 );
nand \U$7260 ( \7507 , \7504 , \7506 );
not \U$7261 ( \7508 , \7507 );
not \U$7262 ( \7509 , \7508 );
or \U$7263 ( \7510 , \7501 , \7509 );
xor \U$7264 ( \7511 , RIbe286d8_26, RIbe29c68_72);
not \U$7265 ( \7512 , \7511 );
not \U$7266 ( \7513 , \4576 );
not \U$7267 ( \7514 , \7513 );
or \U$7268 ( \7515 , \7512 , \7514 );
xor \U$7269 ( \7516 , RIbe27ee0_9, RIbe29c68_72);
nand \U$7270 ( \7517 , \4580 , \7516 );
nand \U$7271 ( \7518 , \7515 , \7517 );
nand \U$7272 ( \7519 , \7510 , \7518 );
not \U$7273 ( \7520 , \7500 );
nand \U$7274 ( \7521 , \7520 , \7507 );
and \U$7275 ( \7522 , \7519 , \7521 );
not \U$7276 ( \7523 , \7522 );
or \U$7277 ( \7524 , \7493 , \7523 );
or \U$7278 ( \7525 , \7492 , \7522 );
nand \U$7279 ( \7526 , \7524 , \7525 );
not \U$7280 ( \7527 , \7526 );
and \U$7281 ( \7528 , RIbe28840_29, RIbe28f48_44);
nor \U$7282 ( \7529 , RIbe28840_29, RIbe28f48_44);
nor \U$7283 ( \7530 , \7528 , \7529 );
not \U$7284 ( \7531 , \7530 );
not \U$7285 ( \7532 , \3256 );
or \U$7286 ( \7533 , \7531 , \7532 );
xor \U$7287 ( \7534 , RIbe28f48_44, RIbe28570_23);
nand \U$7288 ( \7535 , \3249 , \7534 );
nand \U$7289 ( \7536 , \7533 , \7535 );
not \U$7290 ( \7537 , \7536 );
xor \U$7291 ( \7538 , RIbe294e8_56, RIbe28390_19);
not \U$7292 ( \7539 , \7538 );
not \U$7293 ( \7540 , \2639 );
or \U$7294 ( \7541 , \7539 , \7540 );
xor \U$7295 ( \7542 , RIbe28390_19, RIbe288b8_30);
nand \U$7296 ( \7543 , \3714 , \7542 );
nand \U$7297 ( \7544 , \7541 , \7543 );
xor \U$7298 ( \7545 , RIbe28b88_36, RIbe282a0_17);
not \U$7299 ( \7546 , \7545 );
not \U$7300 ( \7547 , \2701 );
or \U$7301 ( \7548 , \7546 , \7547 );
buf \U$7302 ( \7549 , \2557 );
buf \U$7303 ( \7550 , \7549 );
nand \U$7304 ( \7551 , \7550 , \7279 );
nand \U$7305 ( \7552 , \7548 , \7551 );
and \U$7306 ( \7553 , \7544 , \7552 );
not \U$7307 ( \7554 , \7544 );
not \U$7308 ( \7555 , \7552 );
and \U$7309 ( \7556 , \7554 , \7555 );
nor \U$7310 ( \7557 , \7553 , \7556 );
not \U$7311 ( \7558 , \7557 );
or \U$7312 ( \7559 , \7537 , \7558 );
nand \U$7313 ( \7560 , \7552 , \7544 );
nand \U$7314 ( \7561 , \7559 , \7560 );
not \U$7315 ( \7562 , \7561 );
or \U$7316 ( \7563 , \7527 , \7562 );
not \U$7317 ( \7564 , \7522 );
nand \U$7318 ( \7565 , \7564 , \7492 );
nand \U$7319 ( \7566 , \7563 , \7565 );
xor \U$7320 ( \7567 , \7465 , \7566 );
not \U$7321 ( \7568 , \7567 );
not \U$7322 ( \7569 , \7488 );
not \U$7323 ( \7570 , \2519 );
or \U$7324 ( \7571 , \7569 , \7570 );
nand \U$7325 ( \7572 , \3075 , \4860 );
nand \U$7326 ( \7573 , \7571 , \7572 );
not \U$7327 ( \7574 , \7573 );
not \U$7328 ( \7575 , \7473 );
not \U$7329 ( \7576 , \331 );
or \U$7330 ( \7577 , \7575 , \7576 );
nand \U$7331 ( \7578 , \1149 , \4869 );
nand \U$7332 ( \7579 , \7577 , \7578 );
xor \U$7333 ( \7580 , RIbe29f38_78, RIbe27b98_2);
not \U$7334 ( \7581 , \7580 );
not \U$7335 ( \7582 , \1295 );
or \U$7336 ( \7583 , \7581 , \7582 );
buf \U$7337 ( \7584 , \266 );
buf \U$7338 ( \7585 , \7584 );
nand \U$7339 ( \7586 , \7585 , \4825 );
nand \U$7340 ( \7587 , \7583 , \7586 );
and \U$7341 ( \7588 , \7579 , \7587 );
not \U$7342 ( \7589 , \7579 );
not \U$7343 ( \7590 , \7587 );
and \U$7344 ( \7591 , \7589 , \7590 );
nor \U$7345 ( \7592 , \7588 , \7591 );
not \U$7346 ( \7593 , \7592 );
or \U$7347 ( \7594 , \7574 , \7593 );
nand \U$7348 ( \7595 , \7587 , \7579 );
nand \U$7349 ( \7596 , \7594 , \7595 );
not \U$7350 ( \7597 , \7542 );
not \U$7351 ( \7598 , \2639 );
or \U$7352 ( \7599 , \7597 , \7598 );
not \U$7353 ( \7600 , RIbe28390_19);
not \U$7354 ( \7601 , RIbe28a98_34);
and \U$7355 ( \7602 , \7600 , \7601 );
and \U$7356 ( \7603 , RIbe28390_19, RIbe28a98_34);
nor \U$7357 ( \7604 , \7602 , \7603 );
nand \U$7358 ( \7605 , \3714 , \7604 );
nand \U$7359 ( \7606 , \7599 , \7605 );
not \U$7360 ( \7607 , \7606 );
not \U$7361 ( \7608 , \7534 );
not \U$7362 ( \7609 , \3255 );
not \U$7363 ( \7610 , \7609 );
or \U$7364 ( \7611 , \7608 , \7610 );
and \U$7365 ( \7612 , RIbe286d8_26, RIbe28f48_44);
nor \U$7366 ( \7613 , RIbe286d8_26, RIbe28f48_44);
nor \U$7367 ( \7614 , \7612 , \7613 );
nand \U$7368 ( \7615 , \4181 , \7614 );
nand \U$7369 ( \7616 , \7611 , \7615 );
not \U$7370 ( \7617 , \7396 );
not \U$7371 ( \7618 , \2617 );
not \U$7372 ( \7619 , \7618 );
or \U$7373 ( \7620 , \7617 , \7619 );
nand \U$7374 ( \7621 , \2625 , \4800 );
nand \U$7375 ( \7622 , \7620 , \7621 );
and \U$7376 ( \7623 , \7616 , \7622 );
not \U$7377 ( \7624 , \7616 );
not \U$7378 ( \7625 , \7622 );
and \U$7379 ( \7626 , \7624 , \7625 );
nor \U$7380 ( \7627 , \7623 , \7626 );
not \U$7381 ( \7628 , \7627 );
or \U$7382 ( \7629 , \7607 , \7628 );
not \U$7383 ( \7630 , \7625 );
nand \U$7384 ( \7631 , \7630 , \7616 );
nand \U$7385 ( \7632 , \7629 , \7631 );
xor \U$7386 ( \7633 , \7596 , \7632 );
and \U$7387 ( \7634 , \2600 , \7354 );
and \U$7388 ( \7635 , \2603 , \4819 );
nor \U$7389 ( \7636 , \7634 , \7635 );
not \U$7390 ( \7637 , \7636 );
not \U$7391 ( \7638 , \7637 );
not \U$7392 ( \7639 , \7516 );
not \U$7393 ( \7640 , \4578 );
or \U$7394 ( \7641 , \7639 , \7640 );
buf \U$7395 ( \7642 , \4580 );
nand \U$7396 ( \7643 , \7642 , \7232 );
nand \U$7397 ( \7644 , \7641 , \7643 );
not \U$7398 ( \7645 , \7644 );
not \U$7399 ( \7646 , \1516 );
not \U$7400 ( \7647 , \4809 );
and \U$7401 ( \7648 , \7646 , \7647 );
and \U$7402 ( \7649 , \2380 , \7413 );
nor \U$7403 ( \7650 , \7648 , \7649 );
not \U$7404 ( \7651 , \7650 );
or \U$7405 ( \7652 , \7645 , \7651 );
or \U$7406 ( \7653 , \7644 , \7650 );
nand \U$7407 ( \7654 , \7652 , \7653 );
not \U$7408 ( \7655 , \7654 );
or \U$7409 ( \7656 , \7638 , \7655 );
not \U$7410 ( \7657 , \7650 );
nand \U$7411 ( \7658 , \7657 , \7644 );
nand \U$7412 ( \7659 , \7656 , \7658 );
xnor \U$7413 ( \7660 , \7633 , \7659 );
not \U$7414 ( \7661 , \7660 );
not \U$7415 ( \7662 , \7661 );
or \U$7416 ( \7663 , \7568 , \7662 );
nand \U$7417 ( \7664 , \7465 , \7566 );
nand \U$7418 ( \7665 , \7663 , \7664 );
not \U$7419 ( \7666 , \7665 );
and \U$7420 ( \7667 , \5048 , \5057 );
not \U$7421 ( \7668 , \5048 );
not \U$7422 ( \7669 , \5057 );
and \U$7423 ( \7670 , \7668 , \7669 );
nor \U$7424 ( \7671 , \7667 , \7670 );
xnor \U$7425 ( \7672 , \7671 , \5071 );
not \U$7426 ( \7673 , \7672 );
not \U$7427 ( \7674 , \4411 );
not \U$7428 ( \7675 , \4425 );
or \U$7429 ( \7676 , \7674 , \7675 );
or \U$7430 ( \7677 , \4425 , \4411 );
nand \U$7431 ( \7678 , \7676 , \7677 );
not \U$7432 ( \7679 , \7678 );
or \U$7433 ( \7680 , \7673 , \7679 );
or \U$7434 ( \7681 , \7678 , \7672 );
nand \U$7435 ( \7682 , \7680 , \7681 );
xor \U$7436 ( \7683 , \4379 , \4391 );
xor \U$7437 ( \7684 , \7683 , \4401 );
xnor \U$7438 ( \7685 , \7682 , \7684 );
not \U$7439 ( \7686 , \7685 );
not \U$7440 ( \7687 , \7659 );
not \U$7441 ( \7688 , \7633 );
or \U$7442 ( \7689 , \7687 , \7688 );
nand \U$7443 ( \7690 , \7596 , \7632 );
nand \U$7444 ( \7691 , \7689 , \7690 );
not \U$7445 ( \7692 , \4936 );
not \U$7446 ( \7693 , \4927 );
not \U$7447 ( \7694 , \7693 );
or \U$7448 ( \7695 , \7692 , \7694 );
or \U$7449 ( \7696 , \4936 , \7693 );
nand \U$7450 ( \7697 , \7695 , \7696 );
not \U$7451 ( \7698 , \7505 );
not \U$7452 ( \7699 , \281 );
or \U$7453 ( \7700 , \7698 , \7699 );
xor \U$7454 ( \7701 , RIbe29038_46, RIbe27df0_7);
nand \U$7455 ( \7702 , \287 , \7701 );
nand \U$7456 ( \7703 , \7700 , \7702 );
not \U$7457 ( \7704 , \7703 );
xor \U$7458 ( \7705 , RIbe27fd0_11, RIbe28750_27);
not \U$7459 ( \7706 , \7705 );
not \U$7460 ( \7707 , \3377 );
or \U$7461 ( \7708 , \7706 , \7707 );
not \U$7462 ( \7709 , \4896 );
nand \U$7463 ( \7710 , \7709 , \4891 );
nand \U$7464 ( \7711 , \7708 , \7710 );
not \U$7465 ( \7712 , \7711 );
or \U$7466 ( \7713 , \7704 , \7712 );
or \U$7467 ( \7714 , \7711 , \7703 );
not \U$7468 ( \7715 , \7369 );
not \U$7469 ( \7716 , \4841 );
not \U$7470 ( \7717 , \7716 );
or \U$7471 ( \7718 , \7715 , \7717 );
nand \U$7472 ( \7719 , \4850 , RIbe29e48_76);
nand \U$7473 ( \7720 , \7718 , \7719 );
nand \U$7474 ( \7721 , \7714 , \7720 );
nand \U$7475 ( \7722 , \7713 , \7721 );
not \U$7476 ( \7723 , \7722 );
nand \U$7477 ( \7724 , \7723 , \7285 );
not \U$7478 ( \7725 , \7724 );
not \U$7479 ( \7726 , \7434 );
not \U$7480 ( \7727 , \966 );
or \U$7481 ( \7728 , \7726 , \7727 );
nand \U$7482 ( \7729 , \1797 , \4905 );
nand \U$7483 ( \7730 , \7728 , \7729 );
not \U$7484 ( \7731 , \7730 );
xor \U$7485 ( \7732 , RIbe28cf0_39, RIbe27d78_6);
not \U$7486 ( \7733 , \7732 );
not \U$7487 ( \7734 , \1164 );
or \U$7488 ( \7735 , \7733 , \7734 );
nand \U$7489 ( \7736 , \314 , \4919 );
nand \U$7490 ( \7737 , \7735 , \7736 );
not \U$7491 ( \7738 , \7404 );
not \U$7492 ( \7739 , \2730 );
or \U$7493 ( \7740 , \7738 , \7739 );
xor \U$7494 ( \7741 , RIbe28d68_40, RIbe290b0_47);
nand \U$7495 ( \7742 , \398 , \7741 );
nand \U$7496 ( \7743 , \7740 , \7742 );
xor \U$7497 ( \7744 , \7737 , \7743 );
not \U$7498 ( \7745 , \7744 );
or \U$7499 ( \7746 , \7731 , \7745 );
nand \U$7500 ( \7747 , \7737 , \7743 );
nand \U$7501 ( \7748 , \7746 , \7747 );
not \U$7502 ( \7749 , \7748 );
or \U$7503 ( \7750 , \7725 , \7749 );
not \U$7504 ( \7751 , \7285 );
nand \U$7505 ( \7752 , \7722 , \7751 );
nand \U$7506 ( \7753 , \7750 , \7752 );
and \U$7507 ( \7754 , \7697 , \7753 );
not \U$7508 ( \7755 , \7697 );
not \U$7509 ( \7756 , \7753 );
and \U$7510 ( \7757 , \7755 , \7756 );
nor \U$7511 ( \7758 , \7754 , \7757 );
xor \U$7512 ( \7759 , \7691 , \7758 );
not \U$7513 ( \7760 , \7759 );
not \U$7514 ( \7761 , \7760 );
or \U$7515 ( \7762 , \7686 , \7761 );
not \U$7516 ( \7763 , \7685 );
nand \U$7517 ( \7764 , \7763 , \7759 );
nand \U$7518 ( \7765 , \7762 , \7764 );
not \U$7519 ( \7766 , \7765 );
or \U$7520 ( \7767 , \7666 , \7766 );
nand \U$7521 ( \7768 , \7759 , \7685 );
nand \U$7522 ( \7769 , \7767 , \7768 );
xor \U$7523 ( \7770 , \7345 , \7769 );
not \U$7524 ( \7771 , \7770 );
not \U$7525 ( \7772 , \7604 );
not \U$7526 ( \7773 , \2640 );
or \U$7527 ( \7774 , \7772 , \7773 );
nand \U$7528 ( \7775 , \5831 , \5005 );
nand \U$7529 ( \7776 , \7774 , \7775 );
not \U$7530 ( \7777 , \7701 );
not \U$7531 ( \7778 , \979 );
or \U$7532 ( \7779 , \7777 , \7778 );
nand \U$7533 ( \7780 , \1805 , \4393 );
nand \U$7534 ( \7781 , \7779 , \7780 );
xor \U$7535 ( \7782 , \7776 , \7781 );
not \U$7536 ( \7783 , \7614 );
not \U$7537 ( \7784 , \3256 );
or \U$7538 ( \7785 , \7783 , \7784 );
nand \U$7539 ( \7786 , \4181 , \4384 );
nand \U$7540 ( \7787 , \7785 , \7786 );
not \U$7541 ( \7788 , \7787 );
and \U$7542 ( \7789 , \7782 , \7788 );
not \U$7543 ( \7790 , \7782 );
and \U$7544 ( \7791 , \7790 , \7787 );
nor \U$7545 ( \7792 , \7789 , \7791 );
not \U$7546 ( \7793 , \7272 );
not \U$7547 ( \7794 , \1779 );
not \U$7548 ( \7795 , \7794 );
not \U$7549 ( \7796 , \7795 );
or \U$7550 ( \7797 , \7793 , \7796 );
nand \U$7551 ( \7798 , \2475 , \5050 );
nand \U$7552 ( \7799 , \7797 , \7798 );
not \U$7553 ( \7800 , \7313 );
not \U$7554 ( \7801 , \1103 );
or \U$7555 ( \7802 , \7800 , \7801 );
nand \U$7556 ( \7803 , \369 , \4929 );
nand \U$7557 ( \7804 , \7802 , \7803 );
xor \U$7558 ( \7805 , \7799 , \7804 );
not \U$7559 ( \7806 , \7741 );
not \U$7560 ( \7807 , \466 );
or \U$7561 ( \7808 , \7806 , \7807 );
nand \U$7562 ( \7809 , \2071 , \5065 );
nand \U$7563 ( \7810 , \7808 , \7809 );
xnor \U$7564 ( \7811 , \7805 , \7810 );
and \U$7565 ( \7812 , \7792 , \7811 );
xor \U$7566 ( \7813 , \4925 , \4899 );
not \U$7567 ( \7814 , \4915 );
xor \U$7568 ( \7815 , \7813 , \7814 );
nor \U$7569 ( \7816 , \7812 , \7815 );
nor \U$7570 ( \7817 , \7792 , \7811 );
nor \U$7571 ( \7818 , \7816 , \7817 );
not \U$7572 ( \7819 , \7818 );
not \U$7573 ( \7820 , \7819 );
xor \U$7574 ( \7821 , \4884 , \4816 );
not \U$7575 ( \7822 , \7821 );
not \U$7576 ( \7823 , \7776 );
not \U$7577 ( \7824 , \7781 );
or \U$7578 ( \7825 , \7823 , \7824 );
nand \U$7579 ( \7826 , \7782 , \7787 );
nand \U$7580 ( \7827 , \7825 , \7826 );
not \U$7581 ( \7828 , \7810 );
xor \U$7582 ( \7829 , \7799 , \7804 );
not \U$7583 ( \7830 , \7829 );
or \U$7584 ( \7831 , \7828 , \7830 );
nand \U$7585 ( \7832 , \7799 , \7804 );
nand \U$7586 ( \7833 , \7831 , \7832 );
not \U$7587 ( \7834 , \7260 );
or \U$7588 ( \7835 , \7834 , \7246 );
nand \U$7589 ( \7836 , \7835 , \7248 );
xor \U$7590 ( \7837 , \7833 , \7836 );
xor \U$7591 ( \7838 , \7827 , \7837 );
not \U$7592 ( \7839 , \7838 );
or \U$7593 ( \7840 , \7822 , \7839 );
or \U$7594 ( \7841 , \7838 , \7821 );
nand \U$7595 ( \7842 , \7840 , \7841 );
not \U$7596 ( \7843 , \7842 );
or \U$7597 ( \7844 , \7820 , \7843 );
not \U$7598 ( \7845 , \7821 );
nand \U$7599 ( \7846 , \7845 , \7838 );
nand \U$7600 ( \7847 , \7844 , \7846 );
nand \U$7601 ( \7848 , \7758 , \7691 );
nand \U$7602 ( \7849 , \7753 , \7697 );
and \U$7603 ( \7850 , \7848 , \7849 );
xor \U$7604 ( \7851 , \4772 , \4775 );
xor \U$7605 ( \7852 , \7851 , \4779 );
xnor \U$7606 ( \7853 , \7850 , \7852 );
xor \U$7607 ( \7854 , \7847 , \7853 );
not \U$7608 ( \7855 , \7854 );
not \U$7609 ( \7856 , \7855 );
or \U$7610 ( \7857 , \7771 , \7856 );
nand \U$7611 ( \7858 , \7769 , \7345 );
nand \U$7612 ( \7859 , \7857 , \7858 );
not \U$7613 ( \7860 , \7859 );
xnor \U$7614 ( \7861 , \4463 , \4404 );
not \U$7615 ( \7862 , \7684 );
not \U$7616 ( \7863 , \7862 );
not \U$7617 ( \7864 , \7682 );
or \U$7618 ( \7865 , \7863 , \7864 );
not \U$7619 ( \7866 , \7672 );
nand \U$7620 ( \7867 , \7866 , \7678 );
nand \U$7621 ( \7868 , \7865 , \7867 );
xor \U$7622 ( \7869 , \7861 , \7868 );
not \U$7623 ( \7870 , \7869 );
xor \U$7624 ( \7871 , \4761 , \4763 );
xor \U$7625 ( \7872 , \7871 , \4768 );
not \U$7626 ( \7873 , \7872 );
and \U$7627 ( \7874 , \7870 , \7873 );
and \U$7628 ( \7875 , \7869 , \7872 );
nor \U$7629 ( \7876 , \7874 , \7875 );
not \U$7630 ( \7877 , \7876 );
not \U$7631 ( \7878 , \7877 );
not \U$7632 ( \7879 , \4889 );
not \U$7633 ( \7880 , \4943 );
and \U$7634 ( \7881 , \7879 , \7880 );
and \U$7635 ( \7882 , \4889 , \4943 );
nor \U$7636 ( \7883 , \7881 , \7882 );
not \U$7637 ( \7884 , \7883 );
not \U$7638 ( \7885 , \7213 );
not \U$7639 ( \7886 , \7211 );
or \U$7640 ( \7887 , \7885 , \7886 );
not \U$7641 ( \7888 , \7204 );
nand \U$7642 ( \7889 , \7888 , \7207 );
nand \U$7643 ( \7890 , \7887 , \7889 );
not \U$7644 ( \7891 , \7890 );
not \U$7645 ( \7892 , \7827 );
not \U$7646 ( \7893 , \7837 );
or \U$7647 ( \7894 , \7892 , \7893 );
nand \U$7648 ( \7895 , \7833 , \7836 );
nand \U$7649 ( \7896 , \7894 , \7895 );
not \U$7650 ( \7897 , \7896 );
xor \U$7651 ( \7898 , \5073 , \5042 );
xor \U$7652 ( \7899 , \7897 , \7898 );
not \U$7653 ( \7900 , \7899 );
or \U$7654 ( \7901 , \7891 , \7900 );
or \U$7655 ( \7902 , \7890 , \7899 );
nand \U$7656 ( \7903 , \7901 , \7902 );
not \U$7657 ( \7904 , \7903 );
or \U$7658 ( \7905 , \7884 , \7904 );
or \U$7659 ( \7906 , \7903 , \7883 );
nand \U$7660 ( \7907 , \7905 , \7906 );
not \U$7661 ( \7908 , \7907 );
or \U$7662 ( \7909 , \7878 , \7908 );
not \U$7663 ( \7910 , \7883 );
nand \U$7664 ( \7911 , \7910 , \7903 );
nand \U$7665 ( \7912 , \7909 , \7911 );
not \U$7666 ( \7913 , \7912 );
xnor \U$7667 ( \7914 , \4771 , \4783 );
xor \U$7668 ( \7915 , \4786 , \7914 );
not \U$7669 ( \7916 , \4984 );
not \U$7670 ( \7917 , \5082 );
or \U$7671 ( \7918 , \7916 , \7917 );
or \U$7672 ( \7919 , \5082 , \4984 );
nand \U$7673 ( \7920 , \7918 , \7919 );
not \U$7674 ( \7921 , \7890 );
not \U$7675 ( \7922 , \7899 );
not \U$7676 ( \7923 , \7922 );
or \U$7677 ( \7924 , \7921 , \7923 );
not \U$7678 ( \7925 , \7897 );
nand \U$7679 ( \7926 , \7925 , \7898 );
nand \U$7680 ( \7927 , \7924 , \7926 );
not \U$7681 ( \7928 , \7927 );
and \U$7682 ( \7929 , \7920 , \7928 );
not \U$7683 ( \7930 , \7920 );
and \U$7684 ( \7931 , \7930 , \7927 );
or \U$7685 ( \7932 , \7929 , \7931 );
xor \U$7686 ( \7933 , \7915 , \7932 );
not \U$7687 ( \7934 , \7933 );
not \U$7688 ( \7935 , \7934 );
or \U$7689 ( \7936 , \7913 , \7935 );
not \U$7690 ( \7937 , \7912 );
nand \U$7691 ( \7938 , \7933 , \7937 );
nand \U$7692 ( \7939 , \7936 , \7938 );
not \U$7693 ( \7940 , \7939 );
or \U$7694 ( \7941 , \7860 , \7940 );
nand \U$7695 ( \7942 , \7933 , \7912 );
nand \U$7696 ( \7943 , \7941 , \7942 );
xor \U$7697 ( \7944 , \7203 , \7943 );
not \U$7698 ( \7945 , \7915 );
not \U$7699 ( \7946 , \7932 );
or \U$7700 ( \7947 , \7945 , \7946 );
nand \U$7701 ( \7948 , \7920 , \7927 );
nand \U$7702 ( \7949 , \7947 , \7948 );
not \U$7703 ( \7950 , \5092 );
not \U$7704 ( \7951 , \4975 );
and \U$7705 ( \7952 , \7950 , \7951 );
and \U$7706 ( \7953 , \5092 , \4975 );
nor \U$7707 ( \7954 , \7952 , \7953 );
and \U$7708 ( \7955 , \7949 , \7954 );
not \U$7709 ( \7956 , \7949 );
not \U$7710 ( \7957 , \7954 );
and \U$7711 ( \7958 , \7956 , \7957 );
or \U$7712 ( \7959 , \7955 , \7958 );
not \U$7713 ( \7960 , \7847 );
or \U$7714 ( \7961 , \7960 , \7853 );
or \U$7715 ( \7962 , \7850 , \7852 );
nand \U$7716 ( \7963 , \7961 , \7962 );
not \U$7717 ( \7964 , \7963 );
not \U$7718 ( \7965 , \7868 );
not \U$7719 ( \7966 , \7861 );
or \U$7720 ( \7967 , \7965 , \7966 );
not \U$7721 ( \7968 , \7872 );
nand \U$7722 ( \7969 , \7968 , \7869 );
nand \U$7723 ( \7970 , \7967 , \7969 );
not \U$7724 ( \7971 , \4947 );
and \U$7725 ( \7972 , \4957 , \7971 );
not \U$7726 ( \7973 , \4957 );
and \U$7727 ( \7974 , \7973 , \4947 );
nor \U$7728 ( \7975 , \7972 , \7974 );
xnor \U$7729 ( \7976 , \7970 , \7975 );
not \U$7730 ( \7977 , \7976 );
or \U$7731 ( \7978 , \7964 , \7977 );
not \U$7732 ( \7979 , \7975 );
nand \U$7733 ( \7980 , \7979 , \7970 );
nand \U$7734 ( \7981 , \7978 , \7980 );
and \U$7735 ( \7982 , \7959 , \7981 );
not \U$7736 ( \7983 , \7959 );
not \U$7737 ( \7984 , \7981 );
and \U$7738 ( \7985 , \7983 , \7984 );
nor \U$7739 ( \7986 , \7982 , \7985 );
xnor \U$7740 ( \7987 , \7944 , \7986 );
not \U$7741 ( \7988 , \7876 );
not \U$7742 ( \7989 , \7907 );
or \U$7743 ( \7990 , \7988 , \7989 );
or \U$7744 ( \7991 , \7907 , \7876 );
nand \U$7745 ( \7992 , \7990 , \7991 );
not \U$7746 ( \7993 , \7992 );
xnor \U$7747 ( \7994 , \7324 , \7307 );
not \U$7748 ( \7995 , \7994 );
not \U$7749 ( \7996 , \7995 );
xnor \U$7750 ( \7997 , \7627 , \7606 );
not \U$7751 ( \7998 , \7997 );
and \U$7752 ( \7999 , \7744 , \7730 );
not \U$7753 ( \8000 , \7744 );
not \U$7754 ( \8001 , \7730 );
and \U$7755 ( \8002 , \8000 , \8001 );
nor \U$7756 ( \8003 , \7999 , \8002 );
not \U$7757 ( \8004 , \8003 );
or \U$7758 ( \8005 , \7998 , \8004 );
or \U$7759 ( \8006 , \8003 , \7997 );
nand \U$7760 ( \8007 , \8005 , \8006 );
not \U$7761 ( \8008 , \8007 );
or \U$7762 ( \8009 , \7996 , \8008 );
not \U$7763 ( \8010 , \7997 );
nand \U$7764 ( \8011 , \8010 , \8003 );
nand \U$7765 ( \8012 , \8009 , \8011 );
not \U$7766 ( \8013 , \8012 );
xnor \U$7767 ( \8014 , RIbe284f8_22, RIbe27fd0_11);
or \U$7768 ( \8015 , \2717 , \8014 );
not \U$7769 ( \8016 , \7705 );
or \U$7770 ( \8017 , \2708 , \8016 );
nand \U$7771 ( \8018 , \8015 , \8017 );
xor \U$7772 ( \8019 , RIbe27d78_6, RIbe27b20_1);
not \U$7773 ( \8020 , \8019 );
not \U$7774 ( \8021 , \1164 );
or \U$7775 ( \8022 , \8020 , \8021 );
nand \U$7776 ( \8023 , \315 , \7732 );
nand \U$7777 ( \8024 , \8022 , \8023 );
xor \U$7778 ( \8025 , \8018 , \8024 );
not \U$7779 ( \8026 , \7580 );
not \U$7780 ( \8027 , \1298 );
or \U$7781 ( \8028 , \8026 , \8027 );
xnor \U$7782 ( \8029 , RIbe27b98_2, RIbe2b6a8_128);
or \U$7783 ( \8030 , \257 , \8029 );
nand \U$7784 ( \8031 , \8028 , \8030 );
and \U$7785 ( \8032 , \8025 , \8031 );
and \U$7786 ( \8033 , \8018 , \8024 );
or \U$7787 ( \8034 , \8032 , \8033 );
not \U$7788 ( \8035 , \8034 );
xor \U$7789 ( \8036 , \7592 , \7573 );
not \U$7790 ( \8037 , \8036 );
or \U$7791 ( \8038 , \8035 , \8037 );
or \U$7792 ( \8039 , \8034 , \8036 );
xor \U$7793 ( \8040 , \7720 , \7711 );
xor \U$7794 ( \8041 , \8040 , \7703 );
nand \U$7795 ( \8042 , \8039 , \8041 );
nand \U$7796 ( \8043 , \8038 , \8042 );
not \U$7797 ( \8044 , \8043 );
xor \U$7798 ( \8045 , \7751 , \7722 );
xnor \U$7799 ( \8046 , \8045 , \7748 );
not \U$7800 ( \8047 , \8046 );
or \U$7801 ( \8048 , \8044 , \8047 );
or \U$7802 ( \8049 , \8043 , \8046 );
nand \U$7803 ( \8050 , \8048 , \8049 );
not \U$7804 ( \8051 , \8050 );
or \U$7805 ( \8052 , \8013 , \8051 );
not \U$7806 ( \8053 , \8046 );
nand \U$7807 ( \8054 , \8053 , \8043 );
nand \U$7808 ( \8055 , \8052 , \8054 );
not \U$7809 ( \8056 , \8055 );
not \U$7810 ( \8057 , \8056 );
xor \U$7811 ( \8058 , \7818 , \7821 );
xnor \U$7812 ( \8059 , \8058 , \7838 );
not \U$7813 ( \8060 , \8059 );
or \U$7814 ( \8061 , \8057 , \8060 );
xor \U$7815 ( \8062 , \7792 , \7815 );
xnor \U$7816 ( \8063 , \8062 , \7811 );
not \U$7817 ( \8064 , \8063 );
xor \U$7818 ( \8065 , \7336 , \7329 );
xor \U$7819 ( \8066 , \7230 , \7298 );
xnor \U$7820 ( \8067 , \8066 , \7291 );
and \U$7821 ( \8068 , \8065 , \8067 );
not \U$7822 ( \8069 , \8065 );
not \U$7823 ( \8070 , \8067 );
and \U$7824 ( \8071 , \8069 , \8070 );
or \U$7825 ( \8072 , \8068 , \8071 );
not \U$7826 ( \8073 , \8072 );
or \U$7827 ( \8074 , \8064 , \8073 );
nand \U$7828 ( \8075 , \8070 , \8065 );
nand \U$7829 ( \8076 , \8074 , \8075 );
nand \U$7830 ( \8077 , \8061 , \8076 );
or \U$7831 ( \8078 , \8056 , \8059 );
and \U$7832 ( \8079 , \8077 , \8078 );
nand \U$7833 ( \8080 , \7993 , \8079 );
not \U$7834 ( \8081 , \8080 );
xor \U$7835 ( \8082 , \7345 , \7769 );
xor \U$7836 ( \8083 , \8082 , \7854 );
not \U$7837 ( \8084 , \8083 );
not \U$7838 ( \8085 , \8084 );
or \U$7839 ( \8086 , \8081 , \8085 );
not \U$7840 ( \8087 , \8079 );
nand \U$7841 ( \8088 , \8087 , \7992 );
nand \U$7842 ( \8089 , \8086 , \8088 );
not \U$7843 ( \8090 , \8089 );
not \U$7844 ( \8091 , \8090 );
xnor \U$7845 ( \8092 , \7976 , \7963 );
not \U$7846 ( \8093 , \8092 );
xor \U$7847 ( \8094 , \7859 , \7939 );
not \U$7848 ( \8095 , \8094 );
or \U$7849 ( \8096 , \8093 , \8095 );
or \U$7850 ( \8097 , \8094 , \8092 );
nand \U$7851 ( \8098 , \8096 , \8097 );
nand \U$7852 ( \8099 , \8091 , \8098 );
not \U$7853 ( \8100 , \8092 );
nand \U$7854 ( \8101 , \8100 , \8094 );
and \U$7855 ( \8102 , \8099 , \8101 );
nand \U$7856 ( \8103 , \7987 , \8102 );
xor \U$7857 ( \8104 , \4320 , \4496 );
not \U$7858 ( \8105 , \7981 );
not \U$7859 ( \8106 , \7959 );
or \U$7860 ( \8107 , \8105 , \8106 );
nand \U$7861 ( \8108 , \7957 , \7949 );
nand \U$7862 ( \8109 , \8107 , \8108 );
xor \U$7863 ( \8110 , \8104 , \8109 );
not \U$7864 ( \8111 , \8110 );
not \U$7865 ( \8112 , \5098 );
nand \U$7866 ( \8113 , \8112 , \5102 );
and \U$7867 ( \8114 , \8113 , \4967 );
not \U$7868 ( \8115 , \8113 );
not \U$7869 ( \8116 , \4967 );
and \U$7870 ( \8117 , \8115 , \8116 );
nor \U$7871 ( \8118 , \8114 , \8117 );
not \U$7872 ( \8119 , \8118 );
and \U$7873 ( \8120 , \8111 , \8119 );
and \U$7874 ( \8121 , \8110 , \8118 );
nor \U$7875 ( \8122 , \8120 , \8121 );
buf \U$7876 ( \8123 , \7203 );
xor \U$7877 ( \8124 , \8123 , \7943 );
and \U$7878 ( \8125 , \8124 , \7986 );
and \U$7879 ( \8126 , \8123 , \7943 );
nor \U$7880 ( \8127 , \8125 , \8126 );
nand \U$7881 ( \8128 , \8122 , \8127 );
xor \U$7882 ( \8129 , \8056 , \8059 );
xnor \U$7883 ( \8130 , \8129 , \8076 );
xnor \U$7884 ( \8131 , \8050 , \8012 );
not \U$7885 ( \8132 , \8131 );
and \U$7886 ( \8133 , \7382 , \7357 );
not \U$7887 ( \8134 , \7382 );
and \U$7888 ( \8135 , \8134 , \7356 );
or \U$7889 ( \8136 , \8133 , \8135 );
not \U$7890 ( \8137 , \8136 );
not \U$7891 ( \8138 , \8137 );
xor \U$7892 ( \8139 , \8018 , \8024 );
xor \U$7893 ( \8140 , \8139 , \8031 );
not \U$7894 ( \8141 , \8140 );
not \U$7895 ( \8142 , \7536 );
buf \U$7896 ( \8143 , \7557 );
xor \U$7897 ( \8144 , \8142 , \8143 );
not \U$7898 ( \8145 , \8144 );
or \U$7899 ( \8146 , \8141 , \8145 );
or \U$7900 ( \8147 , \8144 , \8140 );
nand \U$7901 ( \8148 , \8146 , \8147 );
not \U$7902 ( \8149 , \8148 );
or \U$7903 ( \8150 , \8138 , \8149 );
not \U$7904 ( \8151 , \8144 );
nand \U$7905 ( \8152 , \8151 , \8140 );
nand \U$7906 ( \8153 , \8150 , \8152 );
not \U$7907 ( \8154 , \8153 );
xor \U$7908 ( \8155 , RIbe28b88_36, RIbe28138_14);
not \U$7909 ( \8156 , \8155 );
not \U$7910 ( \8157 , \2554 );
or \U$7911 ( \8158 , \8156 , \8157 );
nand \U$7912 ( \8159 , \2691 , \7545 );
nand \U$7913 ( \8160 , \8158 , \8159 );
not \U$7914 ( \8161 , RIbe2a028_80);
nor \U$7915 ( \8162 , RIbe2a2f8_86, RIbe2acd0_107);
not \U$7916 ( \8163 , \8162 );
or \U$7917 ( \8164 , \8161 , \8163 );
not \U$7918 ( \8165 , RIbe2a028_80);
nand \U$7919 ( \8166 , \8165 , RIbe2a2f8_86, RIbe2acd0_107);
nand \U$7920 ( \8167 , \8164 , \8166 );
buf \U$7921 ( \8168 , \8167 );
buf \U$7922 ( \8169 , \8168 );
buf \U$7923 ( \8170 , \8169 );
xor \U$7924 ( \8171 , RIbe2a2f8_86, RIbe2acd0_107);
buf \U$7925 ( \8172 , \8171 );
or \U$7926 ( \8173 , \8170 , \8172 );
nand \U$7927 ( \8174 , \8173 , RIbe2a028_80);
nor \U$7928 ( \8175 , \8160 , \8174 );
not \U$7929 ( \8176 , \8175 );
not \U$7930 ( \8177 , \8176 );
not \U$7931 ( \8178 , RIbe27e68_8);
not \U$7932 ( \8179 , RIbe28c00_37);
and \U$7933 ( \8180 , \8178 , \8179 );
and \U$7934 ( \8181 , RIbe27e68_8, RIbe28c00_37);
nor \U$7935 ( \8182 , \8180 , \8181 );
not \U$7936 ( \8183 , \8182 );
not \U$7937 ( \8184 , \2600 );
or \U$7938 ( \8185 , \8183 , \8184 );
nand \U$7939 ( \8186 , \2464 , \7350 );
nand \U$7940 ( \8187 , \8185 , \8186 );
not \U$7941 ( \8188 , \8187 );
and \U$7942 ( \8189 , RIbe2aa00_101, RIbe27b98_2);
xor \U$7943 ( \8190 , RIbe28a20_33, RIbe29740_61);
not \U$7944 ( \8191 , \8190 );
not \U$7945 ( \8192 , \1781 );
or \U$7946 ( \8193 , \8191 , \8192 );
nand \U$7947 ( \8194 , \5055 , \7445 );
nand \U$7948 ( \8195 , \8193 , \8194 );
xor \U$7949 ( \8196 , \8189 , \8195 );
not \U$7950 ( \8197 , \8196 );
or \U$7951 ( \8198 , \8188 , \8197 );
nand \U$7952 ( \8199 , \8195 , \8189 );
nand \U$7953 ( \8200 , \8198 , \8199 );
not \U$7954 ( \8201 , \8200 );
or \U$7955 ( \8202 , \8177 , \8201 );
nand \U$7956 ( \8203 , \8160 , \8174 );
nand \U$7957 ( \8204 , \8202 , \8203 );
not \U$7958 ( \8205 , \8204 );
xor \U$7959 ( \8206 , RIbe29470_55, RIbe28390_19);
not \U$7960 ( \8207 , \8206 );
or \U$7961 ( \8208 , \2774 , \8207 );
not \U$7962 ( \8209 , \7538 );
or \U$7963 ( \8210 , \2778 , \8209 );
nand \U$7964 ( \8211 , \8208 , \8210 );
not \U$7965 ( \8212 , \8211 );
xor \U$7966 ( \8213 , RIbe29998_66, RIbe29038_46);
not \U$7967 ( \8214 , \8213 );
or \U$7968 ( \8215 , \2388 , \8214 );
not \U$7969 ( \8216 , \7502 );
or \U$7970 ( \8217 , \1465 , \8216 );
nand \U$7971 ( \8218 , \8215 , \8217 );
xor \U$7972 ( \8219 , RIbe28f48_44, RIbe28750_27);
not \U$7973 ( \8220 , \8219 );
not \U$7974 ( \8221 , \3255 );
not \U$7975 ( \8222 , \8221 );
or \U$7976 ( \8223 , \8220 , \8222 );
nand \U$7977 ( \8224 , \3249 , \7530 );
nand \U$7978 ( \8225 , \8223 , \8224 );
xor \U$7979 ( \8226 , \8218 , \8225 );
not \U$7980 ( \8227 , \8226 );
or \U$7981 ( \8228 , \8212 , \8227 );
nand \U$7982 ( \8229 , \8225 , \8218 );
nand \U$7983 ( \8230 , \8228 , \8229 );
not \U$7984 ( \8231 , \8230 );
xor \U$7985 ( \8232 , RIbe27d78_6, RIbe29b78_70);
not \U$7986 ( \8233 , \8232 );
not \U$7987 ( \8234 , \1043 );
or \U$7988 ( \8235 , \8233 , \8234 );
nand \U$7989 ( \8236 , \314 , \8019 );
nand \U$7990 ( \8237 , \8235 , \8236 );
and \U$7991 ( \8238 , RIbe29e48_76, RIbe27ee0_9);
not \U$7992 ( \8239 , RIbe29e48_76);
and \U$7993 ( \8240 , \8239 , \317 );
nor \U$7994 ( \8241 , \8238 , \8240 );
not \U$7995 ( \8242 , \8241 );
not \U$7996 ( \8243 , \7372 );
or \U$7997 ( \8244 , \8242 , \8243 );
buf \U$7998 ( \8245 , \4849 );
nand \U$7999 ( \8246 , \8245 , \7376 );
nand \U$8000 ( \8247 , \8244 , \8246 );
xor \U$8001 ( \8248 , \8237 , \8247 );
xnor \U$8002 ( \8249 , RIbe28318_18, RIbe27fd0_11);
or \U$8003 ( \8250 , \2718 , \8249 );
or \U$8004 ( \8251 , \2708 , \8014 );
nand \U$8005 ( \8252 , \8250 , \8251 );
and \U$8006 ( \8253 , \8248 , \8252 );
and \U$8007 ( \8254 , \8237 , \8247 );
nor \U$8008 ( \8255 , \8253 , \8254 );
not \U$8009 ( \8256 , \8255 );
xor \U$8010 ( \8257 , RIbe29c68_72, RIbe28570_23);
not \U$8011 ( \8258 , \8257 );
not \U$8012 ( \8259 , \4576 );
not \U$8013 ( \8260 , \8259 );
or \U$8014 ( \8261 , \8258 , \8260 );
nand \U$8015 ( \8262 , \4580 , \7511 );
nand \U$8016 ( \8263 , \8261 , \8262 );
not \U$8017 ( \8264 , \8263 );
xor \U$8018 ( \8265 , RIbe293f8_54, RIbe285e8_24);
not \U$8019 ( \8266 , \8265 );
not \U$8020 ( \8267 , \2617 );
not \U$8021 ( \8268 , \8267 );
or \U$8022 ( \8269 , \8266 , \8268 );
buf \U$8023 ( \8270 , \2623 );
nand \U$8024 ( \8271 , \8270 , \7392 );
nand \U$8025 ( \8272 , \8269 , \8271 );
not \U$8026 ( \8273 , \8272 );
not \U$8027 ( \8274 , \8273 );
xor \U$8028 ( \8275 , RIbe29218_50, RIbe280c0_13);
not \U$8029 ( \8276 , \8275 );
not \U$8030 ( \8277 , \1053 );
or \U$8031 ( \8278 , \8276 , \8277 );
nand \U$8032 ( \8279 , \869 , \7407 );
nand \U$8033 ( \8280 , \8278 , \8279 );
not \U$8034 ( \8281 , \8280 );
or \U$8035 ( \8282 , \8274 , \8281 );
or \U$8036 ( \8283 , \8280 , \8273 );
nand \U$8037 ( \8284 , \8282 , \8283 );
not \U$8038 ( \8285 , \8284 );
or \U$8039 ( \8286 , \8264 , \8285 );
nand \U$8040 ( \8287 , \8272 , \8280 );
nand \U$8041 ( \8288 , \8286 , \8287 );
not \U$8042 ( \8289 , \8288 );
or \U$8043 ( \8290 , \8256 , \8289 );
or \U$8044 ( \8291 , \8255 , \8288 );
nand \U$8045 ( \8292 , \8290 , \8291 );
not \U$8046 ( \8293 , \8292 );
or \U$8047 ( \8294 , \8231 , \8293 );
not \U$8048 ( \8295 , \8255 );
nand \U$8049 ( \8296 , \8295 , \8288 );
nand \U$8050 ( \8297 , \8294 , \8296 );
xnor \U$8051 ( \8298 , \8205 , \8297 );
not \U$8052 ( \8299 , \8298 );
or \U$8053 ( \8300 , \8154 , \8299 );
not \U$8054 ( \8301 , \8205 );
nand \U$8055 ( \8302 , \8301 , \8297 );
nand \U$8056 ( \8303 , \8300 , \8302 );
not \U$8057 ( \8304 , \8303 );
or \U$8058 ( \8305 , \8132 , \8304 );
or \U$8059 ( \8306 , \8303 , \8131 );
nand \U$8060 ( \8307 , \8305 , \8306 );
not \U$8061 ( \8308 , \8307 );
xor \U$8062 ( \8309 , \8063 , \8072 );
not \U$8063 ( \8310 , \8309 );
or \U$8064 ( \8311 , \8308 , \8310 );
not \U$8065 ( \8312 , \8131 );
nand \U$8066 ( \8313 , \8312 , \8303 );
nand \U$8067 ( \8314 , \8311 , \8313 );
not \U$8068 ( \8315 , \8314 );
xor \U$8069 ( \8316 , \8130 , \8315 );
not \U$8070 ( \8317 , \7340 );
not \U$8071 ( \8318 , \7218 );
and \U$8072 ( \8319 , \8317 , \8318 );
and \U$8073 ( \8320 , \7340 , \7218 );
nor \U$8074 ( \8321 , \8319 , \8320 );
not \U$8075 ( \8322 , \7660 );
not \U$8076 ( \8323 , \7567 );
or \U$8077 ( \8324 , \8322 , \8323 );
or \U$8078 ( \8325 , \7660 , \7567 );
nand \U$8079 ( \8326 , \8324 , \8325 );
not \U$8080 ( \8327 , \8326 );
xnor \U$8081 ( \8328 , \7286 , \7274 );
not \U$8082 ( \8329 , \8328 );
not \U$8083 ( \8330 , \7637 );
not \U$8084 ( \8331 , \7654 );
not \U$8085 ( \8332 , \8331 );
or \U$8086 ( \8333 , \8330 , \8332 );
nand \U$8087 ( \8334 , \7654 , \7636 );
nand \U$8088 ( \8335 , \8333 , \8334 );
not \U$8089 ( \8336 , \8335 );
or \U$8090 ( \8337 , \8329 , \8336 );
or \U$8091 ( \8338 , \8328 , \8335 );
nand \U$8092 ( \8339 , \8337 , \8338 );
not \U$8093 ( \8340 , \8339 );
xor \U$8094 ( \8341 , RIbe296c8_60, RIbe27c88_4);
not \U$8095 ( \8342 , \8341 );
not \U$8096 ( \8343 , \1130 );
or \U$8097 ( \8344 , \8342 , \8343 );
nand \U$8098 ( \8345 , \1137 , \7494 );
nand \U$8099 ( \8346 , \8344 , \8345 );
xor \U$8100 ( \8347 , RIbe29b00_69, RIbe28228_16);
not \U$8101 ( \8348 , \8347 );
not \U$8102 ( \8349 , \879 );
or \U$8103 ( \8350 , \8348 , \8349 );
nand \U$8104 ( \8351 , \885 , \7361 );
nand \U$8105 ( \8352 , \8350 , \8351 );
or \U$8106 ( \8353 , \8346 , \8352 );
not \U$8107 ( \8354 , \7438 );
not \U$8108 ( \8355 , \370 );
or \U$8109 ( \8356 , \8354 , \8355 );
xnor \U$8110 ( \8357 , RIbe29d58_74, RIbe27c10_3);
not \U$8111 ( \8358 , \8357 );
nand \U$8112 ( \8359 , \8358 , \1103 );
nand \U$8113 ( \8360 , \8356 , \8359 );
nand \U$8114 ( \8361 , \8353 , \8360 );
nand \U$8115 ( \8362 , \8352 , \8346 );
and \U$8116 ( \8363 , \8361 , \8362 );
not \U$8117 ( \8364 , \8363 );
not \U$8118 ( \8365 , \8364 );
xnor \U$8119 ( \8366 , RIbe288b8_30, RIbe28480_21);
or \U$8120 ( \8367 , \3345 , \8366 );
not \U$8121 ( \8368 , \7479 );
or \U$8122 ( \8369 , \2672 , \8368 );
nand \U$8123 ( \8370 , \8367 , \8369 );
not \U$8124 ( \8371 , \8370 );
xor \U$8125 ( \8372 , RIbe28de0_41, RIbe29f38_78);
not \U$8126 ( \8373 , \8372 );
not \U$8127 ( \8374 , \331 );
or \U$8128 ( \8375 , \8373 , \8374 );
nand \U$8129 ( \8376 , \346 , \7468 );
nand \U$8130 ( \8377 , \8375 , \8376 );
xor \U$8131 ( \8378 , RIbe2aa78_102, RIbe27b98_2);
not \U$8132 ( \8379 , \8378 );
not \U$8133 ( \8380 , \255 );
not \U$8134 ( \8381 , \8380 );
or \U$8135 ( \8382 , \8379 , \8381 );
not \U$8136 ( \8383 , \8029 );
nand \U$8137 ( \8384 , \8383 , \7585 );
nand \U$8138 ( \8385 , \8382 , \8384 );
xor \U$8139 ( \8386 , \8377 , \8385 );
not \U$8140 ( \8387 , \8386 );
or \U$8141 ( \8388 , \8371 , \8387 );
nand \U$8142 ( \8389 , \8385 , \8377 );
nand \U$8143 ( \8390 , \8388 , \8389 );
xor \U$8144 ( \8391 , RIbe290b0_47, RIbe28cf0_39);
not \U$8145 ( \8392 , \8391 );
not \U$8146 ( \8393 , \386 );
or \U$8147 ( \8394 , \8392 , \8393 );
nand \U$8148 ( \8395 , \399 , \7400 );
nand \U$8149 ( \8396 , \8394 , \8395 );
not \U$8150 ( \8397 , \8396 );
xor \U$8151 ( \8398 , RIbe29380_53, RIbe2a028_80);
not \U$8152 ( \8399 , \8398 );
buf \U$8153 ( \8400 , \8167 );
buf \U$8154 ( \8401 , \8400 );
not \U$8155 ( \8402 , \8401 );
or \U$8156 ( \8403 , \8399 , \8402 );
nand \U$8157 ( \8404 , \8172 , RIbe2a028_80);
nand \U$8158 ( \8405 , \8403 , \8404 );
not \U$8159 ( \8406 , \8405 );
or \U$8160 ( \8407 , \8397 , \8406 );
or \U$8161 ( \8408 , \8396 , \8405 );
and \U$8162 ( \8409 , RIbe28930_31, RIbe291a0_49);
nor \U$8163 ( \8410 , RIbe28930_31, RIbe291a0_49);
nor \U$8164 ( \8411 , \8409 , \8410 );
not \U$8165 ( \8412 , \8411 );
not \U$8166 ( \8413 , \1793 );
or \U$8167 ( \8414 , \8412 , \8413 );
nand \U$8168 ( \8415 , \1199 , \7426 );
nand \U$8169 ( \8416 , \8414 , \8415 );
nand \U$8170 ( \8417 , \8408 , \8416 );
nand \U$8171 ( \8418 , \8407 , \8417 );
xor \U$8172 ( \8419 , \8390 , \8418 );
not \U$8173 ( \8420 , \8419 );
or \U$8174 ( \8421 , \8365 , \8420 );
nand \U$8175 ( \8422 , \8390 , \8418 );
nand \U$8176 ( \8423 , \8421 , \8422 );
not \U$8177 ( \8424 , \8423 );
or \U$8178 ( \8425 , \8340 , \8424 );
not \U$8179 ( \8426 , \8328 );
nand \U$8180 ( \8427 , \8426 , \8335 );
nand \U$8181 ( \8428 , \8425 , \8427 );
xor \U$8182 ( \8429 , \7461 , \7387 );
not \U$8183 ( \8430 , \8429 );
not \U$8184 ( \8431 , \7526 );
not \U$8185 ( \8432 , \7561 );
not \U$8186 ( \8433 , \8432 );
or \U$8187 ( \8434 , \8431 , \8433 );
or \U$8188 ( \8435 , \8432 , \7526 );
nand \U$8189 ( \8436 , \8434 , \8435 );
not \U$8190 ( \8437 , \7507 );
not \U$8191 ( \8438 , \7500 );
or \U$8192 ( \8439 , \8437 , \8438 );
nand \U$8193 ( \8440 , \7520 , \7508 );
nand \U$8194 ( \8441 , \8439 , \8440 );
not \U$8195 ( \8442 , \7518 );
and \U$8196 ( \8443 , \8441 , \8442 );
not \U$8197 ( \8444 , \8441 );
and \U$8198 ( \8445 , \8444 , \7518 );
nor \U$8199 ( \8446 , \8443 , \8445 );
xor \U$8200 ( \8447 , \7466 , \7475 );
xnor \U$8201 ( \8448 , \8447 , \7490 );
nand \U$8202 ( \8449 , \8446 , \8448 );
not \U$8203 ( \8450 , \8449 );
and \U$8204 ( \8451 , \7416 , \7398 );
not \U$8205 ( \8452 , \7416 );
not \U$8206 ( \8453 , \7398 );
and \U$8207 ( \8454 , \8452 , \8453 );
nor \U$8208 ( \8455 , \8451 , \8454 );
not \U$8209 ( \8456 , \8455 );
or \U$8210 ( \8457 , \8450 , \8456 );
not \U$8211 ( \8458 , \8448 );
not \U$8212 ( \8459 , \8446 );
nand \U$8213 ( \8460 , \8458 , \8459 );
nand \U$8214 ( \8461 , \8457 , \8460 );
and \U$8215 ( \8462 , \8436 , \8461 );
not \U$8216 ( \8463 , \8436 );
not \U$8217 ( \8464 , \8461 );
and \U$8218 ( \8465 , \8463 , \8464 );
nor \U$8219 ( \8466 , \8462 , \8465 );
not \U$8220 ( \8467 , \8466 );
or \U$8221 ( \8468 , \8430 , \8467 );
nand \U$8222 ( \8469 , \8436 , \8461 );
nand \U$8223 ( \8470 , \8468 , \8469 );
and \U$8224 ( \8471 , \8428 , \8470 );
not \U$8225 ( \8472 , \8428 );
not \U$8226 ( \8473 , \8470 );
and \U$8227 ( \8474 , \8472 , \8473 );
nor \U$8228 ( \8475 , \8471 , \8474 );
not \U$8229 ( \8476 , \8475 );
or \U$8230 ( \8477 , \8327 , \8476 );
not \U$8231 ( \8478 , \8473 );
nand \U$8232 ( \8479 , \8478 , \8428 );
nand \U$8233 ( \8480 , \8477 , \8479 );
xor \U$8234 ( \8481 , \8321 , \8480 );
not \U$8235 ( \8482 , \7665 );
not \U$8236 ( \8483 , \8482 );
not \U$8237 ( \8484 , \7765 );
or \U$8238 ( \8485 , \8483 , \8484 );
or \U$8239 ( \8486 , \8482 , \7765 );
nand \U$8240 ( \8487 , \8485 , \8486 );
xor \U$8241 ( \8488 , \8481 , \8487 );
and \U$8242 ( \8489 , \8316 , \8488 );
and \U$8243 ( \8490 , \8130 , \8315 );
or \U$8244 ( \8491 , \8489 , \8490 );
not \U$8245 ( \8492 , \8491 );
not \U$8246 ( \8493 , \8084 );
xor \U$8247 ( \8494 , \7992 , \8079 );
not \U$8248 ( \8495 , \8494 );
not \U$8249 ( \8496 , \8495 );
or \U$8250 ( \8497 , \8493 , \8496 );
nand \U$8251 ( \8498 , \8494 , \8083 );
nand \U$8252 ( \8499 , \8497 , \8498 );
not \U$8253 ( \8500 , \8499 );
not \U$8254 ( \8501 , \8487 );
nand \U$8255 ( \8502 , \8501 , \8321 );
nand \U$8256 ( \8503 , \8502 , \8480 );
not \U$8257 ( \8504 , \8321 );
not \U$8258 ( \8505 , \8501 );
nand \U$8259 ( \8506 , \8504 , \8505 );
nand \U$8260 ( \8507 , \8503 , \8506 );
nand \U$8261 ( \8508 , \8500 , \8507 );
not \U$8262 ( \8509 , \8508 );
or \U$8263 ( \8510 , \8492 , \8509 );
not \U$8264 ( \8511 , \8507 );
nand \U$8265 ( \8512 , \8511 , \8499 );
nand \U$8266 ( \8513 , \8510 , \8512 );
not \U$8267 ( \8514 , \8090 );
not \U$8268 ( \8515 , \8098 );
not \U$8269 ( \8516 , \8515 );
or \U$8270 ( \8517 , \8514 , \8516 );
nand \U$8271 ( \8518 , \8517 , \8099 );
nand \U$8272 ( \8519 , \8513 , \8518 );
and \U$8273 ( \8520 , \8103 , \8128 , \8519 );
not \U$8274 ( \8521 , \8520 );
xor \U$8275 ( \8522 , RIbe29a10_67, RIbe28228_16);
not \U$8276 ( \8523 , \8522 );
not \U$8277 ( \8524 , \885 );
or \U$8278 ( \8525 , \8523 , \8524 );
xor \U$8279 ( \8526 , RIbe29218_50, RIbe28228_16);
nand \U$8280 ( \8527 , \879 , \8526 );
nand \U$8281 ( \8528 , \8525 , \8527 );
xor \U$8282 ( \8529 , RIbe296c8_60, RIbe29998_66);
not \U$8283 ( \8530 , \8529 );
not \U$8284 ( \8531 , \899 );
not \U$8285 ( \8532 , \8531 );
or \U$8286 ( \8533 , \8530 , \8532 );
buf \U$8287 ( \8534 , \1937 );
xor \U$8288 ( \8535 , RIbe28d68_40, RIbe296c8_60);
nand \U$8289 ( \8536 , \8534 , \8535 );
nand \U$8290 ( \8537 , \8533 , \8536 );
or \U$8291 ( \8538 , \8528 , \8537 );
xor \U$8292 ( \8539 , RIbe29f38_78, RIbe27c10_3);
not \U$8293 ( \8540 , \8539 );
not \U$8294 ( \8541 , \1493 );
or \U$8295 ( \8542 , \8540 , \8541 );
xor \U$8296 ( \8543 , RIbe29ec0_77, RIbe27c10_3);
nand \U$8297 ( \8544 , \1173 , \8543 );
nand \U$8298 ( \8545 , \8542 , \8544 );
nand \U$8299 ( \8546 , \8538 , \8545 );
nand \U$8300 ( \8547 , \8528 , \8537 );
and \U$8301 ( \8548 , \8546 , \8547 );
xor \U$8302 ( \8549 , RIbe280c0_13, RIbe27c88_4);
not \U$8303 ( \8550 , \8549 );
not \U$8304 ( \8551 , \859 );
not \U$8305 ( \8552 , \8551 );
or \U$8306 ( \8553 , \8550 , \8552 );
xor \U$8307 ( \8554 , RIbe280c0_13, RIbe27df0_7);
nand \U$8308 ( \8555 , \2369 , \8554 );
nand \U$8309 ( \8556 , \8553 , \8555 );
xor \U$8310 ( \8557 , RIbe285e8_24, RIbe288b8_30);
not \U$8311 ( \8558 , \8557 );
not \U$8312 ( \8559 , \2618 );
or \U$8313 ( \8560 , \8558 , \8559 );
xnor \U$8314 ( \8561 , RIbe285e8_24, RIbe28a98_34);
not \U$8315 ( \8562 , \8561 );
nand \U$8316 ( \8563 , \8562 , \2625 );
nand \U$8317 ( \8564 , \8560 , \8563 );
or \U$8318 ( \8565 , \8556 , \8564 );
xor \U$8319 ( \8566 , RIbe28390_19, RIbe28138_14);
not \U$8320 ( \8567 , \8566 );
not \U$8321 ( \8568 , \3408 );
or \U$8322 ( \8569 , \8567 , \8568 );
xor \U$8323 ( \8570 , RIbe28390_19, RIbe282a0_17);
nand \U$8324 ( \8571 , \2648 , \8570 );
nand \U$8325 ( \8572 , \8569 , \8571 );
nand \U$8326 ( \8573 , \8565 , \8572 );
nand \U$8327 ( \8574 , \8556 , \8564 );
nand \U$8328 ( \8575 , \8573 , \8574 );
not \U$8329 ( \8576 , \8575 );
and \U$8330 ( \8577 , \8548 , \8576 );
not \U$8331 ( \8578 , \8548 );
and \U$8332 ( \8579 , \8578 , \8575 );
nor \U$8333 ( \8580 , \8577 , \8579 );
not \U$8334 ( \8581 , \4843 );
xnor \U$8335 ( \8582 , RIbe29e48_76, RIbe28570_23);
or \U$8336 ( \8583 , \8581 , \8582 );
not \U$8337 ( \8584 , \8245 );
and \U$8338 ( \8585 , RIbe29e48_76, \304 );
not \U$8339 ( \8586 , RIbe29e48_76);
and \U$8340 ( \8587 , \8586 , RIbe286d8_26);
nor \U$8341 ( \8588 , \8585 , \8587 );
or \U$8342 ( \8589 , \8584 , \8588 );
nand \U$8343 ( \8590 , \8583 , \8589 );
not \U$8344 ( \8591 , \8590 );
xor \U$8345 ( \8592 , RIbe29c68_72, RIbe28750_27);
not \U$8346 ( \8593 , \8592 );
not \U$8347 ( \8594 , \4576 );
buf \U$8348 ( \8595 , \8594 );
not \U$8349 ( \8596 , \8595 );
or \U$8350 ( \8597 , \8593 , \8596 );
xor \U$8351 ( \8598 , RIbe29c68_72, RIbe28840_29);
nand \U$8352 ( \8599 , \4580 , \8598 );
nand \U$8353 ( \8600 , \8597 , \8599 );
not \U$8354 ( \8601 , \8600 );
xor \U$8355 ( \8602 , RIbe293f8_54, RIbe27e68_8);
and \U$8356 ( \8603 , \8602 , \2600 );
xor \U$8357 ( \8604 , RIbe29308_52, RIbe27e68_8);
and \U$8358 ( \8605 , \2603 , \8604 );
nor \U$8359 ( \8606 , \8603 , \8605 );
not \U$8360 ( \8607 , \8606 );
or \U$8361 ( \8608 , \8601 , \8607 );
or \U$8362 ( \8609 , \8606 , \8600 );
nand \U$8363 ( \8610 , \8608 , \8609 );
not \U$8364 ( \8611 , \8610 );
or \U$8365 ( \8612 , \8591 , \8611 );
not \U$8366 ( \8613 , \8606 );
nand \U$8367 ( \8614 , \8613 , \8600 );
nand \U$8368 ( \8615 , \8612 , \8614 );
xor \U$8369 ( \8616 , \8580 , \8615 );
not \U$8370 ( \8617 , \2762 );
not \U$8371 ( \8618 , \8561 );
and \U$8372 ( \8619 , \8617 , \8618 );
and \U$8373 ( \8620 , \8270 , \8265 );
nor \U$8374 ( \8621 , \8619 , \8620 );
not \U$8375 ( \8622 , \8621 );
not \U$8376 ( \8623 , \8554 );
buf \U$8377 ( \8624 , \858 );
not \U$8378 ( \8625 , \8624 );
or \U$8379 ( \8626 , \8623 , \8625 );
nand \U$8380 ( \8627 , \1263 , \8275 );
nand \U$8381 ( \8628 , \8626 , \8627 );
not \U$8382 ( \8629 , \8628 );
xor \U$8383 ( \8630 , RIbe28a20_33, RIbe295d8_58);
not \U$8384 ( \8631 , \8630 );
not \U$8385 ( \8632 , \1780 );
or \U$8386 ( \8633 , \8631 , \8632 );
nand \U$8387 ( \8634 , \5055 , \8190 );
nand \U$8388 ( \8635 , \8633 , \8634 );
not \U$8389 ( \8636 , \8635 );
not \U$8390 ( \8637 , \8636 );
or \U$8391 ( \8638 , \8629 , \8637 );
or \U$8392 ( \8639 , \8628 , \8636 );
nand \U$8393 ( \8640 , \8638 , \8639 );
not \U$8394 ( \8641 , \8640 );
or \U$8395 ( \8642 , \8622 , \8641 );
or \U$8396 ( \8643 , \8640 , \8621 );
nand \U$8397 ( \8644 , \8642 , \8643 );
not \U$8398 ( \8645 , \8535 );
not \U$8399 ( \8646 , \2875 );
or \U$8400 ( \8647 , \8645 , \8646 );
nand \U$8401 ( \8648 , \1137 , \8341 );
nand \U$8402 ( \8649 , \8647 , \8648 );
not \U$8403 ( \8650 , \8570 );
not \U$8404 ( \8651 , \2638 );
not \U$8405 ( \8652 , \8651 );
or \U$8406 ( \8653 , \8650 , \8652 );
not \U$8407 ( \8654 , \2646 );
nand \U$8408 ( \8655 , \8654 , \8206 );
nand \U$8409 ( \8656 , \8653 , \8655 );
xor \U$8410 ( \8657 , \8649 , \8656 );
xor \U$8411 ( \8658 , RIbe29038_46, RIbe298a8_64);
not \U$8412 ( \8659 , \8658 );
not \U$8413 ( \8660 , \282 );
or \U$8414 ( \8661 , \8659 , \8660 );
nand \U$8415 ( \8662 , \287 , \8213 );
nand \U$8416 ( \8663 , \8661 , \8662 );
xor \U$8417 ( \8664 , \8657 , \8663 );
xor \U$8418 ( \8665 , \8644 , \8664 );
not \U$8419 ( \8666 , \8604 );
not \U$8420 ( \8667 , \2600 );
or \U$8421 ( \8668 , \8666 , \8667 );
nand \U$8422 ( \8669 , \2464 , \8182 );
nand \U$8423 ( \8670 , \8668 , \8669 );
not \U$8424 ( \8671 , \8598 );
not \U$8425 ( \8672 , \8259 );
or \U$8426 ( \8673 , \8671 , \8672 );
nand \U$8427 ( \8674 , \4580 , \8257 );
nand \U$8428 ( \8675 , \8673 , \8674 );
not \U$8429 ( \8676 , \8522 );
not \U$8430 ( \8677 , \879 );
or \U$8431 ( \8678 , \8676 , \8677 );
buf \U$8432 ( \8679 , \877 );
buf \U$8433 ( \8680 , \8679 );
nand \U$8434 ( \8681 , \8680 , \8347 );
nand \U$8435 ( \8682 , \8678 , \8681 );
xor \U$8436 ( \8683 , \8675 , \8682 );
xor \U$8437 ( \8684 , \8670 , \8683 );
xor \U$8438 ( \8685 , \8665 , \8684 );
xor \U$8439 ( \8686 , \8616 , \8685 );
xor \U$8440 ( \8687 , RIbe2a2f8_86, RIbe29380_53);
not \U$8441 ( \8688 , \8687 );
and \U$8442 ( \8689 , RIbe2a370_87, RIbe2a2f8_86);
not \U$8443 ( \8690 , RIbe2a370_87);
and \U$8444 ( \8691 , \8690 , RIbe2a3e8_88);
nor \U$8445 ( \8692 , \8689 , \8691 );
nor \U$8446 ( \8693 , RIbe2a2f8_86, RIbe2a3e8_88);
not \U$8447 ( \8694 , \8693 );
nand \U$8448 ( \8695 , \8692 , \8694 );
buf \U$8449 ( \8696 , \8695 );
not \U$8450 ( \8697 , \8696 );
not \U$8451 ( \8698 , \8697 );
or \U$8452 ( \8699 , \8688 , \8698 );
not \U$8453 ( \8700 , RIbe2a370_87);
not \U$8454 ( \8701 , RIbe2a3e8_88);
and \U$8455 ( \8702 , \8700 , \8701 );
and \U$8456 ( \8703 , RIbe2a370_87, RIbe2a3e8_88);
nor \U$8457 ( \8704 , \8702 , \8703 );
buf \U$8458 ( \8705 , \8704 );
buf \U$8459 ( \8706 , \8705 );
nand \U$8460 ( \8707 , \8706 , RIbe2a2f8_86);
nand \U$8461 ( \8708 , \8699 , \8707 );
not \U$8462 ( \8709 , \8708 );
not \U$8463 ( \8710 , \8709 );
not \U$8464 ( \8711 , \2700 );
not \U$8465 ( \8712 , \8711 );
not \U$8466 ( \8713 , \8712 );
xnor \U$8467 ( \8714 , RIbe29740_61, RIbe28b88_36);
not \U$8468 ( \8715 , \8714 );
and \U$8469 ( \8716 , \8713 , \8715 );
xor \U$8470 ( \8717 , RIbe297b8_62, RIbe28b88_36);
and \U$8471 ( \8718 , \2560 , \8717 );
nor \U$8472 ( \8719 , \8716 , \8718 );
not \U$8473 ( \8720 , \8719 );
or \U$8474 ( \8721 , \8710 , \8720 );
xor \U$8475 ( \8722 , RIbe29b78_70, RIbe290b0_47);
not \U$8476 ( \8723 , \8722 );
not \U$8477 ( \8724 , \2730 );
or \U$8478 ( \8725 , \8723 , \8724 );
xor \U$8479 ( \8726 , RIbe27b20_1, RIbe290b0_47);
nand \U$8480 ( \8727 , \399 , \8726 );
nand \U$8481 ( \8728 , \8725 , \8727 );
nand \U$8482 ( \8729 , \8721 , \8728 );
not \U$8483 ( \8730 , \8719 );
nand \U$8484 ( \8731 , \8730 , \8708 );
nand \U$8485 ( \8732 , \8729 , \8731 );
not \U$8486 ( \8733 , \8732 );
xor \U$8487 ( \8734 , RIbe294e8_56, RIbe28480_21);
not \U$8488 ( \8735 , \8734 );
not \U$8489 ( \8736 , \2519 );
or \U$8490 ( \8737 , \8735 , \8736 );
not \U$8491 ( \8738 , \8366 );
nand \U$8492 ( \8739 , \8738 , \2527 );
nand \U$8493 ( \8740 , \8737 , \8739 );
and \U$8494 ( \8741 , RIbe2a898_98, RIbe27b98_2);
xor \U$8495 ( \8742 , RIbe28de0_41, RIbe2b6a8_128);
not \U$8496 ( \8743 , \8742 );
not \U$8497 ( \8744 , \331 );
or \U$8498 ( \8745 , \8743 , \8744 );
nand \U$8499 ( \8746 , \347 , \8372 );
nand \U$8500 ( \8747 , \8745 , \8746 );
xor \U$8501 ( \8748 , \8741 , \8747 );
xnor \U$8502 ( \8749 , \8740 , \8748 );
not \U$8503 ( \8750 , \8749 );
or \U$8504 ( \8751 , \8733 , \8750 );
not \U$8505 ( \8752 , \8740 );
not \U$8506 ( \8753 , \8752 );
not \U$8507 ( \8754 , \8748 );
or \U$8508 ( \8755 , \8753 , \8754 );
or \U$8509 ( \8756 , \8748 , \8752 );
nand \U$8510 ( \8757 , \8755 , \8756 );
nand \U$8511 ( \8758 , \8729 , \8731 , \8757 );
nand \U$8512 ( \8759 , \8751 , \8758 );
xor \U$8513 ( \8760 , RIbe2aa00_101, RIbe27b98_2);
not \U$8514 ( \8761 , \8760 );
not \U$8515 ( \8762 , \8380 );
or \U$8516 ( \8763 , \8761 , \8762 );
nand \U$8517 ( \8764 , \7585 , \8378 );
nand \U$8518 ( \8765 , \8763 , \8764 );
xor \U$8519 ( \8766 , RIbe27d78_6, RIbe29ce0_73);
not \U$8520 ( \8767 , \8766 );
not \U$8521 ( \8768 , \300 );
not \U$8522 ( \8769 , \8768 );
or \U$8523 ( \8770 , \8767 , \8769 );
nand \U$8524 ( \8771 , \314 , \8232 );
nand \U$8525 ( \8772 , \8770 , \8771 );
xor \U$8526 ( \8773 , \8765 , \8772 );
xor \U$8527 ( \8774 , RIbe28c78_38, RIbe27fd0_11);
not \U$8528 ( \8775 , \8774 );
not \U$8529 ( \8776 , \3378 );
or \U$8530 ( \8777 , \8775 , \8776 );
not \U$8531 ( \8778 , \8249 );
nand \U$8532 ( \8779 , \8778 , \2707 );
nand \U$8533 ( \8780 , \8777 , \8779 );
xor \U$8534 ( \8781 , \8773 , \8780 );
xor \U$8535 ( \8782 , \8759 , \8781 );
xor \U$8536 ( \8783 , \8686 , \8782 );
not \U$8537 ( \8784 , \8783 );
xor \U$8538 ( \8785 , RIbe28d68_40, RIbe280c0_13);
not \U$8539 ( \8786 , \8785 );
not \U$8540 ( \8787 , \861 );
or \U$8541 ( \8788 , \8786 , \8787 );
nand \U$8542 ( \8789 , \1263 , \8549 );
nand \U$8543 ( \8790 , \8788 , \8789 );
not \U$8544 ( \8791 , \8790 );
xor \U$8545 ( \8792 , RIbe2a910_99, RIbe2b5b8_126);
buf \U$8546 ( \8793 , \8792 );
buf \U$8547 ( \8794 , \8793 );
not \U$8548 ( \8795 , \8794 );
not \U$8549 ( \8796 , \8795 );
and \U$8550 ( \8797 , RIbe2a910_99, RIbe2a3e8_88);
not \U$8551 ( \8798 , RIbe2a910_99);
and \U$8552 ( \8799 , \8798 , RIbe2b5b8_126);
nor \U$8553 ( \8800 , \8797 , \8799 );
nor \U$8554 ( \8801 , RIbe2a3e8_88, RIbe2b5b8_126);
not \U$8555 ( \8802 , \8801 );
nand \U$8556 ( \8803 , \8800 , \8802 );
not \U$8557 ( \8804 , \8803 );
buf \U$8558 ( \8805 , \8804 );
buf \U$8559 ( \8806 , \8805 );
not \U$8560 ( \8807 , \8806 );
not \U$8561 ( \8808 , \8807 );
or \U$8562 ( \8809 , \8796 , \8808 );
nand \U$8563 ( \8810 , \8809 , RIbe2a3e8_88);
xor \U$8564 ( \8811 , RIbe294e8_56, RIbe285e8_24);
not \U$8565 ( \8812 , \8811 );
not \U$8566 ( \8813 , \2617 );
not \U$8567 ( \8814 , \8813 );
or \U$8568 ( \8815 , \8812 , \8814 );
nand \U$8569 ( \8816 , \8270 , \8557 );
nand \U$8570 ( \8817 , \8815 , \8816 );
nand \U$8571 ( \8818 , \8810 , \8817 );
nand \U$8572 ( \8819 , \8791 , \8818 );
not \U$8573 ( \8820 , \8810 );
not \U$8574 ( \8821 , \8817 );
nand \U$8575 ( \8822 , \8820 , \8821 );
and \U$8576 ( \8823 , \8819 , \8822 );
xor \U$8577 ( \8824 , RIbe27e68_8, RIbe28a98_34);
not \U$8578 ( \8825 , \8824 );
not \U$8579 ( \8826 , \2600 );
or \U$8580 ( \8827 , \8825 , \8826 );
nand \U$8581 ( \8828 , \2464 , \8602 );
nand \U$8582 ( \8829 , \8827 , \8828 );
not \U$8583 ( \8830 , \8829 );
xor \U$8584 ( \8831 , RIbe286d8_26, RIbe2a028_80);
not \U$8585 ( \8832 , \8831 );
not \U$8586 ( \8833 , \8401 );
or \U$8587 ( \8834 , \8832 , \8833 );
xor \U$8588 ( \8835 , RIbe2a028_80, RIbe27ee0_9);
nand \U$8589 ( \8836 , \8172 , \8835 );
nand \U$8590 ( \8837 , \8834 , \8836 );
not \U$8591 ( \8838 , \8837 );
or \U$8592 ( \8839 , \8830 , \8838 );
or \U$8593 ( \8840 , \8829 , \8837 );
xor \U$8594 ( \8841 , RIbe29e48_76, RIbe28840_29);
not \U$8595 ( \8842 , \8841 );
not \U$8596 ( \8843 , \4842 );
or \U$8597 ( \8844 , \8842 , \8843 );
not \U$8598 ( \8845 , \8582 );
nand \U$8599 ( \8846 , \8845 , \7368 );
nand \U$8600 ( \8847 , \8844 , \8846 );
nand \U$8601 ( \8848 , \8840 , \8847 );
nand \U$8602 ( \8849 , \8839 , \8848 );
xor \U$8603 ( \8850 , \8823 , \8849 );
xor \U$8604 ( \8851 , RIbe27df0_7, RIbe28228_16);
not \U$8605 ( \8852 , \8851 );
not \U$8606 ( \8853 , \3056 );
or \U$8607 ( \8854 , \8852 , \8853 );
nand \U$8608 ( \8855 , \885 , \8526 );
nand \U$8609 ( \8856 , \8854 , \8855 );
not \U$8610 ( \8857 , \8856 );
xor \U$8611 ( \8858 , RIbe29c68_72, RIbe284f8_22);
not \U$8612 ( \8859 , \8858 );
not \U$8613 ( \8860 , \8259 );
or \U$8614 ( \8861 , \8859 , \8860 );
nand \U$8615 ( \8862 , \7237 , \8592 );
nand \U$8616 ( \8863 , \8861 , \8862 );
xor \U$8617 ( \8864 , RIbe297b8_62, RIbe28390_19);
not \U$8618 ( \8865 , \8864 );
not \U$8619 ( \8866 , \3712 );
or \U$8620 ( \8867 , \8865 , \8866 );
buf \U$8621 ( \8868 , \2647 );
nand \U$8622 ( \8869 , \8868 , \8566 );
nand \U$8623 ( \8870 , \8867 , \8869 );
xor \U$8624 ( \8871 , \8863 , \8870 );
not \U$8625 ( \8872 , \8871 );
or \U$8626 ( \8873 , \8857 , \8872 );
nand \U$8627 ( \8874 , \8863 , \8870 );
nand \U$8628 ( \8875 , \8873 , \8874 );
xor \U$8629 ( \8876 , \8850 , \8875 );
not \U$8630 ( \8877 , \2718 );
xor \U$8631 ( \8878 , RIbe28c00_37, RIbe27fd0_11);
not \U$8632 ( \8879 , \8878 );
not \U$8633 ( \8880 , \8879 );
and \U$8634 ( \8881 , \8877 , \8880 );
and \U$8635 ( \8882 , \2707 , \8774 );
nor \U$8636 ( \8883 , \8881 , \8882 );
xor \U$8637 ( \8884 , RIbe28930_31, RIbe29b00_69);
not \U$8638 ( \8885 , \8884 );
not \U$8639 ( \8886 , \961 );
nor \U$8640 ( \8887 , \8886 , \963 );
not \U$8641 ( \8888 , \8887 );
or \U$8642 ( \8889 , \8885 , \8888 );
xor \U$8643 ( \8890 , RIbe28930_31, RIbe29128_48);
nand \U$8644 ( \8891 , \1797 , \8890 );
nand \U$8645 ( \8892 , \8889 , \8891 );
not \U$8646 ( \8893 , \8892 );
not \U$8647 ( \8894 , \8893 );
xor \U$8648 ( \8895 , RIbe27d78_6, RIbe29d58_74);
not \U$8649 ( \8896 , \8895 );
nand \U$8650 ( \8897 , \297 , \298 );
not \U$8651 ( \8898 , \8897 );
not \U$8652 ( \8899 , \8898 );
or \U$8653 ( \8900 , \8896 , \8899 );
nand \U$8654 ( \8901 , \314 , \8766 );
nand \U$8655 ( \8902 , \8900 , \8901 );
not \U$8656 ( \8903 , \8902 );
or \U$8657 ( \8904 , \8894 , \8903 );
or \U$8658 ( \8905 , \8893 , \8902 );
nand \U$8659 ( \8906 , \8904 , \8905 );
xnor \U$8660 ( \8907 , \8883 , \8906 );
not \U$8661 ( \8908 , \8907 );
not \U$8662 ( \8909 , \8908 );
xor \U$8663 ( \8910 , RIbe28cf0_39, RIbe29038_46);
not \U$8664 ( \8911 , \8910 );
not \U$8665 ( \8912 , \281 );
or \U$8666 ( \8913 , \8911 , \8912 );
nand \U$8667 ( \8914 , \1583 , \8658 );
nand \U$8668 ( \8915 , \8913 , \8914 );
xor \U$8669 ( \8916 , RIbe28a20_33, RIbe291a0_49);
not \U$8670 ( \8917 , \8916 );
not \U$8671 ( \8918 , \1780 );
or \U$8672 ( \8919 , \8917 , \8918 );
nand \U$8673 ( \8920 , \5055 , \8630 );
nand \U$8674 ( \8921 , \8919 , \8920 );
and \U$8675 ( \8922 , \8915 , \8921 );
not \U$8676 ( \8923 , \8915 );
not \U$8677 ( \8924 , \8921 );
and \U$8678 ( \8925 , \8923 , \8924 );
nor \U$8679 ( \8926 , \8922 , \8925 );
not \U$8680 ( \8927 , \8835 );
not \U$8681 ( \8928 , \8401 );
or \U$8682 ( \8929 , \8927 , \8928 );
buf \U$8683 ( \8930 , \8171 );
xor \U$8684 ( \8931 , RIbe28048_12, RIbe2a028_80);
nand \U$8685 ( \8932 , \8930 , \8931 );
nand \U$8686 ( \8933 , \8929 , \8932 );
xor \U$8687 ( \8934 , \8926 , \8933 );
not \U$8688 ( \8935 , \8934 );
or \U$8689 ( \8936 , \8909 , \8935 );
not \U$8690 ( \8937 , \8934 );
nand \U$8691 ( \8938 , \8937 , \8907 );
nand \U$8692 ( \8939 , \8936 , \8938 );
not \U$8693 ( \8940 , \8590 );
not \U$8694 ( \8941 , \8610 );
not \U$8695 ( \8942 , \8941 );
or \U$8696 ( \8943 , \8940 , \8942 );
not \U$8697 ( \8944 , \8590 );
nand \U$8698 ( \8945 , \8944 , \8610 );
nand \U$8699 ( \8946 , \8943 , \8945 );
and \U$8700 ( \8947 , \8939 , \8946 );
not \U$8701 ( \8948 , \8939 );
not \U$8702 ( \8949 , \8946 );
and \U$8703 ( \8950 , \8948 , \8949 );
nor \U$8704 ( \8951 , \8947 , \8950 );
xor \U$8705 ( \8952 , \8876 , \8951 );
xor \U$8706 ( \8953 , RIbe29470_55, RIbe28480_21);
not \U$8707 ( \8954 , \8953 );
not \U$8708 ( \8955 , \3483 );
or \U$8709 ( \8956 , \8954 , \8955 );
nand \U$8710 ( \8957 , \2527 , \8734 );
nand \U$8711 ( \8958 , \8956 , \8957 );
xor \U$8712 ( \8959 , RIbe2aa78_102, RIbe28de0_41);
not \U$8713 ( \8960 , \8959 );
not \U$8714 ( \8961 , \332 );
or \U$8715 ( \8962 , \8960 , \8961 );
nand \U$8716 ( \8963 , \514 , \8742 );
nand \U$8717 ( \8964 , \8962 , \8963 );
xor \U$8718 ( \8965 , \8958 , \8964 );
xor \U$8719 ( \8966 , RIbe2a898_98, RIbe27b98_2);
not \U$8720 ( \8967 , \8966 );
not \U$8721 ( \8968 , \256 );
or \U$8722 ( \8969 , \8967 , \8968 );
nand \U$8723 ( \8970 , \269 , \8760 );
nand \U$8724 ( \8971 , \8969 , \8970 );
xor \U$8725 ( \8972 , \8965 , \8971 );
xor \U$8726 ( \8973 , RIbe2b6a8_128, RIbe27c10_3);
not \U$8727 ( \8974 , \8973 );
not \U$8728 ( \8975 , \1493 );
or \U$8729 ( \8976 , \8974 , \8975 );
nand \U$8730 ( \8977 , \1173 , \8539 );
nand \U$8731 ( \8978 , \8976 , \8977 );
xor \U$8732 ( \8979 , RIbe29a10_67, RIbe28930_31);
not \U$8733 ( \8980 , \8979 );
not \U$8734 ( \8981 , \966 );
or \U$8735 ( \8982 , \8980 , \8981 );
nand \U$8736 ( \8983 , \1797 , \8884 );
nand \U$8737 ( \8984 , \8982 , \8983 );
xor \U$8738 ( \8985 , \8978 , \8984 );
xor \U$8739 ( \8986 , RIbe2a2f8_86, RIbe28048_12);
not \U$8740 ( \8987 , \8986 );
buf \U$8741 ( \8988 , \8696 );
not \U$8742 ( \8989 , \8988 );
not \U$8743 ( \8990 , \8989 );
or \U$8744 ( \8991 , \8987 , \8990 );
nand \U$8745 ( \8992 , \8706 , \8687 );
nand \U$8746 ( \8993 , \8991 , \8992 );
and \U$8747 ( \8994 , \8985 , \8993 );
and \U$8748 ( \8995 , \8978 , \8984 );
or \U$8749 ( \8996 , \8994 , \8995 );
xor \U$8750 ( \8997 , \8972 , \8996 );
xor \U$8751 ( \8998 , \8556 , \8564 );
xor \U$8752 ( \8999 , \8998 , \8572 );
and \U$8753 ( \9000 , \8997 , \8999 );
not \U$8754 ( \9001 , \8997 );
not \U$8755 ( \9002 , \8999 );
and \U$8756 ( \9003 , \9001 , \9002 );
nor \U$8757 ( \9004 , \9000 , \9003 );
and \U$8758 ( \9005 , \8952 , \9004 );
and \U$8759 ( \9006 , \8876 , \8951 );
or \U$8760 ( \9007 , \9005 , \9006 );
not \U$8761 ( \9008 , \9007 );
nand \U$8762 ( \9009 , \8784 , \9008 );
not \U$8763 ( \9010 , \9009 );
not \U$8764 ( \9011 , RIbe28318_18);
not \U$8765 ( \9012 , RIbe29c68_72);
and \U$8766 ( \9013 , \9011 , \9012 );
and \U$8767 ( \9014 , RIbe28318_18, RIbe29c68_72);
nor \U$8768 ( \9015 , \9013 , \9014 );
not \U$8769 ( \9016 , \9015 );
not \U$8770 ( \9017 , \8595 );
or \U$8771 ( \9018 , \9016 , \9017 );
nand \U$8772 ( \9019 , \4580 , \8858 );
nand \U$8773 ( \9020 , \9018 , \9019 );
not \U$8774 ( \9021 , \9020 );
xor \U$8775 ( \9022 , RIbe28228_16, RIbe27c88_4);
not \U$8776 ( \9023 , \9022 );
not \U$8777 ( \9024 , \879 );
or \U$8778 ( \9025 , \9023 , \9024 );
nand \U$8779 ( \9026 , \885 , \8851 );
nand \U$8780 ( \9027 , \9025 , \9026 );
not \U$8781 ( \9028 , \9027 );
not \U$8782 ( \9029 , \9028 );
xor \U$8783 ( \9030 , RIbe28cf0_39, RIbe296c8_60);
not \U$8784 ( \9031 , \9030 );
not \U$8785 ( \9032 , \2875 );
or \U$8786 ( \9033 , \9031 , \9032 );
xor \U$8787 ( \9034 , RIbe296c8_60, RIbe298a8_64);
nand \U$8788 ( \9035 , \8534 , \9034 );
nand \U$8789 ( \9036 , \9033 , \9035 );
not \U$8790 ( \9037 , \9036 );
not \U$8791 ( \9038 , \9037 );
or \U$8792 ( \9039 , \9029 , \9038 );
xor \U$8793 ( \9040 , RIbe27c10_3, RIbe2aa78_102);
not \U$8794 ( \9041 , \9040 );
not \U$8795 ( \9042 , \1103 );
or \U$8796 ( \9043 , \9041 , \9042 );
nand \U$8797 ( \9044 , \369 , \8973 );
nand \U$8798 ( \9045 , \9043 , \9044 );
nand \U$8799 ( \9046 , \9039 , \9045 );
nand \U$8800 ( \9047 , \9027 , \9036 );
nand \U$8801 ( \9048 , \9046 , \9047 );
xor \U$8802 ( \9049 , \9021 , \9048 );
xor \U$8803 ( \9050 , RIbe28b88_36, RIbe291a0_49);
not \U$8804 ( \9051 , \9050 );
buf \U$8805 ( \9052 , \2552 );
not \U$8806 ( \9053 , \9052 );
or \U$8807 ( \9054 , \9051 , \9053 );
and \U$8808 ( \9055 , RIbe28b88_36, RIbe295d8_58);
not \U$8809 ( \9056 , RIbe28b88_36);
and \U$8810 ( \9057 , \9056 , \2995 );
nor \U$8811 ( \9058 , \9055 , \9057 );
nand \U$8812 ( \9059 , \9058 , \2559 );
nand \U$8813 ( \9060 , \9054 , \9059 );
xor \U$8814 ( \9061 , RIbe28570_23, RIbe2a028_80);
not \U$8815 ( \9062 , \9061 );
not \U$8816 ( \9063 , \8168 );
or \U$8817 ( \9064 , \9062 , \9063 );
buf \U$8818 ( \9065 , \8172 );
nand \U$8819 ( \9066 , \9065 , \8831 );
nand \U$8820 ( \9067 , \9064 , \9066 );
xor \U$8821 ( \9068 , \9060 , \9067 );
xor \U$8822 ( \9069 , RIbe29038_46, RIbe29b78_70);
not \U$8823 ( \9070 , \9069 );
not \U$8824 ( \9071 , \281 );
or \U$8825 ( \9072 , \9070 , \9071 );
xor \U$8826 ( \9073 , RIbe27b20_1, RIbe29038_46);
nand \U$8827 ( \9074 , \287 , \9073 );
nand \U$8828 ( \9075 , \9072 , \9074 );
and \U$8829 ( \9076 , \9068 , \9075 );
and \U$8830 ( \9077 , \9060 , \9067 );
or \U$8831 ( \9078 , \9076 , \9077 );
xnor \U$8832 ( \9079 , \9049 , \9078 );
xor \U$8833 ( \9080 , RIbe27fd0_11, RIbe293f8_54);
nand \U$8834 ( \9081 , \2713 , \2715 );
not \U$8835 ( \9082 , \9081 );
and \U$8836 ( \9083 , \9080 , \9082 );
xor \U$8837 ( \9084 , RIbe27fd0_11, RIbe29308_52);
and \U$8838 ( \9085 , \7709 , \9084 );
nor \U$8839 ( \9086 , \9083 , \9085 );
not \U$8840 ( \9087 , \9086 );
not \U$8841 ( \9088 , \9087 );
buf \U$8842 ( \9089 , \8792 );
not \U$8843 ( \9090 , \9089 );
not \U$8844 ( \9091 , RIbe2a3e8_88);
or \U$8845 ( \9092 , \9090 , \9091 );
xnor \U$8846 ( \9093 , RIbe29380_53, RIbe2a3e8_88);
not \U$8847 ( \9094 , \9093 );
not \U$8848 ( \9095 , \8804 );
not \U$8849 ( \9096 , \9095 );
nand \U$8850 ( \9097 , \9094 , \9096 );
nand \U$8851 ( \9098 , \9092 , \9097 );
not \U$8852 ( \9099 , \9098 );
or \U$8853 ( \9100 , \9088 , \9099 );
and \U$8854 ( \9101 , \1199 , \8979 );
xor \U$8855 ( \9102 , RIbe28930_31, RIbe29218_50);
not \U$8856 ( \9103 , \9102 );
not \U$8857 ( \9104 , \965 );
nor \U$8858 ( \9105 , \9103 , \9104 );
nor \U$8859 ( \9106 , \9101 , \9105 );
not \U$8860 ( \9107 , \9106 );
not \U$8861 ( \9108 , \9098 );
nand \U$8862 ( \9109 , \9108 , \9086 );
nand \U$8863 ( \9110 , \9107 , \9109 );
nand \U$8864 ( \9111 , \9100 , \9110 );
xor \U$8865 ( \9112 , RIbe29d58_74, RIbe290b0_47);
not \U$8866 ( \9113 , \9112 );
not \U$8867 ( \9114 , \385 );
not \U$8868 ( \9115 , \9114 );
or \U$8869 ( \9116 , \9113 , \9115 );
xor \U$8870 ( \9117 , RIbe29ce0_73, RIbe290b0_47);
nand \U$8871 ( \9118 , \399 , \9117 );
nand \U$8872 ( \9119 , \9116 , \9118 );
xor \U$8873 ( \9120 , RIbe28138_14, RIbe28480_21);
not \U$8874 ( \9121 , \9120 );
not \U$8875 ( \9122 , \2519 );
or \U$8876 ( \9123 , \9121 , \9122 );
xor \U$8877 ( \9124 , RIbe28480_21, RIbe282a0_17);
nand \U$8878 ( \9125 , \2527 , \9124 );
nand \U$8879 ( \9126 , \9123 , \9125 );
xor \U$8880 ( \9127 , \9119 , \9126 );
xor \U$8881 ( \9128 , RIbe2a898_98, RIbe28de0_41);
not \U$8882 ( \9129 , \9128 );
not \U$8883 ( \9130 , \3103 );
or \U$8884 ( \9131 , \9129 , \9130 );
xor \U$8885 ( \9132 , RIbe2aa00_101, RIbe28de0_41);
nand \U$8886 ( \9133 , \514 , \9132 );
nand \U$8887 ( \9134 , \9131 , \9133 );
and \U$8888 ( \9135 , \9127 , \9134 );
and \U$8889 ( \9136 , \9119 , \9126 );
or \U$8890 ( \9137 , \9135 , \9136 );
xor \U$8891 ( \9138 , \9111 , \9137 );
not \U$8892 ( \9139 , \9084 );
not \U$8893 ( \9140 , \4893 );
or \U$8894 ( \9141 , \9139 , \9140 );
nand \U$8895 ( \9142 , \2707 , \8878 );
nand \U$8896 ( \9143 , \9141 , \9142 );
not \U$8897 ( \9144 , \9143 );
not \U$8898 ( \9145 , \269 );
not \U$8899 ( \9146 , \8966 );
or \U$8900 ( \9147 , \9145 , \9146 );
xnor \U$8901 ( \9148 , RIbe27b98_2, RIbe2a820_97);
or \U$8902 ( \9149 , \1566 , \9148 );
nand \U$8903 ( \9150 , \9147 , \9149 );
not \U$8904 ( \9151 , \9150 );
not \U$8905 ( \9152 , \9151 );
or \U$8906 ( \9153 , \9144 , \9152 );
not \U$8907 ( \9154 , \9143 );
nand \U$8908 ( \9155 , \9150 , \9154 );
nand \U$8909 ( \9156 , \9153 , \9155 );
xor \U$8910 ( \9157 , RIbe29ec0_77, RIbe27d78_6);
not \U$8911 ( \9158 , \9157 );
not \U$8912 ( \9159 , \1164 );
or \U$8913 ( \9160 , \9158 , \9159 );
nand \U$8914 ( \9161 , \315 , \8895 );
nand \U$8915 ( \9162 , \9160 , \9161 );
and \U$8916 ( \9163 , \9156 , \9162 );
not \U$8917 ( \9164 , \9156 );
not \U$8918 ( \9165 , \9162 );
and \U$8919 ( \9166 , \9164 , \9165 );
nor \U$8920 ( \9167 , \9163 , \9166 );
xor \U$8921 ( \9168 , \9138 , \9167 );
xor \U$8922 ( \9169 , \9079 , \9168 );
xor \U$8923 ( \9170 , \9119 , \9126 );
xor \U$8924 ( \9171 , \9170 , \9134 );
xor \U$8925 ( \9172 , RIbe28f48_44, RIbe28c00_37);
not \U$8926 ( \9173 , \9172 );
not \U$8927 ( \9174 , \3256 );
or \U$8928 ( \9175 , \9173 , \9174 );
xor \U$8929 ( \9176 , RIbe28f48_44, RIbe28c78_38);
nand \U$8930 ( \9177 , \4181 , \9176 );
nand \U$8931 ( \9178 , \9175 , \9177 );
xor \U$8932 ( \9179 , RIbe29f38_78, RIbe27d78_6);
not \U$8933 ( \9180 , \9179 );
not \U$8934 ( \9181 , \1164 );
or \U$8935 ( \9182 , \9180 , \9181 );
nand \U$8936 ( \9183 , \314 , \9157 );
nand \U$8937 ( \9184 , \9182 , \9183 );
nor \U$8938 ( \9185 , \9178 , \9184 );
not \U$8939 ( \9186 , \9185 );
nand \U$8940 ( \9187 , \9178 , \9184 );
nand \U$8941 ( \9188 , \9186 , \9187 );
not \U$8942 ( \9189 , \9188 );
xor \U$8943 ( \9190 , RIbe29128_48, RIbe28a20_33);
and \U$8944 ( \9191 , \2475 , \9190 );
buf \U$8945 ( \9192 , \1779 );
not \U$8946 ( \9193 , \9192 );
not \U$8947 ( \9194 , \9193 );
xor \U$8948 ( \9195 , RIbe29b00_69, RIbe28a20_33);
and \U$8949 ( \9196 , \9194 , \9195 );
nor \U$8950 ( \9197 , \9191 , \9196 );
buf \U$8951 ( \9198 , \9197 );
not \U$8952 ( \9199 , \9198 );
and \U$8953 ( \9200 , \9189 , \9199 );
and \U$8954 ( \9201 , \9188 , \9198 );
nor \U$8955 ( \9202 , \9200 , \9201 );
xor \U$8956 ( \9203 , \9171 , \9202 );
xor \U$8957 ( \9204 , RIbe29740_61, RIbe28390_19);
not \U$8958 ( \9205 , \9204 );
not \U$8959 ( \9206 , \2639 );
or \U$8960 ( \9207 , \9205 , \9206 );
nand \U$8961 ( \9208 , \5831 , \8864 );
nand \U$8962 ( \9209 , \9207 , \9208 );
xor \U$8963 ( \9210 , RIbe27b98_2, RIbe2a118_82);
not \U$8964 ( \9211 , \9210 );
not \U$8965 ( \9212 , \4828 );
or \U$8966 ( \9213 , \9211 , \9212 );
not \U$8967 ( \9214 , \9148 );
nand \U$8968 ( \9215 , \9214 , \1734 );
nand \U$8969 ( \9216 , \9213 , \9215 );
nor \U$8970 ( \9217 , \9209 , \9216 );
not \U$8971 ( \9218 , \9217 );
nand \U$8972 ( \9219 , \9216 , \9209 );
nand \U$8973 ( \9220 , \9218 , \9219 );
xor \U$8974 ( \9221 , RIbe285e8_24, RIbe29470_55);
and \U$8975 ( \9222 , \2890 , \9221 );
and \U$8976 ( \9223 , \2626 , \8811 );
nor \U$8977 ( \9224 , \9222 , \9223 );
xor \U$8978 ( \9225 , \9220 , \9224 );
and \U$8979 ( \9226 , \9203 , \9225 );
and \U$8980 ( \9227 , \9171 , \9202 );
or \U$8981 ( \9228 , \9226 , \9227 );
and \U$8982 ( \9229 , \9169 , \9228 );
and \U$8983 ( \9230 , \9079 , \9168 );
or \U$8984 ( \9231 , \9229 , \9230 );
not \U$8985 ( \9232 , \9231 );
xor \U$8986 ( \9233 , RIbe294e8_56, RIbe27e68_8);
not \U$8987 ( \9234 , \9233 );
not \U$8988 ( \9235 , \4443 );
or \U$8989 ( \9236 , \9234 , \9235 );
xor \U$8990 ( \9237 , RIbe288b8_30, RIbe27e68_8);
nand \U$8991 ( \9238 , \2603 , \9237 );
nand \U$8992 ( \9239 , \9236 , \9238 );
not \U$8993 ( \9240 , \9239 );
xor \U$8994 ( \9241 , RIbe28d68_40, RIbe28228_16);
not \U$8995 ( \9242 , \9241 );
not \U$8996 ( \9243 , \879 );
or \U$8997 ( \9244 , \9242 , \9243 );
nand \U$8998 ( \9245 , \8680 , \9022 );
nand \U$8999 ( \9246 , \9244 , \9245 );
not \U$9000 ( \9247 , \9246 );
or \U$9001 ( \9248 , \9240 , \9247 );
or \U$9002 ( \9249 , \9246 , \9239 );
xor \U$9003 ( \9250 , RIbe284f8_22, RIbe29e48_76);
not \U$9004 ( \9251 , \9250 );
not \U$9005 ( \9252 , \7371 );
not \U$9006 ( \9253 , \9252 );
or \U$9007 ( \9254 , \9251 , \9253 );
xor \U$9008 ( \9255 , RIbe29e48_76, RIbe28750_27);
nand \U$9009 ( \9256 , \4851 , \9255 );
nand \U$9010 ( \9257 , \9254 , \9256 );
nand \U$9011 ( \9258 , \9249 , \9257 );
nand \U$9012 ( \9259 , \9248 , \9258 );
xor \U$9013 ( \9260 , RIbe2a3e8_88, RIbe28048_12);
not \U$9014 ( \9261 , \9260 );
buf \U$9015 ( \9262 , \8804 );
buf \U$9016 ( \9263 , \9262 );
buf \U$9017 ( \9264 , \9263 );
not \U$9018 ( \9265 , \9264 );
or \U$9019 ( \9266 , \9261 , \9265 );
not \U$9020 ( \9267 , \9093 );
buf \U$9021 ( \9268 , \9089 );
nand \U$9022 ( \9269 , \9267 , \9268 );
nand \U$9023 ( \9270 , \9266 , \9269 );
not \U$9024 ( \9271 , \9270 );
xor \U$9025 ( \9272 , RIbe280c0_13, RIbe298a8_64);
not \U$9026 ( \9273 , \9272 );
xnor \U$9027 ( \9274 , RIbe280c0_13, RIbe281b0_15);
nor \U$9028 ( \9275 , \9273 , \9274 );
not \U$9029 ( \9276 , \9275 );
not \U$9030 ( \9277 , \1516 );
or \U$9031 ( \9278 , \9276 , \9277 );
xor \U$9032 ( \9279 , RIbe29998_66, RIbe280c0_13);
nand \U$9033 ( \9280 , \1263 , \9279 );
nand \U$9034 ( \9281 , \9278 , \9280 );
xor \U$9035 ( \9282 , RIbe285e8_24, RIbe282a0_17);
not \U$9036 ( \9283 , \9282 );
not \U$9037 ( \9284 , \8267 );
or \U$9038 ( \9285 , \9283 , \9284 );
nand \U$9039 ( \9286 , \2758 , \9221 );
nand \U$9040 ( \9287 , \9285 , \9286 );
and \U$9041 ( \9288 , \9281 , \9287 );
not \U$9042 ( \9289 , \9281 );
not \U$9043 ( \9290 , \9287 );
and \U$9044 ( \9291 , \9289 , \9290 );
nor \U$9045 ( \9292 , \9288 , \9291 );
not \U$9046 ( \9293 , \9292 );
or \U$9047 ( \9294 , \9271 , \9293 );
nand \U$9048 ( \9295 , \9287 , \9281 );
nand \U$9049 ( \9296 , \9294 , \9295 );
xor \U$9050 ( \9297 , \9259 , \9296 );
not \U$9051 ( \9298 , RIbe28b88_36);
not \U$9052 ( \9299 , RIbe29128_48);
and \U$9053 ( \9300 , \9298 , \9299 );
and \U$9054 ( \9301 , RIbe28b88_36, RIbe29128_48);
nor \U$9055 ( \9302 , \9300 , \9301 );
not \U$9056 ( \9303 , \9302 );
not \U$9057 ( \9304 , \2554 );
or \U$9058 ( \9305 , \9303 , \9304 );
nand \U$9059 ( \9306 , \2560 , \9050 );
nand \U$9060 ( \9307 , \9305 , \9306 );
not \U$9061 ( \9308 , \9307 );
xor \U$9062 ( \9309 , RIbe28c78_38, RIbe29c68_72);
not \U$9063 ( \9310 , \9309 );
not \U$9064 ( \9311 , \8595 );
or \U$9065 ( \9312 , \9310 , \9311 );
nand \U$9066 ( \9313 , \4580 , \9015 );
nand \U$9067 ( \9314 , \9312 , \9313 );
not \U$9068 ( \9315 , \9314 );
or \U$9069 ( \9316 , \9308 , \9315 );
xor \U$9070 ( \9317 , \9314 , \9307 );
not \U$9071 ( \9318 , \9317 );
not \U$9072 ( \9319 , RIbe28390_19);
not \U$9073 ( \9320 , RIbe295d8_58);
and \U$9074 ( \9321 , \9319 , \9320 );
and \U$9075 ( \9322 , RIbe28390_19, RIbe295d8_58);
nor \U$9076 ( \9323 , \9321 , \9322 );
and \U$9077 ( \9324 , \3408 , \9323 );
and \U$9078 ( \9325 , \3714 , \9204 );
nor \U$9079 ( \9326 , \9324 , \9325 );
or \U$9080 ( \9327 , \9318 , \9326 );
nand \U$9081 ( \9328 , \9316 , \9327 );
and \U$9082 ( \9329 , \9297 , \9328 );
and \U$9083 ( \9330 , \9259 , \9296 );
or \U$9084 ( \9331 , \9329 , \9330 );
not \U$9085 ( \9332 , \9331 );
not \U$9086 ( \9333 , \8820 );
not \U$9087 ( \9334 , \8821 );
or \U$9088 ( \9335 , \9333 , \9334 );
nand \U$9089 ( \9336 , \9335 , \8818 );
xnor \U$9090 ( \9337 , \8790 , \9336 );
not \U$9091 ( \9338 , \9021 );
nand \U$9092 ( \9339 , RIbe27b98_2, RIbe2a0a0_81);
not \U$9093 ( \9340 , \9255 );
not \U$9094 ( \9341 , \7716 );
or \U$9095 ( \9342 , \9340 , \9341 );
nand \U$9096 ( \9343 , \7368 , \8841 );
nand \U$9097 ( \9344 , \9342 , \9343 );
not \U$9098 ( \9345 , \9344 );
xor \U$9099 ( \9346 , \9339 , \9345 );
not \U$9100 ( \9347 , \9346 );
or \U$9101 ( \9348 , \9338 , \9347 );
not \U$9102 ( \9349 , \9339 );
nand \U$9103 ( \9350 , \9349 , \9344 );
nand \U$9104 ( \9351 , \9348 , \9350 );
and \U$9105 ( \9352 , \9337 , \9351 );
not \U$9106 ( \9353 , \9337 );
not \U$9107 ( \9354 , \9351 );
and \U$9108 ( \9355 , \9353 , \9354 );
nor \U$9109 ( \9356 , \9352 , \9355 );
not \U$9110 ( \9357 , \9356 );
or \U$9111 ( \9358 , \9332 , \9357 );
nand \U$9112 ( \9359 , \9351 , \9337 );
nand \U$9113 ( \9360 , \9358 , \9359 );
not \U$9114 ( \9361 , \8824 );
not \U$9115 ( \9362 , \2464 );
or \U$9116 ( \9363 , \9361 , \9362 );
nand \U$9117 ( \9364 , \9237 , \2600 );
nand \U$9118 ( \9365 , \9363 , \9364 );
not \U$9119 ( \9366 , \9365 );
not \U$9120 ( \9367 , \9279 );
not \U$9121 ( \9368 , \861 );
or \U$9122 ( \9369 , \9367 , \9368 );
nand \U$9123 ( \9370 , \869 , \8785 );
nand \U$9124 ( \9371 , \9369 , \9370 );
xor \U$9125 ( \9372 , RIbe2a2f8_86, RIbe27ee0_9);
not \U$9126 ( \9373 , \9372 );
not \U$9127 ( \9374 , \8696 );
buf \U$9128 ( \9375 , \9374 );
not \U$9129 ( \9376 , \9375 );
or \U$9130 ( \9377 , \9373 , \9376 );
not \U$9131 ( \9378 , \8705 );
not \U$9132 ( \9379 , \9378 );
nand \U$9133 ( \9380 , \9379 , \8986 );
nand \U$9134 ( \9381 , \9377 , \9380 );
xor \U$9135 ( \9382 , \9371 , \9381 );
not \U$9136 ( \9383 , \9382 );
or \U$9137 ( \9384 , \9366 , \9383 );
nand \U$9138 ( \9385 , \9371 , \9381 );
nand \U$9139 ( \9386 , \9384 , \9385 );
not \U$9140 ( \9387 , \9386 );
or \U$9141 ( \9388 , \9185 , \9197 );
nand \U$9142 ( \9389 , \9388 , \9187 );
or \U$9143 ( \9390 , \9217 , \9224 );
nand \U$9144 ( \9391 , \9390 , \9219 );
xor \U$9145 ( \9392 , \9389 , \9391 );
not \U$9146 ( \9393 , \9392 );
or \U$9147 ( \9394 , \9387 , \9393 );
nand \U$9148 ( \9395 , \9391 , \9389 );
nand \U$9149 ( \9396 , \9394 , \9395 );
xor \U$9150 ( \9397 , \8708 , \8728 );
xor \U$9151 ( \9398 , \9397 , \8730 );
xor \U$9152 ( \9399 , \8537 , \8528 );
xor \U$9153 ( \9400 , \9399 , \8545 );
xor \U$9154 ( \9401 , \9398 , \9400 );
xor \U$9155 ( \9402 , \9396 , \9401 );
xor \U$9156 ( \9403 , \9360 , \9402 );
not \U$9157 ( \9404 , \9403 );
or \U$9158 ( \9405 , \9232 , \9404 );
nand \U$9159 ( \9406 , \9402 , \9360 );
nand \U$9160 ( \9407 , \9405 , \9406 );
not \U$9161 ( \9408 , \9407 );
or \U$9162 ( \9409 , \9010 , \9408 );
nand \U$9163 ( \9410 , \8783 , \9007 );
nand \U$9164 ( \9411 , \9409 , \9410 );
xnor \U$9165 ( \9412 , \8386 , \8370 );
not \U$9166 ( \9413 , \9412 );
not \U$9167 ( \9414 , \8890 );
not \U$9168 ( \9415 , \1793 );
or \U$9169 ( \9416 , \9414 , \9415 );
nand \U$9170 ( \9417 , \1199 , \8411 );
nand \U$9171 ( \9418 , \9416 , \9417 );
not \U$9172 ( \9419 , \9378 );
not \U$9173 ( \9420 , \8988 );
or \U$9174 ( \9421 , \9419 , \9420 );
nand \U$9175 ( \9422 , \9421 , RIbe2a2f8_86);
or \U$9176 ( \9423 , \9418 , \9422 );
not \U$9177 ( \9424 , \8543 );
not \U$9178 ( \9425 , \936 );
or \U$9179 ( \9426 , \9424 , \9425 );
not \U$9180 ( \9427 , \8357 );
nand \U$9181 ( \9428 , \9427 , \370 );
nand \U$9182 ( \9429 , \9426 , \9428 );
nand \U$9183 ( \9430 , \9423 , \9429 );
nand \U$9184 ( \9431 , \9418 , \9422 );
nand \U$9185 ( \9432 , \9430 , \9431 );
not \U$9186 ( \9433 , \8780 );
not \U$9187 ( \9434 , \8773 );
or \U$9188 ( \9435 , \9433 , \9434 );
nand \U$9189 ( \9436 , \8772 , \8765 );
nand \U$9190 ( \9437 , \9435 , \9436 );
xor \U$9191 ( \9438 , \9432 , \9437 );
not \U$9192 ( \9439 , \9438 );
or \U$9193 ( \9440 , \9413 , \9439 );
or \U$9194 ( \9441 , \9438 , \9412 );
nand \U$9195 ( \9442 , \9440 , \9441 );
not \U$9196 ( \9443 , \9442 );
not \U$9197 ( \9444 , \8781 );
not \U$9198 ( \9445 , \8759 );
or \U$9199 ( \9446 , \9444 , \9445 );
not \U$9200 ( \9447 , \8749 );
nand \U$9201 ( \9448 , \9447 , \8732 );
nand \U$9202 ( \9449 , \9446 , \9448 );
not \U$9203 ( \9450 , \9449 );
not \U$9204 ( \9451 , \9450 );
or \U$9205 ( \9452 , \9443 , \9451 );
not \U$9206 ( \9453 , \9442 );
nand \U$9207 ( \9454 , \9453 , \9449 );
nand \U$9208 ( \9455 , \9452 , \9454 );
not \U$9209 ( \9456 , \8160 );
not \U$9210 ( \9457 , \8621 );
not \U$9211 ( \9458 , \9457 );
not \U$9212 ( \9459 , \8640 );
or \U$9213 ( \9460 , \9458 , \9459 );
nand \U$9214 ( \9461 , \8635 , \8628 );
nand \U$9215 ( \9462 , \9460 , \9461 );
xor \U$9216 ( \9463 , \9456 , \9462 );
not \U$9217 ( \9464 , \8670 );
not \U$9218 ( \9465 , \8683 );
or \U$9219 ( \9466 , \9464 , \9465 );
nand \U$9220 ( \9467 , \8675 , \8682 );
nand \U$9221 ( \9468 , \9466 , \9467 );
xor \U$9222 ( \9469 , \9463 , \9468 );
xor \U$9223 ( \9470 , \9455 , \9469 );
not \U$9224 ( \9471 , \9470 );
xor \U$9225 ( \9472 , \8649 , \8656 );
and \U$9226 ( \9473 , \9472 , \8663 );
and \U$9227 ( \9474 , \8649 , \8656 );
or \U$9228 ( \9475 , \9473 , \9474 );
xor \U$9229 ( \9476 , RIbe28f48_44, RIbe284f8_22);
not \U$9230 ( \9477 , \9476 );
not \U$9231 ( \9478 , \8221 );
or \U$9232 ( \9479 , \9477 , \9478 );
nand \U$9233 ( \9480 , \4181 , \8219 );
nand \U$9234 ( \9481 , \9479 , \9480 );
not \U$9235 ( \9482 , \9481 );
not \U$9236 ( \9483 , \8717 );
not \U$9237 ( \9484 , \2554 );
or \U$9238 ( \9485 , \9483 , \9484 );
nand \U$9239 ( \9486 , \2560 , \8155 );
nand \U$9240 ( \9487 , \9485 , \9486 );
not \U$9241 ( \9488 , \9487 );
or \U$9242 ( \9489 , \9482 , \9488 );
or \U$9243 ( \9490 , \9487 , \9481 );
not \U$9244 ( \9491 , \8726 );
not \U$9245 ( \9492 , \2731 );
or \U$9246 ( \9493 , \9491 , \9492 );
nand \U$9247 ( \9494 , \2071 , \8391 );
nand \U$9248 ( \9495 , \9493 , \9494 );
nand \U$9249 ( \9496 , \9490 , \9495 );
nand \U$9250 ( \9497 , \9489 , \9496 );
xor \U$9251 ( \9498 , \9475 , \9497 );
not \U$9252 ( \9499 , \8740 );
not \U$9253 ( \9500 , \8748 );
or \U$9254 ( \9501 , \9499 , \9500 );
nand \U$9255 ( \9502 , \8747 , \8741 );
nand \U$9256 ( \9503 , \9501 , \9502 );
xor \U$9257 ( \9504 , \9498 , \9503 );
xor \U$9258 ( \9505 , \8644 , \8664 );
and \U$9259 ( \9506 , \9505 , \8684 );
and \U$9260 ( \9507 , \8644 , \8664 );
or \U$9261 ( \9508 , \9506 , \9507 );
nand \U$9262 ( \9509 , \9504 , \9508 );
not \U$9263 ( \9510 , \9508 );
not \U$9264 ( \9511 , \9504 );
nand \U$9265 ( \9512 , \9510 , \9511 );
nand \U$9266 ( \9513 , \9509 , \9512 );
xor \U$9267 ( \9514 , \9422 , \9429 );
xor \U$9268 ( \9515 , \9514 , \9418 );
xor \U$9269 ( \9516 , \9487 , \9481 );
xor \U$9270 ( \9517 , \9516 , \9495 );
xor \U$9271 ( \9518 , \9515 , \9517 );
xor \U$9272 ( \9519 , RIbe28f48_44, RIbe28318_18);
not \U$9273 ( \9520 , \9519 );
not \U$9274 ( \9521 , \8221 );
or \U$9275 ( \9522 , \9520 , \9521 );
not \U$9276 ( \9523 , \3252 );
buf \U$9277 ( \9524 , \9523 );
nand \U$9278 ( \9525 , \9524 , \9476 );
nand \U$9279 ( \9526 , \9522 , \9525 );
not \U$9280 ( \9527 , \8931 );
not \U$9281 ( \9528 , \8168 );
buf \U$9282 ( \9529 , \9528 );
not \U$9283 ( \9530 , \9529 );
buf \U$9284 ( \9531 , \9530 );
not \U$9285 ( \9532 , \9531 );
or \U$9286 ( \9533 , \9527 , \9532 );
nand \U$9287 ( \9534 , \8172 , \8398 );
nand \U$9288 ( \9535 , \9533 , \9534 );
xor \U$9289 ( \9536 , \9526 , \9535 );
not \U$9290 ( \9537 , \8241 );
not \U$9291 ( \9538 , \8245 );
or \U$9292 ( \9539 , \9537 , \9538 );
or \U$9293 ( \9540 , \7371 , \8588 );
nand \U$9294 ( \9541 , \9539 , \9540 );
xor \U$9295 ( \9542 , \9536 , \9541 );
and \U$9296 ( \9543 , \9518 , \9542 );
and \U$9297 ( \9544 , \9515 , \9517 );
or \U$9298 ( \9545 , \9543 , \9544 );
not \U$9299 ( \9546 , \9545 );
and \U$9300 ( \9547 , \9513 , \9546 );
not \U$9301 ( \9548 , \9513 );
not \U$9302 ( \9549 , \9546 );
and \U$9303 ( \9550 , \9548 , \9549 );
nor \U$9304 ( \9551 , \9547 , \9550 );
not \U$9305 ( \9552 , \9551 );
or \U$9306 ( \9553 , \9471 , \9552 );
or \U$9307 ( \9554 , \9470 , \9551 );
nand \U$9308 ( \9555 , \9553 , \9554 );
not \U$9309 ( \9556 , \9555 );
xor \U$9310 ( \9557 , \8263 , \8284 );
not \U$9311 ( \9558 , \8252 );
and \U$9312 ( \9559 , \8248 , \9558 );
not \U$9313 ( \9560 , \8248 );
and \U$9314 ( \9561 , \9560 , \8252 );
nor \U$9315 ( \9562 , \9559 , \9561 );
xnor \U$9316 ( \9563 , \9557 , \9562 );
not \U$9317 ( \9564 , \8211 );
and \U$9318 ( \9565 , \8226 , \9564 );
not \U$9319 ( \9566 , \8226 );
and \U$9320 ( \9567 , \9566 , \8211 );
nor \U$9321 ( \9568 , \9565 , \9567 );
xor \U$9322 ( \9569 , \9563 , \9568 );
not \U$9323 ( \9570 , \9569 );
xor \U$9324 ( \9571 , \8396 , \8405 );
xor \U$9325 ( \9572 , \9571 , \8416 );
not \U$9326 ( \9573 , \9572 );
not \U$9327 ( \9574 , \9573 );
xnor \U$9328 ( \9575 , \8196 , \8187 );
not \U$9329 ( \9576 , \9575 );
not \U$9330 ( \9577 , \9576 );
or \U$9331 ( \9578 , \9574 , \9577 );
nand \U$9332 ( \9579 , \9572 , \9575 );
nand \U$9333 ( \9580 , \9578 , \9579 );
xor \U$9334 ( \9581 , \8352 , \8346 );
xor \U$9335 ( \9582 , \9581 , \8360 );
not \U$9336 ( \9583 , \9582 );
and \U$9337 ( \9584 , \9580 , \9583 );
not \U$9338 ( \9585 , \9580 );
and \U$9339 ( \9586 , \9585 , \9582 );
or \U$9340 ( \9587 , \9584 , \9586 );
not \U$9341 ( \9588 , \9587 );
or \U$9342 ( \9589 , \9570 , \9588 );
or \U$9343 ( \9590 , \9587 , \9569 );
nand \U$9344 ( \9591 , \9589 , \9590 );
not \U$9345 ( \9592 , \9591 );
nand \U$9346 ( \9593 , RIbe27b98_2, RIbe2a820_97);
nand \U$9347 ( \9594 , \9526 , \9593 );
not \U$9348 ( \9595 , \9594 );
not \U$9349 ( \9596 , \9154 );
not \U$9350 ( \9597 , \9151 );
or \U$9351 ( \9598 , \9596 , \9597 );
nand \U$9352 ( \9599 , \9598 , \9162 );
nand \U$9353 ( \9600 , \9150 , \9143 );
nand \U$9354 ( \9601 , \9599 , \9600 );
not \U$9355 ( \9602 , \9601 );
or \U$9356 ( \9603 , \9595 , \9602 );
nor \U$9357 ( \9604 , \9526 , \9593 );
not \U$9358 ( \9605 , \9604 );
nand \U$9359 ( \9606 , \9603 , \9605 );
xor \U$9360 ( \9607 , \8823 , \8849 );
and \U$9361 ( \9608 , \9607 , \8875 );
and \U$9362 ( \9609 , \8823 , \8849 );
or \U$9363 ( \9610 , \9608 , \9609 );
xor \U$9364 ( \9611 , \9606 , \9610 );
not \U$9365 ( \9612 , \9190 );
not \U$9366 ( \9613 , \9194 );
or \U$9367 ( \9614 , \9612 , \9613 );
nand \U$9368 ( \9615 , \2475 , \8916 );
nand \U$9369 ( \9616 , \9614 , \9615 );
not \U$9370 ( \9617 , \9176 );
not \U$9371 ( \9618 , \3255 );
not \U$9372 ( \9619 , \9618 );
or \U$9373 ( \9620 , \9617 , \9619 );
nand \U$9374 ( \9621 , \4181 , \9519 );
nand \U$9375 ( \9622 , \9620 , \9621 );
xor \U$9376 ( \9623 , \9616 , \9622 );
not \U$9377 ( \9624 , \9117 );
not \U$9378 ( \9625 , \386 );
or \U$9379 ( \9626 , \9624 , \9625 );
nand \U$9380 ( \9627 , \399 , \8722 );
nand \U$9381 ( \9628 , \9626 , \9627 );
and \U$9382 ( \9629 , \9623 , \9628 );
and \U$9383 ( \9630 , \9616 , \9622 );
or \U$9384 ( \9631 , \9629 , \9630 );
not \U$9385 ( \9632 , \9631 );
not \U$9386 ( \9633 , \9058 );
not \U$9387 ( \9634 , \3401 );
or \U$9388 ( \9635 , \9633 , \9634 );
not \U$9389 ( \9636 , \8714 );
nand \U$9390 ( \9637 , \9636 , \2560 );
nand \U$9391 ( \9638 , \9635 , \9637 );
not \U$9392 ( \9639 , \9638 );
not \U$9393 ( \9640 , \9034 );
not \U$9394 ( \9641 , \8531 );
or \U$9395 ( \9642 , \9640 , \9641 );
nand \U$9396 ( \9643 , \907 , \8529 );
nand \U$9397 ( \9644 , \9642 , \9643 );
not \U$9398 ( \9645 , \9073 );
not \U$9399 ( \9646 , \281 );
or \U$9400 ( \9647 , \9645 , \9646 );
nand \U$9401 ( \9648 , \286 , \8910 );
nand \U$9402 ( \9649 , \9647 , \9648 );
xor \U$9403 ( \9650 , \9644 , \9649 );
not \U$9404 ( \9651 , \9650 );
or \U$9405 ( \9652 , \9639 , \9651 );
nand \U$9406 ( \9653 , \9649 , \9644 );
nand \U$9407 ( \9654 , \9652 , \9653 );
not \U$9408 ( \9655 , \9124 );
not \U$9409 ( \9656 , \2519 );
or \U$9410 ( \9657 , \9655 , \9656 );
nand \U$9411 ( \9658 , \2527 , \8953 );
nand \U$9412 ( \9659 , \9657 , \9658 );
not \U$9413 ( \9660 , \9659 );
and \U$9414 ( \9661 , RIbe27b98_2, RIbe2a118_82);
not \U$9415 ( \9662 , \9132 );
not \U$9416 ( \9663 , \331 );
or \U$9417 ( \9664 , \9662 , \9663 );
nand \U$9418 ( \9665 , \347 , \8959 );
nand \U$9419 ( \9666 , \9664 , \9665 );
xor \U$9420 ( \9667 , \9661 , \9666 );
not \U$9421 ( \9668 , \9667 );
or \U$9422 ( \9669 , \9660 , \9668 );
nand \U$9423 ( \9670 , RIbe27b98_2, RIbe2a118_82, \9666 );
nand \U$9424 ( \9671 , \9669 , \9670 );
and \U$9425 ( \9672 , \9654 , \9671 );
not \U$9426 ( \9673 , \9654 );
not \U$9427 ( \9674 , \9671 );
and \U$9428 ( \9675 , \9673 , \9674 );
nor \U$9429 ( \9676 , \9672 , \9675 );
not \U$9430 ( \9677 , \9676 );
or \U$9431 ( \9678 , \9632 , \9677 );
nand \U$9432 ( \9679 , \9671 , \9654 );
nand \U$9433 ( \9680 , \9678 , \9679 );
and \U$9434 ( \9681 , \9611 , \9680 );
and \U$9435 ( \9682 , \9606 , \9610 );
or \U$9436 ( \9683 , \9681 , \9682 );
not \U$9437 ( \9684 , \9683 );
not \U$9438 ( \9685 , \9684 );
and \U$9439 ( \9686 , \9592 , \9685 );
and \U$9440 ( \9687 , \9591 , \9684 );
nor \U$9441 ( \9688 , \9686 , \9687 );
not \U$9442 ( \9689 , \9688 );
and \U$9443 ( \9690 , \9556 , \9689 );
and \U$9444 ( \9691 , \9555 , \9688 );
nor \U$9445 ( \9692 , \9690 , \9691 );
xor \U$9446 ( \9693 , \9411 , \9692 );
xor \U$9447 ( \9694 , \9111 , \9137 );
and \U$9448 ( \9695 , \9694 , \9167 );
and \U$9449 ( \9696 , \9111 , \9137 );
or \U$9450 ( \9697 , \9695 , \9696 );
and \U$9451 ( \9698 , \9650 , \9638 );
not \U$9452 ( \9699 , \9650 );
not \U$9453 ( \9700 , \9638 );
and \U$9454 ( \9701 , \9699 , \9700 );
nor \U$9455 ( \9702 , \9698 , \9701 );
xor \U$9456 ( \9703 , \9616 , \9622 );
xor \U$9457 ( \9704 , \9703 , \9628 );
xor \U$9458 ( \9705 , \9702 , \9704 );
xor \U$9459 ( \9706 , \8978 , \8984 );
xor \U$9460 ( \9707 , \9706 , \8993 );
and \U$9461 ( \9708 , \9705 , \9707 );
and \U$9462 ( \9709 , \9702 , \9704 );
or \U$9463 ( \9710 , \9708 , \9709 );
xor \U$9464 ( \9711 , \9697 , \9710 );
xor \U$9465 ( \9712 , \9667 , \9659 );
xor \U$9466 ( \9713 , \8847 , \8829 );
xor \U$9467 ( \9714 , \9713 , \8837 );
xor \U$9468 ( \9715 , \9712 , \9714 );
xor \U$9469 ( \9716 , \8871 , \8856 );
and \U$9470 ( \9717 , \9715 , \9716 );
and \U$9471 ( \9718 , \9712 , \9714 );
or \U$9472 ( \9719 , \9717 , \9718 );
xor \U$9473 ( \9720 , \9711 , \9719 );
not \U$9474 ( \9721 , \9720 );
xor \U$9475 ( \9722 , \9365 , \9382 );
not \U$9476 ( \9723 , \9722 );
xor \U$9477 ( \9724 , RIbe2a550_91, RIbe2a988_100);
buf \U$9478 ( \9725 , \9724 );
buf \U$9479 ( \9726 , \9725 );
not \U$9480 ( \9727 , RIbe2a910_99);
not \U$9481 ( \9728 , \9727 );
nand \U$9482 ( \9729 , RIbe2a550_91, RIbe2a988_100);
not \U$9483 ( \9730 , \9729 );
not \U$9484 ( \9731 , \9730 );
or \U$9485 ( \9732 , \9728 , \9731 );
nor \U$9486 ( \9733 , RIbe2a550_91, RIbe2a988_100);
nand \U$9487 ( \9734 , \9733 , RIbe2a910_99);
nand \U$9488 ( \9735 , \9732 , \9734 );
buf \U$9489 ( \9736 , \9735 );
buf \U$9490 ( \9737 , \9736 );
buf \U$9491 ( \9738 , \9737 );
or \U$9492 ( \9739 , \9726 , \9738 );
nand \U$9493 ( \9740 , \9739 , RIbe2a910_99);
not \U$9494 ( \9741 , \9740 );
xor \U$9495 ( \9742 , RIbe29308_52, RIbe28f48_44);
not \U$9496 ( \9743 , \9742 );
not \U$9497 ( \9744 , \9618 );
or \U$9498 ( \9745 , \9743 , \9744 );
nand \U$9499 ( \9746 , \9524 , \9172 );
nand \U$9500 ( \9747 , \9745 , \9746 );
not \U$9501 ( \9748 , \9747 );
xor \U$9502 ( \9749 , RIbe29a10_67, RIbe28a20_33);
not \U$9503 ( \9750 , \9749 );
not \U$9504 ( \9751 , \7795 );
or \U$9505 ( \9752 , \9750 , \9751 );
nand \U$9506 ( \9753 , \5055 , \9195 );
nand \U$9507 ( \9754 , \9752 , \9753 );
not \U$9508 ( \9755 , \9754 );
not \U$9509 ( \9756 , \9755 );
or \U$9510 ( \9757 , \9748 , \9756 );
or \U$9511 ( \9758 , \9747 , \9755 );
nand \U$9512 ( \9759 , \9757 , \9758 );
not \U$9513 ( \9760 , \9759 );
or \U$9514 ( \9761 , \9741 , \9760 );
nand \U$9515 ( \9762 , \9754 , \9747 );
nand \U$9516 ( \9763 , \9761 , \9762 );
nand \U$9517 ( \9764 , RIbe27b98_2, RIbe2b360_121);
not \U$9518 ( \9765 , \9764 );
not \U$9519 ( \9766 , \9765 );
xor \U$9520 ( \9767 , RIbe2a820_97, RIbe28de0_41);
not \U$9521 ( \9768 , \9767 );
not \U$9522 ( \9769 , \331 );
or \U$9523 ( \9770 , \9768 , \9769 );
nand \U$9524 ( \9771 , \347 , \9128 );
nand \U$9525 ( \9772 , \9770 , \9771 );
not \U$9526 ( \9773 , \9772 );
or \U$9527 ( \9774 , \9766 , \9773 );
xor \U$9528 ( \9775 , \9772 , \9764 );
not \U$9529 ( \9776 , \9775 );
xor \U$9530 ( \9777 , RIbe28480_21, RIbe297b8_62);
not \U$9531 ( \9778 , \9777 );
not \U$9532 ( \9779 , \3344 );
or \U$9533 ( \9780 , \9778 , \9779 );
nand \U$9534 ( \9781 , \3075 , \9120 );
nand \U$9535 ( \9782 , \9780 , \9781 );
nand \U$9536 ( \9783 , \9776 , \9782 );
nand \U$9537 ( \9784 , \9774 , \9783 );
xor \U$9538 ( \9785 , \9763 , \9784 );
not \U$9539 ( \9786 , \9785 );
or \U$9540 ( \9787 , \9723 , \9786 );
nand \U$9541 ( \9788 , \9763 , \9784 );
nand \U$9542 ( \9789 , \9787 , \9788 );
not \U$9543 ( \9790 , \9789 );
xor \U$9544 ( \9791 , RIbe27b20_1, RIbe296c8_60);
not \U$9545 ( \9792 , \9791 );
not \U$9546 ( \9793 , \898 );
not \U$9547 ( \9794 , \9793 );
or \U$9548 ( \9795 , \9792 , \9794 );
nand \U$9549 ( \9796 , \907 , \9030 );
nand \U$9550 ( \9797 , \9795 , \9796 );
not \U$9551 ( \9798 , \9797 );
xor \U$9552 ( \9799 , RIbe29038_46, RIbe29ce0_73);
not \U$9553 ( \9800 , \9799 );
not \U$9554 ( \9801 , \281 );
or \U$9555 ( \9802 , \9800 , \9801 );
nand \U$9556 ( \9803 , \1583 , \9069 );
nand \U$9557 ( \9804 , \9802 , \9803 );
not \U$9558 ( \9805 , \9804 );
or \U$9559 ( \9806 , \9798 , \9805 );
or \U$9560 ( \9807 , \9804 , \9797 );
xor \U$9561 ( \9808 , RIbe29ec0_77, RIbe290b0_47);
not \U$9562 ( \9809 , \9808 );
not \U$9563 ( \9810 , \9114 );
or \U$9564 ( \9811 , \9809 , \9810 );
nand \U$9565 ( \9812 , \2071 , \9112 );
nand \U$9566 ( \9813 , \9811 , \9812 );
nand \U$9567 ( \9814 , \9807 , \9813 );
nand \U$9568 ( \9815 , \9806 , \9814 );
xor \U$9569 ( \9816 , RIbe2b6a8_128, RIbe27d78_6);
not \U$9570 ( \9817 , \9816 );
not \U$9571 ( \9818 , \1164 );
or \U$9572 ( \9819 , \9817 , \9818 );
nand \U$9573 ( \9820 , \314 , \9179 );
nand \U$9574 ( \9821 , \9819 , \9820 );
not \U$9575 ( \9822 , \9821 );
xor \U$9576 ( \9823 , RIbe27fd0_11, RIbe28a98_34);
not \U$9577 ( \9824 , \9823 );
not \U$9578 ( \9825 , \2717 );
not \U$9579 ( \9826 , \9825 );
or \U$9580 ( \9827 , \9824 , \9826 );
nand \U$9581 ( \9828 , \4897 , \9080 );
nand \U$9582 ( \9829 , \9827 , \9828 );
not \U$9583 ( \9830 , \9829 );
xor \U$9584 ( \9831 , RIbe27b98_2, RIbe2a0a0_81);
not \U$9585 ( \9832 , \9831 );
and \U$9586 ( \9833 , \252 , \250 , \253 );
not \U$9587 ( \9834 , \9833 );
or \U$9588 ( \9835 , \9832 , \9834 );
nand \U$9589 ( \9836 , \9210 , \267 );
nand \U$9590 ( \9837 , \9835 , \9836 );
not \U$9591 ( \9838 , \9837 );
nand \U$9592 ( \9839 , \9830 , \9838 );
not \U$9593 ( \9840 , \9839 );
or \U$9594 ( \9841 , \9822 , \9840 );
nand \U$9595 ( \9842 , \9829 , \9837 );
nand \U$9596 ( \9843 , \9841 , \9842 );
or \U$9597 ( \9844 , \9815 , \9843 );
xor \U$9598 ( \9845 , RIbe286d8_26, RIbe2a2f8_86);
not \U$9599 ( \9846 , \9845 );
not \U$9600 ( \9847 , \9375 );
or \U$9601 ( \9848 , \9846 , \9847 );
nand \U$9602 ( \9849 , \8706 , \9372 );
nand \U$9603 ( \9850 , \9848 , \9849 );
not \U$9604 ( \9851 , \9850 );
xor \U$9605 ( \9852 , RIbe28930_31, RIbe27df0_7);
and \U$9606 ( \9853 , \9852 , \965 );
and \U$9607 ( \9854 , \1199 , \9102 );
nor \U$9608 ( \9855 , \9853 , \9854 );
xor \U$9609 ( \9856 , RIbe27c10_3, RIbe2aa00_101);
and \U$9610 ( \9857 , \357 , \9856 );
not \U$9611 ( \9858 , \9857 );
not \U$9612 ( \9859 , \1172 );
or \U$9613 ( \9860 , \9858 , \9859 );
nand \U$9614 ( \9861 , \1173 , \9040 );
nand \U$9615 ( \9862 , \9860 , \9861 );
not \U$9616 ( \9863 , \9862 );
and \U$9617 ( \9864 , \9855 , \9863 );
not \U$9618 ( \9865 , \9855 );
and \U$9619 ( \9866 , \9865 , \9862 );
nor \U$9620 ( \9867 , \9864 , \9866 );
not \U$9621 ( \9868 , \9867 );
or \U$9622 ( \9869 , \9851 , \9868 );
not \U$9623 ( \9870 , \9855 );
nand \U$9624 ( \9871 , \9870 , \9862 );
nand \U$9625 ( \9872 , \9869 , \9871 );
nand \U$9626 ( \9873 , \9844 , \9872 );
nand \U$9627 ( \9874 , \9815 , \9843 );
and \U$9628 ( \9875 , \9873 , \9874 );
not \U$9629 ( \9876 , \9875 );
not \U$9630 ( \9877 , \9086 );
not \U$9631 ( \9878 , \9098 );
or \U$9632 ( \9879 , \9877 , \9878 );
or \U$9633 ( \9880 , \9098 , \9086 );
nand \U$9634 ( \9881 , \9879 , \9880 );
not \U$9635 ( \9882 , \9881 );
not \U$9636 ( \9883 , \9106 );
and \U$9637 ( \9884 , \9882 , \9883 );
and \U$9638 ( \9885 , \9881 , \9106 );
nor \U$9639 ( \9886 , \9884 , \9885 );
not \U$9640 ( \9887 , \9886 );
not \U$9641 ( \9888 , \9887 );
xor \U$9642 ( \9889 , \9060 , \9067 );
xor \U$9643 ( \9890 , \9889 , \9075 );
not \U$9644 ( \9891 , \9890 );
or \U$9645 ( \9892 , \9888 , \9891 );
or \U$9646 ( \9893 , \9887 , \9890 );
not \U$9647 ( \9894 , \9027 );
not \U$9648 ( \9895 , \9037 );
or \U$9649 ( \9896 , \9894 , \9895 );
nand \U$9650 ( \9897 , \9028 , \9036 );
nand \U$9651 ( \9898 , \9896 , \9897 );
and \U$9652 ( \9899 , \9898 , \9045 );
not \U$9653 ( \9900 , \9898 );
not \U$9654 ( \9901 , \9045 );
and \U$9655 ( \9902 , \9900 , \9901 );
nor \U$9656 ( \9903 , \9899 , \9902 );
nand \U$9657 ( \9904 , \9893 , \9903 );
nand \U$9658 ( \9905 , \9892 , \9904 );
not \U$9659 ( \9906 , \9905 );
or \U$9660 ( \9907 , \9876 , \9906 );
or \U$9661 ( \9908 , \9905 , \9875 );
nand \U$9662 ( \9909 , \9907 , \9908 );
not \U$9663 ( \9910 , \9909 );
or \U$9664 ( \9911 , \9790 , \9910 );
not \U$9665 ( \9912 , \9875 );
nand \U$9666 ( \9913 , \9912 , \9905 );
nand \U$9667 ( \9914 , \9911 , \9913 );
not \U$9668 ( \9915 , \9914 );
or \U$9669 ( \9916 , \9078 , \9020 );
nand \U$9670 ( \9917 , \9916 , \9048 );
nand \U$9671 ( \9918 , \9078 , \9020 );
nand \U$9672 ( \9919 , \9917 , \9918 );
not \U$9673 ( \9920 , \9919 );
not \U$9674 ( \9921 , \9601 );
not \U$9675 ( \9922 , \9604 );
nand \U$9676 ( \9923 , \9922 , \9594 );
not \U$9677 ( \9924 , \9923 );
and \U$9678 ( \9925 , \9921 , \9924 );
and \U$9679 ( \9926 , \9601 , \9923 );
nor \U$9680 ( \9927 , \9925 , \9926 );
not \U$9681 ( \9928 , \9927 );
or \U$9682 ( \9929 , \9920 , \9928 );
or \U$9683 ( \9930 , \9927 , \9919 );
nand \U$9684 ( \9931 , \9929 , \9930 );
xor \U$9685 ( \9932 , \9676 , \9631 );
xor \U$9686 ( \9933 , \9931 , \9932 );
not \U$9687 ( \9934 , \9933 );
not \U$9688 ( \9935 , \9934 );
or \U$9689 ( \9936 , \9915 , \9935 );
not \U$9690 ( \9937 , \9914 );
nand \U$9691 ( \9938 , \9937 , \9933 );
nand \U$9692 ( \9939 , \9936 , \9938 );
not \U$9693 ( \9940 , \9939 );
or \U$9694 ( \9941 , \9721 , \9940 );
nand \U$9695 ( \9942 , \9933 , \9914 );
nand \U$9696 ( \9943 , \9941 , \9942 );
not \U$9697 ( \9944 , \9931 );
not \U$9698 ( \9945 , \9932 );
or \U$9699 ( \9946 , \9944 , \9945 );
not \U$9700 ( \9947 , \9927 );
nand \U$9701 ( \9948 , \9947 , \9919 );
nand \U$9702 ( \9949 , \9946 , \9948 );
xor \U$9703 ( \9950 , \9606 , \9610 );
xor \U$9704 ( \9951 , \9950 , \9680 );
xor \U$9705 ( \9952 , \9949 , \9951 );
xor \U$9706 ( \9953 , \8958 , \8964 );
and \U$9707 ( \9954 , \9953 , \8971 );
and \U$9708 ( \9955 , \8958 , \8964 );
or \U$9709 ( \9956 , \9954 , \9955 );
not \U$9710 ( \9957 , \8883 );
not \U$9711 ( \9958 , \9957 );
not \U$9712 ( \9959 , \8906 );
or \U$9713 ( \9960 , \9958 , \9959 );
nand \U$9714 ( \9961 , \8902 , \8892 );
nand \U$9715 ( \9962 , \9960 , \9961 );
xor \U$9716 ( \9963 , \9956 , \9962 );
not \U$9717 ( \9964 , \8933 );
not \U$9718 ( \9965 , \8926 );
or \U$9719 ( \9966 , \9964 , \9965 );
nand \U$9720 ( \9967 , \8921 , \8915 );
nand \U$9721 ( \9968 , \9966 , \9967 );
xor \U$9722 ( \9969 , \9963 , \9968 );
not \U$9723 ( \9970 , \8946 );
not \U$9724 ( \9971 , \8939 );
or \U$9725 ( \9972 , \9970 , \9971 );
nand \U$9726 ( \9973 , \8934 , \8907 );
nand \U$9727 ( \9974 , \9972 , \9973 );
xor \U$9728 ( \9975 , \9969 , \9974 );
not \U$9729 ( \9976 , \8999 );
not \U$9730 ( \9977 , \8997 );
or \U$9731 ( \9978 , \9976 , \9977 );
nand \U$9732 ( \9979 , \8972 , \8996 );
nand \U$9733 ( \9980 , \9978 , \9979 );
xor \U$9734 ( \9981 , \9975 , \9980 );
xor \U$9735 ( \9982 , \9952 , \9981 );
nand \U$9736 ( \9983 , \9943 , \9982 );
xor \U$9737 ( \9984 , \9515 , \9517 );
xor \U$9738 ( \9985 , \9984 , \9542 );
not \U$9739 ( \9986 , \9401 );
not \U$9740 ( \9987 , \9396 );
or \U$9741 ( \9988 , \9986 , \9987 );
nand \U$9742 ( \9989 , \9400 , \9398 );
nand \U$9743 ( \9990 , \9988 , \9989 );
xor \U$9744 ( \9991 , \9985 , \9990 );
xor \U$9745 ( \9992 , \9697 , \9710 );
and \U$9746 ( \9993 , \9992 , \9719 );
and \U$9747 ( \9994 , \9697 , \9710 );
or \U$9748 ( \9995 , \9993 , \9994 );
xnor \U$9749 ( \9996 , \9991 , \9995 );
not \U$9750 ( \9997 , \9996 );
nand \U$9751 ( \9998 , \9997 , \9943 );
not \U$9752 ( \9999 , \9996 );
nand \U$9753 ( \10000 , \9999 , \9982 );
nand \U$9754 ( \10001 , \9983 , \9998 , \10000 );
and \U$9755 ( \10002 , \9693 , \10001 );
and \U$9756 ( \10003 , \9411 , \9692 );
or \U$9757 ( \10004 , \10002 , \10003 );
not \U$9758 ( \10005 , \10004 );
xor \U$9759 ( \10006 , \8616 , \8685 );
and \U$9760 ( \10007 , \10006 , \8782 );
and \U$9761 ( \10008 , \8616 , \8685 );
or \U$9762 ( \10009 , \10007 , \10008 );
xor \U$9763 ( \10010 , \9526 , \9535 );
and \U$9764 ( \10011 , \10010 , \9541 );
and \U$9765 ( \10012 , \9526 , \9535 );
or \U$9766 ( \10013 , \10011 , \10012 );
not \U$9767 ( \10014 , \8590 );
not \U$9768 ( \10015 , \8610 );
or \U$9769 ( \10016 , \10014 , \10015 );
nand \U$9770 ( \10017 , \10016 , \8614 );
not \U$9771 ( \10018 , \10017 );
not \U$9772 ( \10019 , \8580 );
or \U$9773 ( \10020 , \10018 , \10019 );
not \U$9774 ( \10021 , \8548 );
nand \U$9775 ( \10022 , \10021 , \8575 );
nand \U$9776 ( \10023 , \10020 , \10022 );
xor \U$9777 ( \10024 , \10013 , \10023 );
xor \U$9778 ( \10025 , \9956 , \9962 );
and \U$9779 ( \10026 , \10025 , \9968 );
and \U$9780 ( \10027 , \9956 , \9962 );
or \U$9781 ( \10028 , \10026 , \10027 );
xor \U$9782 ( \10029 , \10024 , \10028 );
xor \U$9783 ( \10030 , \10009 , \10029 );
xor \U$9784 ( \10031 , \9969 , \9974 );
and \U$9785 ( \10032 , \10031 , \9980 );
and \U$9786 ( \10033 , \9969 , \9974 );
or \U$9787 ( \10034 , \10032 , \10033 );
xor \U$9788 ( \10035 , \10030 , \10034 );
not \U$9789 ( \10036 , \10035 );
not \U$9790 ( \10037 , \9995 );
not \U$9791 ( \10038 , \9991 );
or \U$9792 ( \10039 , \10037 , \10038 );
nand \U$9793 ( \10040 , \9990 , \9985 );
nand \U$9794 ( \10041 , \10039 , \10040 );
xor \U$9795 ( \10042 , \9949 , \9951 );
and \U$9796 ( \10043 , \10042 , \9981 );
and \U$9797 ( \10044 , \9949 , \9951 );
or \U$9798 ( \10045 , \10043 , \10044 );
and \U$9799 ( \10046 , \10041 , \10045 );
not \U$9800 ( \10047 , \10041 );
not \U$9801 ( \10048 , \10045 );
and \U$9802 ( \10049 , \10047 , \10048 );
nor \U$9803 ( \10050 , \10046 , \10049 );
not \U$9804 ( \10051 , \10050 );
or \U$9805 ( \10052 , \10036 , \10051 );
not \U$9806 ( \10053 , \10048 );
nand \U$9807 ( \10054 , \10053 , \10041 );
nand \U$9808 ( \10055 , \10052 , \10054 );
not \U$9809 ( \10056 , \10009 );
not \U$9810 ( \10057 , \10029 );
or \U$9811 ( \10058 , \10056 , \10057 );
or \U$9812 ( \10059 , \10029 , \10009 );
nand \U$9813 ( \10060 , \10059 , \10034 );
nand \U$9814 ( \10061 , \10058 , \10060 );
not \U$9815 ( \10062 , \10061 );
xor \U$9816 ( \10063 , \10013 , \10023 );
and \U$9817 ( \10064 , \10063 , \10028 );
and \U$9818 ( \10065 , \10013 , \10023 );
or \U$9819 ( \10066 , \10064 , \10065 );
not \U$9820 ( \10067 , \8136 );
not \U$9821 ( \10068 , \8148 );
or \U$9822 ( \10069 , \10067 , \10068 );
or \U$9823 ( \10070 , \8148 , \8136 );
nand \U$9824 ( \10071 , \10069 , \10070 );
not \U$9825 ( \10072 , \10071 );
and \U$9826 ( \10073 , \8458 , \8446 );
not \U$9827 ( \10074 , \8458 );
and \U$9828 ( \10075 , \10074 , \8459 );
nor \U$9829 ( \10076 , \10073 , \10075 );
xor \U$9830 ( \10077 , \8455 , \10076 );
not \U$9831 ( \10078 , \10077 );
and \U$9832 ( \10079 , \10072 , \10078 );
and \U$9833 ( \10080 , \10071 , \10077 );
nor \U$9834 ( \10081 , \10079 , \10080 );
not \U$9835 ( \10082 , \10081 );
xor \U$9836 ( \10083 , \10066 , \10082 );
and \U$9837 ( \10084 , \10062 , \10083 );
not \U$9838 ( \10085 , \10062 );
xor \U$9839 ( \10086 , \10066 , \10081 );
and \U$9840 ( \10087 , \10085 , \10086 );
nor \U$9841 ( \10088 , \10084 , \10087 );
xor \U$9842 ( \10089 , \9475 , \9497 );
and \U$9843 ( \10090 , \10089 , \9503 );
and \U$9844 ( \10091 , \9475 , \9497 );
or \U$9845 ( \10092 , \10090 , \10091 );
xor \U$9846 ( \10093 , \7451 , \7436 );
not \U$9847 ( \10094 , \10093 );
not \U$9848 ( \10095 , \8175 );
nand \U$9849 ( \10096 , \10095 , \8203 );
xor \U$9850 ( \10097 , \10096 , \8200 );
not \U$9851 ( \10098 , \10097 );
or \U$9852 ( \10099 , \10094 , \10098 );
or \U$9853 ( \10100 , \10093 , \10097 );
nand \U$9854 ( \10101 , \10099 , \10100 );
xnor \U$9855 ( \10102 , \10092 , \10101 );
not \U$9856 ( \10103 , \10102 );
not \U$9857 ( \10104 , \9469 );
not \U$9858 ( \10105 , \9455 );
or \U$9859 ( \10106 , \10104 , \10105 );
nand \U$9860 ( \10107 , \9449 , \9442 );
nand \U$9861 ( \10108 , \10106 , \10107 );
not \U$9862 ( \10109 , \10108 );
or \U$9863 ( \10110 , \10103 , \10109 );
or \U$9864 ( \10111 , \10108 , \10102 );
nand \U$9865 ( \10112 , \10110 , \10111 );
not \U$9866 ( \10113 , \10112 );
xor \U$9867 ( \10114 , \9456 , \9462 );
and \U$9868 ( \10115 , \10114 , \9468 );
and \U$9869 ( \10116 , \9456 , \9462 );
nor \U$9870 ( \10117 , \10115 , \10116 );
not \U$9871 ( \10118 , \10117 );
not \U$9872 ( \10119 , \8363 );
not \U$9873 ( \10120 , \8419 );
or \U$9874 ( \10121 , \10119 , \10120 );
or \U$9875 ( \10122 , \8363 , \8419 );
nand \U$9876 ( \10123 , \10121 , \10122 );
not \U$9877 ( \10124 , \10123 );
or \U$9878 ( \10125 , \10118 , \10124 );
or \U$9879 ( \10126 , \10123 , \10117 );
nand \U$9880 ( \10127 , \10125 , \10126 );
not \U$9881 ( \10128 , \9563 );
not \U$9882 ( \10129 , \9568 );
not \U$9883 ( \10130 , \10129 );
or \U$9884 ( \10131 , \10128 , \10130 );
not \U$9885 ( \10132 , \9562 );
nand \U$9886 ( \10133 , \10132 , \9557 );
nand \U$9887 ( \10134 , \10131 , \10133 );
xnor \U$9888 ( \10135 , \10127 , \10134 );
not \U$9889 ( \10136 , \10135 );
and \U$9890 ( \10137 , \10113 , \10136 );
and \U$9891 ( \10138 , \10112 , \10135 );
nor \U$9892 ( \10139 , \10137 , \10138 );
xnor \U$9893 ( \10140 , \10088 , \10139 );
xor \U$9894 ( \10141 , \10055 , \10140 );
not \U$9895 ( \10142 , \9683 );
not \U$9896 ( \10143 , \9591 );
or \U$9897 ( \10144 , \10142 , \10143 );
not \U$9898 ( \10145 , \9569 );
nand \U$9899 ( \10146 , \10145 , \9587 );
nand \U$9900 ( \10147 , \10144 , \10146 );
not \U$9901 ( \10148 , \9582 );
not \U$9902 ( \10149 , \9580 );
or \U$9903 ( \10150 , \10148 , \10149 );
nand \U$9904 ( \10151 , \9576 , \9572 );
nand \U$9905 ( \10152 , \10150 , \10151 );
or \U$9906 ( \10153 , \9504 , \9508 );
nand \U$9907 ( \10154 , \10153 , \9545 );
nand \U$9908 ( \10155 , \10154 , \9509 );
xor \U$9909 ( \10156 , \10152 , \10155 );
not \U$9910 ( \10157 , \9438 );
not \U$9911 ( \10158 , \9412 );
not \U$9912 ( \10159 , \10158 );
or \U$9913 ( \10160 , \10157 , \10159 );
nand \U$9914 ( \10161 , \9437 , \9432 );
nand \U$9915 ( \10162 , \10160 , \10161 );
not \U$9916 ( \10163 , \10162 );
xnor \U$9917 ( \10164 , \8292 , \8230 );
not \U$9918 ( \10165 , \10164 );
or \U$9919 ( \10166 , \10163 , \10165 );
or \U$9920 ( \10167 , \10164 , \10162 );
nand \U$9921 ( \10168 , \10166 , \10167 );
not \U$9922 ( \10169 , \10168 );
xnor \U$9923 ( \10170 , \10156 , \10169 );
xor \U$9924 ( \10171 , \10147 , \10170 );
nor \U$9925 ( \10172 , \9470 , \9551 );
or \U$9926 ( \10173 , \10172 , \9688 );
nand \U$9927 ( \10174 , \9470 , \9551 );
nand \U$9928 ( \10175 , \10173 , \10174 );
not \U$9929 ( \10176 , \10175 );
and \U$9930 ( \10177 , \10171 , \10176 );
not \U$9931 ( \10178 , \10171 );
and \U$9932 ( \10179 , \10178 , \10175 );
or \U$9933 ( \10180 , \10177 , \10179 );
xnor \U$9934 ( \10181 , \10141 , \10180 );
not \U$9935 ( \10182 , \10181 );
or \U$9936 ( \10183 , \10005 , \10182 );
not \U$9937 ( \10184 , \10140 );
xor \U$9938 ( \10185 , \10055 , \10180 );
nand \U$9939 ( \10186 , \10184 , \10185 );
nand \U$9940 ( \10187 , \10183 , \10186 );
not \U$9941 ( \10188 , \10187 );
xor \U$9942 ( \10189 , \8298 , \8153 );
not \U$9943 ( \10190 , \10081 );
nand \U$9944 ( \10191 , \10190 , \10066 );
not \U$9945 ( \10192 , \10077 );
nand \U$9946 ( \10193 , \10192 , \10071 );
and \U$9947 ( \10194 , \10191 , \10193 );
xor \U$9948 ( \10195 , \10189 , \10194 );
xnor \U$9949 ( \10196 , \8423 , \8339 );
not \U$9950 ( \10197 , \10152 );
not \U$9951 ( \10198 , \10168 );
or \U$9952 ( \10199 , \10197 , \10198 );
not \U$9953 ( \10200 , \10164 );
nand \U$9954 ( \10201 , \10200 , \10162 );
nand \U$9955 ( \10202 , \10199 , \10201 );
xnor \U$9956 ( \10203 , \10196 , \10202 );
xnor \U$9957 ( \10204 , \10195 , \10203 );
not \U$9958 ( \10205 , \10135 );
not \U$9959 ( \10206 , \10205 );
not \U$9960 ( \10207 , \10112 );
or \U$9961 ( \10208 , \10206 , \10207 );
not \U$9962 ( \10209 , \10102 );
nand \U$9963 ( \10210 , \10209 , \10108 );
nand \U$9964 ( \10211 , \10208 , \10210 );
not \U$9965 ( \10212 , \10211 );
and \U$9966 ( \10213 , \10204 , \10212 );
not \U$9967 ( \10214 , \10204 );
and \U$9968 ( \10215 , \10214 , \10211 );
nor \U$9969 ( \10216 , \10213 , \10215 );
not \U$9970 ( \10217 , \10216 );
not \U$9971 ( \10218 , \10217 );
or \U$9972 ( \10219 , \10139 , \10088 );
not \U$9973 ( \10220 , \10062 );
nand \U$9974 ( \10221 , \10220 , \10083 );
nand \U$9975 ( \10222 , \10219 , \10221 );
not \U$9976 ( \10223 , \10092 );
not \U$9977 ( \10224 , \10101 );
or \U$9978 ( \10225 , \10223 , \10224 );
not \U$9979 ( \10226 , \10097 );
nand \U$9980 ( \10227 , \10226 , \10093 );
nand \U$9981 ( \10228 , \10225 , \10227 );
not \U$9982 ( \10229 , \7994 );
not \U$9983 ( \10230 , \8007 );
or \U$9984 ( \10231 , \10229 , \10230 );
or \U$9985 ( \10232 , \8007 , \7994 );
nand \U$9986 ( \10233 , \10231 , \10232 );
not \U$9987 ( \10234 , \10233 );
xor \U$9988 ( \10235 , \8034 , \8036 );
buf \U$9989 ( \10236 , \8041 );
xnor \U$9990 ( \10237 , \10235 , \10236 );
not \U$9991 ( \10238 , \10237 );
and \U$9992 ( \10239 , \10234 , \10238 );
and \U$9993 ( \10240 , \10233 , \10237 );
nor \U$9994 ( \10241 , \10239 , \10240 );
xor \U$9995 ( \10242 , \10228 , \10241 );
not \U$9996 ( \10243 , \10242 );
buf \U$9997 ( \10244 , \8466 );
not \U$9998 ( \10245 , \8429 );
and \U$9999 ( \10246 , \10244 , \10245 );
not \U$10000 ( \10247 , \10244 );
and \U$10001 ( \10248 , \10247 , \8429 );
nor \U$10002 ( \10249 , \10246 , \10248 );
not \U$10003 ( \10250 , \10249 );
not \U$10004 ( \10251 , \10134 );
not \U$10005 ( \10252 , \10127 );
or \U$10006 ( \10253 , \10251 , \10252 );
not \U$10007 ( \10254 , \10117 );
nand \U$10008 ( \10255 , \10254 , \10123 );
nand \U$10009 ( \10256 , \10253 , \10255 );
not \U$10010 ( \10257 , \10256 );
or \U$10011 ( \10258 , \10250 , \10257 );
or \U$10012 ( \10259 , \10256 , \10249 );
nand \U$10013 ( \10260 , \10258 , \10259 );
not \U$10014 ( \10261 , \10260 );
or \U$10015 ( \10262 , \10243 , \10261 );
or \U$10016 ( \10263 , \10260 , \10242 );
nand \U$10017 ( \10264 , \10262 , \10263 );
not \U$10018 ( \10265 , \10147 );
not \U$10019 ( \10266 , \10170 );
or \U$10020 ( \10267 , \10265 , \10266 );
not \U$10021 ( \10268 , \10152 );
nand \U$10022 ( \10269 , \10268 , \10168 );
not \U$10023 ( \10270 , \10269 );
nand \U$10024 ( \10271 , \10169 , \10152 );
not \U$10025 ( \10272 , \10271 );
or \U$10026 ( \10273 , \10270 , \10272 );
nand \U$10027 ( \10274 , \10273 , \10155 );
nand \U$10028 ( \10275 , \10267 , \10274 );
xor \U$10029 ( \10276 , \10264 , \10275 );
xor \U$10030 ( \10277 , \10222 , \10276 );
not \U$10031 ( \10278 , \10277 );
not \U$10032 ( \10279 , \10278 );
or \U$10033 ( \10280 , \10218 , \10279 );
nand \U$10034 ( \10281 , \10277 , \10216 );
nand \U$10035 ( \10282 , \10280 , \10281 );
not \U$10036 ( \10283 , \10055 );
not \U$10037 ( \10284 , \10180 );
or \U$10038 ( \10285 , \10283 , \10284 );
nand \U$10039 ( \10286 , \10171 , \10175 );
nand \U$10040 ( \10287 , \10285 , \10286 );
xnor \U$10041 ( \10288 , \10282 , \10287 );
nand \U$10042 ( \10289 , \10188 , \10288 );
not \U$10043 ( \10290 , \10287 );
not \U$10044 ( \10291 , \10282 );
or \U$10045 ( \10292 , \10290 , \10291 );
nand \U$10046 ( \10293 , \10277 , \10217 );
nand \U$10047 ( \10294 , \10292 , \10293 );
not \U$10048 ( \10295 , \10294 );
not \U$10049 ( \10296 , \10241 );
nand \U$10050 ( \10297 , \10296 , \10228 );
not \U$10051 ( \10298 , \10237 );
nand \U$10052 ( \10299 , \10298 , \10233 );
and \U$10053 ( \10300 , \10297 , \10299 );
xor \U$10054 ( \10301 , \8326 , \8475 );
xor \U$10055 ( \10302 , \10300 , \10301 );
not \U$10056 ( \10303 , \10189 );
not \U$10057 ( \10304 , \10203 );
or \U$10058 ( \10305 , \10303 , \10304 );
not \U$10059 ( \10306 , \10196 );
nand \U$10060 ( \10307 , \10306 , \10202 );
nand \U$10061 ( \10308 , \10305 , \10307 );
xnor \U$10062 ( \10309 , \10302 , \10308 );
not \U$10063 ( \10310 , \10242 );
not \U$10064 ( \10311 , \10310 );
not \U$10065 ( \10312 , \10260 );
or \U$10066 ( \10313 , \10311 , \10312 );
not \U$10067 ( \10314 , \10249 );
nand \U$10068 ( \10315 , \10314 , \10256 );
nand \U$10069 ( \10316 , \10313 , \10315 );
xor \U$10070 ( \10317 , \8309 , \8307 );
nor \U$10071 ( \10318 , \10316 , \10317 );
not \U$10072 ( \10319 , \10318 );
nand \U$10073 ( \10320 , \10316 , \10317 );
nand \U$10074 ( \10321 , \10319 , \10320 );
not \U$10075 ( \10322 , \10321 );
and \U$10076 ( \10323 , \10309 , \10322 );
not \U$10077 ( \10324 , \10309 );
and \U$10078 ( \10325 , \10324 , \10321 );
nor \U$10079 ( \10326 , \10323 , \10325 );
not \U$10080 ( \10327 , \10326 );
not \U$10081 ( \10328 , \10222 );
not \U$10082 ( \10329 , \10276 );
or \U$10083 ( \10330 , \10328 , \10329 );
nand \U$10084 ( \10331 , \10275 , \10264 );
nand \U$10085 ( \10332 , \10330 , \10331 );
not \U$10086 ( \10333 , \10211 );
not \U$10087 ( \10334 , \10204 );
or \U$10088 ( \10335 , \10333 , \10334 );
not \U$10089 ( \10336 , \10194 );
xor \U$10090 ( \10337 , \10189 , \10203 );
nand \U$10091 ( \10338 , \10336 , \10337 );
nand \U$10092 ( \10339 , \10335 , \10338 );
xor \U$10093 ( \10340 , \10332 , \10339 );
not \U$10094 ( \10341 , \10340 );
or \U$10095 ( \10342 , \10327 , \10341 );
or \U$10096 ( \10343 , \10340 , \10326 );
nand \U$10097 ( \10344 , \10342 , \10343 );
nand \U$10098 ( \10345 , \10295 , \10344 );
nand \U$10099 ( \10346 , \10289 , \10345 );
not \U$10100 ( \10347 , \10318 );
not \U$10101 ( \10348 , \10347 );
not \U$10102 ( \10349 , \10309 );
or \U$10103 ( \10350 , \10348 , \10349 );
nand \U$10104 ( \10351 , \10350 , \10320 );
not \U$10105 ( \10352 , \10351 );
not \U$10106 ( \10353 , \10352 );
xor \U$10107 ( \10354 , \8130 , \8315 );
xor \U$10108 ( \10355 , \10354 , \8488 );
not \U$10109 ( \10356 , \10355 );
not \U$10110 ( \10357 , \10301 );
not \U$10111 ( \10358 , \10300 );
not \U$10112 ( \10359 , \10308 );
or \U$10113 ( \10360 , \10358 , \10359 );
or \U$10114 ( \10361 , \10308 , \10300 );
nand \U$10115 ( \10362 , \10360 , \10361 );
not \U$10116 ( \10363 , \10362 );
or \U$10117 ( \10364 , \10357 , \10363 );
not \U$10118 ( \10365 , \10300 );
nand \U$10119 ( \10366 , \10365 , \10308 );
nand \U$10120 ( \10367 , \10364 , \10366 );
not \U$10121 ( \10368 , \10367 );
and \U$10122 ( \10369 , \10356 , \10368 );
and \U$10123 ( \10370 , \10367 , \10355 );
nor \U$10124 ( \10371 , \10369 , \10370 );
not \U$10125 ( \10372 , \10371 );
or \U$10126 ( \10373 , \10353 , \10372 );
or \U$10127 ( \10374 , \10371 , \10352 );
nand \U$10128 ( \10375 , \10373 , \10374 );
not \U$10129 ( \10376 , \10340 );
not \U$10130 ( \10377 , \10326 );
not \U$10131 ( \10378 , \10377 );
or \U$10132 ( \10379 , \10376 , \10378 );
or \U$10133 ( \10380 , \10332 , \10339 );
nand \U$10134 ( \10381 , \10379 , \10380 );
nand \U$10135 ( \10382 , \10375 , \10381 );
not \U$10136 ( \10383 , \10355 );
not \U$10137 ( \10384 , \10367 );
not \U$10138 ( \10385 , \10384 );
or \U$10139 ( \10386 , \10383 , \10385 );
nand \U$10140 ( \10387 , \10386 , \10351 );
not \U$10141 ( \10388 , \10355 );
nand \U$10142 ( \10389 , \10388 , \10367 );
and \U$10143 ( \10390 , \10387 , \10389 );
xor \U$10144 ( \10391 , \8507 , \8491 );
xnor \U$10145 ( \10392 , \10391 , \8499 );
nand \U$10146 ( \10393 , \10390 , \10392 );
nand \U$10147 ( \10394 , \10382 , \10393 );
nor \U$10148 ( \10395 , \10346 , \10394 );
xor \U$10149 ( \10396 , RIbe28570_23, RIbe2a910_99);
not \U$10150 ( \10397 , \10396 );
not \U$10151 ( \10398 , \9737 );
or \U$10152 ( \10399 , \10397 , \10398 );
buf \U$10153 ( \10400 , \9724 );
buf \U$10154 ( \10401 , \10400 );
xor \U$10155 ( \10402 , RIbe2a910_99, RIbe286d8_26);
nand \U$10156 ( \10403 , \10401 , \10402 );
nand \U$10157 ( \10404 , \10399 , \10403 );
xor \U$10158 ( \10405 , RIbe28f48_44, RIbe29470_55);
not \U$10159 ( \10406 , \10405 );
not \U$10160 ( \10407 , \9618 );
or \U$10161 ( \10408 , \10406 , \10407 );
xor \U$10162 ( \10409 , RIbe294e8_56, RIbe28f48_44);
nand \U$10163 ( \10410 , \9524 , \10409 );
nand \U$10164 ( \10411 , \10408 , \10410 );
or \U$10165 ( \10412 , \10404 , \10411 );
xor \U$10166 ( \10413 , RIbe2a118_82, RIbe27d78_6);
not \U$10167 ( \10414 , \10413 );
not \U$10168 ( \10415 , \1164 );
or \U$10169 ( \10416 , \10414 , \10415 );
xor \U$10170 ( \10417 , RIbe2a820_97, RIbe27d78_6);
nand \U$10171 ( \10418 , \314 , \10417 );
nand \U$10172 ( \10419 , \10416 , \10418 );
nand \U$10173 ( \10420 , \10412 , \10419 );
nand \U$10174 ( \10421 , \10404 , \10411 );
nand \U$10175 ( \10422 , \10420 , \10421 );
xor \U$10176 ( \10423 , RIbe27ee0_9, RIbe2a550_91);
not \U$10177 ( \10424 , \10423 );
and \U$10178 ( \10425 , RIbe2a190_83, RIbe2a5c8_92);
not \U$10179 ( \10426 , RIbe2a190_83);
and \U$10180 ( \10427 , \10426 , RIbe2a550_91);
nor \U$10181 ( \10428 , \10425 , \10427 );
nand \U$10182 ( \10429 , RIbe2a550_91, RIbe2a5c8_92);
not \U$10183 ( \10430 , \10429 );
nor \U$10184 ( \10431 , \10428 , \10430 );
buf \U$10185 ( \10432 , \10431 );
buf \U$10186 ( \10433 , \10432 );
buf \U$10187 ( \10434 , \10433 );
not \U$10188 ( \10435 , \10434 );
or \U$10189 ( \10436 , \10424 , \10435 );
xor \U$10190 ( \10437 , RIbe2a190_83, RIbe2a5c8_92);
not \U$10191 ( \10438 , \10437 );
buf \U$10192 ( \10439 , \10438 );
not \U$10193 ( \10440 , \10439 );
xor \U$10194 ( \10441 , RIbe2a550_91, RIbe28048_12);
nand \U$10195 ( \10442 , \10440 , \10441 );
nand \U$10196 ( \10443 , \10436 , \10442 );
xor \U$10197 ( \10444 , RIbe28318_18, RIbe2a2f8_86);
not \U$10198 ( \10445 , \10444 );
not \U$10199 ( \10446 , \8988 );
not \U$10200 ( \10447 , \10446 );
or \U$10201 ( \10448 , \10445 , \10447 );
xor \U$10202 ( \10449 , RIbe2a2f8_86, RIbe284f8_22);
nand \U$10203 ( \10450 , \9379 , \10449 );
nand \U$10204 ( \10451 , \10448 , \10450 );
or \U$10205 ( \10452 , \10443 , \10451 );
xor \U$10206 ( \10453 , RIbe29038_46, RIbe2aa78_102);
not \U$10207 ( \10454 , \10453 );
not \U$10208 ( \10455 , \282 );
or \U$10209 ( \10456 , \10454 , \10455 );
xor \U$10210 ( \10457 , RIbe2b6a8_128, RIbe29038_46);
nand \U$10211 ( \10458 , \287 , \10457 );
nand \U$10212 ( \10459 , \10456 , \10458 );
nand \U$10213 ( \10460 , \10452 , \10459 );
nand \U$10214 ( \10461 , \10443 , \10451 );
nand \U$10215 ( \10462 , \10460 , \10461 );
xor \U$10216 ( \10463 , \10422 , \10462 );
xor \U$10217 ( \10464 , RIbe27fd0_11, RIbe28138_14);
not \U$10218 ( \10465 , \10464 );
not \U$10219 ( \10466 , \2717 );
not \U$10220 ( \10467 , \10466 );
or \U$10221 ( \10468 , \10465 , \10467 );
xor \U$10222 ( \10469 , RIbe27fd0_11, RIbe282a0_17);
nand \U$10223 ( \10470 , \2707 , \10469 );
nand \U$10224 ( \10471 , \10468 , \10470 );
xor \U$10225 ( \10472 , RIbe28750_27, RIbe2a3e8_88);
not \U$10226 ( \10473 , \10472 );
not \U$10227 ( \10474 , \9096 );
or \U$10228 ( \10475 , \10473 , \10474 );
buf \U$10229 ( \10476 , \9089 );
xor \U$10230 ( \10477 , RIbe28840_29, RIbe2a3e8_88);
nand \U$10231 ( \10478 , \10476 , \10477 );
nand \U$10232 ( \10479 , \10475 , \10478 );
xor \U$10233 ( \10480 , \10471 , \10479 );
xor \U$10234 ( \10481 , RIbe28cf0_39, RIbe28930_31);
not \U$10235 ( \10482 , \10481 );
not \U$10236 ( \10483 , \965 );
or \U$10237 ( \10484 , \10482 , \10483 );
xor \U$10238 ( \10485 , RIbe298a8_64, RIbe28930_31);
nand \U$10239 ( \10486 , \1199 , \10485 );
nand \U$10240 ( \10487 , \10484 , \10486 );
and \U$10241 ( \10488 , \10480 , \10487 );
and \U$10242 ( \10489 , \10471 , \10479 );
or \U$10243 ( \10490 , \10488 , \10489 );
buf \U$10244 ( \10491 , \10490 );
xnor \U$10245 ( \10492 , \10463 , \10491 );
xor \U$10246 ( \10493 , RIbe28228_16, RIbe29b78_70);
not \U$10247 ( \10494 , \10493 );
not \U$10248 ( \10495 , \879 );
or \U$10249 ( \10496 , \10494 , \10495 );
xor \U$10250 ( \10497 , RIbe27b20_1, RIbe28228_16);
nand \U$10251 ( \10498 , \885 , \10497 );
nand \U$10252 ( \10499 , \10496 , \10498 );
not \U$10253 ( \10500 , \10499 );
xor \U$10254 ( \10501 , RIbe27c10_3, RIbe2b360_121);
not \U$10255 ( \10502 , \10501 );
not \U$10256 ( \10503 , \7440 );
or \U$10257 ( \10504 , \10502 , \10503 );
xor \U$10258 ( \10505 , RIbe27c10_3, RIbe2a0a0_81);
nand \U$10259 ( \10506 , \1173 , \10505 );
nand \U$10260 ( \10507 , \10504 , \10506 );
not \U$10261 ( \10508 , \10507 );
and \U$10262 ( \10509 , \10500 , \10508 );
not \U$10263 ( \10510 , \10500 );
and \U$10264 ( \10511 , \10510 , \10507 );
nor \U$10265 ( \10512 , \10509 , \10511 );
xor \U$10266 ( \10513 , RIbe29f38_78, RIbe296c8_60);
not \U$10267 ( \10514 , \10513 );
not \U$10268 ( \10515 , \1452 );
or \U$10269 ( \10516 , \10514 , \10515 );
xor \U$10270 ( \10517 , RIbe29ec0_77, RIbe296c8_60);
nand \U$10271 ( \10518 , \908 , \10517 );
nand \U$10272 ( \10519 , \10516 , \10518 );
and \U$10273 ( \10520 , \10512 , \10519 );
not \U$10274 ( \10521 , \10512 );
not \U$10275 ( \10522 , \10519 );
and \U$10276 ( \10523 , \10521 , \10522 );
nor \U$10277 ( \10524 , \10520 , \10523 );
xor \U$10278 ( \10525 , RIbe29218_50, RIbe28390_19);
not \U$10279 ( \10526 , \10525 );
not \U$10280 ( \10527 , \8651 );
or \U$10281 ( \10528 , \10526 , \10527 );
xor \U$10282 ( \10529 , RIbe28390_19, RIbe29a10_67);
nand \U$10283 ( \10530 , \2648 , \10529 );
nand \U$10284 ( \10531 , \10528 , \10530 );
xor \U$10285 ( \10532 , RIbe27b98_2, RIbe2adc0_109);
not \U$10286 ( \10533 , \10532 );
not \U$10287 ( \10534 , \1295 );
or \U$10288 ( \10535 , \10533 , \10534 );
xor \U$10289 ( \10536 , RIbe2a460_89, RIbe27b98_2);
nand \U$10290 ( \10537 , \1734 , \10536 );
nand \U$10291 ( \10538 , \10535 , \10537 );
xor \U$10292 ( \10539 , \10531 , \10538 );
xor \U$10293 ( \10540 , RIbe29d58_74, RIbe280c0_13);
not \U$10294 ( \10541 , \10540 );
not \U$10295 ( \10542 , \859 );
not \U$10296 ( \10543 , \10542 );
or \U$10297 ( \10544 , \10541 , \10543 );
xor \U$10298 ( \10545 , RIbe29ce0_73, RIbe280c0_13);
nand \U$10299 ( \10546 , \869 , \10545 );
nand \U$10300 ( \10547 , \10544 , \10546 );
xor \U$10301 ( \10548 , \10539 , \10547 );
xor \U$10302 ( \10549 , \10524 , \10548 );
xor \U$10303 ( \10550 , RIbe2a028_80, RIbe28c00_37);
not \U$10304 ( \10551 , \10550 );
not \U$10305 ( \10552 , \8401 );
or \U$10306 ( \10553 , \10551 , \10552 );
xor \U$10307 ( \10554 , RIbe2a028_80, RIbe28c78_38);
nand \U$10308 ( \10555 , \9065 , \10554 );
nand \U$10309 ( \10556 , \10553 , \10555 );
xor \U$10310 ( \10557 , RIbe28de0_41, RIbe2a4d8_90);
not \U$10311 ( \10558 , \10557 );
not \U$10312 ( \10559 , \331 );
or \U$10313 ( \10560 , \10558 , \10559 );
xor \U$10314 ( \10561 , RIbe2b2e8_120, RIbe28de0_41);
nand \U$10315 ( \10562 , \347 , \10561 );
nand \U$10316 ( \10563 , \10560 , \10562 );
xor \U$10317 ( \10564 , \10556 , \10563 );
xor \U$10318 ( \10565 , RIbe290b0_47, RIbe2a898_98);
not \U$10319 ( \10566 , \10565 );
not \U$10320 ( \10567 , \384 );
buf \U$10321 ( \10568 , \10567 );
not \U$10322 ( \10569 , \10568 );
or \U$10323 ( \10570 , \10566 , \10569 );
xor \U$10324 ( \10571 , RIbe2aa00_101, RIbe290b0_47);
nand \U$10325 ( \10572 , \398 , \10571 );
nand \U$10326 ( \10573 , \10570 , \10572 );
xor \U$10327 ( \10574 , \10564 , \10573 );
and \U$10328 ( \10575 , \10549 , \10574 );
and \U$10329 ( \10576 , \10524 , \10548 );
or \U$10330 ( \10577 , \10575 , \10576 );
buf \U$10331 ( \10578 , \10577 );
xor \U$10332 ( \10579 , \10492 , \10578 );
not \U$10333 ( \10580 , \10451 );
xor \U$10334 ( \10581 , \10443 , \10580 );
xor \U$10335 ( \10582 , \10581 , \10459 );
xor \U$10336 ( \10583 , RIbe29b00_69, RIbe28480_21);
not \U$10337 ( \10584 , \10583 );
not \U$10338 ( \10585 , \3344 );
or \U$10339 ( \10586 , \10584 , \10585 );
and \U$10340 ( \10587 , RIbe28480_21, RIbe29128_48);
nor \U$10341 ( \10588 , RIbe28480_21, RIbe29128_48);
nor \U$10342 ( \10589 , \10587 , \10588 );
nand \U$10343 ( \10590 , \7483 , \10589 );
nand \U$10344 ( \10591 , \10586 , \10590 );
xor \U$10345 ( \10592 , RIbe285e8_24, RIbe291a0_49);
not \U$10346 ( \10593 , \10592 );
not \U$10347 ( \10594 , \2618 );
or \U$10348 ( \10595 , \10593 , \10594 );
xor \U$10349 ( \10596 , RIbe285e8_24, RIbe295d8_58);
nand \U$10350 ( \10597 , \8270 , \10596 );
nand \U$10351 ( \10598 , \10595 , \10597 );
xor \U$10352 ( \10599 , \10591 , \10598 );
xor \U$10353 ( \10600 , RIbe28a20_33, RIbe29998_66);
not \U$10354 ( \10601 , \10600 );
not \U$10355 ( \10602 , \2276 );
or \U$10356 ( \10603 , \10601 , \10602 );
not \U$10357 ( \10604 , RIbe28d68_40);
not \U$10358 ( \10605 , RIbe28a20_33);
or \U$10359 ( \10606 , \10604 , \10605 );
or \U$10360 ( \10607 , RIbe28a20_33, RIbe28d68_40);
nand \U$10361 ( \10608 , \10606 , \10607 );
not \U$10362 ( \10609 , \10608 );
nand \U$10363 ( \10610 , \10609 , \1769 );
nand \U$10364 ( \10611 , \10603 , \10610 );
xnor \U$10365 ( \10612 , \10599 , \10611 );
nand \U$10366 ( \10613 , \10582 , \10612 );
not \U$10367 ( \10614 , \10613 );
xor \U$10368 ( \10615 , \10404 , \10419 );
xor \U$10369 ( \10616 , \10615 , \10411 );
not \U$10370 ( \10617 , \10616 );
or \U$10371 ( \10618 , \10614 , \10617 );
not \U$10372 ( \10619 , \10582 );
not \U$10373 ( \10620 , \10612 );
nand \U$10374 ( \10621 , \10619 , \10620 );
nand \U$10375 ( \10622 , \10618 , \10621 );
xnor \U$10376 ( \10623 , \10579 , \10622 );
not \U$10377 ( \10624 , \10623 );
nand \U$10378 ( \10625 , RIbe27b98_2, RIbe2b540_125);
not \U$10379 ( \10626 , \10625 );
xor \U$10380 ( \10627 , RIbe28de0_41, RIbe2a460_89);
not \U$10381 ( \10628 , \10627 );
not \U$10382 ( \10629 , \924 );
or \U$10383 ( \10630 , \10628 , \10629 );
nand \U$10384 ( \10631 , \347 , \10557 );
nand \U$10385 ( \10632 , \10630 , \10631 );
not \U$10386 ( \10633 , \10632 );
or \U$10387 ( \10634 , \10626 , \10633 );
or \U$10388 ( \10635 , \10632 , \10625 );
nand \U$10389 ( \10636 , \10634 , \10635 );
xor \U$10390 ( \10637 , RIbe28480_21, RIbe29a10_67);
not \U$10391 ( \10638 , \10637 );
not \U$10392 ( \10639 , \2519 );
or \U$10393 ( \10640 , \10638 , \10639 );
nand \U$10394 ( \10641 , \3075 , \10583 );
nand \U$10395 ( \10642 , \10640 , \10641 );
xor \U$10396 ( \10643 , \10636 , \10642 );
not \U$10397 ( \10644 , \10643 );
xor \U$10398 ( \10645 , RIbe296c8_60, RIbe2aa78_102);
not \U$10399 ( \10646 , \10645 );
not \U$10400 ( \10647 , \8531 );
or \U$10401 ( \10648 , \10646 , \10647 );
xor \U$10402 ( \10649 , RIbe2b6a8_128, RIbe296c8_60);
nand \U$10403 ( \10650 , \8534 , \10649 );
nand \U$10404 ( \10651 , \10648 , \10650 );
not \U$10405 ( \10652 , \10651 );
xor \U$10406 ( \10653 , RIbe29d58_74, RIbe28228_16);
not \U$10407 ( \10654 , \10653 );
not \U$10408 ( \10655 , \879 );
or \U$10409 ( \10656 , \10654 , \10655 );
xor \U$10410 ( \10657 , RIbe28228_16, RIbe29ce0_73);
nand \U$10411 ( \10658 , \885 , \10657 );
nand \U$10412 ( \10659 , \10656 , \10658 );
not \U$10413 ( \10660 , \10659 );
or \U$10414 ( \10661 , \10652 , \10660 );
or \U$10415 ( \10662 , \10659 , \10651 );
xor \U$10416 ( \10663 , RIbe2a4d8_90, RIbe27c10_3);
not \U$10417 ( \10664 , \10663 );
not \U$10418 ( \10665 , \936 );
or \U$10419 ( \10666 , \10664 , \10665 );
xor \U$10420 ( \10667 , RIbe2b2e8_120, RIbe27c10_3);
nand \U$10421 ( \10668 , \369 , \10667 );
nand \U$10422 ( \10669 , \10666 , \10668 );
nand \U$10423 ( \10670 , \10662 , \10669 );
nand \U$10424 ( \10671 , \10661 , \10670 );
xor \U$10425 ( \10672 , RIbe2a028_80, RIbe293f8_54);
not \U$10426 ( \10673 , \10672 );
not \U$10427 ( \10674 , \9528 );
not \U$10428 ( \10675 , \10674 );
or \U$10429 ( \10676 , \10673 , \10675 );
xor \U$10430 ( \10677 , RIbe29308_52, RIbe2a028_80);
nand \U$10431 ( \10678 , \9065 , \10677 );
nand \U$10432 ( \10679 , \10676 , \10678 );
xor \U$10433 ( \10680 , RIbe27ee0_9, RIbe2a190_83);
not \U$10434 ( \10681 , \10680 );
and \U$10435 ( \10682 , RIbe2a280_85, RIbe2a190_83);
not \U$10436 ( \10683 , RIbe2a280_85);
and \U$10437 ( \10684 , \10683 , RIbe2a208_84);
nor \U$10438 ( \10685 , \10682 , \10684 );
nor \U$10439 ( \10686 , RIbe2a190_83, RIbe2a208_84);
not \U$10440 ( \10687 , \10686 );
nand \U$10441 ( \10688 , \10685 , \10687 );
buf \U$10442 ( \10689 , \10688 );
not \U$10443 ( \10690 , \10689 );
not \U$10444 ( \10691 , \10690 );
or \U$10445 ( \10692 , \10681 , \10691 );
xor \U$10446 ( \10693 , RIbe2a208_84, RIbe2a280_85);
not \U$10447 ( \10694 , \10693 );
not \U$10448 ( \10695 , \10694 );
buf \U$10449 ( \10696 , \10695 );
xor \U$10450 ( \10697 , RIbe28048_12, RIbe2a190_83);
nand \U$10451 ( \10698 , \10696 , \10697 );
nand \U$10452 ( \10699 , \10692 , \10698 );
or \U$10453 ( \10700 , \10679 , \10699 );
xor \U$10454 ( \10701 , RIbe2a898_98, RIbe29038_46);
not \U$10455 ( \10702 , \10701 );
not \U$10456 ( \10703 , \282 );
or \U$10457 ( \10704 , \10702 , \10703 );
xor \U$10458 ( \10705 , RIbe29038_46, RIbe2aa00_101);
nand \U$10459 ( \10706 , \287 , \10705 );
nand \U$10460 ( \10707 , \10704 , \10706 );
nand \U$10461 ( \10708 , \10700 , \10707 );
nand \U$10462 ( \10709 , \10679 , \10699 );
nand \U$10463 ( \10710 , \10708 , \10709 );
xor \U$10464 ( \10711 , \10671 , \10710 );
not \U$10465 ( \10712 , \10711 );
or \U$10466 ( \10713 , \10644 , \10712 );
nand \U$10467 ( \10714 , \10710 , \10671 );
nand \U$10468 ( \10715 , \10713 , \10714 );
not \U$10469 ( \10716 , \10715 );
not \U$10470 ( \10717 , \10716 );
xor \U$10471 ( \10718 , RIbe294e8_56, RIbe29c68_72);
not \U$10472 ( \10719 , \10718 );
not \U$10473 ( \10720 , \4576 );
not \U$10474 ( \10721 , \10720 );
or \U$10475 ( \10722 , \10719 , \10721 );
xor \U$10476 ( \10723 , RIbe288b8_30, RIbe29c68_72);
nand \U$10477 ( \10724 , \4580 , \10723 );
nand \U$10478 ( \10725 , \10722 , \10724 );
xor \U$10479 ( \10726 , RIbe290b0_47, RIbe2a820_97);
not \U$10480 ( \10727 , \10726 );
not \U$10481 ( \10728 , \523 );
or \U$10482 ( \10729 , \10727 , \10728 );
not \U$10483 ( \10730 , \468 );
nand \U$10484 ( \10731 , \10730 , \10565 );
nand \U$10485 ( \10732 , \10729 , \10731 );
xor \U$10486 ( \10733 , \10725 , \10732 );
xor \U$10487 ( \10734 , RIbe28b88_36, RIbe28d68_40);
not \U$10488 ( \10735 , \10734 );
not \U$10489 ( \10736 , \2701 );
or \U$10490 ( \10737 , \10735 , \10736 );
xor \U$10491 ( \10738 , RIbe28b88_36, RIbe27c88_4);
nand \U$10492 ( \10739 , \2691 , \10738 );
nand \U$10493 ( \10740 , \10737 , \10739 );
xor \U$10494 ( \10741 , \10733 , \10740 );
not \U$10495 ( \10742 , \4893 );
xor \U$10496 ( \10743 , RIbe27fd0_11, RIbe297b8_62);
not \U$10497 ( \10744 , \10743 );
or \U$10498 ( \10745 , \10742 , \10744 );
nand \U$10499 ( \10746 , \7709 , \10464 );
nand \U$10500 ( \10747 , \10745 , \10746 );
xor \U$10501 ( \10748 , RIbe2a0a0_81, RIbe27d78_6);
not \U$10502 ( \10749 , \10748 );
not \U$10503 ( \10750 , \8898 );
or \U$10504 ( \10751 , \10749 , \10750 );
xor \U$10505 ( \10752 , RIbe290b0_47, RIbe29a88_68);
nand \U$10506 ( \10753 , \10752 , \10413 );
nand \U$10507 ( \10754 , \10751 , \10753 );
not \U$10508 ( \10755 , \10754 );
xor \U$10509 ( \10756 , RIbe2ad48_108, RIbe27b98_2);
not \U$10510 ( \10757 , \10756 );
not \U$10511 ( \10758 , \9833 );
or \U$10512 ( \10759 , \10757 , \10758 );
nand \U$10513 ( \10760 , \267 , \10532 );
nand \U$10514 ( \10761 , \10759 , \10760 );
not \U$10515 ( \10762 , \10761 );
not \U$10516 ( \10763 , \10762 );
or \U$10517 ( \10764 , \10755 , \10763 );
or \U$10518 ( \10765 , \10762 , \10754 );
nand \U$10519 ( \10766 , \10764 , \10765 );
xor \U$10520 ( \10767 , \10747 , \10766 );
buf \U$10521 ( \10768 , \10767 );
or \U$10522 ( \10769 , \10741 , \10768 );
xor \U$10523 ( \10770 , RIbe28930_31, RIbe27b20_1);
not \U$10524 ( \10771 , \10770 );
not \U$10525 ( \10772 , \1793 );
or \U$10526 ( \10773 , \10771 , \10772 );
nand \U$10527 ( \10774 , \970 , \10481 );
nand \U$10528 ( \10775 , \10773 , \10774 );
not \U$10529 ( \10776 , \10667 );
not \U$10530 ( \10777 , \7440 );
or \U$10531 ( \10778 , \10776 , \10777 );
nand \U$10532 ( \10779 , \1173 , \10501 );
nand \U$10533 ( \10780 , \10778 , \10779 );
and \U$10534 ( \10781 , \10775 , \10780 );
not \U$10535 ( \10782 , \10775 );
not \U$10536 ( \10783 , \10780 );
and \U$10537 ( \10784 , \10782 , \10783 );
nor \U$10538 ( \10785 , \10781 , \10784 );
not \U$10539 ( \10786 , RIbe28c78_38);
not \U$10540 ( \10787 , RIbe2a2f8_86);
and \U$10541 ( \10788 , \10786 , \10787 );
and \U$10542 ( \10789 , RIbe28c78_38, RIbe2a2f8_86);
nor \U$10543 ( \10790 , \10788 , \10789 );
not \U$10544 ( \10791 , \10790 );
not \U$10545 ( \10792 , \8696 );
not \U$10546 ( \10793 , \10792 );
or \U$10547 ( \10794 , \10791 , \10793 );
nand \U$10548 ( \10795 , \8706 , \10444 );
nand \U$10549 ( \10796 , \10794 , \10795 );
xor \U$10550 ( \10797 , \10785 , \10796 );
nand \U$10551 ( \10798 , \10769 , \10797 );
nand \U$10552 ( \10799 , \10768 , \10741 );
nand \U$10553 ( \10800 , \10798 , \10799 );
not \U$10554 ( \10801 , \10800 );
or \U$10555 ( \10802 , \10717 , \10801 );
or \U$10556 ( \10803 , \10800 , \10716 );
nand \U$10557 ( \10804 , \10802 , \10803 );
xor \U$10558 ( \10805 , RIbe286d8_26, RIbe2a550_91);
not \U$10559 ( \10806 , \10805 );
not \U$10560 ( \10807 , \10434 );
or \U$10561 ( \10808 , \10806 , \10807 );
nand \U$10562 ( \10809 , \10440 , \10423 );
nand \U$10563 ( \10810 , \10808 , \10809 );
not \U$10564 ( \10811 , \10649 );
not \U$10565 ( \10812 , \899 );
not \U$10566 ( \10813 , \10812 );
or \U$10567 ( \10814 , \10811 , \10813 );
nand \U$10568 ( \10815 , \8534 , \10513 );
nand \U$10569 ( \10816 , \10814 , \10815 );
not \U$10570 ( \10817 , \10705 );
not \U$10571 ( \10818 , \281 );
or \U$10572 ( \10819 , \10817 , \10818 );
nand \U$10573 ( \10820 , \1583 , \10453 );
nand \U$10574 ( \10821 , \10819 , \10820 );
and \U$10575 ( \10822 , \10816 , \10821 );
not \U$10576 ( \10823 , \10816 );
not \U$10577 ( \10824 , \10821 );
and \U$10578 ( \10825 , \10823 , \10824 );
nor \U$10579 ( \10826 , \10822 , \10825 );
xor \U$10580 ( \10827 , \10810 , \10826 );
not \U$10581 ( \10828 , \10827 );
not \U$10582 ( \10829 , \10697 );
nand \U$10583 ( \10830 , \10685 , \10687 );
not \U$10584 ( \10831 , \10830 );
not \U$10585 ( \10832 , \10831 );
or \U$10586 ( \10833 , \10829 , \10832 );
not \U$10587 ( \10834 , \10694 );
xor \U$10588 ( \10835 , RIbe29380_53, RIbe2a190_83);
nand \U$10589 ( \10836 , \10834 , \10835 );
nand \U$10590 ( \10837 , \10833 , \10836 );
and \U$10591 ( \10838 , RIbe2b108_116, RIbe2b090_115);
not \U$10592 ( \10839 , RIbe2b108_116);
and \U$10593 ( \10840 , \10839 , RIbe2a280_85);
nor \U$10594 ( \10841 , \10838 , \10840 );
not \U$10595 ( \10842 , \10841 );
nand \U$10596 ( \10843 , RIbe2a280_85, RIbe2b090_115);
nand \U$10597 ( \10844 , \10842 , \10843 );
not \U$10598 ( \10845 , \10844 );
buf \U$10599 ( \10846 , \10845 );
xor \U$10600 ( \10847 , RIbe2b090_115, RIbe2b108_116);
not \U$10601 ( \10848 , \10847 );
not \U$10602 ( \10849 , \10848 );
or \U$10603 ( \10850 , \10846 , \10849 );
nand \U$10604 ( \10851 , \10850 , RIbe2a280_85);
xor \U$10605 ( \10852 , \10837 , \10851 );
not \U$10606 ( \10853 , \10657 );
not \U$10607 ( \10854 , \879 );
or \U$10608 ( \10855 , \10853 , \10854 );
nand \U$10609 ( \10856 , \885 , \10493 );
nand \U$10610 ( \10857 , \10855 , \10856 );
xor \U$10611 ( \10858 , \10852 , \10857 );
not \U$10612 ( \10859 , \10858 );
xor \U$10613 ( \10860 , RIbe285e8_24, RIbe29128_48);
not \U$10614 ( \10861 , \10860 );
nand \U$10615 ( \10862 , \2613 , \2615 );
not \U$10616 ( \10863 , \10862 );
not \U$10617 ( \10864 , \10863 );
or \U$10618 ( \10865 , \10861 , \10864 );
nand \U$10619 ( \10866 , \2758 , \10592 );
nand \U$10620 ( \10867 , \10865 , \10866 );
xor \U$10621 ( \10868 , RIbe284f8_22, RIbe2a3e8_88);
not \U$10622 ( \10869 , \10868 );
not \U$10623 ( \10870 , \9262 );
or \U$10624 ( \10871 , \10869 , \10870 );
nand \U$10625 ( \10872 , \8793 , \10472 );
nand \U$10626 ( \10873 , \10871 , \10872 );
xor \U$10627 ( \10874 , \10867 , \10873 );
xor \U$10628 ( \10875 , RIbe29ec0_77, RIbe280c0_13);
not \U$10629 ( \10876 , \10875 );
not \U$10630 ( \10877 , \8551 );
or \U$10631 ( \10878 , \10876 , \10877 );
nand \U$10632 ( \10879 , \2369 , \10540 );
nand \U$10633 ( \10880 , \10878 , \10879 );
not \U$10634 ( \10881 , \10880 );
and \U$10635 ( \10882 , \10874 , \10881 );
not \U$10636 ( \10883 , \10874 );
and \U$10637 ( \10884 , \10883 , \10880 );
nor \U$10638 ( \10885 , \10882 , \10884 );
not \U$10639 ( \10886 , \10885 );
and \U$10640 ( \10887 , \10859 , \10886 );
and \U$10641 ( \10888 , \10858 , \10885 );
nor \U$10642 ( \10889 , \10887 , \10888 );
not \U$10643 ( \10890 , \10889 );
not \U$10644 ( \10891 , \10890 );
or \U$10645 ( \10892 , \10828 , \10891 );
not \U$10646 ( \10893 , \10885 );
nand \U$10647 ( \10894 , \10893 , \10858 );
nand \U$10648 ( \10895 , \10892 , \10894 );
nand \U$10649 ( \10896 , \10804 , \10895 );
nand \U$10650 ( \10897 , \10800 , \10715 );
nand \U$10651 ( \10898 , \10896 , \10897 );
not \U$10652 ( \10899 , \10747 );
not \U$10653 ( \10900 , \10766 );
or \U$10654 ( \10901 , \10899 , \10900 );
nand \U$10655 ( \10902 , \10761 , \10754 );
nand \U$10656 ( \10903 , \10901 , \10902 );
not \U$10657 ( \10904 , \10642 );
not \U$10658 ( \10905 , \10636 );
or \U$10659 ( \10906 , \10904 , \10905 );
not \U$10660 ( \10907 , \10625 );
nand \U$10661 ( \10908 , \10907 , \10632 );
nand \U$10662 ( \10909 , \10906 , \10908 );
xor \U$10663 ( \10910 , \10903 , \10909 );
not \U$10664 ( \10911 , \10796 );
not \U$10665 ( \10912 , \10785 );
or \U$10666 ( \10913 , \10911 , \10912 );
nand \U$10667 ( \10914 , \10775 , \10780 );
nand \U$10668 ( \10915 , \10913 , \10914 );
xnor \U$10669 ( \10916 , \10910 , \10915 );
xor \U$10670 ( \10917 , \10837 , \10851 );
and \U$10671 ( \10918 , \10917 , \10857 );
and \U$10672 ( \10919 , \10837 , \10851 );
or \U$10673 ( \10920 , \10918 , \10919 );
not \U$10674 ( \10921 , \10920 );
xor \U$10675 ( \10922 , \10725 , \10732 );
and \U$10676 ( \10923 , \10922 , \10740 );
and \U$10677 ( \10924 , \10725 , \10732 );
or \U$10678 ( \10925 , \10923 , \10924 );
not \U$10679 ( \10926 , \10925 );
not \U$10680 ( \10927 , \10926 );
or \U$10681 ( \10928 , \10921 , \10927 );
not \U$10682 ( \10929 , \10920 );
nand \U$10683 ( \10930 , \10929 , \10925 );
nand \U$10684 ( \10931 , \10928 , \10930 );
not \U$10685 ( \10932 , RIbe28a98_34);
not \U$10686 ( \10933 , RIbe29e48_76);
and \U$10687 ( \10934 , \10932 , \10933 );
and \U$10688 ( \10935 , RIbe28a98_34, RIbe29e48_76);
nor \U$10689 ( \10936 , \10934 , \10935 );
not \U$10690 ( \10937 , \10936 );
not \U$10691 ( \10938 , \7371 );
not \U$10692 ( \10939 , \10938 );
or \U$10693 ( \10940 , \10937 , \10939 );
xor \U$10694 ( \10941 , RIbe29e48_76, RIbe293f8_54);
nand \U$10695 ( \10942 , \8245 , \10941 );
nand \U$10696 ( \10943 , \10940 , \10942 );
not \U$10697 ( \10944 , \10943 );
xor \U$10698 ( \10945 , RIbe27e68_8, RIbe295d8_58);
not \U$10699 ( \10946 , \10945 );
not \U$10700 ( \10947 , \2600 );
or \U$10701 ( \10948 , \10946 , \10947 );
xor \U$10702 ( \10949 , RIbe29740_61, RIbe27e68_8);
nand \U$10703 ( \10950 , \2603 , \10949 );
nand \U$10704 ( \10951 , \10948 , \10950 );
xor \U$10705 ( \10952 , RIbe27df0_7, RIbe28390_19);
not \U$10706 ( \10953 , \10952 );
not \U$10707 ( \10954 , \2640 );
or \U$10708 ( \10955 , \10953 , \10954 );
nand \U$10709 ( \10956 , \2777 , \10525 );
nand \U$10710 ( \10957 , \10955 , \10956 );
xor \U$10711 ( \10958 , \10951 , \10957 );
not \U$10712 ( \10959 , \10958 );
or \U$10713 ( \10960 , \10944 , \10959 );
nand \U$10714 ( \10961 , \10951 , \10957 );
nand \U$10715 ( \10962 , \10960 , \10961 );
not \U$10716 ( \10963 , \10962 );
and \U$10717 ( \10964 , \10931 , \10963 );
not \U$10718 ( \10965 , \10931 );
and \U$10719 ( \10966 , \10965 , \10962 );
nor \U$10720 ( \10967 , \10964 , \10966 );
or \U$10721 ( \10968 , \10916 , \10967 );
not \U$10722 ( \10969 , \10967 );
not \U$10723 ( \10970 , \10916 );
or \U$10724 ( \10971 , \10969 , \10970 );
not \U$10725 ( \10972 , \10880 );
not \U$10726 ( \10973 , \10874 );
or \U$10727 ( \10974 , \10972 , \10973 );
nand \U$10728 ( \10975 , \10873 , \10867 );
nand \U$10729 ( \10976 , \10974 , \10975 );
not \U$10730 ( \10977 , \10976 );
xor \U$10731 ( \10978 , RIbe28a20_33, RIbe298a8_64);
not \U$10732 ( \10979 , \10978 );
not \U$10733 ( \10980 , \1780 );
or \U$10734 ( \10981 , \10979 , \10980 );
nand \U$10735 ( \10982 , \2475 , \10600 );
nand \U$10736 ( \10983 , \10981 , \10982 );
not \U$10737 ( \10984 , \10983 );
xor \U$10738 ( \10985 , RIbe28840_29, RIbe2a910_99);
not \U$10739 ( \10986 , \10985 );
buf \U$10740 ( \10987 , \9736 );
not \U$10741 ( \10988 , \10987 );
or \U$10742 ( \10989 , \10986 , \10988 );
nand \U$10743 ( \10990 , \9726 , \10396 );
nand \U$10744 ( \10991 , \10989 , \10990 );
not \U$10745 ( \10992 , \10991 );
or \U$10746 ( \10993 , \10984 , \10992 );
or \U$10747 ( \10994 , \10991 , \10983 );
xor \U$10748 ( \10995 , RIbe28f48_44, RIbe282a0_17);
not \U$10749 ( \10996 , \10995 );
not \U$10750 ( \10997 , \7609 );
or \U$10751 ( \10998 , \10996 , \10997 );
nand \U$10752 ( \10999 , \9524 , \10405 );
nand \U$10753 ( \11000 , \10998 , \10999 );
nand \U$10754 ( \11001 , \10994 , \11000 );
nand \U$10755 ( \11002 , \10993 , \11001 );
not \U$10756 ( \11003 , \11002 );
not \U$10757 ( \11004 , \11003 );
and \U$10758 ( \11005 , \10977 , \11004 );
and \U$10759 ( \11006 , \10976 , \11003 );
nor \U$10760 ( \11007 , \11005 , \11006 );
not \U$10761 ( \11008 , \10810 );
not \U$10762 ( \11009 , \10826 );
or \U$10763 ( \11010 , \11008 , \11009 );
nand \U$10764 ( \11011 , \10821 , \10816 );
nand \U$10765 ( \11012 , \11010 , \11011 );
and \U$10766 ( \11013 , \11007 , \11012 );
not \U$10767 ( \11014 , \11007 );
not \U$10768 ( \11015 , \11012 );
and \U$10769 ( \11016 , \11014 , \11015 );
nor \U$10770 ( \11017 , \11013 , \11016 );
not \U$10771 ( \11018 , \11017 );
nand \U$10772 ( \11019 , \10971 , \11018 );
nand \U$10773 ( \11020 , \10968 , \11019 );
xor \U$10774 ( \11021 , \10898 , \11020 );
not \U$10775 ( \11022 , \11021 );
or \U$10776 ( \11023 , \10624 , \11022 );
not \U$10777 ( \11024 , \10897 );
not \U$10778 ( \11025 , \10896 );
or \U$10779 ( \11026 , \11024 , \11025 );
nand \U$10780 ( \11027 , \11026 , \11020 );
nand \U$10781 ( \11028 , \11023 , \11027 );
not \U$10782 ( \11029 , \11028 );
not \U$10783 ( \11030 , \10577 );
nand \U$10784 ( \11031 , \11030 , \10492 );
not \U$10785 ( \11032 , \11031 );
not \U$10786 ( \11033 , \10622 );
or \U$10787 ( \11034 , \11032 , \11033 );
not \U$10788 ( \11035 , \10492 );
nand \U$10789 ( \11036 , \11035 , \10577 );
nand \U$10790 ( \11037 , \11034 , \11036 );
not \U$10791 ( \11038 , \11037 );
not \U$10792 ( \11039 , \4841 );
buf \U$10793 ( \11040 , \11039 );
and \U$10794 ( \11041 , \11040 , \10941 );
xor \U$10795 ( \11042 , RIbe29e48_76, RIbe29308_52);
and \U$10796 ( \11043 , \7368 , \11042 );
nor \U$10797 ( \11044 , \11041 , \11043 );
not \U$10798 ( \11045 , \11044 );
not \U$10799 ( \11046 , \11045 );
and \U$10800 ( \11047 , RIbe2ad48_108, RIbe27b98_2);
not \U$10801 ( \11048 , \11047 );
not \U$10802 ( \11049 , \10738 );
not \U$10803 ( \11050 , \9052 );
or \U$10804 ( \11051 , \11049 , \11050 );
xor \U$10805 ( \11052 , RIbe28b88_36, RIbe27df0_7);
nand \U$10806 ( \11053 , \7549 , \11052 );
nand \U$10807 ( \11054 , \11051 , \11053 );
not \U$10808 ( \11055 , \11054 );
or \U$10809 ( \11056 , \11048 , \11055 );
or \U$10810 ( \11057 , \11054 , \11047 );
nand \U$10811 ( \11058 , \11056 , \11057 );
not \U$10812 ( \11059 , \11058 );
or \U$10813 ( \11060 , \11046 , \11059 );
not \U$10814 ( \11061 , \11054 );
nand \U$10815 ( \11062 , \11061 , \11047 );
nand \U$10816 ( \11063 , \11060 , \11062 );
not \U$10817 ( \11064 , \11063 );
not \U$10818 ( \11065 , \11002 );
not \U$10819 ( \11066 , \10976 );
or \U$10820 ( \11067 , \11065 , \11066 );
or \U$10821 ( \11068 , \10976 , \11002 );
nand \U$10822 ( \11069 , \11068 , \11012 );
nand \U$10823 ( \11070 , \11067 , \11069 );
not \U$10824 ( \11071 , \11070 );
or \U$10825 ( \11072 , \11064 , \11071 );
not \U$10826 ( \11073 , \10962 );
not \U$10827 ( \11074 , \10931 );
or \U$10828 ( \11075 , \11073 , \11074 );
nand \U$10829 ( \11076 , \10925 , \10920 );
nand \U$10830 ( \11077 , \11075 , \11076 );
not \U$10831 ( \11078 , \11070 );
not \U$10832 ( \11079 , \11063 );
nand \U$10833 ( \11080 , \11078 , \11079 );
nand \U$10834 ( \11081 , \11077 , \11080 );
nand \U$10835 ( \11082 , \11072 , \11081 );
xor \U$10836 ( \11083 , RIbe2a028_80, RIbe28318_18);
not \U$10837 ( \11084 , \11083 );
not \U$10838 ( \11085 , \8400 );
or \U$10839 ( \11086 , \11084 , \11085 );
xor \U$10840 ( \11087 , RIbe2a028_80, RIbe284f8_22);
nand \U$10841 ( \11088 , \8930 , \11087 );
nand \U$10842 ( \11089 , \11086 , \11088 );
xor \U$10843 ( \11090 , RIbe28750_27, RIbe2a2f8_86);
not \U$10844 ( \11091 , \11090 );
not \U$10845 ( \11092 , \10792 );
or \U$10846 ( \11093 , \11091 , \11092 );
buf \U$10847 ( \11094 , \8705 );
xor \U$10848 ( \11095 , RIbe28840_29, RIbe2a2f8_86);
nand \U$10849 ( \11096 , \11094 , \11095 );
nand \U$10850 ( \11097 , \11093 , \11096 );
xor \U$10851 ( \11098 , \11089 , \11097 );
xor \U$10852 ( \11099 , RIbe29f38_78, RIbe29038_46);
not \U$10853 ( \11100 , \11099 );
not \U$10854 ( \11101 , \281 );
or \U$10855 ( \11102 , \11100 , \11101 );
xor \U$10856 ( \11103 , RIbe29038_46, RIbe29ec0_77);
nand \U$10857 ( \11104 , \1583 , \11103 );
nand \U$10858 ( \11105 , \11102 , \11104 );
xor \U$10859 ( \11106 , \11098 , \11105 );
and \U$10860 ( \11107 , RIbe29e48_76, RIbe28c00_37);
not \U$10861 ( \11108 , RIbe29e48_76);
and \U$10862 ( \11109 , \11108 , \2479 );
nor \U$10863 ( \11110 , \11107 , \11109 );
not \U$10864 ( \11111 , \11110 );
not \U$10865 ( \11112 , \4842 );
or \U$10866 ( \11113 , \11111 , \11112 );
xor \U$10867 ( \11114 , RIbe28c78_38, RIbe29e48_76);
nand \U$10868 ( \11115 , \8245 , \11114 );
nand \U$10869 ( \11116 , \11113 , \11115 );
xor \U$10870 ( \11117 , RIbe29b78_70, RIbe280c0_13);
not \U$10871 ( \11118 , \11117 );
not \U$10872 ( \11119 , \10542 );
or \U$10873 ( \11120 , \11118 , \11119 );
xor \U$10874 ( \11121 , RIbe27b20_1, RIbe280c0_13);
nand \U$10875 ( \11122 , \869 , \11121 );
nand \U$10876 ( \11123 , \11120 , \11122 );
xor \U$10877 ( \11124 , RIbe2a4d8_90, RIbe27b98_2);
not \U$10878 ( \11125 , \11124 );
not \U$10879 ( \11126 , \1295 );
or \U$10880 ( \11127 , \11125 , \11126 );
xor \U$10881 ( \11128 , RIbe2b2e8_120, RIbe27b98_2);
nand \U$10882 ( \11129 , \267 , \11128 );
nand \U$10883 ( \11130 , \11127 , \11129 );
and \U$10884 ( \11131 , \11123 , \11130 );
not \U$10885 ( \11132 , \11123 );
not \U$10886 ( \11133 , \11130 );
and \U$10887 ( \11134 , \11132 , \11133 );
nor \U$10888 ( \11135 , \11131 , \11134 );
xor \U$10889 ( \11136 , \11116 , \11135 );
xor \U$10890 ( \11137 , \11106 , \11136 );
xor \U$10891 ( \11138 , RIbe28f48_44, RIbe288b8_30);
not \U$10892 ( \11139 , \11138 );
not \U$10893 ( \11140 , \7609 );
or \U$10894 ( \11141 , \11139 , \11140 );
xor \U$10895 ( \11142 , RIbe28f48_44, RIbe28a98_34);
nand \U$10896 ( \11143 , \4180 , \11142 );
nand \U$10897 ( \11144 , \11141 , \11143 );
xor \U$10898 ( \11145 , RIbe28390_19, RIbe29b00_69);
not \U$10899 ( \11146 , \11145 );
not \U$10900 ( \11147 , \8651 );
or \U$10901 ( \11148 , \11146 , \11147 );
xor \U$10902 ( \11149 , RIbe28390_19, RIbe29128_48);
nand \U$10903 ( \11150 , \2777 , \11149 );
nand \U$10904 ( \11151 , \11148 , \11150 );
xor \U$10905 ( \11152 , \11144 , \11151 );
xor \U$10906 ( \11153 , RIbe2a898_98, RIbe27d78_6);
not \U$10907 ( \11154 , \11153 );
not \U$10908 ( \11155 , \1086 );
or \U$10909 ( \11156 , \11154 , \11155 );
xnor \U$10910 ( \11157 , RIbe27d78_6, RIbe2aa00_101);
not \U$10911 ( \11158 , \11157 );
nand \U$10912 ( \11159 , \11158 , \315 );
nand \U$10913 ( \11160 , \11156 , \11159 );
xnor \U$10914 ( \11161 , \11152 , \11160 );
xnor \U$10915 ( \11162 , \11137 , \11161 );
not \U$10916 ( \11163 , \11162 );
and \U$10917 ( \11164 , \11082 , \11163 );
not \U$10918 ( \11165 , \11082 );
and \U$10919 ( \11166 , \11165 , \11162 );
nor \U$10920 ( \11167 , \11164 , \11166 );
not \U$10921 ( \11168 , \11167 );
or \U$10922 ( \11169 , \11038 , \11168 );
or \U$10923 ( \11170 , \11167 , \11037 );
nand \U$10924 ( \11171 , \11169 , \11170 );
xor \U$10925 ( \11172 , RIbe285e8_24, RIbe29b00_69);
not \U$10926 ( \11173 , \11172 );
not \U$10927 ( \11174 , \2617 );
not \U$10928 ( \11175 , \11174 );
or \U$10929 ( \11176 , \11173 , \11175 );
nand \U$10930 ( \11177 , \8270 , \10860 );
nand \U$10931 ( \11178 , \11176 , \11177 );
not \U$10932 ( \11179 , \11178 );
xor \U$10933 ( \11180 , RIbe27b98_2, RIbe2b540_125);
not \U$10934 ( \11181 , \11180 );
not \U$10935 ( \11182 , \8380 );
or \U$10936 ( \11183 , \11181 , \11182 );
nand \U$10937 ( \11184 , \7585 , \10756 );
nand \U$10938 ( \11185 , \11183 , \11184 );
not \U$10939 ( \11186 , \11185 );
or \U$10940 ( \11187 , \11179 , \11186 );
or \U$10941 ( \11188 , \11185 , \11178 );
xor \U$10942 ( \11189 , RIbe29f38_78, RIbe280c0_13);
not \U$10943 ( \11190 , \11189 );
not \U$10944 ( \11191 , \8551 );
or \U$10945 ( \11192 , \11190 , \11191 );
nand \U$10946 ( \11193 , \1265 , \10875 );
nand \U$10947 ( \11194 , \11192 , \11193 );
nand \U$10948 ( \11195 , \11188 , \11194 );
nand \U$10949 ( \11196 , \11187 , \11195 );
xor \U$10950 ( \11197 , RIbe28f48_44, RIbe28138_14);
not \U$10951 ( \11198 , \11197 );
not \U$10952 ( \11199 , \8221 );
or \U$10953 ( \11200 , \11198 , \11199 );
buf \U$10954 ( \11201 , \3248 );
nand \U$10955 ( \11202 , \11201 , \10995 );
nand \U$10956 ( \11203 , \11200 , \11202 );
not \U$10957 ( \11204 , \11203 );
xor \U$10958 ( \11205 , RIbe2a910_99, RIbe28750_27);
not \U$10959 ( \11206 , \11205 );
not \U$10960 ( \11207 , \10987 );
or \U$10961 ( \11208 , \11206 , \11207 );
nand \U$10962 ( \11209 , \10401 , \10985 );
nand \U$10963 ( \11210 , \11208 , \11209 );
not \U$10964 ( \11211 , \11210 );
or \U$10965 ( \11212 , \11204 , \11211 );
or \U$10966 ( \11213 , \11210 , \11203 );
xor \U$10967 ( \11214 , RIbe2b360_121, RIbe27d78_6);
not \U$10968 ( \11215 , \11214 );
not \U$10969 ( \11216 , \1613 );
or \U$10970 ( \11217 , \11215 , \11216 );
nand \U$10971 ( \11218 , \314 , \10748 );
nand \U$10972 ( \11219 , \11217 , \11218 );
nand \U$10973 ( \11220 , \11213 , \11219 );
nand \U$10974 ( \11221 , \11212 , \11220 );
xor \U$10975 ( \11222 , \11196 , \11221 );
xor \U$10976 ( \11223 , RIbe2a550_91, RIbe28570_23);
not \U$10977 ( \11224 , \11223 );
not \U$10978 ( \11225 , \10434 );
or \U$10979 ( \11226 , \11224 , \11225 );
not \U$10980 ( \11227 , \10439 );
buf \U$10981 ( \11228 , \11227 );
nand \U$10982 ( \11229 , \11228 , \10805 );
nand \U$10983 ( \11230 , \11226 , \11229 );
not \U$10984 ( \11231 , \11230 );
xor \U$10985 ( \11232 , RIbe29c68_72, RIbe29470_55);
not \U$10986 ( \11233 , \11232 );
not \U$10987 ( \11234 , \8594 );
or \U$10988 ( \11235 , \11233 , \11234 );
nand \U$10989 ( \11236 , \4580 , \10718 );
nand \U$10990 ( \11237 , \11235 , \11236 );
not \U$10991 ( \11238 , \11237 );
xor \U$10992 ( \11239 , RIbe28cf0_39, RIbe28a20_33);
not \U$10993 ( \11240 , \11239 );
not \U$10994 ( \11241 , \1780 );
or \U$10995 ( \11242 , \11240 , \11241 );
nand \U$10996 ( \11243 , \1769 , \10978 );
nand \U$10997 ( \11244 , \11242 , \11243 );
not \U$10998 ( \11245 , \11244 );
not \U$10999 ( \11246 , \11245 );
or \U$11000 ( \11247 , \11238 , \11246 );
or \U$11001 ( \11248 , \11237 , \11245 );
nand \U$11002 ( \11249 , \11247 , \11248 );
not \U$11003 ( \11250 , \11249 );
or \U$11004 ( \11251 , \11231 , \11250 );
not \U$11005 ( \11252 , \11245 );
nand \U$11006 ( \11253 , \11252 , \11237 );
nand \U$11007 ( \11254 , \11251 , \11253 );
and \U$11008 ( \11255 , \11222 , \11254 );
and \U$11009 ( \11256 , \11196 , \11221 );
or \U$11010 ( \11257 , \11255 , \11256 );
not \U$11011 ( \11258 , \11257 );
xor \U$11012 ( \11259 , RIbe28480_21, RIbe29218_50);
not \U$11013 ( \11260 , \11259 );
not \U$11014 ( \11261 , \2518 );
or \U$11015 ( \11262 , \11260 , \11261 );
not \U$11016 ( \11263 , \2526 );
nand \U$11017 ( \11264 , \11263 , \10637 );
nand \U$11018 ( \11265 , \11262 , \11264 );
not \U$11019 ( \11266 , \11265 );
xor \U$11020 ( \11267 , RIbe28b88_36, RIbe29998_66);
not \U$11021 ( \11268 , \11267 );
not \U$11022 ( \11269 , \3401 );
or \U$11023 ( \11270 , \11268 , \11269 );
nand \U$11024 ( \11271 , \2559 , \10734 );
nand \U$11025 ( \11272 , \11270 , \11271 );
not \U$11026 ( \11273 , \11272 );
or \U$11027 ( \11274 , \11266 , \11273 );
or \U$11028 ( \11275 , \11272 , \11265 );
xor \U$11029 ( \11276 , RIbe27c88_4, RIbe28390_19);
not \U$11030 ( \11277 , \11276 );
not \U$11031 ( \11278 , \3408 );
or \U$11032 ( \11279 , \11277 , \11278 );
nand \U$11033 ( \11280 , \2777 , \10952 );
nand \U$11034 ( \11281 , \11279 , \11280 );
nand \U$11035 ( \11282 , \11275 , \11281 );
nand \U$11036 ( \11283 , \11274 , \11282 );
not \U$11037 ( \11284 , \11283 );
nand \U$11038 ( \11285 , RIbe27b98_2, RIbe2b4c8_124);
not \U$11039 ( \11286 , \11285 );
xor \U$11040 ( \11287 , RIbe27e68_8, RIbe291a0_49);
not \U$11041 ( \11288 , \11287 );
not \U$11042 ( \11289 , \2457 );
or \U$11043 ( \11290 , \11288 , \11289 );
nand \U$11044 ( \11291 , \2463 , \10945 );
nand \U$11045 ( \11292 , \11290 , \11291 );
not \U$11046 ( \11293 , \11292 );
or \U$11047 ( \11294 , \11286 , \11293 );
or \U$11048 ( \11295 , \11292 , \11285 );
nand \U$11049 ( \11296 , \11294 , \11295 );
not \U$11050 ( \11297 , \11296 );
xor \U$11051 ( \11298 , RIbe29e48_76, RIbe288b8_30);
not \U$11052 ( \11299 , \11298 );
not \U$11053 ( \11300 , \10938 );
or \U$11054 ( \11301 , \11299 , \11300 );
nand \U$11055 ( \11302 , \4851 , \10936 );
nand \U$11056 ( \11303 , \11301 , \11302 );
not \U$11057 ( \11304 , \11303 );
or \U$11058 ( \11305 , \11297 , \11304 );
not \U$11059 ( \11306 , \11285 );
nand \U$11060 ( \11307 , \11306 , \11292 );
nand \U$11061 ( \11308 , \11305 , \11307 );
not \U$11062 ( \11309 , \11308 );
or \U$11063 ( \11310 , \11284 , \11309 );
or \U$11064 ( \11311 , \11308 , \11283 );
xor \U$11065 ( \11312 , RIbe2a2f8_86, RIbe28c00_37);
not \U$11066 ( \11313 , \11312 );
not \U$11067 ( \11314 , \9375 );
or \U$11068 ( \11315 , \11313 , \11314 );
nand \U$11069 ( \11316 , \8706 , \10790 );
nand \U$11070 ( \11317 , \11315 , \11316 );
not \U$11071 ( \11318 , \11317 );
xor \U$11072 ( \11319 , RIbe28de0_41, RIbe2adc0_109);
not \U$11073 ( \11320 , \11319 );
nor \U$11074 ( \11321 , \327 , \329 );
not \U$11075 ( \11322 , \11321 );
or \U$11076 ( \11323 , \11320 , \11322 );
nand \U$11077 ( \11324 , \7472 , \10627 );
nand \U$11078 ( \11325 , \11323 , \11324 );
xor \U$11079 ( \11326 , RIbe290b0_47, RIbe2a118_82);
not \U$11080 ( \11327 , \11326 );
not \U$11081 ( \11328 , \10567 );
or \U$11082 ( \11329 , \11327 , \11328 );
nand \U$11083 ( \11330 , \398 , \10726 );
nand \U$11084 ( \11331 , \11329 , \11330 );
xor \U$11085 ( \11332 , \11325 , \11331 );
not \U$11086 ( \11333 , \11332 );
or \U$11087 ( \11334 , \11318 , \11333 );
nand \U$11088 ( \11335 , \11331 , \11325 );
nand \U$11089 ( \11336 , \11334 , \11335 );
nand \U$11090 ( \11337 , \11311 , \11336 );
nand \U$11091 ( \11338 , \11310 , \11337 );
not \U$11092 ( \11339 , \11338 );
xor \U$11093 ( \11340 , RIbe2a280_85, RIbe29380_53);
not \U$11094 ( \11341 , \11340 );
not \U$11095 ( \11342 , \10841 );
nand \U$11096 ( \11343 , \11342 , \10843 );
buf \U$11097 ( \11344 , \11343 );
not \U$11098 ( \11345 , \11344 );
not \U$11099 ( \11346 , \11345 );
or \U$11100 ( \11347 , \11341 , \11346 );
buf \U$11101 ( \11348 , \10847 );
nand \U$11102 ( \11349 , \11348 , RIbe2a280_85);
nand \U$11103 ( \11350 , \11347 , \11349 );
not \U$11104 ( \11351 , \10677 );
not \U$11105 ( \11352 , \8401 );
or \U$11106 ( \11353 , \11351 , \11352 );
nand \U$11107 ( \11354 , \8172 , \10550 );
nand \U$11108 ( \11355 , \11353 , \11354 );
or \U$11109 ( \11356 , \11350 , \11355 );
not \U$11110 ( \11357 , \11356 );
xor \U$11111 ( \11358 , RIbe28318_18, RIbe2a3e8_88);
not \U$11112 ( \11359 , \11358 );
not \U$11113 ( \11360 , \9263 );
or \U$11114 ( \11361 , \11359 , \11360 );
nand \U$11115 ( \11362 , \8794 , \10868 );
nand \U$11116 ( \11363 , \11361 , \11362 );
xor \U$11117 ( \11364 , RIbe27fd0_11, RIbe29740_61);
not \U$11118 ( \11365 , \11364 );
not \U$11119 ( \11366 , \2717 );
not \U$11120 ( \11367 , \11366 );
or \U$11121 ( \11368 , \11365 , \11367 );
nand \U$11122 ( \11369 , \2707 , \10743 );
nand \U$11123 ( \11370 , \11368 , \11369 );
or \U$11124 ( \11371 , \11363 , \11370 );
xor \U$11125 ( \11372 , RIbe29b78_70, RIbe28930_31);
not \U$11126 ( \11373 , \11372 );
not \U$11127 ( \11374 , \9104 );
not \U$11128 ( \11375 , \11374 );
or \U$11129 ( \11376 , \11373 , \11375 );
nand \U$11130 ( \11377 , \1199 , \10770 );
nand \U$11131 ( \11378 , \11376 , \11377 );
nand \U$11132 ( \11379 , \11371 , \11378 );
nand \U$11133 ( \11380 , \11363 , \11370 );
nand \U$11134 ( \11381 , \11379 , \11380 );
not \U$11135 ( \11382 , \11381 );
or \U$11136 ( \11383 , \11357 , \11382 );
nand \U$11137 ( \11384 , \11355 , \11350 );
nand \U$11138 ( \11385 , \11383 , \11384 );
not \U$11139 ( \11386 , \11385 );
not \U$11140 ( \11387 , \11386 );
or \U$11141 ( \11388 , \11339 , \11387 );
or \U$11142 ( \11389 , \11338 , \11386 );
nand \U$11143 ( \11390 , \11388 , \11389 );
not \U$11144 ( \11391 , \11390 );
or \U$11145 ( \11392 , \11258 , \11391 );
nand \U$11146 ( \11393 , \11338 , \11385 );
nand \U$11147 ( \11394 , \11392 , \11393 );
not \U$11148 ( \11395 , \10835 );
not \U$11149 ( \11396 , \10689 );
not \U$11150 ( \11397 , \11396 );
or \U$11151 ( \11398 , \11395 , \11397 );
buf \U$11152 ( \11399 , \10693 );
buf \U$11153 ( \11400 , \11399 );
nand \U$11154 ( \11401 , \11400 , RIbe2a190_83);
nand \U$11155 ( \11402 , \11398 , \11401 );
not \U$11156 ( \11403 , \11402 );
not \U$11157 ( \11404 , \10723 );
not \U$11158 ( \11405 , \8595 );
or \U$11159 ( \11406 , \11404 , \11405 );
xnor \U$11160 ( \11407 , RIbe29c68_72, RIbe28a98_34);
not \U$11161 ( \11408 , \11407 );
nand \U$11162 ( \11409 , \11408 , \4580 );
nand \U$11163 ( \11410 , \11406 , \11409 );
xor \U$11164 ( \11411 , \11403 , \11410 );
not \U$11165 ( \11412 , \10949 );
not \U$11166 ( \11413 , \2459 );
or \U$11167 ( \11414 , \11412 , \11413 );
xor \U$11168 ( \11415 , RIbe297b8_62, RIbe27e68_8);
nand \U$11169 ( \11416 , \4447 , \11415 );
nand \U$11170 ( \11417 , \11414 , \11416 );
not \U$11171 ( \11418 , \11417 );
xor \U$11172 ( \11419 , \11411 , \11418 );
not \U$11173 ( \11420 , \11419 );
xor \U$11174 ( \11421 , \10471 , \10479 );
xor \U$11175 ( \11422 , \11421 , \10487 );
xor \U$11176 ( \11423 , \11044 , \11058 );
xnor \U$11177 ( \11424 , \11422 , \11423 );
not \U$11178 ( \11425 , \11424 );
or \U$11179 ( \11426 , \11420 , \11425 );
not \U$11180 ( \11427 , \11423 );
nand \U$11181 ( \11428 , \11427 , \11422 );
nand \U$11182 ( \11429 , \11426 , \11428 );
and \U$11183 ( \11430 , \11394 , \11429 );
not \U$11184 ( \11431 , \11394 );
not \U$11185 ( \11432 , \11429 );
and \U$11186 ( \11433 , \11431 , \11432 );
nor \U$11187 ( \11434 , \11430 , \11433 );
not \U$11188 ( \11435 , \11434 );
xor \U$11189 ( \11436 , \11079 , \11070 );
xor \U$11190 ( \11437 , \11436 , \11077 );
not \U$11191 ( \11438 , \11437 );
not \U$11192 ( \11439 , \11438 );
or \U$11193 ( \11440 , \11435 , \11439 );
nand \U$11194 ( \11441 , \11394 , \11429 );
nand \U$11195 ( \11442 , \11440 , \11441 );
xor \U$11196 ( \11443 , \11171 , \11442 );
not \U$11197 ( \11444 , \11443 );
or \U$11198 ( \11445 , \11029 , \11444 );
nand \U$11199 ( \11446 , \11171 , \11442 );
nand \U$11200 ( \11447 , \11445 , \11446 );
not \U$11201 ( \11448 , \11447 );
not \U$11202 ( \11449 , \11448 );
xor \U$11203 ( \11450 , RIbe2a910_99, RIbe28048_12);
not \U$11204 ( \11451 , \11450 );
not \U$11205 ( \11452 , \9736 );
not \U$11206 ( \11453 , \11452 );
not \U$11207 ( \11454 , \11453 );
or \U$11208 ( \11455 , \11451 , \11454 );
buf \U$11209 ( \11456 , \10400 );
xor \U$11210 ( \11457 , RIbe2a910_99, RIbe29380_53);
nand \U$11211 ( \11458 , \11456 , \11457 );
nand \U$11212 ( \11459 , \11455 , \11458 );
not \U$11213 ( \11460 , \11142 );
not \U$11214 ( \11461 , \3255 );
not \U$11215 ( \11462 , \11461 );
or \U$11216 ( \11463 , \11460 , \11462 );
xnor \U$11217 ( \11464 , RIbe293f8_54, RIbe28f48_44);
not \U$11218 ( \11465 , \11464 );
nand \U$11219 ( \11466 , \11465 , \11201 );
nand \U$11220 ( \11467 , \11463 , \11466 );
xor \U$11221 ( \11468 , \11459 , \11467 );
xor \U$11222 ( \11469 , RIbe28a20_33, RIbe27df0_7);
not \U$11223 ( \11470 , \11469 );
not \U$11224 ( \11471 , \1781 );
or \U$11225 ( \11472 , \11470 , \11471 );
xor \U$11226 ( \11473 , RIbe29218_50, RIbe28a20_33);
nand \U$11227 ( \11474 , \2476 , \11473 );
nand \U$11228 ( \11475 , \11472 , \11474 );
xor \U$11229 ( \11476 , \11468 , \11475 );
not \U$11230 ( \11477 , \11103 );
not \U$11231 ( \11478 , \281 );
or \U$11232 ( \11479 , \11477 , \11478 );
xor \U$11233 ( \11480 , RIbe29038_46, RIbe29d58_74);
nand \U$11234 ( \11481 , \286 , \11480 );
nand \U$11235 ( \11482 , \11479 , \11481 );
not \U$11236 ( \11483 , \11482 );
not \U$11237 ( \11484 , \10438 );
buf \U$11238 ( \11485 , \11484 );
or \U$11239 ( \11486 , \10433 , \11485 );
nand \U$11240 ( \11487 , \11486 , RIbe2a550_91);
not \U$11241 ( \11488 , \11487 );
not \U$11242 ( \11489 , \11488 );
or \U$11243 ( \11490 , \11483 , \11489 );
or \U$11244 ( \11491 , \11488 , \11482 );
nand \U$11245 ( \11492 , \11490 , \11491 );
xor \U$11246 ( \11493 , RIbe29ce0_73, RIbe296c8_60);
not \U$11247 ( \11494 , \11493 );
not \U$11248 ( \11495 , \1130 );
or \U$11249 ( \11496 , \11494 , \11495 );
xor \U$11250 ( \11497 , RIbe296c8_60, RIbe29b78_70);
nand \U$11251 ( \11498 , \908 , \11497 );
nand \U$11252 ( \11499 , \11496 , \11498 );
xor \U$11253 ( \11500 , \11492 , \11499 );
and \U$11254 ( \11501 , \11476 , \11500 );
not \U$11255 ( \11502 , \11476 );
not \U$11256 ( \11503 , \11500 );
and \U$11257 ( \11504 , \11502 , \11503 );
nor \U$11258 ( \11505 , \11501 , \11504 );
xor \U$11259 ( \11506 , RIbe28d68_40, RIbe28930_31);
not \U$11260 ( \11507 , \11506 );
not \U$11261 ( \11508 , \965 );
or \U$11262 ( \11509 , \11507 , \11508 );
xor \U$11263 ( \11510 , RIbe28930_31, RIbe27c88_4);
nand \U$11264 ( \11511 , \1199 , \11510 );
nand \U$11265 ( \11512 , \11509 , \11511 );
xor \U$11266 ( \11513 , RIbe27c10_3, RIbe2a820_97);
not \U$11267 ( \11514 , \11513 );
not \U$11268 ( \11515 , \1103 );
or \U$11269 ( \11516 , \11514 , \11515 );
xor \U$11270 ( \11517 , RIbe2a898_98, RIbe27c10_3);
nand \U$11271 ( \11518 , \1498 , \11517 );
nand \U$11272 ( \11519 , \11516 , \11518 );
xor \U$11273 ( \11520 , \11512 , \11519 );
not \U$11274 ( \11521 , \11095 );
not \U$11275 ( \11522 , \10792 );
or \U$11276 ( \11523 , \11521 , \11522 );
xor \U$11277 ( \11524 , RIbe2a2f8_86, RIbe28570_23);
nand \U$11278 ( \11525 , \8706 , \11524 );
nand \U$11279 ( \11526 , \11523 , \11525 );
not \U$11280 ( \11527 , \11526 );
and \U$11281 ( \11528 , \11520 , \11527 );
not \U$11282 ( \11529 , \11520 );
and \U$11283 ( \11530 , \11529 , \11526 );
or \U$11284 ( \11531 , \11528 , \11530 );
and \U$11285 ( \11532 , \11505 , \11531 );
not \U$11286 ( \11533 , \11505 );
not \U$11287 ( \11534 , \11531 );
and \U$11288 ( \11535 , \11533 , \11534 );
nor \U$11289 ( \11536 , \11532 , \11535 );
not \U$11290 ( \11537 , \11536 );
xor \U$11291 ( \11538 , RIbe2a3e8_88, RIbe27ee0_9);
not \U$11292 ( \11539 , \11538 );
not \U$11293 ( \11540 , \9268 );
not \U$11294 ( \11541 , \11540 );
not \U$11295 ( \11542 , \11541 );
or \U$11296 ( \11543 , \11539 , \11542 );
not \U$11297 ( \11544 , \9263 );
xor \U$11298 ( \11545 , RIbe2a3e8_88, RIbe286d8_26);
not \U$11299 ( \11546 , \11545 );
or \U$11300 ( \11547 , \11544 , \11546 );
nand \U$11301 ( \11548 , \11543 , \11547 );
not \U$11302 ( \11549 , \11121 );
not \U$11303 ( \11550 , \2379 );
or \U$11304 ( \11551 , \11549 , \11550 );
xor \U$11305 ( \11552 , RIbe28cf0_39, RIbe280c0_13);
nand \U$11306 ( \11553 , \1263 , \11552 );
nand \U$11307 ( \11554 , \11551 , \11553 );
xor \U$11308 ( \11555 , RIbe285e8_24, RIbe297b8_62);
not \U$11309 ( \11556 , \11555 );
not \U$11310 ( \11557 , \8813 );
or \U$11311 ( \11558 , \11556 , \11557 );
xor \U$11312 ( \11559 , RIbe28138_14, RIbe285e8_24);
nand \U$11313 ( \11560 , \2625 , \11559 );
nand \U$11314 ( \11561 , \11558 , \11560 );
and \U$11315 ( \11562 , \11554 , \11561 );
not \U$11316 ( \11563 , \11554 );
not \U$11317 ( \11564 , \11561 );
and \U$11318 ( \11565 , \11563 , \11564 );
nor \U$11319 ( \11566 , \11562 , \11565 );
xor \U$11320 ( \11567 , \11548 , \11566 );
not \U$11321 ( \11568 , \2553 );
not \U$11322 ( \11569 , RIbe28b88_36);
not \U$11323 ( \11570 , RIbe29218_50);
and \U$11324 ( \11571 , \11569 , \11570 );
and \U$11325 ( \11572 , RIbe28b88_36, RIbe29218_50);
nor \U$11326 ( \11573 , \11571 , \11572 );
not \U$11327 ( \11574 , \11573 );
or \U$11328 ( \11575 , \11568 , \11574 );
xor \U$11329 ( \11576 , RIbe29a10_67, RIbe28b88_36);
nand \U$11330 ( \11577 , \2559 , \11576 );
nand \U$11331 ( \11578 , \11575 , \11577 );
not \U$11332 ( \11579 , \11087 );
not \U$11333 ( \11580 , \8169 );
or \U$11334 ( \11581 , \11579 , \11580 );
xor \U$11335 ( \11582 , RIbe2a028_80, RIbe28750_27);
nand \U$11336 ( \11583 , \8930 , \11582 );
nand \U$11337 ( \11584 , \11581 , \11583 );
nor \U$11338 ( \11585 , \11578 , \11584 );
not \U$11339 ( \11586 , \11585 );
nand \U$11340 ( \11587 , \11578 , \11584 );
nand \U$11341 ( \11588 , \11586 , \11587 );
not \U$11342 ( \11589 , \11114 );
not \U$11343 ( \11590 , \4842 );
or \U$11344 ( \11591 , \11589 , \11590 );
and \U$11345 ( \11592 , RIbe29e48_76, RIbe28318_18);
not \U$11346 ( \11593 , RIbe29e48_76);
and \U$11347 ( \11594 , \11593 , \2244 );
nor \U$11348 ( \11595 , \11592 , \11594 );
nand \U$11349 ( \11596 , \8245 , \11595 );
nand \U$11350 ( \11597 , \11591 , \11596 );
xor \U$11351 ( \11598 , \11588 , \11597 );
xor \U$11352 ( \11599 , \11567 , \11598 );
not \U$11353 ( \11600 , \11415 );
not \U$11354 ( \11601 , \2459 );
or \U$11355 ( \11602 , \11600 , \11601 );
xor \U$11356 ( \11603 , RIbe27e68_8, RIbe28138_14);
nand \U$11357 ( \11604 , \2464 , \11603 );
nand \U$11358 ( \11605 , \11602 , \11604 );
not \U$11359 ( \11606 , \11605 );
not \U$11360 ( \11607 , \10554 );
not \U$11361 ( \11608 , \8401 );
or \U$11362 ( \11609 , \11607 , \11608 );
nand \U$11363 ( \11610 , \8172 , \11083 );
nand \U$11364 ( \11611 , \11609 , \11610 );
not \U$11365 ( \11612 , \11611 );
or \U$11366 ( \11613 , \11606 , \11612 );
or \U$11367 ( \11614 , \11611 , \11605 );
not \U$11368 ( \11615 , \11042 );
not \U$11369 ( \11616 , \4842 );
or \U$11370 ( \11617 , \11615 , \11616 );
nand \U$11371 ( \11618 , \7368 , \11110 );
nand \U$11372 ( \11619 , \11617 , \11618 );
nand \U$11373 ( \11620 , \11614 , \11619 );
nand \U$11374 ( \11621 , \11613 , \11620 );
not \U$11375 ( \11622 , \11621 );
nand \U$11376 ( \11623 , RIbe27b98_2, RIbe2a460_89);
not \U$11377 ( \11624 , \11623 );
and \U$11378 ( \11625 , \11578 , \11624 );
not \U$11379 ( \11626 , \11578 );
and \U$11380 ( \11627 , \11626 , \11623 );
or \U$11381 ( \11628 , \11625 , \11627 );
not \U$11382 ( \11629 , \11628 );
or \U$11383 ( \11630 , \11622 , \11629 );
not \U$11384 ( \11631 , \11578 );
nand \U$11385 ( \11632 , \11631 , \11624 );
nand \U$11386 ( \11633 , \11630 , \11632 );
xor \U$11387 ( \11634 , \11599 , \11633 );
not \U$11388 ( \11635 , \11634 );
or \U$11389 ( \11636 , \11537 , \11635 );
or \U$11390 ( \11637 , \11634 , \11536 );
nand \U$11391 ( \11638 , \11636 , \11637 );
not \U$11392 ( \11639 , \11054 );
not \U$11393 ( \11640 , \10611 );
not \U$11394 ( \11641 , \10599 );
or \U$11395 ( \11642 , \11640 , \11641 );
nand \U$11396 ( \11643 , \10598 , \10591 );
nand \U$11397 ( \11644 , \11642 , \11643 );
not \U$11398 ( \11645 , \11644 );
or \U$11399 ( \11646 , \11639 , \11645 );
or \U$11400 ( \11647 , \11644 , \11054 );
not \U$11401 ( \11648 , \10547 );
not \U$11402 ( \11649 , \10538 );
or \U$11403 ( \11650 , \11648 , \11649 );
or \U$11404 ( \11651 , \10538 , \10547 );
nand \U$11405 ( \11652 , \11651 , \10531 );
nand \U$11406 ( \11653 , \11650 , \11652 );
nand \U$11407 ( \11654 , \11647 , \11653 );
nand \U$11408 ( \11655 , \11646 , \11654 );
not \U$11409 ( \11656 , \11655 );
xor \U$11410 ( \11657 , RIbe2a3e8_88, RIbe28570_23);
not \U$11411 ( \11658 , \11657 );
not \U$11412 ( \11659 , \8806 );
or \U$11413 ( \11660 , \11658 , \11659 );
nand \U$11414 ( \11661 , \9268 , \11545 );
nand \U$11415 ( \11662 , \11660 , \11661 );
buf \U$11416 ( \11663 , \11662 );
xor \U$11417 ( \11664 , RIbe29470_55, RIbe27fd0_11);
not \U$11418 ( \11665 , \11664 );
not \U$11419 ( \11666 , \9825 );
or \U$11420 ( \11667 , \11665 , \11666 );
xor \U$11421 ( \11668 , RIbe27fd0_11, RIbe294e8_56);
nand \U$11422 ( \11669 , \7709 , \11668 );
nand \U$11423 ( \11670 , \11667 , \11669 );
xor \U$11424 ( \11671 , \11663 , \11670 );
xor \U$11425 ( \11672 , RIbe29998_66, RIbe28930_31);
not \U$11426 ( \11673 , \11672 );
not \U$11427 ( \11674 , \1793 );
or \U$11428 ( \11675 , \11673 , \11674 );
nand \U$11429 ( \11676 , \1797 , \11506 );
nand \U$11430 ( \11677 , \11675 , \11676 );
xor \U$11431 ( \11678 , \11671 , \11677 );
xor \U$11432 ( \11679 , \11628 , \11621 );
xor \U$11433 ( \11680 , \11678 , \11679 );
not \U$11434 ( \11681 , \11680 );
or \U$11435 ( \11682 , \11656 , \11681 );
nand \U$11436 ( \11683 , \11679 , \11678 );
nand \U$11437 ( \11684 , \11682 , \11683 );
and \U$11438 ( \11685 , \11638 , \11684 );
not \U$11439 ( \11686 , \11638 );
not \U$11440 ( \11687 , \11684 );
and \U$11441 ( \11688 , \11686 , \11687 );
nor \U$11442 ( \11689 , \11685 , \11688 );
not \U$11443 ( \11690 , \10573 );
not \U$11444 ( \11691 , \10556 );
or \U$11445 ( \11692 , \11690 , \11691 );
or \U$11446 ( \11693 , \10573 , \10556 );
nand \U$11447 ( \11694 , \11693 , \10563 );
nand \U$11448 ( \11695 , \11692 , \11694 );
not \U$11449 ( \11696 , \10507 );
not \U$11450 ( \11697 , \10499 );
or \U$11451 ( \11698 , \11696 , \11697 );
not \U$11452 ( \11699 , \10508 );
not \U$11453 ( \11700 , \10500 );
or \U$11454 ( \11701 , \11699 , \11700 );
nand \U$11455 ( \11702 , \11701 , \10519 );
nand \U$11456 ( \11703 , \11698 , \11702 );
not \U$11457 ( \11704 , \11703 );
xor \U$11458 ( \11705 , \11695 , \11704 );
not \U$11459 ( \11706 , \11417 );
nand \U$11460 ( \11707 , \11706 , \11403 );
not \U$11461 ( \11708 , \11707 );
not \U$11462 ( \11709 , \11410 );
or \U$11463 ( \11710 , \11708 , \11709 );
nand \U$11464 ( \11711 , \11402 , \11417 );
nand \U$11465 ( \11712 , \11710 , \11711 );
xor \U$11466 ( \11713 , \11705 , \11712 );
not \U$11467 ( \11714 , \11713 );
not \U$11468 ( \11715 , \11714 );
xor \U$11469 ( \11716 , \11054 , \11653 );
xnor \U$11470 ( \11717 , \11716 , \11644 );
not \U$11471 ( \11718 , \11717 );
not \U$11472 ( \11719 , \11718 );
or \U$11473 ( \11720 , \11715 , \11719 );
not \U$11474 ( \11721 , \11717 );
not \U$11475 ( \11722 , \11713 );
or \U$11476 ( \11723 , \11721 , \11722 );
not \U$11477 ( \11724 , \10903 );
not \U$11478 ( \11725 , \10915 );
or \U$11479 ( \11726 , \11724 , \11725 );
or \U$11480 ( \11727 , \10915 , \10903 );
nand \U$11481 ( \11728 , \11727 , \10909 );
nand \U$11482 ( \11729 , \11726 , \11728 );
nand \U$11483 ( \11730 , \11723 , \11729 );
nand \U$11484 ( \11731 , \11720 , \11730 );
not \U$11485 ( \11732 , \11731 );
not \U$11486 ( \11733 , \11732 );
not \U$11487 ( \11734 , \11695 );
nand \U$11488 ( \11735 , \11734 , \11704 );
not \U$11489 ( \11736 , \11735 );
not \U$11490 ( \11737 , \11712 );
or \U$11491 ( \11738 , \11736 , \11737 );
nand \U$11492 ( \11739 , \11703 , \11695 );
nand \U$11493 ( \11740 , \11738 , \11739 );
or \U$11494 ( \11741 , \10490 , \10422 );
nand \U$11495 ( \11742 , \11741 , \10462 );
nand \U$11496 ( \11743 , \10491 , \10422 );
nand \U$11497 ( \11744 , \11742 , \11743 );
not \U$11498 ( \11745 , \11744 );
xor \U$11499 ( \11746 , \11740 , \11745 );
not \U$11500 ( \11747 , \10449 );
not \U$11501 ( \11748 , \10446 );
or \U$11502 ( \11749 , \11747 , \11748 );
nand \U$11503 ( \11750 , \8706 , \11090 );
nand \U$11504 ( \11751 , \11749 , \11750 );
not \U$11505 ( \11752 , \10485 );
not \U$11506 ( \11753 , \965 );
or \U$11507 ( \11754 , \11752 , \11753 );
nand \U$11508 ( \11755 , \1199 , \11672 );
nand \U$11509 ( \11756 , \11754 , \11755 );
xor \U$11510 ( \11757 , \11751 , \11756 );
not \U$11511 ( \11758 , \10505 );
not \U$11512 ( \11759 , \1103 );
or \U$11513 ( \11760 , \11758 , \11759 );
xor \U$11514 ( \11761 , RIbe27c10_3, RIbe2a118_82);
nand \U$11515 ( \11762 , \1173 , \11761 );
nand \U$11516 ( \11763 , \11760 , \11762 );
and \U$11517 ( \11764 , \11757 , \11763 );
and \U$11518 ( \11765 , \11751 , \11756 );
or \U$11519 ( \11766 , \11764 , \11765 );
not \U$11520 ( \11767 , \10469 );
not \U$11521 ( \11768 , \11366 );
nor \U$11522 ( \11769 , \11767 , \11768 );
and \U$11523 ( \11770 , \2707 , \11664 );
nor \U$11524 ( \11771 , \11769 , \11770 );
not \U$11525 ( \11772 , \11771 );
not \U$11526 ( \11773 , \11772 );
not \U$11527 ( \11774 , \10417 );
not \U$11528 ( \11775 , \1164 );
or \U$11529 ( \11776 , \11774 , \11775 );
nand \U$11530 ( \11777 , \314 , \11153 );
nand \U$11531 ( \11778 , \11776 , \11777 );
not \U$11532 ( \11779 , \10536 );
not \U$11533 ( \11780 , \256 );
or \U$11534 ( \11781 , \11779 , \11780 );
nand \U$11535 ( \11782 , \267 , \11124 );
nand \U$11536 ( \11783 , \11781 , \11782 );
xor \U$11537 ( \11784 , \11778 , \11783 );
not \U$11538 ( \11785 , \11784 );
or \U$11539 ( \11786 , \11773 , \11785 );
nand \U$11540 ( \11787 , \11783 , \11778 );
nand \U$11541 ( \11788 , \11786 , \11787 );
xor \U$11542 ( \11789 , \11766 , \11788 );
nand \U$11543 ( \11790 , RIbe27b98_2, RIbe2adc0_109);
not \U$11544 ( \11791 , \11790 );
not \U$11545 ( \11792 , \11791 );
not \U$11546 ( \11793 , \10561 );
not \U$11547 ( \11794 , \924 );
or \U$11548 ( \11795 , \11793 , \11794 );
xor \U$11549 ( \11796 , RIbe2b360_121, RIbe28de0_41);
nand \U$11550 ( \11797 , \347 , \11796 );
nand \U$11551 ( \11798 , \11795 , \11797 );
not \U$11552 ( \11799 , \11798 );
or \U$11553 ( \11800 , \11792 , \11799 );
xor \U$11554 ( \11801 , \11798 , \11790 );
not \U$11555 ( \11802 , \11801 );
and \U$11556 ( \11803 , \2520 , \10589 );
xor \U$11557 ( \11804 , RIbe28480_21, RIbe291a0_49);
and \U$11558 ( \11805 , \2527 , \11804 );
nor \U$11559 ( \11806 , \11803 , \11805 );
not \U$11560 ( \11807 , \11806 );
nand \U$11561 ( \11808 , \11802 , \11807 );
nand \U$11562 ( \11809 , \11800 , \11808 );
xor \U$11563 ( \11810 , \11789 , \11809 );
xor \U$11564 ( \11811 , \11746 , \11810 );
not \U$11565 ( \11812 , \11811 );
or \U$11566 ( \11813 , \11733 , \11812 );
xor \U$11567 ( \11814 , \11655 , \11680 );
nand \U$11568 ( \11815 , \11813 , \11814 );
not \U$11569 ( \11816 , \11811 );
nand \U$11570 ( \11817 , \11816 , \11731 );
nand \U$11571 ( \11818 , \11815 , \11817 );
not \U$11572 ( \11819 , \11818 );
xor \U$11573 ( \11820 , \11689 , \11819 );
not \U$11574 ( \11821 , \11037 );
not \U$11575 ( \11822 , \11167 );
not \U$11576 ( \11823 , \11822 );
or \U$11577 ( \11824 , \11821 , \11823 );
nand \U$11578 ( \11825 , \11162 , \11082 );
nand \U$11579 ( \11826 , \11824 , \11825 );
not \U$11580 ( \11827 , \11826 );
xor \U$11581 ( \11828 , \11820 , \11827 );
not \U$11582 ( \11829 , \11828 );
not \U$11583 ( \11830 , \11829 );
or \U$11584 ( \11831 , \11449 , \11830 );
not \U$11585 ( \11832 , \11447 );
not \U$11586 ( \11833 , \11828 );
or \U$11587 ( \11834 , \11832 , \11833 );
xor \U$11588 ( \11835 , RIbe285e8_24, RIbe29740_61);
not \U$11589 ( \11836 , \11835 );
not \U$11590 ( \11837 , \2618 );
or \U$11591 ( \11838 , \11836 , \11837 );
nand \U$11592 ( \11839 , \8270 , \11555 );
nand \U$11593 ( \11840 , \11838 , \11839 );
xor \U$11594 ( \11841 , RIbe2a550_91, RIbe29380_53);
not \U$11595 ( \11842 , \11841 );
not \U$11596 ( \11843 , \10433 );
or \U$11597 ( \11844 , \11842 , \11843 );
nand \U$11598 ( \11845 , \11227 , RIbe2a550_91);
nand \U$11599 ( \11846 , \11844 , \11845 );
not \U$11600 ( \11847 , \11846 );
and \U$11601 ( \11848 , \11840 , \11847 );
not \U$11602 ( \11849 , \11840 );
and \U$11603 ( \11850 , \11849 , \11846 );
or \U$11604 ( \11851 , \11848 , \11850 );
xor \U$11605 ( \11852 , RIbe28a20_33, RIbe27c88_4);
not \U$11606 ( \11853 , \11852 );
not \U$11607 ( \11854 , \2276 );
or \U$11608 ( \11855 , \11853 , \11854 );
nand \U$11609 ( \11856 , \5055 , \11469 );
nand \U$11610 ( \11857 , \11855 , \11856 );
not \U$11611 ( \11858 , \11857 );
not \U$11612 ( \11859 , \11858 );
and \U$11613 ( \11860 , \11851 , \11859 );
not \U$11614 ( \11861 , \11851 );
and \U$11615 ( \11862 , \11861 , \11858 );
nor \U$11616 ( \11863 , \11860 , \11862 );
not \U$11617 ( \11864 , \11863 );
xor \U$11618 ( \11865 , RIbe2a910_99, RIbe27ee0_9);
not \U$11619 ( \11866 , \11865 );
not \U$11620 ( \11867 , \9737 );
or \U$11621 ( \11868 , \11866 , \11867 );
nand \U$11622 ( \11869 , \10400 , \11450 );
nand \U$11623 ( \11870 , \11868 , \11869 );
not \U$11624 ( \11871 , \11603 );
not \U$11625 ( \11872 , \2457 );
or \U$11626 ( \11873 , \11871 , \11872 );
xor \U$11627 ( \11874 , RIbe27e68_8, RIbe282a0_17);
nand \U$11628 ( \11875 , \2463 , \11874 );
nand \U$11629 ( \11876 , \11873 , \11875 );
or \U$11630 ( \11877 , \11870 , \11876 );
not \U$11631 ( \11878 , \11865 );
not \U$11632 ( \11879 , \9737 );
or \U$11633 ( \11880 , \11878 , \11879 );
nand \U$11634 ( \11881 , \11880 , \11869 );
nand \U$11635 ( \11882 , \11881 , \11876 );
nand \U$11636 ( \11883 , \11877 , \11882 );
not \U$11637 ( \11884 , \4577 );
xnor \U$11638 ( \11885 , RIbe293f8_54, RIbe29c68_72);
not \U$11639 ( \11886 , \11885 );
and \U$11640 ( \11887 , \11884 , \11886 );
xnor \U$11641 ( \11888 , RIbe29308_52, RIbe29c68_72);
nor \U$11642 ( \11889 , \4581 , \11888 );
nor \U$11643 ( \11890 , \11887 , \11889 );
not \U$11644 ( \11891 , \11890 );
and \U$11645 ( \11892 , \11883 , \11891 );
not \U$11646 ( \11893 , \11883 );
and \U$11647 ( \11894 , \11893 , \11890 );
nor \U$11648 ( \11895 , \11892 , \11894 );
not \U$11649 ( \11896 , \11895 );
or \U$11650 ( \11897 , \11864 , \11896 );
or \U$11651 ( \11898 , \11895 , \11863 );
nand \U$11652 ( \11899 , \11897 , \11898 );
xor \U$11653 ( \11900 , RIbe296c8_60, RIbe29d58_74);
not \U$11654 ( \11901 , \11900 );
not \U$11655 ( \11902 , \2875 );
or \U$11656 ( \11903 , \11901 , \11902 );
nand \U$11657 ( \11904 , \908 , \11493 );
nand \U$11658 ( \11905 , \11903 , \11904 );
not \U$11659 ( \11906 , \11761 );
and \U$11660 ( \11907 , \356 , \357 );
not \U$11661 ( \11908 , \11907 );
or \U$11662 ( \11909 , \11906 , \11908 );
nand \U$11663 ( \11910 , \1173 , \11513 );
nand \U$11664 ( \11911 , \11909 , \11910 );
not \U$11665 ( \11912 , \11911 );
xor \U$11666 ( \11913 , \11905 , \11912 );
xor \U$11667 ( \11914 , RIbe28228_16, RIbe28cf0_39);
not \U$11668 ( \11915 , \11914 );
not \U$11669 ( \11916 , \3056 );
or \U$11670 ( \11917 , \11915 , \11916 );
xor \U$11671 ( \11918 , RIbe28228_16, RIbe298a8_64);
nand \U$11672 ( \11919 , \8679 , \11918 );
nand \U$11673 ( \11920 , \11917 , \11919 );
xor \U$11674 ( \11921 , \11913 , \11920 );
and \U$11675 ( \11922 , \11899 , \11921 );
not \U$11676 ( \11923 , \11899 );
not \U$11677 ( \11924 , \11921 );
and \U$11678 ( \11925 , \11923 , \11924 );
nor \U$11679 ( \11926 , \11922 , \11925 );
not \U$11680 ( \11927 , \11926 );
not \U$11681 ( \11928 , \10571 );
not \U$11682 ( \11929 , \9114 );
or \U$11683 ( \11930 , \11928 , \11929 );
xor \U$11684 ( \11931 , RIbe290b0_47, RIbe2aa78_102);
nand \U$11685 ( \11932 , \2071 , \11931 );
nand \U$11686 ( \11933 , \11930 , \11932 );
or \U$11687 ( \11934 , \4577 , \11407 );
or \U$11688 ( \11935 , \7236 , \11885 );
nand \U$11689 ( \11936 , \11934 , \11935 );
nor \U$11690 ( \11937 , \11933 , \11936 );
not \U$11691 ( \11938 , \3401 );
not \U$11692 ( \11939 , \11938 );
not \U$11693 ( \11940 , \11052 );
not \U$11694 ( \11941 , \11940 );
and \U$11695 ( \11942 , \11939 , \11941 );
and \U$11696 ( \11943 , \2560 , \11573 );
nor \U$11697 ( \11944 , \11942 , \11943 );
or \U$11698 ( \11945 , \11937 , \11944 );
nand \U$11699 ( \11946 , \11936 , \11933 );
nand \U$11700 ( \11947 , \11945 , \11946 );
not \U$11701 ( \11948 , \11931 );
not \U$11702 ( \11949 , \2730 );
or \U$11703 ( \11950 , \11948 , \11949 );
xor \U$11704 ( \11951 , RIbe290b0_47, RIbe2b6a8_128);
nand \U$11705 ( \11952 , \10730 , \11951 );
nand \U$11706 ( \11953 , \11950 , \11952 );
not \U$11707 ( \11954 , \11804 );
not \U$11708 ( \11955 , \2518 );
or \U$11709 ( \11956 , \11954 , \11955 );
xor \U$11710 ( \11957 , RIbe28480_21, RIbe295d8_58);
nand \U$11711 ( \11958 , \3074 , \11957 );
nand \U$11712 ( \11959 , \11956 , \11958 );
not \U$11713 ( \11960 , \11959 );
xor \U$11714 ( \11961 , \11953 , \11960 );
not \U$11715 ( \11962 , \11796 );
not \U$11716 ( \11963 , \924 );
or \U$11717 ( \11964 , \11962 , \11963 );
xor \U$11718 ( \11965 , RIbe28de0_41, RIbe2a0a0_81);
nand \U$11719 ( \11966 , \347 , \11965 );
nand \U$11720 ( \11967 , \11964 , \11966 );
xor \U$11721 ( \11968 , \11961 , \11967 );
not \U$11722 ( \11969 , \11968 );
xor \U$11723 ( \11970 , \11947 , \11969 );
not \U$11724 ( \11971 , \11400 );
not \U$11725 ( \11972 , \11971 );
not \U$11726 ( \11973 , \11396 );
not \U$11727 ( \11974 , \11973 );
or \U$11728 ( \11975 , \11972 , \11974 );
nand \U$11729 ( \11976 , \11975 , RIbe2a190_83);
not \U$11730 ( \11977 , \11976 );
not \U$11731 ( \11978 , \10497 );
not \U$11732 ( \11979 , \879 );
or \U$11733 ( \11980 , \11978 , \11979 );
nand \U$11734 ( \11981 , \885 , \11914 );
nand \U$11735 ( \11982 , \11980 , \11981 );
not \U$11736 ( \11983 , \10529 );
not \U$11737 ( \11984 , \2639 );
or \U$11738 ( \11985 , \11983 , \11984 );
nand \U$11739 ( \11986 , \8654 , \11145 );
nand \U$11740 ( \11987 , \11985 , \11986 );
xor \U$11741 ( \11988 , \11982 , \11987 );
not \U$11742 ( \11989 , \11988 );
or \U$11743 ( \11990 , \11977 , \11989 );
nand \U$11744 ( \11991 , \11982 , \11987 );
nand \U$11745 ( \11992 , \11990 , \11991 );
xnor \U$11746 ( \11993 , \11970 , \11992 );
not \U$11747 ( \11994 , \11993 );
nand \U$11748 ( \11995 , \11927 , \11994 );
nand \U$11749 ( \11996 , \11926 , \11993 );
nand \U$11750 ( \11997 , \11995 , \11996 );
not \U$11751 ( \11998 , \10441 );
buf \U$11752 ( \11999 , \10432 );
buf \U$11753 ( \12000 , \11999 );
not \U$11754 ( \12001 , \12000 );
or \U$11755 ( \12002 , \11998 , \12001 );
not \U$11756 ( \12003 , \11484 );
not \U$11757 ( \12004 , \12003 );
nand \U$11758 ( \12005 , \12004 , \11841 );
nand \U$11759 ( \12006 , \12002 , \12005 );
not \U$11760 ( \12007 , \10457 );
not \U$11761 ( \12008 , \281 );
or \U$11762 ( \12009 , \12007 , \12008 );
nand \U$11763 ( \12010 , \1583 , \11099 );
nand \U$11764 ( \12011 , \12009 , \12010 );
nor \U$11765 ( \12012 , \12006 , \12011 );
not \U$11766 ( \12013 , \2876 );
not \U$11767 ( \12014 , \10517 );
not \U$11768 ( \12015 , \12014 );
and \U$11769 ( \12016 , \12013 , \12015 );
and \U$11770 ( \12017 , \907 , \11900 );
nor \U$11771 ( \12018 , \12016 , \12017 );
or \U$11772 ( \12019 , \12012 , \12018 );
nand \U$11773 ( \12020 , \12011 , \12006 );
nand \U$11774 ( \12021 , \12019 , \12020 );
not \U$11775 ( \12022 , \10402 );
not \U$11776 ( \12023 , \10987 );
or \U$11777 ( \12024 , \12022 , \12023 );
nand \U$11778 ( \12025 , \11456 , \11865 );
nand \U$11779 ( \12026 , \12024 , \12025 );
not \U$11780 ( \12027 , \1780 );
or \U$11781 ( \12028 , \12027 , \10608 );
nand \U$11782 ( \12029 , \5055 , \11852 );
nand \U$11783 ( \12030 , \12028 , \12029 );
nor \U$11784 ( \12031 , \12026 , \12030 );
buf \U$11785 ( \12032 , \12031 );
not \U$11786 ( \12033 , \10409 );
not \U$11787 ( \12034 , \3256 );
or \U$11788 ( \12035 , \12033 , \12034 );
nand \U$11789 ( \12036 , \3249 , \11138 );
nand \U$11790 ( \12037 , \12035 , \12036 );
not \U$11791 ( \12038 , \12037 );
or \U$11792 ( \12039 , \12032 , \12038 );
nand \U$11793 ( \12040 , \12026 , \12030 );
nand \U$11794 ( \12041 , \12039 , \12040 );
xor \U$11795 ( \12042 , \12021 , \12041 );
not \U$11796 ( \12043 , \10545 );
not \U$11797 ( \12044 , \2379 );
or \U$11798 ( \12045 , \12043 , \12044 );
nand \U$11799 ( \12046 , \869 , \11117 );
nand \U$11800 ( \12047 , \12045 , \12046 );
not \U$11801 ( \12048 , \12047 );
not \U$11802 ( \12049 , \10596 );
not \U$11803 ( \12050 , \2761 );
or \U$11804 ( \12051 , \12049 , \12050 );
nand \U$11805 ( \12052 , \8270 , \11835 );
nand \U$11806 ( \12053 , \12051 , \12052 );
not \U$11807 ( \12054 , \12053 );
or \U$11808 ( \12055 , \12048 , \12054 );
xnor \U$11809 ( \12056 , \12047 , \12053 );
not \U$11810 ( \12057 , \10477 );
not \U$11811 ( \12058 , \9264 );
or \U$11812 ( \12059 , \12057 , \12058 );
nand \U$11813 ( \12060 , \8794 , \11657 );
nand \U$11814 ( \12061 , \12059 , \12060 );
not \U$11815 ( \12062 , \12061 );
or \U$11816 ( \12063 , \12056 , \12062 );
nand \U$11817 ( \12064 , \12055 , \12063 );
xor \U$11818 ( \12065 , \12042 , \12064 );
not \U$11819 ( \12066 , \12065 );
and \U$11820 ( \12067 , \11997 , \12066 );
not \U$11821 ( \12068 , \11997 );
and \U$11822 ( \12069 , \12068 , \12065 );
nor \U$11823 ( \12070 , \12067 , \12069 );
not \U$11824 ( \12071 , \12070 );
not \U$11825 ( \12072 , \12071 );
and \U$11826 ( \12073 , \11801 , \11806 );
not \U$11827 ( \12074 , \11801 );
and \U$11828 ( \12075 , \12074 , \11807 );
nor \U$11829 ( \12076 , \12073 , \12075 );
not \U$11830 ( \12077 , \11611 );
not \U$11831 ( \12078 , \11605 );
not \U$11832 ( \12079 , \12078 );
or \U$11833 ( \12080 , \12077 , \12079 );
not \U$11834 ( \12081 , \11611 );
nand \U$11835 ( \12082 , \12081 , \11605 );
nand \U$11836 ( \12083 , \12080 , \12082 );
and \U$11837 ( \12084 , \12083 , \11619 );
not \U$11838 ( \12085 , \12083 );
not \U$11839 ( \12086 , \11619 );
and \U$11840 ( \12087 , \12085 , \12086 );
nor \U$11841 ( \12088 , \12084 , \12087 );
xor \U$11842 ( \12089 , \12076 , \12088 );
not \U$11843 ( \12090 , \11771 );
not \U$11844 ( \12091 , \11784 );
or \U$11845 ( \12092 , \12090 , \12091 );
or \U$11846 ( \12093 , \11784 , \11771 );
nand \U$11847 ( \12094 , \12092 , \12093 );
and \U$11848 ( \12095 , \12089 , \12094 );
and \U$11849 ( \12096 , \12076 , \12088 );
or \U$11850 ( \12097 , \12095 , \12096 );
not \U$11851 ( \12098 , \12097 );
not \U$11852 ( \12099 , RIbe2a190_83);
nor \U$11853 ( \12100 , \11400 , \11396 );
nor \U$11854 ( \12101 , \12099 , \12100 );
not \U$11855 ( \12102 , \12101 );
not \U$11856 ( \12103 , \11988 );
and \U$11857 ( \12104 , \12102 , \12103 );
and \U$11858 ( \12105 , \11988 , \12101 );
nor \U$11859 ( \12106 , \12104 , \12105 );
not \U$11860 ( \12107 , \12106 );
xor \U$11861 ( \12108 , \12011 , \12018 );
xor \U$11862 ( \12109 , \12108 , \12006 );
not \U$11863 ( \12110 , \12109 );
or \U$11864 ( \12111 , \12107 , \12110 );
xor \U$11865 ( \12112 , \11751 , \11756 );
xor \U$11866 ( \12113 , \12112 , \11763 );
nand \U$11867 ( \12114 , \12111 , \12113 );
not \U$11868 ( \12115 , \12106 );
not \U$11869 ( \12116 , \12109 );
nand \U$11870 ( \12117 , \12115 , \12116 );
nand \U$11871 ( \12118 , \12114 , \12117 );
not \U$11872 ( \12119 , \12118 );
not \U$11873 ( \12120 , \12061 );
not \U$11874 ( \12121 , \12056 );
and \U$11875 ( \12122 , \12120 , \12121 );
and \U$11876 ( \12123 , \12056 , \12061 );
nor \U$11877 ( \12124 , \12122 , \12123 );
not \U$11878 ( \12125 , \12124 );
not \U$11879 ( \12126 , \12125 );
not \U$11880 ( \12127 , \12031 );
nand \U$11881 ( \12128 , \12127 , \12040 );
and \U$11882 ( \12129 , \12128 , \12037 );
not \U$11883 ( \12130 , \12128 );
and \U$11884 ( \12131 , \12130 , \12038 );
nor \U$11885 ( \12132 , \12129 , \12131 );
not \U$11886 ( \12133 , \12132 );
not \U$11887 ( \12134 , \12133 );
or \U$11888 ( \12135 , \12126 , \12134 );
not \U$11889 ( \12136 , \12132 );
not \U$11890 ( \12137 , \12124 );
or \U$11891 ( \12138 , \12136 , \12137 );
not \U$11892 ( \12139 , \11937 );
nand \U$11893 ( \12140 , \12139 , \11946 );
and \U$11894 ( \12141 , \12140 , \11944 );
not \U$11895 ( \12142 , \12140 );
not \U$11896 ( \12143 , \11944 );
and \U$11897 ( \12144 , \12142 , \12143 );
nor \U$11898 ( \12145 , \12141 , \12144 );
nand \U$11899 ( \12146 , \12138 , \12145 );
nand \U$11900 ( \12147 , \12135 , \12146 );
not \U$11901 ( \12148 , \12147 );
not \U$11902 ( \12149 , \12148 );
and \U$11903 ( \12150 , \12119 , \12149 );
and \U$11904 ( \12151 , \12118 , \12148 );
nor \U$11905 ( \12152 , \12150 , \12151 );
not \U$11906 ( \12153 , \12152 );
or \U$11907 ( \12154 , \12098 , \12153 );
or \U$11908 ( \12155 , \12097 , \12152 );
nand \U$11909 ( \12156 , \12154 , \12155 );
not \U$11910 ( \12157 , \12156 );
not \U$11911 ( \12158 , \12133 );
not \U$11912 ( \12159 , \12124 );
or \U$11913 ( \12160 , \12158 , \12159 );
nand \U$11914 ( \12161 , \12125 , \12132 );
nand \U$11915 ( \12162 , \12160 , \12161 );
and \U$11916 ( \12163 , \12162 , \12145 );
not \U$11917 ( \12164 , \12162 );
not \U$11918 ( \12165 , \12145 );
and \U$11919 ( \12166 , \12164 , \12165 );
nor \U$11920 ( \12167 , \12163 , \12166 );
not \U$11921 ( \12168 , \12167 );
xor \U$11922 ( \12169 , \12076 , \12088 );
xor \U$11923 ( \12170 , \12169 , \12094 );
not \U$11924 ( \12171 , \12170 );
or \U$11925 ( \12172 , \12168 , \12171 );
or \U$11926 ( \12173 , \12167 , \12170 );
xor \U$11927 ( \12174 , \12113 , \12106 );
xnor \U$11928 ( \12175 , \12174 , \12116 );
nand \U$11929 ( \12176 , \12173 , \12175 );
nand \U$11930 ( \12177 , \12172 , \12176 );
not \U$11931 ( \12178 , \12177 );
not \U$11932 ( \12179 , \12178 );
and \U$11933 ( \12180 , \12157 , \12179 );
and \U$11934 ( \12181 , \12156 , \12178 );
nor \U$11935 ( \12182 , \12180 , \12181 );
not \U$11936 ( \12183 , \12182 );
not \U$11937 ( \12184 , \12183 );
or \U$11938 ( \12185 , \12072 , \12184 );
nand \U$11939 ( \12186 , \12182 , \12070 );
nand \U$11940 ( \12187 , \12185 , \12186 );
not \U$11941 ( \12188 , \11814 );
not \U$11942 ( \12189 , \11731 );
buf \U$11943 ( \12190 , \11811 );
nand \U$11944 ( \12191 , \12189 , \12190 );
nand \U$11945 ( \12192 , \12191 , \11817 );
not \U$11946 ( \12193 , \12192 );
or \U$11947 ( \12194 , \12188 , \12193 );
or \U$11948 ( \12195 , \12192 , \11814 );
nand \U$11949 ( \12196 , \12194 , \12195 );
or \U$11950 ( \12197 , \12187 , \12196 );
buf \U$11951 ( \12198 , \12170 );
not \U$11952 ( \12199 , \12198 );
not \U$11953 ( \12200 , \12167 );
and \U$11954 ( \12201 , \12175 , \12200 );
not \U$11955 ( \12202 , \12175 );
and \U$11956 ( \12203 , \12202 , \12167 );
nor \U$11957 ( \12204 , \12201 , \12203 );
not \U$11958 ( \12205 , \12204 );
or \U$11959 ( \12206 , \12199 , \12205 );
or \U$11960 ( \12207 , \12204 , \12198 );
nand \U$11961 ( \12208 , \12206 , \12207 );
not \U$11962 ( \12209 , \12208 );
xor \U$11963 ( \12210 , \11718 , \11714 );
not \U$11964 ( \12211 , \11729 );
xor \U$11965 ( \12212 , \12210 , \12211 );
not \U$11966 ( \12213 , \12212 );
nand \U$11967 ( \12214 , \10621 , \10613 );
not \U$11968 ( \12215 , \10616 );
and \U$11969 ( \12216 , \12214 , \12215 );
not \U$11970 ( \12217 , \12214 );
and \U$11971 ( \12218 , \12217 , \10616 );
nor \U$11972 ( \12219 , \12216 , \12218 );
not \U$11973 ( \12220 , \12219 );
not \U$11974 ( \12221 , \11419 );
not \U$11975 ( \12222 , \12221 );
not \U$11976 ( \12223 , \11424 );
and \U$11977 ( \12224 , \12222 , \12223 );
and \U$11978 ( \12225 , \11424 , \12221 );
nor \U$11979 ( \12226 , \12224 , \12225 );
not \U$11980 ( \12227 , \12226 );
xor \U$11981 ( \12228 , \10524 , \10548 );
xor \U$11982 ( \12229 , \12228 , \10574 );
not \U$11983 ( \12230 , \12229 );
or \U$11984 ( \12231 , \12227 , \12230 );
or \U$11985 ( \12232 , \12226 , \12229 );
nand \U$11986 ( \12233 , \12231 , \12232 );
not \U$11987 ( \12234 , \12233 );
or \U$11988 ( \12235 , \12220 , \12234 );
not \U$11989 ( \12236 , \12226 );
nand \U$11990 ( \12237 , \12236 , \12229 );
nand \U$11991 ( \12238 , \12235 , \12237 );
not \U$11992 ( \12239 , \12238 );
or \U$11993 ( \12240 , \12213 , \12239 );
or \U$11994 ( \12241 , \12238 , \12212 );
nand \U$11995 ( \12242 , \12240 , \12241 );
not \U$11996 ( \12243 , \12242 );
or \U$11997 ( \12244 , \12209 , \12243 );
not \U$11998 ( \12245 , \12212 );
nand \U$11999 ( \12246 , \12245 , \12238 );
nand \U$12000 ( \12247 , \12244 , \12246 );
nand \U$12001 ( \12248 , \12197 , \12247 );
nand \U$12002 ( \12249 , \12187 , \12196 );
nand \U$12003 ( \12250 , \12248 , \12249 );
not \U$12004 ( \12251 , \12250 );
nand \U$12005 ( \12252 , \11834 , \12251 );
nand \U$12006 ( \12253 , \11831 , \12252 );
not \U$12007 ( \12254 , \12253 );
xor \U$12008 ( \12255 , \12021 , \12041 );
and \U$12009 ( \12256 , \12255 , \12064 );
and \U$12010 ( \12257 , \12021 , \12041 );
or \U$12011 ( \12258 , \12256 , \12257 );
not \U$12012 ( \12259 , \11105 );
not \U$12013 ( \12260 , \11089 );
or \U$12014 ( \12261 , \12259 , \12260 );
or \U$12015 ( \12262 , \11089 , \11105 );
nand \U$12016 ( \12263 , \12262 , \11097 );
nand \U$12017 ( \12264 , \12261 , \12263 );
nor \U$12018 ( \12265 , \11881 , \11876 );
or \U$12019 ( \12266 , \12265 , \11890 );
nand \U$12020 ( \12267 , \12266 , \11882 );
xor \U$12021 ( \12268 , \12264 , \12267 );
nor \U$12022 ( \12269 , \11953 , \11967 );
or \U$12023 ( \12270 , \12269 , \11960 );
nand \U$12024 ( \12271 , \11953 , \11967 );
nand \U$12025 ( \12272 , \12270 , \12271 );
xor \U$12026 ( \12273 , \12268 , \12272 );
nor \U$12027 ( \12274 , \12258 , \12273 );
buf \U$12028 ( \12275 , \12274 );
xor \U$12029 ( \12276 , \11766 , \11788 );
and \U$12030 ( \12277 , \12276 , \11809 );
and \U$12031 ( \12278 , \11766 , \11788 );
or \U$12032 ( \12279 , \12277 , \12278 );
not \U$12033 ( \12280 , \12279 );
or \U$12034 ( \12281 , \12275 , \12280 );
nand \U$12035 ( \12282 , \12258 , \12273 );
nand \U$12036 ( \12283 , \12281 , \12282 );
xor \U$12037 ( \12284 , \12264 , \12267 );
and \U$12038 ( \12285 , \12284 , \12272 );
and \U$12039 ( \12286 , \12264 , \12267 );
or \U$12040 ( \12287 , \12285 , \12286 );
not \U$12041 ( \12288 , \11670 );
not \U$12042 ( \12289 , \11662 );
or \U$12043 ( \12290 , \12288 , \12289 );
or \U$12044 ( \12291 , \11662 , \11670 );
nand \U$12045 ( \12292 , \12291 , \11677 );
nand \U$12046 ( \12293 , \12290 , \12292 );
not \U$12047 ( \12294 , \12293 );
or \U$12048 ( \12295 , \11920 , \11911 );
nand \U$12049 ( \12296 , \12295 , \11905 );
nand \U$12050 ( \12297 , \11920 , \11911 );
and \U$12051 ( \12298 , \12296 , \12297 );
not \U$12052 ( \12299 , \12298 );
not \U$12053 ( \12300 , \12299 );
or \U$12054 ( \12301 , \12294 , \12300 );
not \U$12055 ( \12302 , \12298 );
not \U$12056 ( \12303 , \12293 );
not \U$12057 ( \12304 , \12303 );
or \U$12058 ( \12305 , \12302 , \12304 );
not \U$12059 ( \12306 , \11160 );
not \U$12060 ( \12307 , \11152 );
or \U$12061 ( \12308 , \12306 , \12307 );
nand \U$12062 ( \12309 , \11144 , \11151 );
nand \U$12063 ( \12310 , \12308 , \12309 );
nand \U$12064 ( \12311 , \12305 , \12310 );
nand \U$12065 ( \12312 , \12301 , \12311 );
xor \U$12066 ( \12313 , \12287 , \12312 );
xor \U$12067 ( \12314 , RIbe29b00_69, RIbe28b88_36);
not \U$12068 ( \12315 , \12314 );
not \U$12069 ( \12316 , \2701 );
or \U$12070 ( \12317 , \12315 , \12316 );
nand \U$12071 ( \12318 , \2691 , \9302 );
nand \U$12072 ( \12319 , \12317 , \12318 );
not \U$12073 ( \12320 , \12319 );
and \U$12074 ( \12321 , \4828 , \11128 );
xor \U$12075 ( \12322 , RIbe2b360_121, RIbe27b98_2);
and \U$12076 ( \12323 , \7585 , \12322 );
nor \U$12077 ( \12324 , \12321 , \12323 );
not \U$12078 ( \12325 , \11668 );
not \U$12079 ( \12326 , \3377 );
or \U$12080 ( \12327 , \12325 , \12326 );
xor \U$12081 ( \12328 , RIbe27fd0_11, RIbe288b8_30);
nand \U$12082 ( \12329 , \4897 , \12328 );
nand \U$12083 ( \12330 , \12327 , \12329 );
not \U$12084 ( \12331 , \10752 );
xor \U$12085 ( \12332 , RIbe2aa78_102, RIbe27d78_6);
not \U$12086 ( \12333 , \12332 );
or \U$12087 ( \12334 , \12331 , \12333 );
or \U$12088 ( \12335 , \8897 , \11157 );
nand \U$12089 ( \12336 , \12334 , \12335 );
nor \U$12090 ( \12337 , \12330 , \12336 );
or \U$12091 ( \12338 , \12324 , \12337 );
nand \U$12092 ( \12339 , \12336 , \12330 );
nand \U$12093 ( \12340 , \12338 , \12339 );
not \U$12094 ( \12341 , \12340 );
or \U$12095 ( \12342 , \12320 , \12341 );
or \U$12096 ( \12343 , \12340 , \12319 );
nand \U$12097 ( \12344 , \12342 , \12343 );
buf \U$12098 ( \12345 , \12344 );
not \U$12099 ( \12346 , \11526 );
not \U$12100 ( \12347 , \11520 );
or \U$12101 ( \12348 , \12346 , \12347 );
nand \U$12102 ( \12349 , \11512 , \11519 );
nand \U$12103 ( \12350 , \12348 , \12349 );
and \U$12104 ( \12351 , \12345 , \12350 );
not \U$12105 ( \12352 , \12345 );
not \U$12106 ( \12353 , \12350 );
and \U$12107 ( \12354 , \12352 , \12353 );
nor \U$12108 ( \12355 , \12351 , \12354 );
not \U$12109 ( \12356 , \12355 );
and \U$12110 ( \12357 , \12313 , \12356 );
not \U$12111 ( \12358 , \12313 );
and \U$12112 ( \12359 , \12358 , \12355 );
nor \U$12113 ( \12360 , \12357 , \12359 );
not \U$12114 ( \12361 , \12360 );
not \U$12115 ( \12362 , \12361 );
xor \U$12116 ( \12363 , \12293 , \12299 );
xnor \U$12117 ( \12364 , \12363 , \12310 );
not \U$12118 ( \12365 , \11947 );
nand \U$12119 ( \12366 , \12365 , \11968 );
not \U$12120 ( \12367 , \12366 );
not \U$12121 ( \12368 , \11992 );
or \U$12122 ( \12369 , \12367 , \12368 );
nand \U$12123 ( \12370 , \11969 , \11947 );
nand \U$12124 ( \12371 , \12369 , \12370 );
not \U$12125 ( \12372 , \11921 );
not \U$12126 ( \12373 , \11895 );
or \U$12127 ( \12374 , \12372 , \12373 );
nand \U$12128 ( \12375 , \12374 , \11863 );
not \U$12129 ( \12376 , \11895 );
nand \U$12130 ( \12377 , \12376 , \11924 );
nand \U$12131 ( \12378 , \12375 , \12377 );
nor \U$12132 ( \12379 , \12371 , \12378 );
or \U$12133 ( \12380 , \12364 , \12379 );
nand \U$12134 ( \12381 , \12378 , \12371 );
nand \U$12135 ( \12382 , \12380 , \12381 );
not \U$12136 ( \12383 , \12382 );
not \U$12137 ( \12384 , \12383 );
or \U$12138 ( \12385 , \12362 , \12384 );
nand \U$12139 ( \12386 , \12382 , \12360 );
nand \U$12140 ( \12387 , \12385 , \12386 );
xor \U$12141 ( \12388 , \12283 , \12387 );
not \U$12142 ( \12389 , \11840 );
not \U$12143 ( \12390 , \11857 );
or \U$12144 ( \12391 , \12389 , \12390 );
nand \U$12145 ( \12392 , \12391 , \11847 );
not \U$12146 ( \12393 , \11840 );
nand \U$12147 ( \12394 , \12393 , \11858 );
and \U$12148 ( \12395 , \12392 , \12394 );
not \U$12149 ( \12396 , \12337 );
nand \U$12150 ( \12397 , \12396 , \12339 );
xor \U$12151 ( \12398 , \12397 , \12324 );
xor \U$12152 ( \12399 , \12395 , \12398 );
not \U$12153 ( \12400 , \11116 );
not \U$12154 ( \12401 , \11135 );
or \U$12155 ( \12402 , \12400 , \12401 );
not \U$12156 ( \12403 , \11133 );
nand \U$12157 ( \12404 , \12403 , \11123 );
nand \U$12158 ( \12405 , \12402 , \12404 );
xor \U$12159 ( \12406 , \12399 , \12405 );
and \U$12160 ( \12407 , \2519 , \11957 );
xor \U$12161 ( \12408 , RIbe28480_21, RIbe29740_61);
not \U$12162 ( \12409 , \12408 );
nor \U$12163 ( \12410 , \12409 , \2670 );
nor \U$12164 ( \12411 , \12407 , \12410 );
nand \U$12165 ( \12412 , RIbe27b98_2, RIbe2a4d8_90);
not \U$12166 ( \12413 , \12412 );
not \U$12167 ( \12414 , \11965 );
not \U$12168 ( \12415 , \11321 );
or \U$12169 ( \12416 , \12414 , \12415 );
xor \U$12170 ( \12417 , RIbe28de0_41, RIbe2a118_82);
nand \U$12171 ( \12418 , \346 , \12417 );
nand \U$12172 ( \12419 , \12416 , \12418 );
not \U$12173 ( \12420 , \12419 );
or \U$12174 ( \12421 , \12413 , \12420 );
or \U$12175 ( \12422 , \12419 , \12412 );
nand \U$12176 ( \12423 , \12421 , \12422 );
xnor \U$12177 ( \12424 , \12411 , \12423 );
not \U$12178 ( \12425 , \11888 );
not \U$12179 ( \12426 , \12425 );
not \U$12180 ( \12427 , \4578 );
or \U$12181 ( \12428 , \12426 , \12427 );
and \U$12182 ( \12429 , RIbe29c68_72, RIbe28c00_37);
not \U$12183 ( \12430 , RIbe29c68_72);
and \U$12184 ( \12431 , \12430 , \2479 );
nor \U$12185 ( \12432 , \12429 , \12431 );
nand \U$12186 ( \12433 , \4580 , \12432 );
nand \U$12187 ( \12434 , \12428 , \12433 );
not \U$12188 ( \12435 , \11951 );
not \U$12189 ( \12436 , \2730 );
or \U$12190 ( \12437 , \12435 , \12436 );
xor \U$12191 ( \12438 , RIbe29f38_78, RIbe290b0_47);
nand \U$12192 ( \12439 , \399 , \12438 );
nand \U$12193 ( \12440 , \12437 , \12439 );
not \U$12194 ( \12441 , \11576 );
not \U$12195 ( \12442 , \3401 );
or \U$12196 ( \12443 , \12441 , \12442 );
nand \U$12197 ( \12444 , \2559 , \12314 );
nand \U$12198 ( \12445 , \12443 , \12444 );
xor \U$12199 ( \12446 , \12440 , \12445 );
xor \U$12200 ( \12447 , \12434 , \12446 );
xor \U$12201 ( \12448 , \12424 , \12447 );
not \U$12202 ( \12449 , \11149 );
not \U$12203 ( \12450 , \2639 );
or \U$12204 ( \12451 , \12449 , \12450 );
xor \U$12205 ( \12452 , RIbe28390_19, RIbe291a0_49);
nand \U$12206 ( \12453 , \2647 , \12452 );
nand \U$12207 ( \12454 , \12451 , \12453 );
not \U$12208 ( \12455 , \12454 );
not \U$12209 ( \12456 , \11918 );
not \U$12210 ( \12457 , \879 );
or \U$12211 ( \12458 , \12456 , \12457 );
xor \U$12212 ( \12459 , RIbe29998_66, RIbe28228_16);
nand \U$12213 ( \12460 , \885 , \12459 );
nand \U$12214 ( \12461 , \12458 , \12460 );
not \U$12215 ( \12462 , \12461 );
not \U$12216 ( \12463 , \12462 );
or \U$12217 ( \12464 , \12455 , \12463 );
not \U$12218 ( \12465 , \12454 );
nand \U$12219 ( \12466 , \12465 , \12461 );
nand \U$12220 ( \12467 , \12464 , \12466 );
not \U$12221 ( \12468 , \12467 );
not \U$12222 ( \12469 , \11874 );
not \U$12223 ( \12470 , \2459 );
or \U$12224 ( \12471 , \12469 , \12470 );
xor \U$12225 ( \12472 , RIbe27e68_8, RIbe29470_55);
nand \U$12226 ( \12473 , \2464 , \12472 );
nand \U$12227 ( \12474 , \12471 , \12473 );
not \U$12228 ( \12475 , \12474 );
not \U$12229 ( \12476 , \12475 );
or \U$12230 ( \12477 , \12468 , \12476 );
or \U$12231 ( \12478 , \12475 , \12467 );
nand \U$12232 ( \12479 , \12477 , \12478 );
xor \U$12233 ( \12480 , \12448 , \12479 );
xor \U$12234 ( \12481 , \12406 , \12480 );
not \U$12235 ( \12482 , \11106 );
not \U$12237 ( \12483 , \11136 );
and \U$12238 ( \12484 , \12483 , \11161 );
nor \U$12239 ( \12485 , 1'b0 , \12484 );
not \U$12240 ( \12486 , \12485 );
or \U$12241 ( \12487 , \12482 , \12486 );
not \U$12242 ( \12488 , \11161 );
nand \U$12243 ( \12489 , \12488 , \11136 );
nand \U$12244 ( \12490 , \12487 , \12489 );
xor \U$12245 ( \12491 , \12481 , \12490 );
not \U$12246 ( \12492 , \12491 );
not \U$12247 ( \12493 , \11996 );
not \U$12248 ( \12494 , \12065 );
or \U$12249 ( \12495 , \12493 , \12494 );
nand \U$12250 ( \12496 , \12495 , \11995 );
not \U$12251 ( \12497 , \12496 );
not \U$12252 ( \12498 , \12379 );
nand \U$12253 ( \12499 , \12498 , \12381 );
not \U$12254 ( \12500 , \12364 );
and \U$12255 ( \12501 , \12499 , \12500 );
not \U$12256 ( \12502 , \12499 );
and \U$12257 ( \12503 , \12502 , \12364 );
nor \U$12258 ( \12504 , \12501 , \12503 );
not \U$12259 ( \12505 , \12504 );
or \U$12260 ( \12506 , \12497 , \12505 );
or \U$12261 ( \12507 , \12504 , \12496 );
nand \U$12262 ( \12508 , \12506 , \12507 );
not \U$12263 ( \12509 , \12508 );
or \U$12264 ( \12510 , \12492 , \12509 );
not \U$12265 ( \12511 , \12504 );
nand \U$12266 ( \12512 , \12511 , \12496 );
nand \U$12267 ( \12513 , \12510 , \12512 );
xor \U$12268 ( \12514 , \12388 , \12513 );
not \U$12269 ( \12515 , \11500 );
not \U$12270 ( \12516 , \11531 );
or \U$12271 ( \12517 , \12515 , \12516 );
or \U$12272 ( \12518 , \11531 , \11500 );
nand \U$12273 ( \12519 , \12518 , \11476 );
nand \U$12274 ( \12520 , \12517 , \12519 );
xor \U$12275 ( \12521 , \12424 , \12447 );
and \U$12276 ( \12522 , \12521 , \12479 );
and \U$12277 ( \12523 , \12424 , \12447 );
or \U$12278 ( \12524 , \12522 , \12523 );
xor \U$12279 ( \12525 , \12520 , \12524 );
not \U$12280 ( \12526 , \12474 );
not \U$12281 ( \12527 , \12467 );
or \U$12282 ( \12528 , \12526 , \12527 );
nand \U$12283 ( \12529 , \12461 , \12454 );
nand \U$12284 ( \12530 , \12528 , \12529 );
not \U$12285 ( \12531 , \12434 );
not \U$12286 ( \12532 , \12446 );
or \U$12287 ( \12533 , \12531 , \12532 );
nand \U$12288 ( \12534 , \12445 , \12440 );
nand \U$12289 ( \12535 , \12533 , \12534 );
xor \U$12290 ( \12536 , \12530 , \12535 );
not \U$12291 ( \12537 , \11548 );
not \U$12292 ( \12538 , \11566 );
or \U$12293 ( \12539 , \12537 , \12538 );
nand \U$12294 ( \12540 , \11554 , \11561 );
nand \U$12295 ( \12541 , \12539 , \12540 );
and \U$12296 ( \12542 , \12536 , \12541 );
not \U$12297 ( \12543 , \12536 );
not \U$12298 ( \12544 , \12541 );
and \U$12299 ( \12545 , \12543 , \12544 );
nor \U$12300 ( \12546 , \12542 , \12545 );
xor \U$12301 ( \12547 , \12525 , \12546 );
xor \U$12302 ( \12548 , \12406 , \12480 );
and \U$12303 ( \12549 , \12548 , \12490 );
and \U$12304 ( \12550 , \12406 , \12480 );
or \U$12305 ( \12551 , \12549 , \12550 );
xor \U$12306 ( \12552 , \12547 , \12551 );
not \U$12307 ( \12553 , \12408 );
not \U$12308 ( \12554 , \2518 );
or \U$12309 ( \12555 , \12553 , \12554 );
nand \U$12310 ( \12556 , \3074 , \9777 );
nand \U$12311 ( \12557 , \12555 , \12556 );
not \U$12312 ( \12558 , \12438 );
not \U$12313 ( \12559 , \2730 );
or \U$12314 ( \12560 , \12558 , \12559 );
nand \U$12315 ( \12561 , \398 , \9808 );
nand \U$12316 ( \12562 , \12560 , \12561 );
xor \U$12317 ( \12563 , \12557 , \12562 );
not \U$12318 ( \12564 , \12417 );
not \U$12319 ( \12565 , \332 );
or \U$12320 ( \12566 , \12564 , \12565 );
nand \U$12321 ( \12567 , \347 , \9767 );
nand \U$12322 ( \12568 , \12566 , \12567 );
xnor \U$12323 ( \12569 , \12563 , \12568 );
not \U$12324 ( \12570 , \11552 );
not \U$12325 ( \12571 , \1053 );
or \U$12326 ( \12572 , \12570 , \12571 );
nand \U$12327 ( \12573 , \1263 , \9272 );
nand \U$12328 ( \12574 , \12572 , \12573 );
not \U$12329 ( \12575 , \11473 );
not \U$12330 ( \12576 , \2276 );
or \U$12331 ( \12577 , \12575 , \12576 );
nand \U$12332 ( \12578 , \5055 , \9749 );
nand \U$12333 ( \12579 , \12577 , \12578 );
xor \U$12334 ( \12580 , \12574 , \12579 );
not \U$12335 ( \12581 , \12432 );
not \U$12336 ( \12582 , \4578 );
or \U$12337 ( \12583 , \12581 , \12582 );
nand \U$12338 ( \12584 , \7642 , \9309 );
nand \U$12339 ( \12585 , \12583 , \12584 );
xor \U$12340 ( \12586 , \12580 , \12585 );
xnor \U$12341 ( \12587 , \12569 , \12586 );
and \U$12342 ( \12588 , RIbe2b2e8_120, RIbe27b98_2);
not \U$12343 ( \12589 , \11538 );
not \U$12344 ( \12590 , \8807 );
not \U$12345 ( \12591 , \12590 );
or \U$12346 ( \12592 , \12589 , \12591 );
nand \U$12347 ( \12593 , \10476 , \9260 );
nand \U$12348 ( \12594 , \12592 , \12593 );
xor \U$12349 ( \12595 , \12588 , \12594 );
not \U$12350 ( \12596 , \12472 );
not \U$12351 ( \12597 , \2459 );
or \U$12352 ( \12598 , \12596 , \12597 );
nand \U$12353 ( \12599 , \4447 , \9233 );
nand \U$12354 ( \12600 , \12598 , \12599 );
xor \U$12355 ( \12601 , \12595 , \12600 );
not \U$12356 ( \12602 , \12601 );
xor \U$12357 ( \12603 , \12587 , \12602 );
not \U$12358 ( \12604 , \12603 );
xor \U$12359 ( \12605 , \12395 , \12398 );
and \U$12360 ( \12606 , \12605 , \12405 );
and \U$12361 ( \12607 , \12395 , \12398 );
or \U$12362 ( \12608 , \12606 , \12607 );
not \U$12363 ( \12609 , \12608 );
not \U$12364 ( \12610 , \11499 );
not \U$12365 ( \12611 , \11492 );
or \U$12366 ( \12612 , \12610 , \12611 );
not \U$12367 ( \12613 , \11488 );
nand \U$12368 ( \12614 , \12613 , \11482 );
nand \U$12369 ( \12615 , \12612 , \12614 );
not \U$12370 ( \12616 , \12411 );
not \U$12371 ( \12617 , \12616 );
not \U$12372 ( \12618 , \12423 );
or \U$12373 ( \12619 , \12617 , \12618 );
not \U$12374 ( \12620 , \12412 );
nand \U$12375 ( \12621 , \12620 , \12419 );
nand \U$12376 ( \12622 , \12619 , \12621 );
xor \U$12377 ( \12623 , \12615 , \12622 );
xor \U$12378 ( \12624 , \11459 , \11467 );
and \U$12379 ( \12625 , \12624 , \11475 );
and \U$12380 ( \12626 , \11459 , \11467 );
or \U$12381 ( \12627 , \12625 , \12626 );
xnor \U$12382 ( \12628 , \12623 , \12627 );
not \U$12383 ( \12629 , \12628 );
or \U$12384 ( \12630 , \12609 , \12629 );
or \U$12385 ( \12631 , \12628 , \12608 );
nand \U$12386 ( \12632 , \12630 , \12631 );
not \U$12387 ( \12633 , \12632 );
or \U$12388 ( \12634 , \12604 , \12633 );
or \U$12389 ( \12635 , \12632 , \12603 );
nand \U$12390 ( \12636 , \12634 , \12635 );
xor \U$12391 ( \12637 , \12552 , \12636 );
xor \U$12392 ( \12638 , \12514 , \12637 );
and \U$12393 ( \12639 , \12254 , \12638 );
not \U$12394 ( \12640 , \12254 );
not \U$12395 ( \12641 , \12638 );
and \U$12396 ( \12642 , \12640 , \12641 );
nor \U$12397 ( \12643 , \12639 , \12642 );
not \U$12398 ( \12644 , \12097 );
not \U$12399 ( \12645 , \12152 );
not \U$12400 ( \12646 , \12645 );
or \U$12401 ( \12647 , \12644 , \12646 );
not \U$12402 ( \12648 , \12148 );
nand \U$12403 ( \12649 , \12648 , \12118 );
nand \U$12404 ( \12650 , \12647 , \12649 );
not \U$12405 ( \12651 , \12650 );
not \U$12406 ( \12652 , \12274 );
nand \U$12407 ( \12653 , \12652 , \12282 );
and \U$12408 ( \12654 , \12653 , \12279 );
not \U$12409 ( \12655 , \12653 );
and \U$12410 ( \12656 , \12655 , \12280 );
nor \U$12411 ( \12657 , \12654 , \12656 );
not \U$12412 ( \12658 , \11740 );
nand \U$12413 ( \12659 , \12658 , \11745 );
not \U$12414 ( \12660 , \12659 );
not \U$12415 ( \12661 , \11810 );
or \U$12416 ( \12662 , \12660 , \12661 );
nand \U$12417 ( \12663 , \11740 , \11744 );
nand \U$12418 ( \12664 , \12662 , \12663 );
not \U$12419 ( \12665 , \12664 );
nand \U$12420 ( \12666 , \12657 , \12665 );
not \U$12421 ( \12667 , \12666 );
or \U$12422 ( \12668 , \12651 , \12667 );
not \U$12423 ( \12669 , \12657 );
not \U$12424 ( \12670 , \12665 );
nand \U$12425 ( \12671 , \12669 , \12670 );
nand \U$12426 ( \12672 , \12668 , \12671 );
not \U$12427 ( \12673 , \11684 );
not \U$12428 ( \12674 , \11638 );
or \U$12429 ( \12675 , \12673 , \12674 );
not \U$12430 ( \12676 , \11634 );
nand \U$12431 ( \12677 , \12676 , \11536 );
nand \U$12432 ( \12678 , \12675 , \12677 );
not \U$12433 ( \12679 , \12678 );
not \U$12434 ( \12680 , \12679 );
not \U$12435 ( \12681 , \11567 );
nand \U$12436 ( \12682 , \12681 , \11598 );
not \U$12437 ( \12683 , \12682 );
not \U$12438 ( \12684 , \11633 );
or \U$12439 ( \12685 , \12683 , \12684 );
not \U$12440 ( \12686 , \11598 );
nand \U$12441 ( \12687 , \12686 , \11567 );
nand \U$12442 ( \12688 , \12685 , \12687 );
not \U$12443 ( \12689 , \11597 );
or \U$12444 ( \12690 , \12689 , \11585 );
nand \U$12445 ( \12691 , \12690 , \11587 );
not \U$12446 ( \12692 , \11524 );
not \U$12447 ( \12693 , \8697 );
or \U$12448 ( \12694 , \12692 , \12693 );
nand \U$12449 ( \12695 , \9379 , \9845 );
nand \U$12450 ( \12696 , \12694 , \12695 );
not \U$12451 ( \12697 , \11582 );
not \U$12452 ( \12698 , \8401 );
or \U$12453 ( \12699 , \12697 , \12698 );
xor \U$12454 ( \12700 , RIbe2a028_80, RIbe28840_29);
nand \U$12455 ( \12701 , \8172 , \12700 );
nand \U$12456 ( \12702 , \12699 , \12701 );
xor \U$12457 ( \12703 , \12696 , \12702 );
not \U$12458 ( \12704 , \11480 );
not \U$12459 ( \12705 , \979 );
or \U$12460 ( \12706 , \12704 , \12705 );
nand \U$12461 ( \12707 , \1805 , \9799 );
nand \U$12462 ( \12708 , \12706 , \12707 );
xor \U$12463 ( \12709 , \12703 , \12708 );
nor \U$12464 ( \12710 , \12691 , \12709 );
not \U$12465 ( \12711 , \12710 );
nand \U$12466 ( \12712 , \12709 , \12691 );
nand \U$12467 ( \12713 , \12711 , \12712 );
not \U$12468 ( \12714 , \11457 );
not \U$12469 ( \12715 , \11452 );
buf \U$12470 ( \12716 , \12715 );
not \U$12471 ( \12717 , \12716 );
or \U$12472 ( \12718 , \12714 , \12717 );
nand \U$12473 ( \12719 , \9726 , RIbe2a910_99);
nand \U$12474 ( \12720 , \12718 , \12719 );
not \U$12475 ( \12721 , \3255 );
not \U$12476 ( \12722 , \12721 );
or \U$12477 ( \12723 , \12722 , \11464 );
not \U$12478 ( \12724 , \9742 );
or \U$12479 ( \12725 , \3250 , \12724 );
nand \U$12480 ( \12726 , \12723 , \12725 );
nor \U$12481 ( \12727 , \12720 , \12726 );
not \U$12482 ( \12728 , \12727 );
nand \U$12483 ( \12729 , \12720 , \12726 );
nand \U$12484 ( \12730 , \12728 , \12729 );
not \U$12485 ( \12731 , \315 );
not \U$12486 ( \12732 , \9816 );
or \U$12487 ( \12733 , \12731 , \12732 );
not \U$12488 ( \12734 , \301 );
nand \U$12489 ( \12735 , \12734 , \12332 );
nand \U$12490 ( \12736 , \12733 , \12735 );
and \U$12491 ( \12737 , \12730 , \12736 );
not \U$12492 ( \12738 , \12730 );
and \U$12493 ( \12739 , \1086 , \12332 );
and \U$12494 ( \12740 , \315 , \9816 );
nor \U$12495 ( \12741 , \12739 , \12740 );
and \U$12496 ( \12742 , \12738 , \12741 );
nor \U$12497 ( \12743 , \12737 , \12742 );
not \U$12498 ( \12744 , \12743 );
and \U$12499 ( \12745 , \12713 , \12744 );
not \U$12500 ( \12746 , \12713 );
and \U$12501 ( \12747 , \12746 , \12743 );
nor \U$12502 ( \12748 , \12745 , \12747 );
xor \U$12503 ( \12749 , \12688 , \12748 );
not \U$12504 ( \12750 , \11559 );
not \U$12505 ( \12751 , \2618 );
or \U$12506 ( \12752 , \12750 , \12751 );
nand \U$12507 ( \12753 , \2626 , \9282 );
nand \U$12508 ( \12754 , \12752 , \12753 );
not \U$12509 ( \12755 , \12322 );
not \U$12510 ( \12756 , \256 );
or \U$12511 ( \12757 , \12755 , \12756 );
nand \U$12512 ( \12758 , \1734 , \9831 );
nand \U$12513 ( \12759 , \12757 , \12758 );
xor \U$12514 ( \12760 , \12754 , \12759 );
not \U$12515 ( \12761 , \11595 );
not \U$12516 ( \12762 , \7372 );
or \U$12517 ( \12763 , \12761 , \12762 );
nand \U$12518 ( \12764 , \8245 , \9250 );
nand \U$12519 ( \12765 , \12763 , \12764 );
xor \U$12520 ( \12766 , \12760 , \12765 );
not \U$12521 ( \12767 , \11517 );
not \U$12522 ( \12768 , \1103 );
or \U$12523 ( \12769 , \12767 , \12768 );
nand \U$12524 ( \12770 , \9856 , \1498 );
nand \U$12525 ( \12771 , \12769 , \12770 );
not \U$12526 ( \12772 , \12771 );
not \U$12527 ( \12773 , \12459 );
not \U$12528 ( \12774 , \1061 );
or \U$12529 ( \12775 , \12773 , \12774 );
nand \U$12530 ( \12776 , \885 , \9241 );
nand \U$12531 ( \12777 , \12775 , \12776 );
not \U$12532 ( \12778 , \12777 );
not \U$12533 ( \12779 , \12778 );
or \U$12534 ( \12780 , \12772 , \12779 );
not \U$12535 ( \12781 , \12771 );
nand \U$12536 ( \12782 , \12781 , \12777 );
nand \U$12537 ( \12783 , \12780 , \12782 );
not \U$12538 ( \12784 , \11497 );
not \U$12539 ( \12785 , \1132 );
or \U$12540 ( \12786 , \12784 , \12785 );
nand \U$12541 ( \12787 , \1137 , \9791 );
nand \U$12542 ( \12788 , \12786 , \12787 );
not \U$12543 ( \12789 , \12788 );
and \U$12544 ( \12790 , \12783 , \12789 );
not \U$12545 ( \12791 , \12783 );
and \U$12546 ( \12792 , \12791 , \12788 );
nor \U$12547 ( \12793 , \12790 , \12792 );
not \U$12548 ( \12794 , \12793 );
nand \U$12549 ( \12795 , \12766 , \12794 );
not \U$12550 ( \12796 , \12766 );
nand \U$12551 ( \12797 , \12796 , \12793 );
nand \U$12552 ( \12798 , \12795 , \12797 );
and \U$12553 ( \12799 , \3408 , \12452 );
and \U$12554 ( \12800 , \2777 , \9323 );
nor \U$12555 ( \12801 , \12799 , \12800 );
not \U$12556 ( \12802 , \11510 );
not \U$12557 ( \12803 , \1793 );
or \U$12558 ( \12804 , \12802 , \12803 );
nand \U$12559 ( \12805 , \1797 , \9852 );
nand \U$12560 ( \12806 , \12804 , \12805 );
not \U$12561 ( \12807 , \12328 );
not \U$12562 ( \12808 , \2718 );
not \U$12563 ( \12809 , \12808 );
or \U$12564 ( \12810 , \12807 , \12809 );
nand \U$12565 ( \12811 , \2707 , \9823 );
nand \U$12566 ( \12812 , \12810 , \12811 );
nor \U$12567 ( \12813 , \12806 , \12812 );
not \U$12568 ( \12814 , \12813 );
nand \U$12569 ( \12815 , \12812 , \12806 );
nand \U$12570 ( \12816 , \12814 , \12815 );
xor \U$12571 ( \12817 , \12801 , \12816 );
xor \U$12572 ( \12818 , \12798 , \12817 );
xnor \U$12573 ( \12819 , \12749 , \12818 );
not \U$12574 ( \12820 , \12819 );
not \U$12575 ( \12821 , \12820 );
or \U$12576 ( \12822 , \12680 , \12821 );
nand \U$12577 ( \12823 , \12819 , \12678 );
nand \U$12578 ( \12824 , \12822 , \12823 );
not \U$12579 ( \12825 , \12824 );
xor \U$12580 ( \12826 , \12672 , \12825 );
not \U$12581 ( \12827 , \11689 );
and \U$12582 ( \12828 , \11827 , \11819 );
not \U$12583 ( \12829 , \11827 );
and \U$12584 ( \12830 , \12829 , \11818 );
nor \U$12585 ( \12831 , \12828 , \12830 );
not \U$12586 ( \12832 , \12831 );
or \U$12587 ( \12833 , \12827 , \12832 );
nand \U$12588 ( \12834 , \11826 , \11818 );
nand \U$12589 ( \12835 , \12833 , \12834 );
not \U$12590 ( \12836 , \12835 );
xor \U$12591 ( \12837 , \12826 , \12836 );
not \U$12592 ( \12838 , \12183 );
not \U$12593 ( \12839 , \12070 );
or \U$12594 ( \12840 , \12838 , \12839 );
nand \U$12595 ( \12841 , \12156 , \12177 );
nand \U$12596 ( \12842 , \12840 , \12841 );
not \U$12597 ( \12843 , \12842 );
buf \U$12598 ( \12844 , \12508 );
not \U$12599 ( \12845 , \12491 );
and \U$12600 ( \12846 , \12844 , \12845 );
not \U$12601 ( \12847 , \12844 );
and \U$12602 ( \12848 , \12847 , \12491 );
nor \U$12603 ( \12849 , \12846 , \12848 );
and \U$12604 ( \12850 , \12669 , \12665 );
not \U$12605 ( \12851 , \12669 );
and \U$12606 ( \12852 , \12851 , \12670 );
nor \U$12607 ( \12853 , \12850 , \12852 );
and \U$12608 ( \12854 , \12853 , \12650 );
not \U$12609 ( \12855 , \12853 );
not \U$12610 ( \12856 , \12650 );
and \U$12611 ( \12857 , \12855 , \12856 );
nor \U$12612 ( \12858 , \12854 , \12857 );
nand \U$12613 ( \12859 , \12849 , \12858 );
not \U$12614 ( \12860 , \12859 );
or \U$12615 ( \12861 , \12843 , \12860 );
not \U$12616 ( \12862 , \12849 );
not \U$12617 ( \12863 , \12858 );
nand \U$12618 ( \12864 , \12862 , \12863 );
nand \U$12619 ( \12865 , \12861 , \12864 );
not \U$12620 ( \12866 , \12865 );
xor \U$12621 ( \12867 , \12837 , \12866 );
nand \U$12622 ( \12868 , \12643 , \12867 );
not \U$12623 ( \12869 , \12254 );
nand \U$12624 ( \12870 , \12869 , \12641 );
nand \U$12625 ( \12871 , \12868 , \12870 );
not \U$12626 ( \12872 , \12355 );
not \U$12627 ( \12873 , \12313 );
or \U$12628 ( \12874 , \12872 , \12873 );
nand \U$12629 ( \12875 , \12312 , \12287 );
nand \U$12630 ( \12876 , \12874 , \12875 );
not \U$12631 ( \12877 , \12876 );
not \U$12632 ( \12878 , \12700 );
not \U$12633 ( \12879 , \9530 );
or \U$12634 ( \12880 , \12878 , \12879 );
nand \U$12635 ( \12881 , \9065 , \9061 );
nand \U$12636 ( \12882 , \12880 , \12881 );
not \U$12637 ( \12883 , \12882 );
not \U$12638 ( \12884 , \12319 );
not \U$12639 ( \12885 , \12884 );
or \U$12640 ( \12886 , \12883 , \12885 );
or \U$12641 ( \12887 , \12884 , \12882 );
nand \U$12642 ( \12888 , \12886 , \12887 );
or \U$12643 ( \12889 , \12562 , \12557 );
nand \U$12644 ( \12890 , \12889 , \12568 );
nand \U$12645 ( \12891 , \12562 , \12557 );
nand \U$12646 ( \12892 , \12890 , \12891 );
xor \U$12647 ( \12893 , \12888 , \12892 );
not \U$12648 ( \12894 , \12350 );
not \U$12649 ( \12895 , \12344 );
or \U$12650 ( \12896 , \12894 , \12895 );
nand \U$12651 ( \12897 , \12340 , \12884 );
nand \U$12652 ( \12898 , \12896 , \12897 );
and \U$12653 ( \12899 , \12893 , \12898 );
not \U$12654 ( \12900 , \12893 );
not \U$12655 ( \12901 , \12898 );
and \U$12656 ( \12902 , \12900 , \12901 );
nor \U$12657 ( \12903 , \12899 , \12902 );
not \U$12658 ( \12904 , \12541 );
not \U$12659 ( \12905 , \12536 );
or \U$12660 ( \12906 , \12904 , \12905 );
nand \U$12661 ( \12907 , \12535 , \12530 );
nand \U$12662 ( \12908 , \12906 , \12907 );
xor \U$12663 ( \12909 , \12903 , \12908 );
not \U$12664 ( \12910 , \12909 );
not \U$12665 ( \12911 , \12910 );
or \U$12666 ( \12912 , \12877 , \12911 );
not \U$12667 ( \12913 , \12876 );
nand \U$12668 ( \12914 , \12913 , \12909 );
nand \U$12669 ( \12915 , \12912 , \12914 );
not \U$12670 ( \12916 , \12546 );
not \U$12671 ( \12917 , \12524 );
not \U$12672 ( \12918 , \12520 );
nand \U$12673 ( \12919 , \12917 , \12918 );
not \U$12674 ( \12920 , \12919 );
or \U$12675 ( \12921 , \12916 , \12920 );
or \U$12676 ( \12922 , \12918 , \12917 );
nand \U$12677 ( \12923 , \12921 , \12922 );
xnor \U$12678 ( \12924 , \12915 , \12923 );
not \U$12679 ( \12925 , \12924 );
xor \U$12680 ( \12926 , \12547 , \12551 );
and \U$12681 ( \12927 , \12926 , \12636 );
and \U$12682 ( \12928 , \12547 , \12551 );
or \U$12683 ( \12929 , \12927 , \12928 );
not \U$12684 ( \12930 , \12929 );
or \U$12685 ( \12931 , \12925 , \12930 );
or \U$12686 ( \12932 , \12924 , \12929 );
nand \U$12687 ( \12933 , \12931 , \12932 );
buf \U$12688 ( \12934 , \12933 );
xor \U$12689 ( \12935 , \12588 , \12594 );
and \U$12690 ( \12936 , \12935 , \12600 );
and \U$12691 ( \12937 , \12588 , \12594 );
or \U$12692 ( \12938 , \12936 , \12937 );
and \U$12693 ( \12939 , \9829 , \9838 );
not \U$12694 ( \12940 , \9829 );
and \U$12695 ( \12941 , \12940 , \9837 );
or \U$12696 ( \12942 , \12939 , \12941 );
xor \U$12697 ( \12943 , \12942 , \9821 );
xor \U$12698 ( \12944 , \12938 , \12943 );
xor \U$12699 ( \12945 , \9239 , \9257 );
xor \U$12700 ( \12946 , \12945 , \9246 );
xor \U$12701 ( \12947 , \12944 , \12946 );
or \U$12702 ( \12948 , \12813 , \12801 );
nand \U$12703 ( \12949 , \12948 , \12815 );
xor \U$12704 ( \12950 , \12696 , \12702 );
and \U$12705 ( \12951 , \12950 , \12708 );
and \U$12706 ( \12952 , \12696 , \12702 );
or \U$12707 ( \12953 , \12951 , \12952 );
xor \U$12708 ( \12954 , \12949 , \12953 );
not \U$12709 ( \12955 , \12788 );
not \U$12710 ( \12956 , \12783 );
or \U$12711 ( \12957 , \12955 , \12956 );
nand \U$12712 ( \12958 , \12777 , \12771 );
nand \U$12713 ( \12959 , \12957 , \12958 );
xor \U$12714 ( \12960 , \12954 , \12959 );
xor \U$12715 ( \12961 , \12947 , \12960 );
or \U$12716 ( \12962 , \12727 , \12741 );
nand \U$12717 ( \12963 , \12962 , \12729 );
xor \U$12718 ( \12964 , \12574 , \12579 );
and \U$12719 ( \12965 , \12964 , \12585 );
and \U$12720 ( \12966 , \12574 , \12579 );
or \U$12721 ( \12967 , \12965 , \12966 );
and \U$12722 ( \12968 , \12963 , \12967 );
not \U$12723 ( \12969 , \12963 );
not \U$12724 ( \12970 , \12967 );
and \U$12725 ( \12971 , \12969 , \12970 );
nor \U$12726 ( \12972 , \12968 , \12971 );
xor \U$12727 ( \12973 , \12754 , \12759 );
and \U$12728 ( \12974 , \12973 , \12765 );
and \U$12729 ( \12975 , \12754 , \12759 );
or \U$12730 ( \12976 , \12974 , \12975 );
xor \U$12731 ( \12977 , \12972 , \12976 );
xor \U$12732 ( \12978 , \12961 , \12977 );
not \U$12733 ( \12979 , \12797 );
not \U$12734 ( \12980 , \12817 );
or \U$12735 ( \12981 , \12979 , \12980 );
nand \U$12736 ( \12982 , \12981 , \12795 );
not \U$12737 ( \12983 , \12601 );
not \U$12738 ( \12984 , \12587 );
or \U$12739 ( \12985 , \12983 , \12984 );
not \U$12740 ( \12986 , \12569 );
nand \U$12741 ( \12987 , \12986 , \12586 );
nand \U$12742 ( \12988 , \12985 , \12987 );
not \U$12743 ( \12989 , \12627 );
not \U$12744 ( \12990 , \12623 );
or \U$12745 ( \12991 , \12989 , \12990 );
nand \U$12746 ( \12992 , \12622 , \12615 );
nand \U$12747 ( \12993 , \12991 , \12992 );
xor \U$12748 ( \12994 , \12988 , \12993 );
xor \U$12749 ( \12995 , \12982 , \12994 );
xor \U$12750 ( \12996 , \12978 , \12995 );
not \U$12751 ( \12997 , \12603 );
not \U$12752 ( \12998 , \12997 );
not \U$12753 ( \12999 , \12632 );
or \U$12754 ( \13000 , \12998 , \12999 );
not \U$12755 ( \13001 , \12628 );
nand \U$12756 ( \13002 , \13001 , \12608 );
nand \U$12757 ( \13003 , \13000 , \13002 );
not \U$12758 ( \13004 , \13003 );
xnor \U$12759 ( \13005 , \12996 , \13004 );
not \U$12760 ( \13006 , \13005 );
and \U$12761 ( \13007 , \12934 , \13006 );
not \U$12762 ( \13008 , \12934 );
and \U$12763 ( \13009 , \13008 , \13005 );
nor \U$12764 ( \13010 , \13007 , \13009 );
not \U$12765 ( \13011 , \12820 );
not \U$12766 ( \13012 , \12678 );
or \U$12767 ( \13013 , \13011 , \13012 );
not \U$12768 ( \13014 , \12819 );
not \U$12769 ( \13015 , \12679 );
or \U$12770 ( \13016 , \13014 , \13015 );
nand \U$12771 ( \13017 , \13016 , \12672 );
nand \U$12772 ( \13018 , \13013 , \13017 );
not \U$12773 ( \13019 , \12748 );
nand \U$12774 ( \13020 , \13019 , \12688 );
and \U$12775 ( \13021 , \13020 , \12818 );
nor \U$12776 ( \13022 , \13019 , \12688 );
nor \U$12777 ( \13023 , \13021 , \13022 );
buf \U$12778 ( \13024 , \12710 );
or \U$12779 ( \13025 , \13024 , \12743 );
nand \U$12780 ( \13026 , \13025 , \12712 );
xor \U$12781 ( \13027 , \9797 , \9804 );
xor \U$12782 ( \13028 , \13027 , \9813 );
xor \U$12783 ( \13029 , \9775 , \9782 );
not \U$12784 ( \13030 , \13029 );
xor \U$12785 ( \13031 , \13028 , \13030 );
not \U$12786 ( \13032 , \9326 );
not \U$12787 ( \13033 , \9317 );
or \U$12788 ( \13034 , \13032 , \13033 );
or \U$12789 ( \13035 , \9317 , \9326 );
nand \U$12790 ( \13036 , \13034 , \13035 );
xor \U$12791 ( \13037 , \13031 , \13036 );
xor \U$12792 ( \13038 , \13026 , \13037 );
xor \U$12793 ( \13039 , \9867 , \9850 );
xor \U$12794 ( \13040 , \9292 , \9270 );
xor \U$12795 ( \13041 , \13039 , \13040 );
xnor \U$12796 ( \13042 , \9759 , \9740 );
xnor \U$12797 ( \13043 , \13041 , \13042 );
xor \U$12798 ( \13044 , \13038 , \13043 );
xor \U$12799 ( \13045 , \13023 , \13044 );
not \U$12800 ( \13046 , \12361 );
not \U$12801 ( \13047 , \12382 );
or \U$12802 ( \13048 , \13046 , \13047 );
not \U$12803 ( \13049 , \12360 );
not \U$12804 ( \13050 , \12383 );
or \U$12805 ( \13051 , \13049 , \13050 );
nand \U$12806 ( \13052 , \13051 , \12283 );
nand \U$12807 ( \13053 , \13048 , \13052 );
xor \U$12808 ( \13054 , \13045 , \13053 );
xor \U$12809 ( \13055 , \13018 , \13054 );
xor \U$12810 ( \13056 , \12388 , \12513 );
and \U$12811 ( \13057 , \13056 , \12637 );
and \U$12812 ( \13058 , \12388 , \12513 );
or \U$12813 ( \13059 , \13057 , \13058 );
and \U$12814 ( \13060 , \13055 , \13059 );
not \U$12815 ( \13061 , \13055 );
not \U$12816 ( \13062 , \13059 );
and \U$12817 ( \13063 , \13061 , \13062 );
or \U$12818 ( \13064 , \13060 , \13063 );
xor \U$12819 ( \13065 , \13010 , \13064 );
xor \U$12820 ( \13066 , \12826 , \12836 );
and \U$12821 ( \13067 , \13066 , \12866 );
and \U$12822 ( \13068 , \12826 , \12836 );
or \U$12823 ( \13069 , \13067 , \13068 );
xor \U$12824 ( \13070 , \13065 , \13069 );
nand \U$12825 ( \13071 , \12871 , \13070 );
not \U$12826 ( \13072 , \13071 );
xnor \U$12827 ( \13073 , \12867 , \12643 );
not \U$12828 ( \13074 , \12849 );
xor \U$12829 ( \13075 , \12863 , \13074 );
xnor \U$12830 ( \13076 , \13075 , \12842 );
not \U$12831 ( \13077 , \13076 );
not \U$12832 ( \13078 , \11828 );
not \U$12833 ( \13079 , \11448 );
or \U$12834 ( \13080 , \13078 , \13079 );
nand \U$12835 ( \13081 , \11829 , \11447 );
nand \U$12836 ( \13082 , \13080 , \13081 );
buf \U$12837 ( \13083 , \12250 );
not \U$12838 ( \13084 , \13083 );
and \U$12839 ( \13085 , \13082 , \13084 );
not \U$12840 ( \13086 , \13082 );
and \U$12841 ( \13087 , \13086 , \13083 );
nor \U$12842 ( \13088 , \13085 , \13087 );
not \U$12843 ( \13089 , \13088 );
or \U$12844 ( \13090 , \13077 , \13089 );
xnor \U$12845 ( \13091 , \11443 , \11028 );
not \U$12846 ( \13092 , \13091 );
not \U$12847 ( \13093 , \13092 );
xor \U$12848 ( \13094 , \10804 , \10895 );
not \U$12849 ( \13095 , \13094 );
not \U$12850 ( \13096 , \11257 );
not \U$12851 ( \13097 , \13096 );
buf \U$12852 ( \13098 , \11390 );
not \U$12853 ( \13099 , \13098 );
or \U$12854 ( \13100 , \13097 , \13099 );
or \U$12855 ( \13101 , \13098 , \13096 );
nand \U$12856 ( \13102 , \13100 , \13101 );
and \U$12857 ( \13103 , \10711 , \10643 );
not \U$12858 ( \13104 , \10711 );
not \U$12859 ( \13105 , \10643 );
and \U$12860 ( \13106 , \13104 , \13105 );
nor \U$12861 ( \13107 , \13103 , \13106 );
not \U$12862 ( \13108 , \13107 );
xor \U$12863 ( \13109 , \11296 , \11303 );
not \U$12864 ( \13110 , \13109 );
not \U$12865 ( \13111 , \9263 );
xor \U$12866 ( \13112 , RIbe28c78_38, RIbe2a3e8_88);
not \U$12867 ( \13113 , \13112 );
or \U$12868 ( \13114 , \13111 , \13113 );
nand \U$12869 ( \13115 , \9268 , \11358 );
nand \U$12870 ( \13116 , \13114 , \13115 );
buf \U$12871 ( \13117 , \13116 );
not \U$12872 ( \13118 , \13117 );
xor \U$12873 ( \13119 , RIbe285e8_24, RIbe29a10_67);
not \U$12874 ( \13120 , \13119 );
not \U$12875 ( \13121 , \7618 );
or \U$12876 ( \13122 , \13120 , \13121 );
nand \U$12877 ( \13123 , \8270 , \11172 );
nand \U$12878 ( \13124 , \13122 , \13123 );
not \U$12879 ( \13125 , \13124 );
or \U$12880 ( \13126 , \13118 , \13125 );
or \U$12881 ( \13127 , \13124 , \13117 );
xor \U$12882 ( \13128 , RIbe2b6a8_128, RIbe280c0_13);
not \U$12883 ( \13129 , \13128 );
not \U$12884 ( \13130 , \1053 );
or \U$12885 ( \13131 , \13129 , \13130 );
nand \U$12886 ( \13132 , \869 , \11189 );
nand \U$12887 ( \13133 , \13131 , \13132 );
nand \U$12888 ( \13134 , \13127 , \13133 );
nand \U$12889 ( \13135 , \13126 , \13134 );
not \U$12890 ( \13136 , \13135 );
buf \U$12891 ( \13137 , \11332 );
not \U$12892 ( \13138 , \11317 );
and \U$12893 ( \13139 , \13137 , \13138 );
not \U$12894 ( \13140 , \13137 );
and \U$12895 ( \13141 , \13140 , \11317 );
nor \U$12896 ( \13142 , \13139 , \13141 );
not \U$12897 ( \13143 , \13142 );
or \U$12898 ( \13144 , \13136 , \13143 );
or \U$12899 ( \13145 , \13135 , \13142 );
nand \U$12900 ( \13146 , \13144 , \13145 );
not \U$12901 ( \13147 , \13146 );
or \U$12902 ( \13148 , \13110 , \13147 );
not \U$12903 ( \13149 , \13142 );
nand \U$12904 ( \13150 , \13149 , \13135 );
nand \U$12905 ( \13151 , \13148 , \13150 );
not \U$12906 ( \13152 , \13151 );
or \U$12907 ( \13153 , \13108 , \13152 );
or \U$12908 ( \13154 , \13151 , \13107 );
xor \U$12909 ( \13155 , \10679 , \10699 );
not \U$12910 ( \13156 , \10707 );
xor \U$12911 ( \13157 , \13155 , \13156 );
xor \U$12912 ( \13158 , \11185 , \11178 );
not \U$12913 ( \13159 , \13158 );
xor \U$12914 ( \13160 , \11194 , \13159 );
nand \U$12915 ( \13161 , \13157 , \13160 );
not \U$12916 ( \13162 , \13161 );
xor \U$12917 ( \13163 , \11249 , \11230 );
not \U$12918 ( \13164 , \13163 );
or \U$12919 ( \13165 , \13162 , \13164 );
not \U$12920 ( \13166 , \13157 );
not \U$12921 ( \13167 , \13160 );
nand \U$12922 ( \13168 , \13166 , \13167 );
nand \U$12923 ( \13169 , \13165 , \13168 );
nand \U$12924 ( \13170 , \13154 , \13169 );
nand \U$12925 ( \13171 , \13153 , \13170 );
xor \U$12926 ( \13172 , \13102 , \13171 );
not \U$12927 ( \13173 , \13172 );
or \U$12928 ( \13174 , \13095 , \13173 );
nand \U$12929 ( \13175 , \13171 , \13102 );
nand \U$12930 ( \13176 , \13174 , \13175 );
not \U$12931 ( \13177 , \13176 );
xor \U$12932 ( \13178 , \10983 , \10991 );
xor \U$12933 ( \13179 , \13178 , \11000 );
not \U$12934 ( \13180 , \13179 );
not \U$12935 ( \13181 , \10943 );
and \U$12936 ( \13182 , \10958 , \13181 );
not \U$12937 ( \13183 , \10958 );
and \U$12938 ( \13184 , \13183 , \10943 );
nor \U$12939 ( \13185 , \13182 , \13184 );
not \U$12940 ( \13186 , \13185 );
not \U$12941 ( \13187 , \13186 );
or \U$12942 ( \13188 , \13180 , \13187 );
not \U$12943 ( \13189 , \13179 );
not \U$12944 ( \13190 , \13189 );
not \U$12945 ( \13191 , \13185 );
or \U$12946 ( \13192 , \13190 , \13191 );
and \U$12947 ( \13193 , \11384 , \11356 );
buf \U$12948 ( \13194 , \11381 );
xor \U$12949 ( \13195 , \13193 , \13194 );
nand \U$12950 ( \13196 , \13192 , \13195 );
nand \U$12951 ( \13197 , \13188 , \13196 );
xor \U$12952 ( \13198 , \11272 , \11265 );
xnor \U$12953 ( \13199 , \13198 , \11281 );
not \U$12954 ( \13200 , \13199 );
xor \U$12955 ( \13201 , \11363 , \11370 );
buf \U$12956 ( \13202 , \11378 );
not \U$12957 ( \13203 , \13202 );
and \U$12958 ( \13204 , \13201 , \13203 );
not \U$12959 ( \13205 , \13201 );
and \U$12960 ( \13206 , \13205 , \13202 );
nor \U$12961 ( \13207 , \13204 , \13206 );
not \U$12962 ( \13208 , \13207 );
or \U$12963 ( \13209 , \13200 , \13208 );
not \U$12964 ( \13210 , \10669 );
not \U$12965 ( \13211 , \13210 );
xor \U$12966 ( \13212 , \10659 , \10651 );
not \U$12967 ( \13213 , \13212 );
or \U$12968 ( \13214 , \13211 , \13213 );
or \U$12969 ( \13215 , \13212 , \13210 );
nand \U$12970 ( \13216 , \13214 , \13215 );
nand \U$12971 ( \13217 , \13209 , \13216 );
not \U$12972 ( \13218 , \13207 );
not \U$12973 ( \13219 , \13199 );
nand \U$12974 ( \13220 , \13218 , \13219 );
nand \U$12975 ( \13221 , \13217 , \13220 );
xor \U$12976 ( \13222 , \11196 , \11221 );
xor \U$12977 ( \13223 , \13222 , \11254 );
nor \U$12978 ( \13224 , \13221 , \13223 );
xor \U$12979 ( \13225 , \11308 , \11283 );
not \U$12980 ( \13226 , \11336 );
and \U$12981 ( \13227 , \13225 , \13226 );
not \U$12982 ( \13228 , \13225 );
and \U$12983 ( \13229 , \13228 , \11336 );
nor \U$12984 ( \13230 , \13227 , \13229 );
or \U$12985 ( \13231 , \13224 , \13230 );
not \U$12986 ( \13232 , \13217 );
not \U$12987 ( \13233 , \13220 );
or \U$12988 ( \13234 , \13232 , \13233 );
nand \U$12989 ( \13235 , \13234 , \13223 );
nand \U$12990 ( \13236 , \13231 , \13235 );
xor \U$12991 ( \13237 , \13197 , \13236 );
xor \U$12992 ( \13238 , RIbe290b0_47, RIbe2a0a0_81);
not \U$12993 ( \13239 , \13238 );
not \U$12994 ( \13240 , \523 );
or \U$12995 ( \13241 , \13239 , \13240 );
nand \U$12996 ( \13242 , \10730 , \11326 );
nand \U$12997 ( \13243 , \13241 , \13242 );
not \U$12998 ( \13244 , \13243 );
xor \U$12999 ( \13245 , RIbe28b88_36, RIbe298a8_64);
not \U$13000 ( \13246 , \13245 );
not \U$13001 ( \13247 , \9052 );
or \U$13002 ( \13248 , \13246 , \13247 );
not \U$13003 ( \13249 , \7549 );
not \U$13004 ( \13250 , \13249 );
nand \U$13005 ( \13251 , \13250 , \11267 );
nand \U$13006 ( \13252 , \13248 , \13251 );
not \U$13007 ( \13253 , \13252 );
nand \U$13008 ( \13254 , \13244 , \13253 );
not \U$13009 ( \13255 , \13254 );
xor \U$13010 ( \13256 , RIbe282a0_17, RIbe29c68_72);
not \U$13011 ( \13257 , \13256 );
not \U$13012 ( \13258 , \8595 );
or \U$13013 ( \13259 , \13257 , \13258 );
nand \U$13014 ( \13260 , \4580 , \11232 );
nand \U$13015 ( \13261 , \13259 , \13260 );
not \U$13016 ( \13262 , \13261 );
or \U$13017 ( \13263 , \13255 , \13262 );
nand \U$13018 ( \13264 , \13252 , \13243 );
nand \U$13019 ( \13265 , \13263 , \13264 );
xor \U$13020 ( \13266 , RIbe2a280_85, RIbe28048_12);
not \U$13021 ( \13267 , \13266 );
not \U$13022 ( \13268 , \11344 );
not \U$13023 ( \13269 , \13268 );
or \U$13024 ( \13270 , \13267 , \13269 );
nand \U$13025 ( \13271 , \10849 , \11340 );
nand \U$13026 ( \13272 , \13270 , \13271 );
not \U$13027 ( \13273 , \13272 );
not \U$13028 ( \13274 , \10689 );
xnor \U$13029 ( \13275 , RIbe286d8_26, RIbe2a190_83);
not \U$13030 ( \13276 , \13275 );
and \U$13031 ( \13277 , \13274 , \13276 );
buf \U$13032 ( \13278 , \11399 );
and \U$13033 ( \13279 , \13278 , \10680 );
nor \U$13034 ( \13280 , \13277 , \13279 );
nand \U$13035 ( \13281 , \13273 , \13280 );
not \U$13036 ( \13282 , \13281 );
xor \U$13037 ( \13283 , RIbe29ec0_77, RIbe28228_16);
not \U$13038 ( \13284 , \13283 );
not \U$13039 ( \13285 , \3056 );
or \U$13040 ( \13286 , \13284 , \13285 );
nand \U$13041 ( \13287 , \8680 , \10653 );
nand \U$13042 ( \13288 , \13286 , \13287 );
not \U$13043 ( \13289 , \13288 );
or \U$13044 ( \13290 , \13282 , \13289 );
not \U$13045 ( \13291 , \13280 );
nand \U$13046 ( \13292 , \13272 , \13291 );
nand \U$13047 ( \13293 , \13290 , \13292 );
nor \U$13048 ( \13294 , \13265 , \13293 );
xor \U$13049 ( \13295 , RIbe28d68_40, RIbe28390_19);
not \U$13050 ( \13296 , \13295 );
not \U$13051 ( \13297 , \8651 );
or \U$13052 ( \13298 , \13296 , \13297 );
nand \U$13053 ( \13299 , \8654 , \11276 );
nand \U$13054 ( \13300 , \13298 , \13299 );
xor \U$13055 ( \13301 , RIbe29128_48, RIbe27e68_8);
not \U$13056 ( \13302 , \13301 );
not \U$13057 ( \13303 , \4443 );
or \U$13058 ( \13304 , \13302 , \13303 );
not \U$13059 ( \13305 , \2463 );
not \U$13060 ( \13306 , \13305 );
nand \U$13061 ( \13307 , \13306 , \11287 );
nand \U$13062 ( \13308 , \13304 , \13307 );
or \U$13063 ( \13309 , \13300 , \13308 );
xor \U$13064 ( \13310 , RIbe29e48_76, RIbe294e8_56);
not \U$13065 ( \13311 , \13310 );
not \U$13066 ( \13312 , \10938 );
or \U$13067 ( \13313 , \13311 , \13312 );
nand \U$13068 ( \13314 , \4851 , \11298 );
nand \U$13069 ( \13315 , \13313 , \13314 );
nand \U$13070 ( \13316 , \13309 , \13315 );
nand \U$13071 ( \13317 , \13300 , \13308 );
and \U$13072 ( \13318 , \13316 , \13317 );
or \U$13073 ( \13319 , \13294 , \13318 );
nand \U$13074 ( \13320 , \13265 , \13293 );
nand \U$13075 ( \13321 , \13319 , \13320 );
not \U$13076 ( \13322 , \13321 );
xor \U$13077 ( \13323 , RIbe2a910_99, RIbe284f8_22);
not \U$13078 ( \13324 , \13323 );
buf \U$13079 ( \13325 , \9737 );
not \U$13080 ( \13326 , \13325 );
or \U$13081 ( \13327 , \13324 , \13326 );
nand \U$13082 ( \13328 , \11456 , \11205 );
nand \U$13083 ( \13329 , \13327 , \13328 );
not \U$13084 ( \13330 , \13329 );
xor \U$13085 ( \13331 , RIbe297b8_62, RIbe28f48_44);
not \U$13086 ( \13332 , \13331 );
not \U$13087 ( \13333 , \11461 );
or \U$13088 ( \13334 , \13332 , \13333 );
nand \U$13089 ( \13335 , \11201 , \11197 );
nand \U$13090 ( \13336 , \13334 , \13335 );
not \U$13091 ( \13337 , \13336 );
not \U$13092 ( \13338 , \9193 );
xnor \U$13093 ( \13339 , RIbe27b20_1, RIbe28a20_33);
not \U$13094 ( \13340 , \13339 );
and \U$13095 ( \13341 , \13338 , \13340 );
and \U$13096 ( \13342 , \2475 , \11239 );
nor \U$13097 ( \13343 , \13341 , \13342 );
not \U$13098 ( \13344 , \13343 );
or \U$13099 ( \13345 , \13337 , \13344 );
or \U$13100 ( \13346 , \13343 , \13336 );
nand \U$13101 ( \13347 , \13345 , \13346 );
not \U$13102 ( \13348 , \13347 );
or \U$13103 ( \13349 , \13330 , \13348 );
not \U$13104 ( \13350 , \13343 );
nand \U$13105 ( \13351 , \13350 , \13336 );
nand \U$13106 ( \13352 , \13349 , \13351 );
not \U$13107 ( \13353 , \11350 );
or \U$13108 ( \13354 , \13352 , \13353 );
xor \U$13109 ( \13355 , RIbe296c8_60, RIbe2aa00_101);
not \U$13110 ( \13356 , \13355 );
not \U$13111 ( \13357 , \1129 );
or \U$13112 ( \13358 , \13356 , \13357 );
nand \U$13113 ( \13359 , \1939 , \10645 );
nand \U$13114 ( \13360 , \13358 , \13359 );
not \U$13115 ( \13361 , \13360 );
xor \U$13116 ( \13362 , RIbe2a550_91, RIbe28840_29);
not \U$13117 ( \13363 , \13362 );
not \U$13118 ( \13364 , \11999 );
or \U$13119 ( \13365 , \13363 , \13364 );
nand \U$13120 ( \13366 , \11485 , \11223 );
nand \U$13121 ( \13367 , \13365 , \13366 );
not \U$13122 ( \13368 , \13367 );
or \U$13123 ( \13369 , \13361 , \13368 );
or \U$13124 ( \13370 , \13367 , \13360 );
xor \U$13125 ( \13371 , RIbe2a820_97, RIbe29038_46);
not \U$13126 ( \13372 , \13371 );
not \U$13127 ( \13373 , \979 );
or \U$13128 ( \13374 , \13372 , \13373 );
nand \U$13129 ( \13375 , \287 , \10701 );
nand \U$13130 ( \13376 , \13374 , \13375 );
nand \U$13131 ( \13377 , \13370 , \13376 );
nand \U$13132 ( \13378 , \13369 , \13377 );
nand \U$13133 ( \13379 , \13354 , \13378 );
nand \U$13134 ( \13380 , \13352 , \13353 );
and \U$13135 ( \13381 , \13379 , \13380 );
xor \U$13136 ( \13382 , \13322 , \13381 );
not \U$13137 ( \13383 , \9375 );
not \U$13138 ( \13384 , \13383 );
xnor \U$13139 ( \13385 , RIbe29308_52, RIbe2a2f8_86);
not \U$13140 ( \13386 , \13385 );
and \U$13141 ( \13387 , \13384 , \13386 );
and \U$13142 ( \13388 , \8706 , \11312 );
nor \U$13143 ( \13389 , \13387 , \13388 );
not \U$13144 ( \13390 , \13389 );
not \U$13145 ( \13391 , \13390 );
xor \U$13146 ( \13392 , RIbe2a460_89, RIbe27c10_3);
not \U$13147 ( \13393 , \13392 );
not \U$13148 ( \13394 , \936 );
or \U$13149 ( \13395 , \13393 , \13394 );
nand \U$13150 ( \13396 , \1174 , \10663 );
nand \U$13151 ( \13397 , \13395 , \13396 );
not \U$13152 ( \13398 , \13397 );
not \U$13153 ( \13399 , \13398 );
xor \U$13154 ( \13400 , RIbe29ce0_73, RIbe28930_31);
not \U$13155 ( \13401 , \13400 );
not \U$13156 ( \13402 , \11374 );
or \U$13157 ( \13403 , \13401 , \13402 );
nand \U$13158 ( \13404 , \1797 , \11372 );
nand \U$13159 ( \13405 , \13403 , \13404 );
not \U$13160 ( \13406 , \13405 );
or \U$13161 ( \13407 , \13399 , \13406 );
or \U$13162 ( \13408 , \13405 , \13398 );
nand \U$13163 ( \13409 , \13407 , \13408 );
not \U$13164 ( \13410 , \13409 );
or \U$13165 ( \13411 , \13391 , \13410 );
nand \U$13166 ( \13412 , \13397 , \13405 );
nand \U$13167 ( \13413 , \13411 , \13412 );
not \U$13168 ( \13414 , \13413 );
nand \U$13169 ( \13415 , RIbe27b98_2, RIbe2a6b8_94);
not \U$13170 ( \13416 , \13415 );
xor \U$13171 ( \13417 , RIbe28de0_41, RIbe2ad48_108);
not \U$13172 ( \13418 , \13417 );
not \U$13173 ( \13419 , \331 );
or \U$13174 ( \13420 , \13418 , \13419 );
nand \U$13175 ( \13421 , \346 , \11319 );
nand \U$13176 ( \13422 , \13420 , \13421 );
not \U$13177 ( \13423 , \13422 );
or \U$13178 ( \13424 , \13416 , \13423 );
or \U$13179 ( \13425 , \13422 , \13415 );
nand \U$13180 ( \13426 , \13424 , \13425 );
and \U$13181 ( \13427 , RIbe27df0_7, RIbe28480_21);
nor \U$13182 ( \13428 , RIbe27df0_7, RIbe28480_21);
nor \U$13183 ( \13429 , \13427 , \13428 );
not \U$13184 ( \13430 , \13429 );
not \U$13185 ( \13431 , \3344 );
or \U$13186 ( \13432 , \13430 , \13431 );
nand \U$13187 ( \13433 , \3075 , \11259 );
nand \U$13188 ( \13434 , \13432 , \13433 );
and \U$13189 ( \13435 , \13426 , \13434 );
not \U$13190 ( \13436 , \13422 );
nor \U$13191 ( \13437 , \13436 , \13415 );
nor \U$13192 ( \13438 , \13435 , \13437 );
not \U$13193 ( \13439 , \13438 );
not \U$13194 ( \13440 , RIbe27fd0_11);
not \U$13195 ( \13441 , RIbe295d8_58);
and \U$13196 ( \13442 , \13440 , \13441 );
and \U$13197 ( \13443 , RIbe27fd0_11, RIbe295d8_58);
nor \U$13198 ( \13444 , \13442 , \13443 );
not \U$13199 ( \13445 , \13444 );
not \U$13200 ( \13446 , \11366 );
or \U$13201 ( \13447 , \13445 , \13446 );
nand \U$13202 ( \13448 , \2707 , \11364 );
nand \U$13203 ( \13449 , \13447 , \13448 );
not \U$13204 ( \13450 , \13449 );
xor \U$13205 ( \13451 , RIbe2b2e8_120, RIbe27d78_6);
not \U$13206 ( \13452 , \13451 );
not \U$13207 ( \13453 , \8898 );
or \U$13208 ( \13454 , \13452 , \13453 );
nand \U$13209 ( \13455 , \10752 , \11214 );
nand \U$13210 ( \13456 , \13454 , \13455 );
not \U$13211 ( \13457 , \13456 );
xor \U$13212 ( \13458 , RIbe27b98_2, RIbe2b4c8_124);
not \U$13213 ( \13459 , \13458 );
not \U$13214 ( \13460 , \4827 );
or \U$13215 ( \13461 , \13459 , \13460 );
nand \U$13216 ( \13462 , \267 , \11180 );
nand \U$13217 ( \13463 , \13461 , \13462 );
not \U$13218 ( \13464 , \13463 );
not \U$13219 ( \13465 , \13464 );
or \U$13220 ( \13466 , \13457 , \13465 );
or \U$13221 ( \13467 , \13464 , \13456 );
nand \U$13222 ( \13468 , \13466 , \13467 );
not \U$13223 ( \13469 , \13468 );
or \U$13224 ( \13470 , \13450 , \13469 );
nand \U$13225 ( \13471 , \13463 , \13456 );
nand \U$13226 ( \13472 , \13470 , \13471 );
not \U$13227 ( \13473 , \13472 );
or \U$13228 ( \13474 , \13439 , \13473 );
or \U$13229 ( \13475 , \13472 , \13438 );
nand \U$13230 ( \13476 , \13474 , \13475 );
not \U$13231 ( \13477 , \13476 );
or \U$13232 ( \13478 , \13414 , \13477 );
not \U$13233 ( \13479 , \13438 );
nand \U$13234 ( \13480 , \13479 , \13472 );
nand \U$13235 ( \13481 , \13478 , \13480 );
not \U$13236 ( \13482 , \13481 );
and \U$13237 ( \13483 , \13382 , \13482 );
and \U$13238 ( \13484 , \13322 , \13381 );
or \U$13239 ( \13485 , \13483 , \13484 );
not \U$13240 ( \13486 , \13485 );
and \U$13241 ( \13487 , \13237 , \13486 );
and \U$13242 ( \13488 , \13197 , \13236 );
or \U$13243 ( \13489 , \13487 , \13488 );
not \U$13244 ( \13490 , \11437 );
not \U$13245 ( \13491 , \11434 );
or \U$13246 ( \13492 , \13490 , \13491 );
or \U$13247 ( \13493 , \11434 , \11437 );
nand \U$13248 ( \13494 , \13492 , \13493 );
nor \U$13249 ( \13495 , \13489 , \13494 );
or \U$13250 ( \13496 , \13177 , \13495 );
nand \U$13251 ( \13497 , \13489 , \13494 );
nand \U$13252 ( \13498 , \13496 , \13497 );
not \U$13253 ( \13499 , \13498 );
or \U$13254 ( \13500 , \13093 , \13499 );
not \U$13255 ( \13501 , \13091 );
not \U$13256 ( \13502 , \13498 );
not \U$13257 ( \13503 , \13502 );
or \U$13258 ( \13504 , \13501 , \13503 );
xor \U$13259 ( \13505 , \12242 , \12208 );
not \U$13260 ( \13506 , \13505 );
xor \U$13261 ( \13507 , \12233 , \12219 );
not \U$13262 ( \13508 , \13507 );
xor \U$13263 ( \13509 , \11017 , \10967 );
xor \U$13264 ( \13510 , \13509 , \10916 );
not \U$13265 ( \13511 , \13510 );
xor \U$13266 ( \13512 , RIbe2a028_80, RIbe28a98_34);
not \U$13267 ( \13513 , \13512 );
not \U$13268 ( \13514 , \9531 );
or \U$13269 ( \13515 , \13513 , \13514 );
nand \U$13270 ( \13516 , \9065 , \10672 );
nand \U$13271 ( \13517 , \13515 , \13516 );
xor \U$13272 ( \13518 , RIbe2b108_116, RIbe29380_53);
not \U$13273 ( \13519 , \13518 );
and \U$13274 ( \13520 , RIbe2b180_117, RIbe2b270_119);
not \U$13275 ( \13521 , RIbe2b180_117);
and \U$13276 ( \13522 , \13521 , RIbe2b108_116);
nor \U$13277 ( \13523 , \13520 , \13522 );
nand \U$13278 ( \13524 , RIbe2b108_116, RIbe2b270_119);
not \U$13279 ( \13525 , \13524 );
nor \U$13280 ( \13526 , \13523 , \13525 );
buf \U$13281 ( \13527 , \13526 );
not \U$13282 ( \13528 , \13527 );
not \U$13283 ( \13529 , \13528 );
not \U$13284 ( \13530 , \13529 );
or \U$13285 ( \13531 , \13519 , \13530 );
xor \U$13286 ( \13532 , RIbe2b180_117, RIbe2b270_119);
buf \U$13287 ( \13533 , \13532 );
buf \U$13288 ( \13534 , \13533 );
nand \U$13289 ( \13535 , \13534 , RIbe2b108_116);
nand \U$13290 ( \13536 , \13531 , \13535 );
or \U$13291 ( \13537 , \13517 , \13536 );
not \U$13292 ( \13538 , \13534 );
not \U$13293 ( \13539 , \13538 );
not \U$13294 ( \13540 , \13527 );
not \U$13295 ( \13541 , \13540 );
buf \U$13296 ( \13542 , \13541 );
buf \U$13297 ( \13543 , \13542 );
not \U$13298 ( \13544 , \13543 );
not \U$13299 ( \13545 , \13544 );
or \U$13300 ( \13546 , \13539 , \13545 );
nand \U$13301 ( \13547 , \13546 , RIbe2b108_116);
nand \U$13302 ( \13548 , \13537 , \13547 );
nand \U$13303 ( \13549 , \13536 , \13517 );
nand \U$13304 ( \13550 , \13548 , \13549 );
xor \U$13305 ( \13551 , \11210 , \11219 );
xor \U$13306 ( \13552 , \13551 , \11203 );
xor \U$13307 ( \13553 , \13550 , \13552 );
not \U$13308 ( \13554 , \13553 );
xor \U$13309 ( \13555 , RIbe28750_27, RIbe2a550_91);
not \U$13310 ( \13556 , \13555 );
not \U$13311 ( \13557 , \10434 );
or \U$13312 ( \13558 , \13556 , \13557 );
nand \U$13313 ( \13559 , \11228 , \13362 );
nand \U$13314 ( \13560 , \13558 , \13559 );
not \U$13315 ( \13561 , \13560 );
xor \U$13316 ( \13562 , RIbe28a20_33, RIbe29b78_70);
not \U$13317 ( \13563 , \13562 );
not \U$13318 ( \13564 , \2276 );
or \U$13319 ( \13565 , \13563 , \13564 );
not \U$13320 ( \13566 , \13339 );
nand \U$13321 ( \13567 , \13566 , \2476 );
nand \U$13322 ( \13568 , \13565 , \13567 );
not \U$13323 ( \13569 , \13568 );
or \U$13324 ( \13570 , \13561 , \13569 );
or \U$13325 ( \13571 , \13568 , \13560 );
xor \U$13326 ( \13572 , RIbe29c68_72, RIbe28138_14);
not \U$13327 ( \13573 , \13572 );
not \U$13328 ( \13574 , \4578 );
or \U$13329 ( \13575 , \13573 , \13574 );
nand \U$13330 ( \13576 , \4580 , \13256 );
nand \U$13331 ( \13577 , \13575 , \13576 );
nand \U$13332 ( \13578 , \13571 , \13577 );
nand \U$13333 ( \13579 , \13570 , \13578 );
not \U$13334 ( \13580 , \13579 );
xor \U$13335 ( \13581 , RIbe2a910_99, RIbe28318_18);
not \U$13336 ( \13582 , \13581 );
not \U$13337 ( \13583 , \10987 );
or \U$13338 ( \13584 , \13582 , \13583 );
nand \U$13339 ( \13585 , \9726 , \13323 );
nand \U$13340 ( \13586 , \13584 , \13585 );
xor \U$13341 ( \13587 , RIbe27d78_6, RIbe2a4d8_90);
not \U$13342 ( \13588 , \13587 );
not \U$13343 ( \13589 , \5739 );
or \U$13344 ( \13590 , \13588 , \13589 );
nand \U$13345 ( \13591 , \10752 , \13451 );
nand \U$13346 ( \13592 , \13590 , \13591 );
nor \U$13347 ( \13593 , \13586 , \13592 );
not \U$13348 ( \13594 , \9618 );
not \U$13349 ( \13595 , \13594 );
xor \U$13350 ( \13596 , RIbe29740_61, RIbe28f48_44);
not \U$13351 ( \13597 , \13596 );
not \U$13352 ( \13598 , \13597 );
and \U$13353 ( \13599 , \13595 , \13598 );
not \U$13354 ( \13600 , \13331 );
nor \U$13355 ( \13601 , \13600 , \3250 );
nor \U$13356 ( \13602 , \13599 , \13601 );
or \U$13357 ( \13603 , \13593 , \13602 );
nand \U$13358 ( \13604 , \13586 , \13592 );
nand \U$13359 ( \13605 , \13603 , \13604 );
not \U$13360 ( \13606 , \13605 );
xor \U$13361 ( \13607 , RIbe28c00_37, RIbe2a3e8_88);
not \U$13362 ( \13608 , \13607 );
not \U$13363 ( \13609 , \8806 );
or \U$13364 ( \13610 , \13608 , \13609 );
nand \U$13365 ( \13611 , \8794 , \13112 );
nand \U$13366 ( \13612 , \13610 , \13611 );
not \U$13367 ( \13613 , \13612 );
not \U$13368 ( \13614 , \13613 );
xor \U$13369 ( \13615 , RIbe27b98_2, RIbe2a6b8_94);
not \U$13370 ( \13616 , \13615 );
not \U$13371 ( \13617 , \8380 );
or \U$13372 ( \13618 , \13616 , \13617 );
nand \U$13373 ( \13619 , \7585 , \13458 );
nand \U$13374 ( \13620 , \13618 , \13619 );
not \U$13375 ( \13621 , \13620 );
not \U$13376 ( \13622 , \13621 );
or \U$13377 ( \13623 , \13614 , \13622 );
xor \U$13378 ( \13624 , RIbe280c0_13, RIbe2aa78_102);
not \U$13379 ( \13625 , \13624 );
not \U$13380 ( \13626 , \2380 );
or \U$13381 ( \13627 , \13625 , \13626 );
nand \U$13382 ( \13628 , \1265 , \13128 );
nand \U$13383 ( \13629 , \13627 , \13628 );
nand \U$13384 ( \13630 , \13623 , \13629 );
nand \U$13385 ( \13631 , \13620 , \13612 );
nand \U$13386 ( \13632 , \13630 , \13631 );
not \U$13387 ( \13633 , \13632 );
not \U$13388 ( \13634 , \13633 );
or \U$13389 ( \13635 , \13606 , \13634 );
not \U$13390 ( \13636 , \13605 );
nand \U$13391 ( \13637 , \13636 , \13632 );
nand \U$13392 ( \13638 , \13635 , \13637 );
not \U$13393 ( \13639 , \13638 );
or \U$13394 ( \13640 , \13580 , \13639 );
nand \U$13395 ( \13641 , \13605 , \13632 );
nand \U$13396 ( \13642 , \13640 , \13641 );
not \U$13397 ( \13643 , \13642 );
or \U$13398 ( \13644 , \13554 , \13643 );
nand \U$13399 ( \13645 , \13552 , \13550 );
nand \U$13400 ( \13646 , \13644 , \13645 );
not \U$13401 ( \13647 , \13646 );
not \U$13402 ( \13648 , \10741 );
not \U$13403 ( \13649 , \10767 );
or \U$13404 ( \13650 , \13648 , \13649 );
or \U$13405 ( \13651 , \10767 , \10741 );
nand \U$13406 ( \13652 , \13650 , \13651 );
and \U$13407 ( \13653 , \13652 , \10797 );
not \U$13408 ( \13654 , \13652 );
not \U$13409 ( \13655 , \10797 );
and \U$13410 ( \13656 , \13654 , \13655 );
nor \U$13411 ( \13657 , \13653 , \13656 );
not \U$13412 ( \13658 , \13657 );
not \U$13413 ( \13659 , \13658 );
not \U$13414 ( \13660 , \10827 );
not \U$13415 ( \13661 , \10889 );
or \U$13416 ( \13662 , \13660 , \13661 );
or \U$13417 ( \13663 , \10889 , \10827 );
nand \U$13418 ( \13664 , \13662 , \13663 );
not \U$13419 ( \13665 , \13664 );
not \U$13420 ( \13666 , \13665 );
or \U$13421 ( \13667 , \13659 , \13666 );
nand \U$13422 ( \13668 , \13657 , \13664 );
nand \U$13423 ( \13669 , \13667 , \13668 );
not \U$13424 ( \13670 , \13669 );
or \U$13425 ( \13671 , \13647 , \13670 );
nand \U$13426 ( \13672 , \13658 , \13664 );
nand \U$13427 ( \13673 , \13671 , \13672 );
not \U$13428 ( \13674 , \13673 );
or \U$13429 ( \13675 , \13511 , \13674 );
or \U$13430 ( \13676 , \13673 , \13510 );
nand \U$13431 ( \13677 , \13675 , \13676 );
not \U$13432 ( \13678 , \13677 );
or \U$13433 ( \13679 , \13508 , \13678 );
not \U$13434 ( \13680 , \13510 );
nand \U$13435 ( \13681 , \13680 , \13673 );
nand \U$13436 ( \13682 , \13679 , \13681 );
not \U$13437 ( \13683 , \10623 );
and \U$13438 ( \13684 , \11021 , \13683 );
not \U$13439 ( \13685 , \11021 );
and \U$13440 ( \13686 , \13685 , \10623 );
nor \U$13441 ( \13687 , \13684 , \13686 );
xnor \U$13442 ( \13688 , \13682 , \13687 );
not \U$13443 ( \13689 , \13688 );
or \U$13444 ( \13690 , \13506 , \13689 );
not \U$13445 ( \13691 , \13687 );
nand \U$13446 ( \13692 , \13691 , \13682 );
nand \U$13447 ( \13693 , \13690 , \13692 );
nand \U$13448 ( \13694 , \13504 , \13693 );
nand \U$13449 ( \13695 , \13500 , \13694 );
nand \U$13450 ( \13696 , \13090 , \13695 );
not \U$13451 ( \13697 , \13088 );
not \U$13452 ( \13698 , \13076 );
nand \U$13453 ( \13699 , \13697 , \13698 );
nand \U$13454 ( \13700 , \13696 , \13699 );
nand \U$13455 ( \13701 , \13073 , \13700 );
or \U$13456 ( \13702 , \13072 , \13701 );
not \U$13457 ( \13703 , \13070 );
buf \U$13458 ( \13704 , \12868 );
buf \U$13459 ( \13705 , \12870 );
nand \U$13460 ( \13706 , \13703 , \13704 , \13705 );
nand \U$13461 ( \13707 , \13702 , \13706 );
not \U$13462 ( \13708 , \12982 );
not \U$13463 ( \13709 , \12994 );
or \U$13464 ( \13710 , \13708 , \13709 );
nand \U$13465 ( \13711 , \12993 , \12988 );
nand \U$13466 ( \13712 , \13710 , \13711 );
not \U$13467 ( \13713 , \13712 );
not \U$13468 ( \13714 , \13713 );
not \U$13469 ( \13715 , \12976 );
not \U$13470 ( \13716 , \12972 );
or \U$13471 ( \13717 , \13715 , \13716 );
not \U$13472 ( \13718 , \12970 );
nand \U$13473 ( \13719 , \13718 , \12963 );
nand \U$13474 ( \13720 , \13717 , \13719 );
not \U$13475 ( \13721 , \12892 );
not \U$13476 ( \13722 , \12888 );
or \U$13477 ( \13723 , \13721 , \13722 );
nand \U$13478 ( \13724 , \12319 , \12882 );
nand \U$13479 ( \13725 , \13723 , \13724 );
and \U$13480 ( \13726 , \9346 , \9020 );
not \U$13481 ( \13727 , \9346 );
and \U$13482 ( \13728 , \13727 , \9021 );
nor \U$13483 ( \13729 , \13726 , \13728 );
xnor \U$13484 ( \13730 , \13725 , \13729 );
xor \U$13485 ( \13731 , \13720 , \13730 );
not \U$13486 ( \13732 , \12908 );
not \U$13487 ( \13733 , \12903 );
or \U$13488 ( \13734 , \13732 , \13733 );
nand \U$13489 ( \13735 , \12898 , \12893 );
nand \U$13490 ( \13736 , \13734 , \13735 );
xor \U$13491 ( \13737 , \13731 , \13736 );
not \U$13492 ( \13738 , \13737 );
and \U$13493 ( \13739 , \13714 , \13738 );
and \U$13494 ( \13740 , \13713 , \13737 );
nor \U$13495 ( \13741 , \13739 , \13740 );
xor \U$13496 ( \13742 , \12947 , \12960 );
and \U$13497 ( \13743 , \13742 , \12977 );
and \U$13498 ( \13744 , \12947 , \12960 );
or \U$13499 ( \13745 , \13743 , \13744 );
not \U$13500 ( \13746 , \13745 );
xor \U$13501 ( \13747 , \12938 , \12943 );
and \U$13502 ( \13748 , \13747 , \12946 );
and \U$13503 ( \13749 , \12938 , \12943 );
or \U$13504 ( \13750 , \13748 , \13749 );
xor \U$13505 ( \13751 , \9259 , \9296 );
xor \U$13506 ( \13752 , \13751 , \9328 );
xor \U$13507 ( \13753 , \13750 , \13752 );
not \U$13508 ( \13754 , \13039 );
not \U$13509 ( \13755 , \13040 );
not \U$13510 ( \13756 , \13042 );
or \U$13511 ( \13757 , \13755 , \13756 );
or \U$13512 ( \13758 , \13042 , \13040 );
nand \U$13513 ( \13759 , \13757 , \13758 );
not \U$13514 ( \13760 , \13759 );
or \U$13515 ( \13761 , \13754 , \13760 );
not \U$13516 ( \13762 , \13042 );
nand \U$13517 ( \13763 , \13762 , \13040 );
nand \U$13518 ( \13764 , \13761 , \13763 );
xor \U$13519 ( \13765 , \13753 , \13764 );
xor \U$13520 ( \13766 , \13746 , \13765 );
not \U$13521 ( \13767 , \13037 );
and \U$13522 ( \13768 , \13043 , \13026 );
not \U$13523 ( \13769 , \13043 );
not \U$13524 ( \13770 , \13026 );
and \U$13525 ( \13771 , \13769 , \13770 );
nor \U$13526 ( \13772 , \13768 , \13771 );
not \U$13527 ( \13773 , \13772 );
or \U$13528 ( \13774 , \13767 , \13773 );
nand \U$13529 ( \13775 , \13043 , \13026 );
nand \U$13530 ( \13776 , \13774 , \13775 );
xnor \U$13531 ( \13777 , \13766 , \13776 );
xor \U$13532 ( \13778 , \13741 , \13777 );
not \U$13533 ( \13779 , \12978 );
not \U$13534 ( \13780 , \12995 );
not \U$13535 ( \13781 , \13004 );
or \U$13536 ( \13782 , \13780 , \13781 );
or \U$13537 ( \13783 , \13004 , \12995 );
nand \U$13538 ( \13784 , \13782 , \13783 );
not \U$13539 ( \13785 , \13784 );
or \U$13540 ( \13786 , \13779 , \13785 );
nand \U$13541 ( \13787 , \13003 , \12995 );
nand \U$13542 ( \13788 , \13786 , \13787 );
not \U$13543 ( \13789 , \13788 );
xnor \U$13544 ( \13790 , \13778 , \13789 );
not \U$13545 ( \13791 , \13790 );
not \U$13546 ( \13792 , \13791 );
not \U$13547 ( \13793 , \13005 );
not \U$13548 ( \13794 , \12933 );
or \U$13549 ( \13795 , \13793 , \13794 );
not \U$13550 ( \13796 , \12924 );
nand \U$13551 ( \13797 , \13796 , \12929 );
nand \U$13552 ( \13798 , \13795 , \13797 );
xor \U$13553 ( \13799 , \9815 , \9843 );
xor \U$13554 ( \13800 , \9872 , \13799 );
not \U$13555 ( \13801 , \9886 );
not \U$13556 ( \13802 , \9890 );
or \U$13557 ( \13803 , \13801 , \13802 );
or \U$13558 ( \13804 , \9886 , \9890 );
nand \U$13559 ( \13805 , \13803 , \13804 );
xor \U$13560 ( \13806 , \9903 , \13805 );
xor \U$13561 ( \13807 , \13800 , \13806 );
xor \U$13562 ( \13808 , \9171 , \9202 );
xor \U$13563 ( \13809 , \13808 , \9225 );
xor \U$13564 ( \13810 , \13807 , \13809 );
not \U$13565 ( \13811 , \13810 );
not \U$13566 ( \13812 , \13028 );
nand \U$13567 ( \13813 , \13812 , \13029 );
not \U$13568 ( \13814 , \13813 );
not \U$13569 ( \13815 , \13036 );
or \U$13570 ( \13816 , \13814 , \13815 );
nand \U$13571 ( \13817 , \13030 , \13028 );
nand \U$13572 ( \13818 , \13816 , \13817 );
xor \U$13573 ( \13819 , \12949 , \12953 );
and \U$13574 ( \13820 , \13819 , \12959 );
and \U$13575 ( \13821 , \12949 , \12953 );
or \U$13576 ( \13822 , \13820 , \13821 );
xor \U$13577 ( \13823 , \13818 , \13822 );
and \U$13578 ( \13824 , \9785 , \9722 );
not \U$13579 ( \13825 , \9785 );
not \U$13580 ( \13826 , \9722 );
and \U$13581 ( \13827 , \13825 , \13826 );
nor \U$13582 ( \13828 , \13824 , \13827 );
and \U$13583 ( \13829 , \13823 , \13828 );
not \U$13584 ( \13830 , \13823 );
not \U$13585 ( \13831 , \13828 );
and \U$13586 ( \13832 , \13830 , \13831 );
nor \U$13587 ( \13833 , \13829 , \13832 );
not \U$13588 ( \13834 , \13833 );
not \U$13589 ( \13835 , \13834 );
or \U$13590 ( \13836 , \13811 , \13835 );
not \U$13591 ( \13837 , \13810 );
nand \U$13592 ( \13838 , \13837 , \13833 );
nand \U$13593 ( \13839 , \13836 , \13838 );
not \U$13594 ( \13840 , \12923 );
not \U$13595 ( \13841 , \12915 );
or \U$13596 ( \13842 , \13840 , \13841 );
nand \U$13597 ( \13843 , \12909 , \12876 );
nand \U$13598 ( \13844 , \13842 , \13843 );
not \U$13599 ( \13845 , \13844 );
xor \U$13600 ( \13846 , \13839 , \13845 );
xor \U$13601 ( \13847 , \13023 , \13044 );
and \U$13602 ( \13848 , \13847 , \13053 );
and \U$13603 ( \13849 , \13023 , \13044 );
or \U$13604 ( \13850 , \13848 , \13849 );
xnor \U$13605 ( \13851 , \13846 , \13850 );
xor \U$13606 ( \13852 , \13798 , \13851 );
not \U$13607 ( \13853 , \13852 );
or \U$13608 ( \13854 , \13792 , \13853 );
not \U$13609 ( \13855 , \13852 );
not \U$13610 ( \13856 , \13855 );
not \U$13611 ( \13857 , \13790 );
or \U$13612 ( \13858 , \13856 , \13857 );
or \U$13613 ( \13859 , \13054 , \13018 );
not \U$13614 ( \13860 , \13859 );
not \U$13615 ( \13861 , \13059 );
or \U$13616 ( \13862 , \13860 , \13861 );
nand \U$13617 ( \13863 , \13054 , \13018 );
nand \U$13618 ( \13864 , \13862 , \13863 );
nand \U$13619 ( \13865 , \13858 , \13864 );
nand \U$13620 ( \13866 , \13854 , \13865 );
not \U$13621 ( \13867 , \13866 );
not \U$13622 ( \13868 , \13777 );
not \U$13623 ( \13869 , \13741 );
not \U$13624 ( \13870 , \13788 );
or \U$13625 ( \13871 , \13869 , \13870 );
or \U$13626 ( \13872 , \13788 , \13741 );
nand \U$13627 ( \13873 , \13871 , \13872 );
not \U$13628 ( \13874 , \13873 );
or \U$13629 ( \13875 , \13868 , \13874 );
not \U$13630 ( \13876 , \13741 );
nand \U$13631 ( \13877 , \13876 , \13788 );
nand \U$13632 ( \13878 , \13875 , \13877 );
not \U$13633 ( \13879 , \13878 );
not \U$13634 ( \13880 , \13798 );
not \U$13635 ( \13881 , \13851 );
or \U$13636 ( \13882 , \13880 , \13881 );
xor \U$13637 ( \13883 , \13839 , \13844 );
nand \U$13638 ( \13884 , \13883 , \13850 );
nand \U$13639 ( \13885 , \13882 , \13884 );
not \U$13640 ( \13886 , \13885 );
xor \U$13641 ( \13887 , \13879 , \13886 );
not \U$13642 ( \13888 , \13737 );
not \U$13643 ( \13889 , \13712 );
or \U$13644 ( \13890 , \13888 , \13889 );
nand \U$13645 ( \13891 , \13736 , \13731 );
nand \U$13646 ( \13892 , \13890 , \13891 );
xor \U$13647 ( \13893 , \13800 , \13806 );
and \U$13648 ( \13894 , \13893 , \13809 );
and \U$13649 ( \13895 , \13800 , \13806 );
or \U$13650 ( \13896 , \13894 , \13895 );
xor \U$13651 ( \13897 , \9079 , \9168 );
xor \U$13652 ( \13898 , \13897 , \9228 );
xor \U$13653 ( \13899 , \13896 , \13898 );
xor \U$13654 ( \13900 , \13750 , \13752 );
and \U$13655 ( \13901 , \13900 , \13764 );
and \U$13656 ( \13902 , \13750 , \13752 );
or \U$13657 ( \13903 , \13901 , \13902 );
xnor \U$13658 ( \13904 , \13899 , \13903 );
xor \U$13659 ( \13905 , \13892 , \13904 );
not \U$13660 ( \13906 , \13765 );
xnor \U$13661 ( \13907 , \13746 , \13776 );
not \U$13662 ( \13908 , \13907 );
or \U$13663 ( \13909 , \13906 , \13908 );
not \U$13664 ( \13910 , \13746 );
nand \U$13665 ( \13911 , \13910 , \13776 );
nand \U$13666 ( \13912 , \13909 , \13911 );
not \U$13667 ( \13913 , \13912 );
xnor \U$13668 ( \13914 , \13905 , \13913 );
not \U$13669 ( \13915 , \13914 );
not \U$13670 ( \13916 , \13839 );
not \U$13671 ( \13917 , \13844 );
or \U$13672 ( \13918 , \13916 , \13917 );
nand \U$13673 ( \13919 , \13810 , \13833 );
nand \U$13674 ( \13920 , \13918 , \13919 );
not \U$13675 ( \13921 , \13920 );
not \U$13676 ( \13922 , \13730 );
not \U$13677 ( \13923 , \13720 );
or \U$13678 ( \13924 , \13922 , \13923 );
not \U$13679 ( \13925 , \13729 );
nand \U$13680 ( \13926 , \13925 , \13725 );
nand \U$13681 ( \13927 , \13924 , \13926 );
xor \U$13682 ( \13928 , \9331 , \9356 );
xor \U$13683 ( \13929 , \13927 , \13928 );
not \U$13684 ( \13930 , \13828 );
not \U$13685 ( \13931 , \13823 );
or \U$13686 ( \13932 , \13930 , \13931 );
nand \U$13687 ( \13933 , \13822 , \13818 );
nand \U$13688 ( \13934 , \13932 , \13933 );
not \U$13689 ( \13935 , \13934 );
and \U$13690 ( \13936 , \13929 , \13935 );
not \U$13691 ( \13937 , \13929 );
and \U$13692 ( \13938 , \13937 , \13934 );
or \U$13693 ( \13939 , \13936 , \13938 );
xor \U$13694 ( \13940 , \9712 , \9714 );
xor \U$13695 ( \13941 , \13940 , \9716 );
xnor \U$13696 ( \13942 , \9392 , \9386 );
xor \U$13697 ( \13943 , \9702 , \9704 );
xor \U$13698 ( \13944 , \13943 , \9707 );
and \U$13699 ( \13945 , \13942 , \13944 );
not \U$13700 ( \13946 , \13942 );
not \U$13701 ( \13947 , \13944 );
and \U$13702 ( \13948 , \13946 , \13947 );
or \U$13703 ( \13949 , \13945 , \13948 );
xor \U$13704 ( \13950 , \13941 , \13949 );
not \U$13705 ( \13951 , \9789 );
and \U$13706 ( \13952 , \9909 , \13951 );
not \U$13707 ( \13953 , \9909 );
and \U$13708 ( \13954 , \13953 , \9789 );
nor \U$13709 ( \13955 , \13952 , \13954 );
xnor \U$13710 ( \13956 , \13950 , \13955 );
not \U$13711 ( \13957 , \13956 );
xor \U$13712 ( \13958 , \13939 , \13957 );
not \U$13713 ( \13959 , \13958 );
or \U$13714 ( \13960 , \13921 , \13959 );
or \U$13715 ( \13961 , \13920 , \13958 );
nand \U$13716 ( \13962 , \13960 , \13961 );
not \U$13717 ( \13963 , \13962 );
and \U$13718 ( \13964 , \13915 , \13963 );
and \U$13719 ( \13965 , \13914 , \13962 );
nor \U$13720 ( \13966 , \13964 , \13965 );
xor \U$13721 ( \13967 , \13887 , \13966 );
nand \U$13722 ( \13968 , \13867 , \13967 );
xor \U$13723 ( \13969 , \13864 , \13790 );
xor \U$13724 ( \13970 , \13969 , \13852 );
xor \U$13725 ( \13971 , \13010 , \13064 );
and \U$13726 ( \13972 , \13971 , \13069 );
and \U$13727 ( \13973 , \13010 , \13064 );
or \U$13728 ( \13974 , \13972 , \13973 );
nand \U$13729 ( \13975 , \13970 , \13974 );
nand \U$13730 ( \13976 , \13968 , \13975 );
not \U$13731 ( \13977 , \13976 );
and \U$13732 ( \13978 , \13707 , \13977 );
not \U$13733 ( \13979 , \13956 );
not \U$13734 ( \13980 , \13939 );
or \U$13735 ( \13981 , \13979 , \13980 );
not \U$13736 ( \13982 , \13955 );
xor \U$13737 ( \13983 , \13949 , \13941 );
nand \U$13738 ( \13984 , \13982 , \13983 );
nand \U$13739 ( \13985 , \13981 , \13984 );
not \U$13740 ( \13986 , \13985 );
xor \U$13741 ( \13987 , \8876 , \8951 );
xor \U$13742 ( \13988 , \13987 , \9004 );
not \U$13743 ( \13989 , \13941 );
not \U$13744 ( \13990 , \13949 );
or \U$13745 ( \13991 , \13989 , \13990 );
not \U$13746 ( \13992 , \13942 );
nand \U$13747 ( \13993 , \13992 , \13944 );
nand \U$13748 ( \13994 , \13991 , \13993 );
and \U$13749 ( \13995 , \13988 , \13994 );
not \U$13750 ( \13996 , \13988 );
not \U$13751 ( \13997 , \13994 );
and \U$13752 ( \13998 , \13996 , \13997 );
nor \U$13753 ( \13999 , \13995 , \13998 );
not \U$13754 ( \14000 , \13999 );
xor \U$13755 ( \14001 , \9231 , \9403 );
not \U$13756 ( \14002 , \14001 );
or \U$13757 ( \14003 , \14000 , \14002 );
not \U$13758 ( \14004 , \13999 );
not \U$13759 ( \14005 , \14001 );
nand \U$13760 ( \14006 , \14004 , \14005 );
nand \U$13761 ( \14007 , \14003 , \14006 );
nand \U$13762 ( \14008 , \13986 , \14007 );
not \U$13763 ( \14009 , \14008 );
not \U$13764 ( \14010 , \13912 );
not \U$13765 ( \14011 , \13892 );
nand \U$13766 ( \14012 , \14011 , \13904 );
not \U$13767 ( \14013 , \14012 );
or \U$13768 ( \14014 , \14010 , \14013 );
xor \U$13769 ( \14015 , \13896 , \13898 );
xor \U$13770 ( \14016 , \14015 , \13903 );
nand \U$13771 ( \14017 , \14016 , \13892 );
nand \U$13772 ( \14018 , \14014 , \14017 );
not \U$13773 ( \14019 , \14018 );
not \U$13774 ( \14020 , \14019 );
not \U$13775 ( \14021 , \14020 );
or \U$13776 ( \14022 , \14009 , \14021 );
or \U$13777 ( \14023 , \13986 , \14007 );
nand \U$13778 ( \14024 , \14022 , \14023 );
not \U$13779 ( \14025 , \14024 );
not \U$13780 ( \14026 , \14025 );
not \U$13781 ( \14027 , \13988 );
nand \U$13782 ( \14028 , \14027 , \13997 );
not \U$13783 ( \14029 , \14028 );
not \U$13784 ( \14030 , \14001 );
or \U$13785 ( \14031 , \14029 , \14030 );
nand \U$13786 ( \14032 , \13994 , \13988 );
nand \U$13787 ( \14033 , \14031 , \14032 );
not \U$13788 ( \14034 , \14033 );
not \U$13789 ( \14035 , \14034 );
nand \U$13790 ( \14036 , \9009 , \9410 );
xor \U$13791 ( \14037 , \14036 , \9407 );
not \U$13792 ( \14038 , \14037 );
not \U$13793 ( \14039 , \14038 );
or \U$13794 ( \14040 , \14035 , \14039 );
nand \U$13795 ( \14041 , \14037 , \14033 );
nand \U$13796 ( \14042 , \14040 , \14041 );
not \U$13797 ( \14043 , \9982 );
xor \U$13798 ( \14044 , \9996 , \14043 );
xnor \U$13799 ( \14045 , \14044 , \9943 );
xor \U$13800 ( \14046 , \14042 , \14045 );
not \U$13801 ( \14047 , \13934 );
not \U$13802 ( \14048 , \13929 );
or \U$13803 ( \14049 , \14047 , \14048 );
nand \U$13804 ( \14050 , \13928 , \13927 );
nand \U$13805 ( \14051 , \14049 , \14050 );
not \U$13806 ( \14052 , \14051 );
not \U$13807 ( \14053 , \14052 );
xor \U$13808 ( \14054 , \9939 , \9720 );
not \U$13809 ( \14055 , \14054 );
or \U$13810 ( \14056 , \14053 , \14055 );
or \U$13811 ( \14057 , \14054 , \14052 );
nand \U$13812 ( \14058 , \14056 , \14057 );
not \U$13813 ( \14059 , \14058 );
xor \U$13814 ( \14060 , \13903 , \13896 );
and \U$13815 ( \14061 , \14060 , \13898 );
and \U$13816 ( \14062 , \13903 , \13896 );
or \U$13817 ( \14063 , \14061 , \14062 );
not \U$13818 ( \14064 , \14063 );
or \U$13819 ( \14065 , \14059 , \14064 );
not \U$13820 ( \14066 , \14052 );
nand \U$13821 ( \14067 , \14066 , \14054 );
nand \U$13822 ( \14068 , \14065 , \14067 );
xor \U$13823 ( \14069 , \14046 , \14068 );
not \U$13824 ( \14070 , \14069 );
or \U$13825 ( \14071 , \14026 , \14070 );
or \U$13826 ( \14072 , \14069 , \14025 );
nand \U$13827 ( \14073 , \14071 , \14072 );
not \U$13828 ( \14074 , \13962 );
not \U$13829 ( \14075 , \13914 );
not \U$13830 ( \14076 , \14075 );
or \U$13831 ( \14077 , \14074 , \14076 );
not \U$13832 ( \14078 , \13958 );
nand \U$13833 ( \14079 , \14078 , \13920 );
nand \U$13834 ( \14080 , \14077 , \14079 );
not \U$13835 ( \14081 , \14007 );
not \U$13836 ( \14082 , \13986 );
or \U$13837 ( \14083 , \14081 , \14082 );
or \U$13838 ( \14084 , \14007 , \13986 );
nand \U$13839 ( \14085 , \14083 , \14084 );
not \U$13840 ( \14086 , \14085 );
and \U$13841 ( \14087 , \14019 , \14086 );
not \U$13842 ( \14088 , \14019 );
and \U$13843 ( \14089 , \14088 , \14085 );
nor \U$13844 ( \14090 , \14087 , \14089 );
xnor \U$13845 ( \14091 , \14058 , \14063 );
nand \U$13846 ( \14092 , \14090 , \14091 );
nand \U$13847 ( \14093 , \14080 , \14092 );
not \U$13848 ( \14094 , \14090 );
not \U$13849 ( \14095 , \14091 );
nand \U$13850 ( \14096 , \14094 , \14095 );
and \U$13851 ( \14097 , \14093 , \14096 );
nand \U$13852 ( \14098 , \14073 , \14097 );
nand \U$13853 ( \14099 , \14096 , \14092 );
and \U$13854 ( \14100 , \14099 , \14080 );
not \U$13855 ( \14101 , \14099 );
not \U$13856 ( \14102 , \14080 );
and \U$13857 ( \14103 , \14101 , \14102 );
nor \U$13858 ( \14104 , \14100 , \14103 );
xor \U$13859 ( \14105 , \13879 , \13886 );
and \U$13860 ( \14106 , \14105 , \13966 );
and \U$13861 ( \14107 , \13879 , \13886 );
or \U$13862 ( \14108 , \14106 , \14107 );
nand \U$13863 ( \14109 , \14104 , \14108 );
nand \U$13864 ( \14110 , \14098 , \14109 );
xnor \U$13865 ( \14111 , \10035 , \10050 );
not \U$13866 ( \14112 , \14111 );
xor \U$13867 ( \14113 , \9411 , \9692 );
xor \U$13868 ( \14114 , \14113 , \10001 );
nand \U$13869 ( \14115 , \14112 , \14114 );
buf \U$13870 ( \14116 , \14115 );
not \U$13871 ( \14117 , \14114 );
nand \U$13872 ( \14118 , \14117 , \14111 );
nand \U$13873 ( \14119 , \14034 , \14037 );
not \U$13874 ( \14120 , \14119 );
not \U$13875 ( \14121 , \14068 );
or \U$13876 ( \14122 , \14120 , \14121 );
nand \U$13877 ( \14123 , \14038 , \14033 );
nand \U$13878 ( \14124 , \14122 , \14123 );
nand \U$13879 ( \14125 , \14118 , \14124 );
nand \U$13880 ( \14126 , \14116 , \14125 );
not \U$13881 ( \14127 , \14126 );
not \U$13882 ( \14128 , \10004 );
xor \U$13883 ( \14129 , \10140 , \14128 );
xnor \U$13884 ( \14130 , \14129 , \10185 );
nand \U$13885 ( \14131 , \14127 , \14130 );
not \U$13886 ( \14132 , \14045 );
not \U$13887 ( \14133 , \14042 );
not \U$13888 ( \14134 , \14068 );
or \U$13889 ( \14135 , \14133 , \14134 );
or \U$13890 ( \14136 , \14068 , \14042 );
nand \U$13891 ( \14137 , \14135 , \14136 );
not \U$13892 ( \14138 , \14137 );
or \U$13893 ( \14139 , \14132 , \14138 );
nand \U$13894 ( \14140 , \14139 , \14024 );
not \U$13895 ( \14141 , \14137 );
not \U$13896 ( \14142 , \14045 );
nand \U$13897 ( \14143 , \14141 , \14142 );
nand \U$13898 ( \14144 , \14140 , \14143 );
not \U$13899 ( \14145 , \14144 );
nand \U$13900 ( \14146 , \14118 , \14115 );
and \U$13901 ( \14147 , \14146 , \14124 );
not \U$13902 ( \14148 , \14146 );
not \U$13903 ( \14149 , \14124 );
and \U$13904 ( \14150 , \14148 , \14149 );
nor \U$13905 ( \14151 , \14147 , \14150 );
nand \U$13906 ( \14152 , \14145 , \14151 );
nand \U$13907 ( \14153 , \14131 , \14152 );
nor \U$13908 ( \14154 , \14110 , \14153 );
nand \U$13909 ( \14155 , \10395 , \13978 , \14154 );
nor \U$13910 ( \14156 , \10381 , \10375 );
buf \U$13911 ( \14157 , \10393 );
and \U$13912 ( \14158 , \14156 , \14157 );
nor \U$13913 ( \14159 , \10390 , \10392 );
nor \U$13914 ( \14160 , \14158 , \14159 );
nand \U$13915 ( \14161 , \14155 , \14160 );
not \U$13916 ( \14162 , \14161 );
or \U$13917 ( \14163 , \8521 , \14162 );
not \U$13918 ( \14164 , \8103 );
not \U$13919 ( \14165 , \8513 );
not \U$13920 ( \14166 , \8518 );
nand \U$13921 ( \14167 , \14165 , \14166 );
or \U$13922 ( \14168 , \14164 , \14167 );
or \U$13923 ( \14169 , \8102 , \7987 );
nand \U$13924 ( \14170 , \14168 , \14169 );
and \U$13925 ( \14171 , \14170 , \8128 );
nor \U$13926 ( \14172 , \8127 , \8122 );
nor \U$13927 ( \14173 , \14171 , \14172 );
nand \U$13928 ( \14174 , \14163 , \14173 );
not \U$13929 ( \14175 , \8118 );
and \U$13930 ( \14176 , \14175 , \8110 );
and \U$13931 ( \14177 , \8104 , \8109 );
nor \U$13932 ( \14178 , \14176 , \14177 );
not \U$13933 ( \14179 , \4755 );
and \U$13934 ( \14180 , \5104 , \14179 );
not \U$13935 ( \14181 , \5104 );
and \U$13936 ( \14182 , \14181 , \4755 );
nor \U$13937 ( \14183 , \14180 , \14182 );
nand \U$13938 ( \14184 , \14178 , \14183 );
nand \U$13939 ( \14185 , \14174 , \14184 );
not \U$13940 ( \14186 , \13967 );
nand \U$13941 ( \14187 , \14186 , \13866 );
not \U$13942 ( \14188 , \14187 );
buf \U$13943 ( \14189 , \13968 );
nor \U$13944 ( \14190 , \13970 , \13974 );
nand \U$13945 ( \14191 , \14189 , \14190 );
not \U$13946 ( \14192 , \14191 );
or \U$13947 ( \14193 , \14188 , \14192 );
nand \U$13948 ( \14194 , \14193 , \14154 );
not \U$13949 ( \14195 , \14194 );
not \U$13950 ( \14196 , \14153 );
not \U$13951 ( \14197 , \14196 );
not \U$13952 ( \14198 , \14104 );
not \U$13953 ( \14199 , \14108 );
nand \U$13954 ( \14200 , \14198 , \14199 );
not \U$13955 ( \14201 , \14098 );
or \U$13956 ( \14202 , \14200 , \14201 );
or \U$13957 ( \14203 , \14097 , \14073 );
nand \U$13958 ( \14204 , \14202 , \14203 );
not \U$13959 ( \14205 , \14204 );
or \U$13960 ( \14206 , \14197 , \14205 );
not \U$13961 ( \14207 , \14151 );
nand \U$13962 ( \14208 , \14207 , \14144 );
not \U$13963 ( \14209 , \14208 );
nand \U$13964 ( \14210 , \14209 , \14131 );
not \U$13965 ( \14211 , \14130 );
nand \U$13966 ( \14212 , \14211 , \14126 );
and \U$13967 ( \14213 , \14210 , \14212 );
nand \U$13968 ( \14214 , \14206 , \14213 );
or \U$13969 ( \14215 , \14195 , \14214 );
buf \U$13970 ( \14216 , \10395 );
nand \U$13971 ( \14217 , \14215 , \14216 );
not \U$13972 ( \14218 , \10394 );
not \U$13973 ( \14219 , \10345 );
not \U$13974 ( \14220 , \10288 );
not \U$13975 ( \14221 , \10187 );
not \U$13976 ( \14222 , \14221 );
nand \U$13977 ( \14223 , \14220 , \14222 );
or \U$13978 ( \14224 , \14219 , \14223 );
not \U$13979 ( \14225 , \10344 );
buf \U$13980 ( \14226 , \10294 );
nand \U$13981 ( \14227 , \14225 , \14226 );
nand \U$13982 ( \14228 , \14224 , \14227 );
nand \U$13983 ( \14229 , \14218 , \14228 );
nand \U$13984 ( \14230 , \14217 , \14229 );
and \U$13985 ( \14231 , \8519 , \8128 , \8103 , \14184 );
nand \U$13986 ( \14232 , \14230 , \14231 );
or \U$13987 ( \14233 , \14178 , \14183 );
and \U$13988 ( \14234 , \14185 , \14232 , \14233 );
xor \U$13989 ( \14235 , RIbe2a910_99, RIbe28c78_38);
not \U$13990 ( \14236 , \14235 );
not \U$13991 ( \14237 , \9736 );
or \U$13992 ( \14238 , \14236 , \14237 );
nand \U$13993 ( \14239 , \10400 , \13581 );
nand \U$13994 ( \14240 , \14238 , \14239 );
xor \U$13995 ( \14241 , RIbe28a20_33, RIbe29ce0_73);
not \U$13996 ( \14242 , \14241 );
not \U$13997 ( \14243 , \1779 );
or \U$13998 ( \14244 , \14242 , \14243 );
nand \U$13999 ( \14245 , \1768 , \13562 );
nand \U$14000 ( \14246 , \14244 , \14245 );
xor \U$14001 ( \14247 , \14240 , \14246 );
buf \U$14002 ( \14248 , \14247 );
xor \U$14003 ( \14249 , RIbe295d8_58, RIbe28f48_44);
not \U$14004 ( \14250 , \14249 );
not \U$14005 ( \14251 , \9618 );
or \U$14006 ( \14252 , \14250 , \14251 );
nand \U$14007 ( \14253 , \11201 , \13596 );
nand \U$14008 ( \14254 , \14252 , \14253 );
xnor \U$14009 ( \14255 , \14248 , \14254 );
not \U$14010 ( \14256 , \14255 );
not \U$14011 ( \14257 , \14256 );
xor \U$14012 ( \14258 , RIbe284f8_22, RIbe2a550_91);
not \U$14013 ( \14259 , \14258 );
not \U$14014 ( \14260 , \10432 );
or \U$14015 ( \14261 , \14259 , \14260 );
nand \U$14016 ( \14262 , \11484 , \13555 );
nand \U$14017 ( \14263 , \14261 , \14262 );
xor \U$14018 ( \14264 , RIbe29038_46, RIbe2a0a0_81);
not \U$14019 ( \14265 , \14264 );
not \U$14020 ( \14266 , \280 );
or \U$14021 ( \14267 , \14265 , \14266 );
xor \U$14022 ( \14268 , RIbe29038_46, RIbe2a118_82);
nand \U$14023 ( \14269 , \284 , \14268 );
nand \U$14024 ( \14270 , \14267 , \14269 );
and \U$14025 ( \14271 , \14263 , \14270 );
not \U$14026 ( \14272 , \14263 );
not \U$14027 ( \14273 , \14270 );
and \U$14028 ( \14274 , \14272 , \14273 );
nor \U$14029 ( \14275 , \14271 , \14274 );
xor \U$14030 ( \14276 , RIbe2a820_97, RIbe296c8_60);
not \U$14031 ( \14277 , \14276 );
not \U$14032 ( \14278 , \1129 );
or \U$14033 ( \14279 , \14277 , \14278 );
xor \U$14034 ( \14280 , RIbe296c8_60, RIbe2a898_98);
nand \U$14035 ( \14281 , \8534 , \14280 );
nand \U$14036 ( \14282 , \14279 , \14281 );
xor \U$14037 ( \14283 , \14275 , \14282 );
not \U$14038 ( \14284 , \14283 );
xor \U$14039 ( \14285 , RIbe293f8_54, RIbe2a3e8_88);
not \U$14040 ( \14286 , \14285 );
not \U$14041 ( \14287 , \9262 );
or \U$14042 ( \14288 , \14286 , \14287 );
xor \U$14043 ( \14289 , RIbe29308_52, RIbe2a3e8_88);
nand \U$14044 ( \14290 , \9089 , \14289 );
nand \U$14045 ( \14291 , \14288 , \14290 );
not \U$14046 ( \14292 , \14291 );
not \U$14047 ( \14293 , \14292 );
xor \U$14048 ( \14294 , RIbe27ee0_9, RIbe2b108_116);
not \U$14049 ( \14295 , \14294 );
buf \U$14050 ( \14296 , \13526 );
buf \U$14051 ( \14297 , \14296 );
not \U$14052 ( \14298 , \14297 );
or \U$14053 ( \14299 , \14295 , \14298 );
xor \U$14054 ( \14300 , RIbe2b108_116, RIbe28048_12);
nand \U$14055 ( \14301 , \13534 , \14300 );
nand \U$14056 ( \14302 , \14299 , \14301 );
not \U$14057 ( \14303 , \14302 );
or \U$14058 ( \14304 , \14293 , \14303 );
xor \U$14059 ( \14305 , RIbe28138_14, RIbe29e48_76);
not \U$14060 ( \14306 , \14305 );
and \U$14061 ( \14307 , \4838 , \4839 );
not \U$14062 ( \14308 , \14307 );
or \U$14063 ( \14309 , \14306 , \14308 );
xor \U$14064 ( \14310 , RIbe282a0_17, RIbe29e48_76);
nand \U$14065 ( \14311 , \4849 , \14310 );
nand \U$14066 ( \14312 , \14309 , \14311 );
nand \U$14067 ( \14313 , \14304 , \14312 );
not \U$14068 ( \14314 , \14302 );
nand \U$14069 ( \14315 , \14314 , \14291 );
and \U$14070 ( \14316 , \14313 , \14315 );
not \U$14071 ( \14317 , \14316 );
or \U$14072 ( \14318 , \14284 , \14317 );
or \U$14073 ( \14319 , \14283 , \14316 );
nand \U$14074 ( \14320 , \14318 , \14319 );
not \U$14075 ( \14321 , \14320 );
or \U$14076 ( \14322 , \14257 , \14321 );
not \U$14077 ( \14323 , \14316 );
nand \U$14078 ( \14324 , \14323 , \14283 );
nand \U$14079 ( \14325 , \14322 , \14324 );
not \U$14080 ( \14326 , \14325 );
not \U$14081 ( \14327 , \14326 );
not \U$14082 ( \14328 , \14280 );
not \U$14083 ( \14329 , \2877 );
or \U$14084 ( \14330 , \14328 , \14329 );
nand \U$14085 ( \14331 , \908 , \13355 );
nand \U$14086 ( \14332 , \14330 , \14331 );
xor \U$14087 ( \14333 , RIbe29f38_78, RIbe28228_16);
not \U$14088 ( \14334 , \14333 );
not \U$14089 ( \14335 , \879 );
or \U$14090 ( \14336 , \14334 , \14335 );
nand \U$14091 ( \14337 , \885 , \13283 );
nand \U$14092 ( \14338 , \14336 , \14337 );
xor \U$14093 ( \14339 , RIbe27c10_3, RIbe2adc0_109);
not \U$14094 ( \14340 , \14339 );
not \U$14095 ( \14341 , \7440 );
or \U$14096 ( \14342 , \14340 , \14341 );
nand \U$14097 ( \14343 , \1173 , \13392 );
nand \U$14098 ( \14344 , \14342 , \14343 );
xor \U$14099 ( \14345 , \14338 , \14344 );
xor \U$14100 ( \14346 , \14332 , \14345 );
not \U$14101 ( \14347 , \14346 );
xor \U$14102 ( \14348 , RIbe28de0_41, RIbe2b540_125);
not \U$14103 ( \14349 , \14348 );
not \U$14104 ( \14350 , \924 );
or \U$14105 ( \14351 , \14349 , \14350 );
nand \U$14106 ( \14352 , \1149 , \13417 );
nand \U$14107 ( \14353 , \14351 , \14352 );
xor \U$14108 ( \14354 , RIbe290b0_47, RIbe2b360_121);
not \U$14109 ( \14355 , \14354 );
not \U$14110 ( \14356 , \9114 );
or \U$14111 ( \14357 , \14355 , \14356 );
nand \U$14112 ( \14358 , \399 , \13238 );
nand \U$14113 ( \14359 , \14357 , \14358 );
xor \U$14114 ( \14360 , \14353 , \14359 );
not \U$14115 ( \14361 , \14360 );
xor \U$14116 ( \14362 , RIbe27c88_4, RIbe28480_21);
and \U$14117 ( \14363 , \2520 , \14362 );
and \U$14118 ( \14364 , \11263 , \13429 );
nor \U$14119 ( \14365 , \14363 , \14364 );
not \U$14120 ( \14366 , \14365 );
and \U$14121 ( \14367 , \14361 , \14366 );
and \U$14122 ( \14368 , \14360 , \14365 );
nor \U$14123 ( \14369 , \14367 , \14368 );
not \U$14124 ( \14370 , \14369 );
or \U$14125 ( \14371 , \14347 , \14370 );
or \U$14126 ( \14372 , \14369 , \14346 );
nand \U$14127 ( \14373 , \14371 , \14372 );
xor \U$14128 ( \14374 , RIbe27fd0_11, RIbe291a0_49);
not \U$14129 ( \14375 , \14374 );
not \U$14130 ( \14376 , \12808 );
or \U$14131 ( \14377 , \14375 , \14376 );
nand \U$14132 ( \14378 , \2707 , \13444 );
nand \U$14133 ( \14379 , \14377 , \14378 );
xor \U$14134 ( \14380 , RIbe2a280_85, RIbe27ee0_9);
not \U$14135 ( \14381 , \14380 );
not \U$14136 ( \14382 , \11344 );
buf \U$14137 ( \14383 , \14382 );
not \U$14138 ( \14384 , \14383 );
or \U$14139 ( \14385 , \14381 , \14384 );
nand \U$14140 ( \14386 , \11348 , \13266 );
nand \U$14141 ( \14387 , \14385 , \14386 );
xor \U$14142 ( \14388 , \14379 , \14387 );
xor \U$14143 ( \14389 , RIbe28930_31, RIbe29d58_74);
not \U$14144 ( \14390 , \14389 );
or \U$14145 ( \14391 , \967 , \14390 );
not \U$14146 ( \14392 , \13400 );
or \U$14147 ( \14393 , \972 , \14392 );
nand \U$14148 ( \14394 , \14391 , \14393 );
xor \U$14149 ( \14395 , \14388 , \14394 );
xnor \U$14150 ( \14396 , \14373 , \14395 );
not \U$14151 ( \14397 , \14396 );
not \U$14152 ( \14398 , \14397 );
or \U$14153 ( \14399 , \14327 , \14398 );
nand \U$14154 ( \14400 , \14396 , \14325 );
nand \U$14155 ( \14401 , \14399 , \14400 );
not \U$14156 ( \14402 , \14401 );
xor \U$14157 ( \14403 , RIbe294e8_56, RIbe2a2f8_86);
not \U$14158 ( \14404 , \14403 );
not \U$14159 ( \14405 , \10792 );
or \U$14160 ( \14406 , \14404 , \14405 );
xor \U$14161 ( \14407 , RIbe288b8_30, RIbe2a2f8_86);
nand \U$14162 ( \14408 , \8706 , \14407 );
nand \U$14163 ( \14409 , \14406 , \14408 );
not \U$14164 ( \14410 , \14409 );
xor \U$14165 ( \14411 , RIbe2afa0_113, RIbe2b018_114);
not \U$14166 ( \14412 , \14411 );
not \U$14167 ( \14413 , \14412 );
not \U$14168 ( \14414 , \14413 );
not \U$14169 ( \14415 , \14414 );
not \U$14170 ( \14416 , RIbe2af28_112);
nor \U$14171 ( \14417 , RIbe2afa0_113, RIbe2b018_114);
not \U$14172 ( \14418 , \14417 );
or \U$14173 ( \14419 , \14416 , \14418 );
not \U$14174 ( \14420 , RIbe2af28_112);
nand \U$14175 ( \14421 , \14420 , RIbe2b018_114, RIbe2afa0_113);
nand \U$14176 ( \14422 , \14419 , \14421 );
buf \U$14177 ( \14423 , \14422 );
not \U$14178 ( \14424 , \14423 );
not \U$14179 ( \14425 , \14424 );
or \U$14180 ( \14426 , \14415 , \14425 );
nand \U$14181 ( \14427 , \14426 , RIbe2af28_112);
not \U$14182 ( \14428 , \14427 );
not \U$14183 ( \14429 , \14428 );
xor \U$14184 ( \14430 , RIbe27c10_3, RIbe2b4c8_124);
not \U$14185 ( \14431 , \14430 );
not \U$14186 ( \14432 , \7440 );
or \U$14187 ( \14433 , \14431 , \14432 );
xor \U$14188 ( \14434 , RIbe27c10_3, RIbe2b540_125);
nand \U$14189 ( \14435 , \369 , \14434 );
nand \U$14190 ( \14436 , \14433 , \14435 );
not \U$14191 ( \14437 , \14436 );
and \U$14192 ( \14438 , \14429 , \14437 );
and \U$14193 ( \14439 , \14428 , \14436 );
nor \U$14194 ( \14440 , \14438 , \14439 );
not \U$14195 ( \14441 , \14440 );
not \U$14196 ( \14442 , \14441 );
or \U$14197 ( \14443 , \14410 , \14442 );
nand \U$14198 ( \14444 , \14427 , \14436 );
nand \U$14199 ( \14445 , \14443 , \14444 );
not \U$14200 ( \14446 , \14445 );
xnor \U$14201 ( \14447 , RIbe285e8_24, RIbe28d68_40);
or \U$14202 ( \14448 , \2762 , \14447 );
xor \U$14203 ( \14449 , RIbe285e8_24, RIbe27c88_4);
not \U$14204 ( \14450 , \14449 );
or \U$14205 ( \14451 , \3502 , \14450 );
nand \U$14206 ( \14452 , \14448 , \14451 );
not \U$14207 ( \14453 , \14452 );
xor \U$14208 ( \14454 , RIbe2a910_99, RIbe29308_52);
not \U$14209 ( \14455 , \14454 );
not \U$14210 ( \14456 , \11453 );
or \U$14211 ( \14457 , \14455 , \14456 );
xor \U$14212 ( \14458 , RIbe2a910_99, RIbe28c00_37);
nand \U$14213 ( \14459 , \9726 , \14458 );
nand \U$14214 ( \14460 , \14457 , \14459 );
xor \U$14215 ( \14461 , RIbe29038_46, RIbe2b2e8_120);
not \U$14216 ( \14462 , \14461 );
not \U$14217 ( \14463 , \281 );
or \U$14218 ( \14464 , \14462 , \14463 );
xor \U$14219 ( \14465 , RIbe2b360_121, RIbe29038_46);
nand \U$14220 ( \14466 , \1583 , \14465 );
nand \U$14221 ( \14467 , \14464 , \14466 );
xor \U$14222 ( \14468 , \14460 , \14467 );
not \U$14223 ( \14469 , \14468 );
or \U$14224 ( \14470 , \14453 , \14469 );
nand \U$14225 ( \14471 , \14460 , \14467 );
nand \U$14226 ( \14472 , \14470 , \14471 );
xor \U$14227 ( \14473 , RIbe2a3e8_88, RIbe28a98_34);
not \U$14228 ( \14474 , \14473 );
not \U$14229 ( \14475 , \9263 );
or \U$14230 ( \14476 , \14474 , \14475 );
nand \U$14231 ( \14477 , \9268 , \14285 );
nand \U$14232 ( \14478 , \14476 , \14477 );
not \U$14233 ( \14479 , \14478 );
xor \U$14234 ( \14480 , RIbe2a820_97, RIbe280c0_13);
not \U$14235 ( \14481 , \14480 );
not \U$14236 ( \14482 , \8624 );
or \U$14237 ( \14483 , \14481 , \14482 );
xor \U$14238 ( \14484 , RIbe2a898_98, RIbe280c0_13);
nand \U$14239 ( \14485 , \1263 , \14484 );
nand \U$14240 ( \14486 , \14483 , \14485 );
not \U$14241 ( \14487 , \14486 );
xor \U$14242 ( \14488 , RIbe28a20_33, RIbe29ec0_77);
not \U$14243 ( \14489 , \14488 );
not \U$14244 ( \14490 , \1780 );
or \U$14245 ( \14491 , \14489 , \14490 );
xor \U$14246 ( \14492 , RIbe28a20_33, RIbe29d58_74);
nand \U$14247 ( \14493 , \1768 , \14492 );
nand \U$14248 ( \14494 , \14491 , \14493 );
not \U$14249 ( \14495 , \14494 );
not \U$14250 ( \14496 , \14495 );
or \U$14251 ( \14497 , \14487 , \14496 );
or \U$14252 ( \14498 , \14495 , \14486 );
nand \U$14253 ( \14499 , \14497 , \14498 );
not \U$14254 ( \14500 , \14499 );
or \U$14255 ( \14501 , \14479 , \14500 );
not \U$14256 ( \14502 , \14495 );
nand \U$14257 ( \14503 , \14502 , \14486 );
nand \U$14258 ( \14504 , \14501 , \14503 );
xor \U$14259 ( \14505 , \14472 , \14504 );
not \U$14260 ( \14506 , \14505 );
or \U$14261 ( \14507 , \14446 , \14506 );
nand \U$14262 ( \14508 , \14472 , \14504 );
nand \U$14263 ( \14509 , \14507 , \14508 );
not \U$14264 ( \14510 , \14509 );
xor \U$14265 ( \14511 , RIbe2a028_80, RIbe282a0_17);
not \U$14266 ( \14512 , \14511 );
buf \U$14267 ( \14513 , \8168 );
not \U$14268 ( \14514 , \14513 );
or \U$14269 ( \14515 , \14512 , \14514 );
xor \U$14270 ( \14516 , RIbe29470_55, RIbe2a028_80);
nand \U$14271 ( \14517 , \8172 , \14516 );
nand \U$14272 ( \14518 , \14515 , \14517 );
not \U$14273 ( \14519 , \14518 );
xor \U$14274 ( \14520 , RIbe27b98_2, RIbe2abe0_105);
not \U$14275 ( \14521 , \14520 );
not \U$14276 ( \14522 , \9833 );
or \U$14277 ( \14523 , \14521 , \14522 );
xor \U$14278 ( \14524 , RIbe2ac58_106, RIbe27b98_2);
nand \U$14279 ( \14525 , \14524 , \267 );
nand \U$14280 ( \14526 , \14523 , \14525 );
not \U$14281 ( \14527 , \14526 );
xor \U$14282 ( \14528 , RIbe27e68_8, RIbe27df0_7);
not \U$14283 ( \14529 , \14528 );
not \U$14284 ( \14530 , \2457 );
or \U$14285 ( \14531 , \14529 , \14530 );
xor \U$14286 ( \14532 , RIbe27e68_8, RIbe29218_50);
nand \U$14287 ( \14533 , \2463 , \14532 );
nand \U$14288 ( \14534 , \14531 , \14533 );
not \U$14289 ( \14535 , \14534 );
nand \U$14290 ( \14536 , \14527 , \14535 );
not \U$14291 ( \14537 , \14536 );
or \U$14292 ( \14538 , \14519 , \14537 );
not \U$14293 ( \14539 , \14535 );
nand \U$14294 ( \14540 , \14539 , \14526 );
nand \U$14295 ( \14541 , \14538 , \14540 );
not \U$14296 ( \14542 , \14541 );
xor \U$14297 ( \14543 , RIbe2b6a8_128, RIbe28930_31);
not \U$14298 ( \14544 , \14543 );
not \U$14299 ( \14545 , \965 );
or \U$14300 ( \14546 , \14544 , \14545 );
xor \U$14301 ( \14547 , RIbe29f38_78, RIbe28930_31);
nand \U$14302 ( \14548 , \970 , \14547 );
nand \U$14303 ( \14549 , \14546 , \14548 );
not \U$14304 ( \14550 , \14549 );
not \U$14305 ( \14551 , \4897 );
xor \U$14306 ( \14552 , RIbe29b00_69, RIbe27fd0_11);
not \U$14307 ( \14553 , \14552 );
or \U$14308 ( \14554 , \14551 , \14553 );
xor \U$14309 ( \14555 , RIbe27fd0_11, RIbe29a10_67);
not \U$14310 ( \14556 , \14555 );
or \U$14311 ( \14557 , \2717 , \14556 );
nand \U$14312 ( \14558 , \14554 , \14557 );
not \U$14313 ( \14559 , \14558 );
or \U$14314 ( \14560 , \14550 , \14559 );
or \U$14315 ( \14561 , \14558 , \14549 );
xor \U$14316 ( \14562 , RIbe2ad48_108, RIbe27d78_6);
not \U$14317 ( \14563 , \14562 );
not \U$14318 ( \14564 , \8768 );
or \U$14319 ( \14565 , \14563 , \14564 );
xor \U$14320 ( \14566 , RIbe27d78_6, RIbe2adc0_109);
nand \U$14321 ( \14567 , \314 , \14566 );
nand \U$14322 ( \14568 , \14565 , \14567 );
nand \U$14323 ( \14569 , \14561 , \14568 );
nand \U$14324 ( \14570 , \14560 , \14569 );
xor \U$14325 ( \14571 , RIbe286d8_26, RIbe2b108_116);
not \U$14326 ( \14572 , \14571 );
not \U$14327 ( \14573 , \14296 );
or \U$14328 ( \14574 , \14572 , \14573 );
nand \U$14329 ( \14575 , \13534 , \14294 );
nand \U$14330 ( \14576 , \14574 , \14575 );
xor \U$14331 ( \14577 , RIbe27b20_1, RIbe28390_19);
not \U$14332 ( \14578 , \14577 );
not \U$14333 ( \14579 , \2638 );
not \U$14334 ( \14580 , \14579 );
or \U$14335 ( \14581 , \14578 , \14580 );
xor \U$14336 ( \14582 , RIbe28390_19, RIbe28cf0_39);
nand \U$14337 ( \14583 , \2647 , \14582 );
nand \U$14338 ( \14584 , \14581 , \14583 );
or \U$14339 ( \14585 , \14576 , \14584 );
xor \U$14340 ( \14586 , RIbe297b8_62, RIbe29e48_76);
not \U$14341 ( \14587 , \14586 );
not \U$14342 ( \14588 , \11039 );
or \U$14343 ( \14589 , \14587 , \14588 );
nand \U$14344 ( \14590 , \4850 , \14305 );
nand \U$14345 ( \14591 , \14589 , \14590 );
nand \U$14346 ( \14592 , \14585 , \14591 );
nand \U$14347 ( \14593 , \14576 , \14584 );
nand \U$14348 ( \14594 , \14592 , \14593 );
xor \U$14349 ( \14595 , \14570 , \14594 );
not \U$14350 ( \14596 , \14595 );
or \U$14351 ( \14597 , \14542 , \14596 );
nand \U$14352 ( \14598 , \14594 , \14570 );
nand \U$14353 ( \14599 , \14597 , \14598 );
xor \U$14354 ( \14600 , RIbe28f48_44, RIbe29128_48);
not \U$14355 ( \14601 , \14600 );
not \U$14356 ( \14602 , \3256 );
or \U$14357 ( \14603 , \14601 , \14602 );
xor \U$14358 ( \14604 , RIbe28f48_44, RIbe291a0_49);
nand \U$14359 ( \14605 , \3249 , \14604 );
nand \U$14360 ( \14606 , \14603 , \14605 );
not \U$14361 ( \14607 , \14606 );
xor \U$14362 ( \14608 , RIbe28c78_38, RIbe2a550_91);
not \U$14363 ( \14609 , \14608 );
not \U$14364 ( \14610 , \11999 );
or \U$14365 ( \14611 , \14609 , \14610 );
not \U$14366 ( \14612 , \10439 );
xor \U$14367 ( \14613 , RIbe28318_18, RIbe2a550_91);
nand \U$14368 ( \14614 , \14612 , \14613 );
nand \U$14369 ( \14615 , \14611 , \14614 );
xor \U$14370 ( \14616 , RIbe290b0_47, RIbe2a460_89);
not \U$14371 ( \14617 , \14616 );
not \U$14372 ( \14618 , \2730 );
or \U$14373 ( \14619 , \14617 , \14618 );
xor \U$14374 ( \14620 , RIbe290b0_47, RIbe2a4d8_90);
nand \U$14375 ( \14621 , \10730 , \14620 );
nand \U$14376 ( \14622 , \14619 , \14621 );
xor \U$14377 ( \14623 , \14615 , \14622 );
not \U$14378 ( \14624 , \14623 );
or \U$14379 ( \14625 , \14607 , \14624 );
nand \U$14380 ( \14626 , \14615 , \14622 );
nand \U$14381 ( \14627 , \14625 , \14626 );
not \U$14382 ( \14628 , \14627 );
xor \U$14383 ( \14629 , RIbe296c8_60, RIbe2a0a0_81);
not \U$14384 ( \14630 , \14629 );
not \U$14385 ( \14631 , \900 );
or \U$14386 ( \14632 , \14630 , \14631 );
xor \U$14387 ( \14633 , RIbe296c8_60, RIbe2a118_82);
nand \U$14388 ( \14634 , \907 , \14633 );
nand \U$14389 ( \14635 , \14632 , \14634 );
xor \U$14390 ( \14636 , RIbe28228_16, RIbe2aa00_101);
not \U$14391 ( \14637 , \14636 );
buf \U$14392 ( \14638 , \878 );
not \U$14393 ( \14639 , \14638 );
or \U$14394 ( \14640 , \14637 , \14639 );
xor \U$14395 ( \14641 , RIbe28228_16, RIbe2aa78_102);
nand \U$14396 ( \14642 , \885 , \14641 );
nand \U$14397 ( \14643 , \14640 , \14642 );
or \U$14398 ( \14644 , \14635 , \14643 );
xor \U$14399 ( \14645 , RIbe28840_29, RIbe2a280_85);
not \U$14400 ( \14646 , \14645 );
not \U$14401 ( \14647 , \11345 );
or \U$14402 ( \14648 , \14646 , \14647 );
not \U$14403 ( \14649 , \10848 );
not \U$14404 ( \14650 , RIbe28570_23);
not \U$14405 ( \14651 , RIbe2a280_85);
and \U$14406 ( \14652 , \14650 , \14651 );
and \U$14407 ( \14653 , RIbe28570_23, RIbe2a280_85);
nor \U$14408 ( \14654 , \14652 , \14653 );
nand \U$14409 ( \14655 , \14649 , \14654 );
nand \U$14410 ( \14656 , \14648 , \14655 );
nand \U$14411 ( \14657 , \14644 , \14656 );
nand \U$14412 ( \14658 , \14643 , \14635 );
nand \U$14413 ( \14659 , \14657 , \14658 );
xor \U$14414 ( \14660 , RIbe295d8_58, RIbe29c68_72);
not \U$14415 ( \14661 , \14660 );
not \U$14416 ( \14662 , \5024 );
or \U$14417 ( \14663 , \14661 , \14662 );
xor \U$14418 ( \14664 , RIbe29740_61, RIbe29c68_72);
nand \U$14419 ( \14665 , \4580 , \14664 );
nand \U$14420 ( \14666 , \14663 , \14665 );
not \U$14421 ( \14667 , \14666 );
xor \U$14422 ( \14668 , RIbe28b88_36, RIbe29ce0_73);
not \U$14423 ( \14669 , \14668 );
not \U$14424 ( \14670 , \2552 );
or \U$14425 ( \14671 , \14669 , \14670 );
xor \U$14426 ( \14672 , RIbe28b88_36, RIbe29b78_70);
nand \U$14427 ( \14673 , \2558 , \14672 );
nand \U$14428 ( \14674 , \14671 , \14673 );
xor \U$14429 ( \14675 , RIbe284f8_22, RIbe2a190_83);
not \U$14430 ( \14676 , \14675 );
not \U$14431 ( \14677 , \10831 );
or \U$14432 ( \14678 , \14676 , \14677 );
xor \U$14433 ( \14679 , RIbe28750_27, RIbe2a190_83);
nand \U$14434 ( \14680 , \11399 , \14679 );
nand \U$14435 ( \14681 , \14678 , \14680 );
xor \U$14436 ( \14682 , \14674 , \14681 );
not \U$14437 ( \14683 , \14682 );
or \U$14438 ( \14684 , \14667 , \14683 );
nand \U$14439 ( \14685 , \14681 , \14674 );
nand \U$14440 ( \14686 , \14684 , \14685 );
and \U$14441 ( \14687 , \14659 , \14686 );
not \U$14442 ( \14688 , \14659 );
not \U$14443 ( \14689 , \14686 );
and \U$14444 ( \14690 , \14688 , \14689 );
nor \U$14445 ( \14691 , \14687 , \14690 );
not \U$14446 ( \14692 , \14691 );
or \U$14447 ( \14693 , \14628 , \14692 );
nand \U$14448 ( \14694 , \14686 , \14659 );
nand \U$14449 ( \14695 , \14693 , \14694 );
xor \U$14450 ( \14696 , \14599 , \14695 );
not \U$14451 ( \14697 , \14696 );
or \U$14452 ( \14698 , \14510 , \14697 );
nand \U$14453 ( \14699 , \14695 , \14599 );
nand \U$14454 ( \14700 , \14698 , \14699 );
not \U$14455 ( \14701 , \14700 );
or \U$14456 ( \14702 , \14402 , \14701 );
not \U$14457 ( \14703 , \14326 );
nand \U$14458 ( \14704 , \14703 , \14397 );
nand \U$14459 ( \14705 , \14702 , \14704 );
not \U$14460 ( \14706 , \14705 );
xor \U$14461 ( \14707 , \13612 , \13621 );
xor \U$14462 ( \14708 , \14707 , \13629 );
not \U$14463 ( \14709 , \14708 );
not \U$14464 ( \14710 , \14709 );
not \U$14465 ( \14711 , \13593 );
nand \U$14466 ( \14712 , \14711 , \13604 );
xor \U$14467 ( \14713 , \14712 , \13602 );
not \U$14468 ( \14714 , \14713 );
not \U$14469 ( \14715 , \14714 );
or \U$14470 ( \14716 , \14710 , \14715 );
nand \U$14471 ( \14717 , \14713 , \14708 );
nand \U$14472 ( \14718 , \14716 , \14717 );
xor \U$14473 ( \14719 , \13560 , \13568 );
xor \U$14474 ( \14720 , \14719 , \13577 );
not \U$14475 ( \14721 , \14720 );
and \U$14476 ( \14722 , \14718 , \14721 );
not \U$14477 ( \14723 , \14718 );
and \U$14478 ( \14724 , \14723 , \14720 );
nor \U$14479 ( \14725 , \14722 , \14724 );
not \U$14480 ( \14726 , \14725 );
not \U$14481 ( \14727 , \14726 );
xor \U$14482 ( \14728 , RIbe28570_23, RIbe2a190_83);
not \U$14483 ( \14729 , \14728 );
not \U$14484 ( \14730 , \10689 );
not \U$14485 ( \14731 , \14730 );
or \U$14486 ( \14732 , \14729 , \14731 );
not \U$14487 ( \14733 , \13275 );
nand \U$14488 ( \14734 , \14733 , \13278 );
nand \U$14489 ( \14735 , \14732 , \14734 );
xor \U$14490 ( \14736 , RIbe28cf0_39, RIbe28b88_36);
not \U$14491 ( \14737 , \14736 );
not \U$14492 ( \14738 , \8711 );
or \U$14493 ( \14739 , \14737 , \14738 );
nand \U$14494 ( \14740 , \2691 , \13245 );
nand \U$14495 ( \14741 , \14739 , \14740 );
xor \U$14496 ( \14742 , \14735 , \14741 );
xor \U$14497 ( \14743 , RIbe28390_19, RIbe29998_66);
not \U$14498 ( \14744 , \14743 );
not \U$14499 ( \14745 , \2640 );
or \U$14500 ( \14746 , \14744 , \14745 );
nand \U$14501 ( \14747 , \2777 , \13295 );
nand \U$14502 ( \14748 , \14746 , \14747 );
xor \U$14503 ( \14749 , \14742 , \14748 );
xor \U$14504 ( \14750 , RIbe29e48_76, RIbe29470_55);
not \U$14505 ( \14751 , \14750 );
not \U$14506 ( \14752 , \4842 );
or \U$14507 ( \14753 , \14751 , \14752 );
nand \U$14508 ( \14754 , \4851 , \13310 );
nand \U$14509 ( \14755 , \14753 , \14754 );
xor \U$14510 ( \14756 , RIbe285e8_24, RIbe29218_50);
not \U$14511 ( \14757 , \14756 );
not \U$14512 ( \14758 , \7618 );
or \U$14513 ( \14759 , \14757 , \14758 );
nand \U$14514 ( \14760 , \2625 , \13119 );
nand \U$14515 ( \14761 , \14759 , \14760 );
xor \U$14516 ( \14762 , \14755 , \14761 );
xor \U$14517 ( \14763 , RIbe27e68_8, RIbe29b00_69);
not \U$14518 ( \14764 , \14763 );
not \U$14519 ( \14765 , \2459 );
or \U$14520 ( \14766 , \14764 , \14765 );
nand \U$14521 ( \14767 , \4447 , \13301 );
nand \U$14522 ( \14768 , \14766 , \14767 );
xor \U$14523 ( \14769 , \14762 , \14768 );
xor \U$14524 ( \14770 , \14749 , \14769 );
xor \U$14525 ( \14771 , RIbe293f8_54, RIbe2a2f8_86);
not \U$14526 ( \14772 , \14771 );
not \U$14527 ( \14773 , \10792 );
or \U$14528 ( \14774 , \14772 , \14773 );
not \U$14529 ( \14775 , \13385 );
nand \U$14530 ( \14776 , \14775 , \8706 );
nand \U$14531 ( \14777 , \14774 , \14776 );
xor \U$14532 ( \14778 , RIbe2a028_80, RIbe288b8_30);
not \U$14533 ( \14779 , \14778 );
not \U$14534 ( \14780 , \9530 );
or \U$14535 ( \14781 , \14779 , \14780 );
nand \U$14536 ( \14782 , \8930 , \13512 );
nand \U$14537 ( \14783 , \14781 , \14782 );
not \U$14538 ( \14784 , \14268 );
not \U$14539 ( \14785 , \979 );
or \U$14540 ( \14786 , \14784 , \14785 );
nand \U$14541 ( \14787 , \1805 , \13371 );
nand \U$14542 ( \14788 , \14786 , \14787 );
xor \U$14543 ( \14789 , \14783 , \14788 );
xor \U$14544 ( \14790 , \14777 , \14789 );
xor \U$14545 ( \14791 , \14770 , \14790 );
not \U$14546 ( \14792 , \14791 );
not \U$14547 ( \14793 , \14310 );
not \U$14548 ( \14794 , \10938 );
or \U$14549 ( \14795 , \14793 , \14794 );
nand \U$14550 ( \14796 , \8245 , \14750 );
nand \U$14551 ( \14797 , \14795 , \14796 );
xor \U$14552 ( \14798 , RIbe27e68_8, RIbe29a10_67);
not \U$14553 ( \14799 , \14798 );
not \U$14554 ( \14800 , \2458 );
or \U$14555 ( \14801 , \14799 , \14800 );
nand \U$14556 ( \14802 , \13306 , \14763 );
nand \U$14557 ( \14803 , \14801 , \14802 );
xor \U$14558 ( \14804 , RIbe28390_19, RIbe298a8_64);
not \U$14559 ( \14805 , \14804 );
not \U$14560 ( \14806 , \2638 );
not \U$14561 ( \14807 , \14806 );
or \U$14562 ( \14808 , \14805 , \14807 );
nand \U$14563 ( \14809 , \2777 , \14743 );
nand \U$14564 ( \14810 , \14808 , \14809 );
and \U$14565 ( \14811 , \14803 , \14810 );
not \U$14566 ( \14812 , \14803 );
not \U$14567 ( \14813 , \14810 );
and \U$14568 ( \14814 , \14812 , \14813 );
nor \U$14569 ( \14815 , \14811 , \14814 );
xor \U$14570 ( \14816 , \14797 , \14815 );
not \U$14571 ( \14817 , \14816 );
xor \U$14572 ( \14818 , RIbe29ec0_77, RIbe28930_31);
not \U$14573 ( \14819 , \14818 );
not \U$14574 ( \14820 , \8887 );
or \U$14575 ( \14821 , \14819 , \14820 );
nand \U$14576 ( \14822 , \1199 , \14389 );
nand \U$14577 ( \14823 , \14821 , \14822 );
xor \U$14578 ( \14824 , RIbe28a98_34, RIbe2a2f8_86);
not \U$14579 ( \14825 , \14824 );
not \U$14580 ( \14826 , \8695 );
buf \U$14581 ( \14827 , \14826 );
not \U$14582 ( \14828 , \14827 );
or \U$14583 ( \14829 , \14825 , \14828 );
nand \U$14584 ( \14830 , \8705 , \14771 );
nand \U$14585 ( \14831 , \14829 , \14830 );
nor \U$14586 ( \14832 , \14823 , \14831 );
not \U$14587 ( \14833 , \14832 );
nand \U$14588 ( \14834 , \14823 , \14831 );
nand \U$14589 ( \14835 , \14833 , \14834 );
xor \U$14590 ( \14836 , RIbe27c10_3, RIbe2ad48_108);
and \U$14591 ( \14837 , \936 , \14836 );
and \U$14592 ( \14838 , \370 , \14339 );
nor \U$14593 ( \14839 , \14837 , \14838 );
not \U$14594 ( \14840 , \14839 );
and \U$14595 ( \14841 , \14835 , \14840 );
not \U$14596 ( \14842 , \14835 );
and \U$14597 ( \14843 , \14842 , \14839 );
nor \U$14598 ( \14844 , \14841 , \14843 );
xor \U$14599 ( \14845 , RIbe2af28_112, RIbe2b1f8_118);
not \U$14600 ( \14846 , \14845 );
not \U$14601 ( \14847 , \14846 );
xnor \U$14602 ( \14848 , RIbe2af28_112, RIbe2b1f8_118);
xor \U$14603 ( \14849 , RIbe2b1f8_118, RIbe2b180_117);
nand \U$14604 ( \14850 , \14848 , \14849 );
not \U$14605 ( \14851 , \14850 );
buf \U$14606 ( \14852 , \14851 );
not \U$14607 ( \14853 , \14852 );
not \U$14608 ( \14854 , \14853 );
or \U$14609 ( \14855 , \14847 , \14854 );
nand \U$14610 ( \14856 , \14855 , RIbe2b180_117);
xor \U$14611 ( \14857 , RIbe294e8_56, RIbe2a028_80);
not \U$14612 ( \14858 , \14857 );
not \U$14613 ( \14859 , \14513 );
or \U$14614 ( \14860 , \14858 , \14859 );
nand \U$14615 ( \14861 , \8172 , \14778 );
nand \U$14616 ( \14862 , \14860 , \14861 );
not \U$14617 ( \14863 , \14300 );
not \U$14618 ( \14864 , \14297 );
or \U$14619 ( \14865 , \14863 , \14864 );
nand \U$14620 ( \14866 , \13534 , \13518 );
nand \U$14621 ( \14867 , \14865 , \14866 );
xor \U$14622 ( \14868 , \14862 , \14867 );
xor \U$14623 ( \14869 , \14856 , \14868 );
xnor \U$14624 ( \14870 , \14844 , \14869 );
not \U$14625 ( \14871 , \14870 );
or \U$14626 ( \14872 , \14817 , \14871 );
not \U$14627 ( \14873 , \14844 );
nand \U$14628 ( \14874 , \14873 , \14869 );
nand \U$14629 ( \14875 , \14872 , \14874 );
not \U$14630 ( \14876 , \14875 );
nand \U$14631 ( \14877 , \14792 , \14876 );
not \U$14632 ( \14878 , \14877 );
or \U$14633 ( \14879 , \14727 , \14878 );
nand \U$14634 ( \14880 , \14875 , \14791 );
nand \U$14635 ( \14881 , \14879 , \14880 );
not \U$14636 ( \14882 , \14881 );
xnor \U$14637 ( \14883 , \13468 , \13449 );
not \U$14638 ( \14884 , \13434 );
and \U$14639 ( \14885 , \13426 , \14884 );
not \U$14640 ( \14886 , \13426 );
and \U$14641 ( \14887 , \14886 , \13434 );
nor \U$14642 ( \14888 , \14885 , \14887 );
buf \U$14643 ( \14889 , \14888 );
xor \U$14644 ( \14890 , \14883 , \14889 );
not \U$14645 ( \14891 , \13389 );
not \U$14646 ( \14892 , \13409 );
or \U$14647 ( \14893 , \14891 , \14892 );
or \U$14648 ( \14894 , \13409 , \13389 );
nand \U$14649 ( \14895 , \14893 , \14894 );
buf \U$14650 ( \14896 , \14895 );
xor \U$14651 ( \14897 , \14890 , \14896 );
not \U$14652 ( \14898 , \14897 );
not \U$14653 ( \14899 , \14898 );
xor \U$14654 ( \14900 , \13308 , \13315 );
not \U$14655 ( \14901 , \13300 );
and \U$14656 ( \14902 , \14900 , \14901 );
not \U$14657 ( \14903 , \14900 );
and \U$14658 ( \14904 , \14903 , \13300 );
nor \U$14659 ( \14905 , \14902 , \14904 );
not \U$14660 ( \14906 , \14905 );
xor \U$14661 ( \14907 , \13116 , \13124 );
xnor \U$14662 ( \14908 , \14907 , \13133 );
not \U$14663 ( \14909 , \14908 );
nand \U$14664 ( \14910 , \14906 , \14909 );
nand \U$14665 ( \14911 , \14908 , \14905 );
nand \U$14666 ( \14912 , \14910 , \14911 );
or \U$14667 ( \14913 , \13291 , \13272 );
nand \U$14668 ( \14914 , \14913 , \13292 );
not \U$14669 ( \14915 , \13288 );
and \U$14670 ( \14916 , \14914 , \14915 );
not \U$14671 ( \14917 , \14914 );
and \U$14672 ( \14918 , \14917 , \13288 );
nor \U$14673 ( \14919 , \14916 , \14918 );
xor \U$14674 ( \14920 , \14912 , \14919 );
not \U$14675 ( \14921 , \14920 );
not \U$14676 ( \14922 , \14921 );
or \U$14677 ( \14923 , \14899 , \14922 );
nand \U$14678 ( \14924 , \14897 , \14920 );
nand \U$14679 ( \14925 , \14923 , \14924 );
not \U$14680 ( \14926 , \13536 );
and \U$14681 ( \14927 , RIbe2a640_93, RIbe27b98_2);
not \U$14682 ( \14928 , \14927 );
and \U$14683 ( \14929 , \14926 , \14928 );
and \U$14684 ( \14930 , \13536 , \14927 );
nor \U$14685 ( \14931 , \14929 , \14930 );
not \U$14686 ( \14932 , \14931 );
xor \U$14687 ( \14933 , RIbe28840_29, RIbe2a190_83);
not \U$14688 ( \14934 , \14933 );
not \U$14689 ( \14935 , \14730 );
or \U$14690 ( \14936 , \14934 , \14935 );
nand \U$14691 ( \14937 , \13278 , \14728 );
nand \U$14692 ( \14938 , \14936 , \14937 );
not \U$14693 ( \14939 , \14938 );
xor \U$14694 ( \14940 , RIbe2a280_85, RIbe286d8_26);
not \U$14695 ( \14941 , \14940 );
not \U$14696 ( \14942 , \11344 );
not \U$14697 ( \14943 , \14942 );
or \U$14698 ( \14944 , \14941 , \14943 );
nand \U$14699 ( \14945 , \14649 , \14380 );
nand \U$14700 ( \14946 , \14944 , \14945 );
not \U$14701 ( \14947 , \14946 );
or \U$14702 ( \14948 , \14939 , \14947 );
or \U$14703 ( \14949 , \14946 , \14938 );
xor \U$14704 ( \14950 , RIbe28228_16, RIbe2b6a8_128);
not \U$14705 ( \14951 , \14950 );
not \U$14706 ( \14952 , \879 );
or \U$14707 ( \14953 , \14951 , \14952 );
nand \U$14708 ( \14954 , \885 , \14333 );
nand \U$14709 ( \14955 , \14953 , \14954 );
nand \U$14710 ( \14956 , \14949 , \14955 );
nand \U$14711 ( \14957 , \14948 , \14956 );
not \U$14712 ( \14958 , \14957 );
or \U$14713 ( \14959 , \14932 , \14958 );
or \U$14714 ( \14960 , \14931 , \14957 );
nand \U$14715 ( \14961 , \14959 , \14960 );
xor \U$14716 ( \14962 , RIbe29380_53, RIbe2b180_117);
not \U$14717 ( \14963 , \14962 );
not \U$14718 ( \14964 , \14852 );
or \U$14719 ( \14965 , \14963 , \14964 );
buf \U$14720 ( \14966 , \14845 );
nand \U$14721 ( \14967 , \14966 , RIbe2b180_117);
nand \U$14722 ( \14968 , \14965 , \14967 );
not \U$14723 ( \14969 , \14968 );
not \U$14724 ( \14970 , \14664 );
and \U$14725 ( \14971 , \4573 , \4574 );
not \U$14726 ( \14972 , \14971 );
or \U$14727 ( \14973 , \14970 , \14972 );
xor \U$14728 ( \14974 , RIbe29c68_72, RIbe297b8_62);
nand \U$14729 ( \14975 , \4580 , \14974 );
nand \U$14730 ( \14976 , \14973 , \14975 );
not \U$14731 ( \14977 , \14672 );
not \U$14732 ( \14978 , \2552 );
or \U$14733 ( \14979 , \14977 , \14978 );
xor \U$14734 ( \14980 , RIbe27b20_1, RIbe28b88_36);
nand \U$14735 ( \14981 , \2559 , \14980 );
nand \U$14736 ( \14982 , \14979 , \14981 );
and \U$14737 ( \14983 , \14976 , \14982 );
not \U$14738 ( \14984 , \14976 );
not \U$14739 ( \14985 , \14982 );
and \U$14740 ( \14986 , \14984 , \14985 );
nor \U$14741 ( \14987 , \14983 , \14986 );
not \U$14742 ( \14988 , \14987 );
or \U$14743 ( \14989 , \14969 , \14988 );
nand \U$14744 ( \14990 , \14982 , \14976 );
nand \U$14745 ( \14991 , \14989 , \14990 );
not \U$14746 ( \14992 , \14991 );
not \U$14747 ( \14993 , \14449 );
not \U$14748 ( \14994 , \8813 );
or \U$14749 ( \14995 , \14993 , \14994 );
not \U$14750 ( \14996 , RIbe27df0_7);
not \U$14751 ( \14997 , RIbe285e8_24);
and \U$14752 ( \14998 , \14996 , \14997 );
and \U$14753 ( \14999 , RIbe27df0_7, RIbe285e8_24);
nor \U$14754 ( \15000 , \14998 , \14999 );
nand \U$14755 ( \15001 , \8270 , \15000 );
nand \U$14756 ( \15002 , \14995 , \15001 );
not \U$14757 ( \15003 , \15002 );
not \U$14758 ( \15004 , \14532 );
not \U$14759 ( \15005 , \2457 );
or \U$14760 ( \15006 , \15004 , \15005 );
nand \U$14761 ( \15007 , \2463 , \14798 );
nand \U$14762 ( \15008 , \15006 , \15007 );
buf \U$14763 ( \15009 , \382 );
nand \U$14764 ( \15010 , \15009 , \14620 );
or \U$14765 ( \15011 , \15010 , \398 );
xor \U$14766 ( \15012 , RIbe290b0_47, RIbe2b2e8_120);
nand \U$14767 ( \15013 , \398 , \15012 );
nand \U$14768 ( \15014 , \15011 , \15013 );
xor \U$14769 ( \15015 , \15008 , \15014 );
not \U$14770 ( \15016 , \15015 );
or \U$14771 ( \15017 , \15003 , \15016 );
nand \U$14772 ( \15018 , \15008 , \15014 );
nand \U$14773 ( \15019 , \15017 , \15018 );
xor \U$14774 ( \15020 , \14302 , \15019 );
not \U$14775 ( \15021 , \15020 );
or \U$14776 ( \15022 , \14992 , \15021 );
nand \U$14777 ( \15023 , \15019 , \14302 );
nand \U$14778 ( \15024 , \15022 , \15023 );
xor \U$14779 ( \15025 , \14961 , \15024 );
not \U$14780 ( \15026 , \14633 );
nor \U$14781 ( \15027 , \15026 , \1254 );
and \U$14782 ( \15028 , \1937 , \14276 );
nor \U$14783 ( \15029 , \15027 , \15028 );
not \U$14784 ( \15030 , \15029 );
not \U$14785 ( \15031 , \15030 );
not \U$14786 ( \15032 , \14547 );
not \U$14787 ( \15033 , \8887 );
or \U$14788 ( \15034 , \15032 , \15033 );
nand \U$14789 ( \15035 , \970 , \14818 );
nand \U$14790 ( \15036 , \15034 , \15035 );
not \U$14791 ( \15037 , \14407 );
not \U$14792 ( \15038 , \14826 );
or \U$14793 ( \15039 , \15037 , \15038 );
nand \U$14794 ( \15040 , \8705 , \14824 );
nand \U$14795 ( \15041 , \15039 , \15040 );
xor \U$14796 ( \15042 , \15036 , \15041 );
not \U$14797 ( \15043 , \15042 );
or \U$14798 ( \15044 , \15031 , \15043 );
nand \U$14799 ( \15045 , \15041 , \15036 );
nand \U$14800 ( \15046 , \15044 , \15045 );
not \U$14801 ( \15047 , \15046 );
not \U$14802 ( \15048 , \2518 );
xnor \U$14803 ( \15049 , RIbe28480_21, RIbe29998_66);
or \U$14804 ( \15050 , \15048 , \15049 );
xor \U$14805 ( \15051 , RIbe28480_21, RIbe28d68_40);
not \U$14806 ( \15052 , \15051 );
or \U$14807 ( \15053 , \2670 , \15052 );
nand \U$14808 ( \15054 , \15050 , \15053 );
not \U$14809 ( \15055 , \15054 );
not \U$14810 ( \15056 , \14641 );
not \U$14811 ( \15057 , RIbe29560_57);
xor \U$14812 ( \15058 , RIbe28228_16, \15057 );
nor \U$14813 ( \15059 , \15058 , \877 );
not \U$14814 ( \15060 , \15059 );
or \U$14815 ( \15061 , \15056 , \15060 );
nand \U$14816 ( \15062 , \885 , \14950 );
nand \U$14817 ( \15063 , \15061 , \15062 );
not \U$14818 ( \15064 , \14516 );
not \U$14819 ( \15065 , \8400 );
or \U$14820 ( \15066 , \15064 , \15065 );
nand \U$14821 ( \15067 , \8930 , \14857 );
nand \U$14822 ( \15068 , \15066 , \15067 );
not \U$14823 ( \15069 , \15068 );
xnor \U$14824 ( \15070 , \15063 , \15069 );
not \U$14825 ( \15071 , \15070 );
or \U$14826 ( \15072 , \15055 , \15071 );
not \U$14827 ( \15073 , \15069 );
nand \U$14828 ( \15074 , \15073 , \15063 );
nand \U$14829 ( \15075 , \15072 , \15074 );
xor \U$14830 ( \15076 , RIbe28de0_41, RIbe2a6b8_94);
not \U$14831 ( \15077 , \15076 );
not \U$14832 ( \15078 , \331 );
or \U$14833 ( \15079 , \15077 , \15078 );
xor \U$14834 ( \15080 , RIbe28de0_41, RIbe2b4c8_124);
nand \U$14835 ( \15081 , \347 , \15080 );
nand \U$14836 ( \15082 , \15079 , \15081 );
not \U$14837 ( \15083 , \15082 );
not \U$14838 ( \15084 , \14434 );
not \U$14839 ( \15085 , \11907 );
or \U$14840 ( \15086 , \15084 , \15085 );
nand \U$14841 ( \15087 , \1173 , \14836 );
nand \U$14842 ( \15088 , \15086 , \15087 );
nand \U$14843 ( \15089 , RIbe27b98_2, RIbe2abe0_105);
and \U$14844 ( \15090 , \15088 , \15089 );
not \U$14845 ( \15091 , \15088 );
not \U$14846 ( \15092 , \15089 );
and \U$14847 ( \15093 , \15091 , \15092 );
or \U$14848 ( \15094 , \15090 , \15093 );
not \U$14849 ( \15095 , \15094 );
or \U$14850 ( \15096 , \15083 , \15095 );
nand \U$14851 ( \15097 , \15088 , \15092 );
nand \U$14852 ( \15098 , \15096 , \15097 );
or \U$14853 ( \15099 , \15075 , \15098 );
not \U$14854 ( \15100 , \15099 );
or \U$14855 ( \15101 , \15047 , \15100 );
nand \U$14856 ( \15102 , \15075 , \15098 );
nand \U$14857 ( \15103 , \15101 , \15102 );
and \U$14858 ( \15104 , \15025 , \15103 );
and \U$14859 ( \15105 , \14961 , \15024 );
or \U$14860 ( \15106 , \15104 , \15105 );
xnor \U$14861 ( \15107 , \14925 , \15106 );
not \U$14862 ( \15108 , \15107 );
or \U$14863 ( \15109 , \14882 , \15108 );
or \U$14864 ( \15110 , \14881 , \15107 );
nand \U$14865 ( \15111 , \15109 , \15110 );
not \U$14866 ( \15112 , \15111 );
or \U$14867 ( \15113 , \14706 , \15112 );
not \U$14868 ( \15114 , \15107 );
nand \U$14869 ( \15115 , \15114 , \14881 );
nand \U$14870 ( \15116 , \15113 , \15115 );
not \U$14871 ( \15117 , \15116 );
not \U$14872 ( \15118 , \14911 );
not \U$14873 ( \15119 , \14919 );
or \U$14874 ( \15120 , \15118 , \15119 );
nand \U$14875 ( \15121 , \15120 , \14910 );
not \U$14876 ( \15122 , \14888 );
not \U$14877 ( \15123 , \14883 );
or \U$14878 ( \15124 , \15122 , \15123 );
nand \U$14879 ( \15125 , \15124 , \14895 );
or \U$14880 ( \15126 , \14888 , \14883 );
nand \U$14881 ( \15127 , \15125 , \15126 );
and \U$14882 ( \15128 , \15121 , \15127 );
not \U$14883 ( \15129 , \15121 );
not \U$14884 ( \15130 , \15127 );
and \U$14885 ( \15131 , \15129 , \15130 );
nor \U$14886 ( \15132 , \15128 , \15131 );
nand \U$14887 ( \15133 , \13161 , \13168 );
not \U$14888 ( \15134 , \13163 );
and \U$14889 ( \15135 , \15133 , \15134 );
not \U$14890 ( \15136 , \15133 );
and \U$14891 ( \15137 , \15136 , \13163 );
nor \U$14892 ( \15138 , \15135 , \15137 );
xor \U$14893 ( \15139 , \15132 , \15138 );
not \U$14894 ( \15140 , \14761 );
not \U$14895 ( \15141 , \14768 );
or \U$14896 ( \15142 , \15140 , \15141 );
or \U$14897 ( \15143 , \14768 , \14761 );
nand \U$14898 ( \15144 , \15143 , \14755 );
nand \U$14899 ( \15145 , \15142 , \15144 );
xor \U$14900 ( \15146 , \14735 , \14741 );
and \U$14901 ( \15147 , \15146 , \14748 );
and \U$14902 ( \15148 , \14735 , \14741 );
or \U$14903 ( \15149 , \15147 , \15148 );
xor \U$14904 ( \15150 , \15145 , \15149 );
not \U$14905 ( \15151 , \14365 );
not \U$14906 ( \15152 , \15151 );
not \U$14907 ( \15153 , \14360 );
or \U$14908 ( \15154 , \15152 , \15153 );
nand \U$14909 ( \15155 , \14353 , \14359 );
nand \U$14910 ( \15156 , \15154 , \15155 );
xor \U$14911 ( \15157 , \15150 , \15156 );
not \U$14912 ( \15158 , \14720 );
not \U$14913 ( \15159 , \14718 );
or \U$14914 ( \15160 , \15158 , \15159 );
nand \U$14915 ( \15161 , \14713 , \14709 );
nand \U$14916 ( \15162 , \15160 , \15161 );
xor \U$14917 ( \15163 , \15157 , \15162 );
xor \U$14918 ( \15164 , \14379 , \14387 );
and \U$14919 ( \15165 , \15164 , \14394 );
and \U$14920 ( \15166 , \14379 , \14387 );
or \U$14921 ( \15167 , \15165 , \15166 );
not \U$14922 ( \15168 , \14777 );
not \U$14923 ( \15169 , \14789 );
or \U$14924 ( \15170 , \15168 , \15169 );
nand \U$14925 ( \15171 , \14783 , \14788 );
nand \U$14926 ( \15172 , \15170 , \15171 );
not \U$14927 ( \15173 , \14332 );
not \U$14928 ( \15174 , \14345 );
or \U$14929 ( \15175 , \15173 , \15174 );
nand \U$14930 ( \15176 , \14338 , \14344 );
nand \U$14931 ( \15177 , \15175 , \15176 );
xor \U$14932 ( \15178 , \15172 , \15177 );
xor \U$14933 ( \15179 , \15167 , \15178 );
and \U$14934 ( \15180 , \15163 , \15179 );
and \U$14935 ( \15181 , \15157 , \15162 );
or \U$14936 ( \15182 , \15180 , \15181 );
xor \U$14937 ( \15183 , \15139 , \15182 );
xor \U$14938 ( \15184 , \13329 , \13347 );
xor \U$14939 ( \15185 , \13367 , \13360 );
xnor \U$14940 ( \15186 , \15185 , \13376 );
not \U$14941 ( \15187 , \15186 );
xor \U$14942 ( \15188 , \15184 , \15187 );
not \U$14943 ( \15189 , \13261 );
not \U$14944 ( \15190 , \13243 );
not \U$14945 ( \15191 , \13253 );
or \U$14946 ( \15192 , \15190 , \15191 );
or \U$14947 ( \15193 , \13253 , \13243 );
nand \U$14948 ( \15194 , \15192 , \15193 );
not \U$14949 ( \15195 , \15194 );
or \U$14950 ( \15196 , \15189 , \15195 );
or \U$14951 ( \15197 , \15194 , \13261 );
nand \U$14952 ( \15198 , \15196 , \15197 );
not \U$14953 ( \15199 , \15198 );
xor \U$14954 ( \15200 , \15188 , \15199 );
not \U$14955 ( \15201 , \15200 );
xor \U$14956 ( \15202 , \14749 , \14769 );
and \U$14957 ( \15203 , \15202 , \14790 );
and \U$14958 ( \15204 , \14749 , \14769 );
or \U$14959 ( \15205 , \15203 , \15204 );
not \U$14960 ( \15206 , \14395 );
not \U$14961 ( \15207 , \14373 );
or \U$14962 ( \15208 , \15206 , \15207 );
not \U$14963 ( \15209 , \14369 );
nand \U$14964 ( \15210 , \15209 , \14346 );
nand \U$14965 ( \15211 , \15208 , \15210 );
xor \U$14966 ( \15212 , \15205 , \15211 );
not \U$14967 ( \15213 , \15212 );
or \U$14968 ( \15214 , \15201 , \15213 );
nand \U$14969 ( \15215 , \15211 , \15205 );
nand \U$14970 ( \15216 , \15214 , \15215 );
xnor \U$14971 ( \15217 , \15183 , \15216 );
not \U$14972 ( \15218 , \15217 );
and \U$14973 ( \15219 , \15117 , \15218 );
and \U$14974 ( \15220 , \15116 , \15217 );
nor \U$14975 ( \15221 , \15219 , \15220 );
not \U$14976 ( \15222 , \13318 );
xnor \U$14977 ( \15223 , \13293 , \13265 );
not \U$14978 ( \15224 , \15223 );
or \U$14979 ( \15225 , \15222 , \15224 );
or \U$14980 ( \15226 , \13318 , \15223 );
nand \U$14981 ( \15227 , \15225 , \15226 );
xor \U$14982 ( \15228 , \11350 , \13378 );
xnor \U$14983 ( \15229 , \15228 , \13352 );
not \U$14984 ( \15230 , \15199 );
not \U$14985 ( \15231 , \15187 );
or \U$14986 ( \15232 , \15230 , \15231 );
not \U$14987 ( \15233 , \15186 );
not \U$14988 ( \15234 , \15198 );
or \U$14989 ( \15235 , \15233 , \15234 );
nand \U$14990 ( \15236 , \15235 , \15184 );
nand \U$14991 ( \15237 , \15232 , \15236 );
nor \U$14992 ( \15238 , \15229 , \15237 );
not \U$14993 ( \15239 , \15238 );
nand \U$14994 ( \15240 , \15229 , \15237 );
nand \U$14995 ( \15241 , \15239 , \15240 );
xor \U$14996 ( \15242 , \15227 , \15241 );
not \U$14997 ( \15243 , \15106 );
not \U$14998 ( \15244 , \14925 );
or \U$14999 ( \15245 , \15243 , \15244 );
nand \U$15000 ( \15246 , \14897 , \14921 );
nand \U$15001 ( \15247 , \15245 , \15246 );
xor \U$15002 ( \15248 , \15242 , \15247 );
not \U$15003 ( \15249 , \15248 );
not \U$15004 ( \15250 , \14931 );
nand \U$15005 ( \15251 , \15250 , \14957 );
not \U$15006 ( \15252 , \13536 );
nand \U$15007 ( \15253 , \15252 , \14927 );
and \U$15008 ( \15254 , \15251 , \15253 );
xor \U$15009 ( \15255 , \13547 , \13517 );
and \U$15010 ( \15256 , \15255 , \13536 );
not \U$15011 ( \15257 , \15255 );
and \U$15012 ( \15258 , \15257 , \15252 );
nor \U$15013 ( \15259 , \15256 , \15258 );
not \U$15014 ( \15260 , \15259 );
nand \U$15015 ( \15261 , \15254 , \15260 );
not \U$15016 ( \15262 , \15261 );
not \U$15017 ( \15263 , \14856 );
not \U$15018 ( \15264 , \14868 );
or \U$15019 ( \15265 , \15263 , \15264 );
nand \U$15020 ( \15266 , \14867 , \14862 );
nand \U$15021 ( \15267 , \15265 , \15266 );
not \U$15022 ( \15268 , \15267 );
xor \U$15023 ( \15269 , RIbe29128_48, RIbe27fd0_11);
not \U$15024 ( \15270 , \15269 );
not \U$15025 ( \15271 , \12808 );
or \U$15026 ( \15272 , \15270 , \15271 );
nand \U$15027 ( \15273 , \2707 , \14374 );
nand \U$15028 ( \15274 , \15272 , \15273 );
not \U$15029 ( \15275 , \15274 );
xor \U$15030 ( \15276 , RIbe27d78_6, RIbe2a460_89);
not \U$15031 ( \15277 , \15276 );
not \U$15032 ( \15278 , \8768 );
or \U$15033 ( \15279 , \15277 , \15278 );
nand \U$15034 ( \15280 , \314 , \13587 );
nand \U$15035 ( \15281 , \15279 , \15280 );
xor \U$15036 ( \15282 , RIbe2a640_93, RIbe27b98_2);
not \U$15037 ( \15283 , \15282 );
not \U$15038 ( \15284 , \8380 );
or \U$15039 ( \15285 , \15283 , \15284 );
nand \U$15040 ( \15286 , \7585 , \13615 );
nand \U$15041 ( \15287 , \15285 , \15286 );
xor \U$15042 ( \15288 , \15281 , \15287 );
not \U$15043 ( \15289 , \15288 );
or \U$15044 ( \15290 , \15275 , \15289 );
nand \U$15045 ( \15291 , \15287 , \15281 );
nand \U$15046 ( \15292 , \15290 , \15291 );
not \U$15047 ( \15293 , \15051 );
not \U$15048 ( \15294 , \3483 );
or \U$15049 ( \15295 , \15293 , \15294 );
nand \U$15050 ( \15296 , \2527 , \14362 );
nand \U$15051 ( \15297 , \15295 , \15296 );
not \U$15052 ( \15298 , \15297 );
and \U$15053 ( \15299 , RIbe2ac58_106, RIbe27b98_2);
not \U$15054 ( \15300 , \15299 );
not \U$15055 ( \15301 , \15080 );
not \U$15056 ( \15302 , \11321 );
or \U$15057 ( \15303 , \15301 , \15302 );
nand \U$15058 ( \15304 , \346 , \14348 );
nand \U$15059 ( \15305 , \15303 , \15304 );
not \U$15060 ( \15306 , \15305 );
nand \U$15061 ( \15307 , \15300 , \15306 );
not \U$15062 ( \15308 , \15307 );
or \U$15063 ( \15309 , \15298 , \15308 );
nand \U$15064 ( \15310 , \15305 , \15299 );
nand \U$15065 ( \15311 , \15309 , \15310 );
xor \U$15066 ( \15312 , \15292 , \15311 );
not \U$15067 ( \15313 , \15312 );
or \U$15068 ( \15314 , \15268 , \15313 );
nand \U$15069 ( \15315 , \15292 , \15311 );
nand \U$15070 ( \15316 , \15314 , \15315 );
not \U$15071 ( \15317 , \15316 );
or \U$15072 ( \15318 , \15262 , \15317 );
or \U$15073 ( \15319 , \15254 , \15260 );
nand \U$15074 ( \15320 , \15318 , \15319 );
and \U$15075 ( \15321 , \13216 , \13207 );
not \U$15076 ( \15322 , \13216 );
and \U$15077 ( \15323 , \15322 , \13218 );
or \U$15078 ( \15324 , \15321 , \15323 );
and \U$15079 ( \15325 , \15324 , \13219 );
not \U$15080 ( \15326 , \15324 );
and \U$15081 ( \15327 , \15326 , \13199 );
nor \U$15082 ( \15328 , \15325 , \15327 );
not \U$15083 ( \15329 , \15328 );
xnor \U$15084 ( \15330 , \13146 , \13109 );
not \U$15085 ( \15331 , \15330 );
or \U$15086 ( \15332 , \15329 , \15331 );
or \U$15087 ( \15333 , \15328 , \15330 );
nand \U$15088 ( \15334 , \15332 , \15333 );
xnor \U$15089 ( \15335 , \15320 , \15334 );
not \U$15090 ( \15336 , \15335 );
and \U$15091 ( \15337 , \15249 , \15336 );
and \U$15092 ( \15338 , \15248 , \15335 );
nor \U$15093 ( \15339 , \15337 , \15338 );
not \U$15094 ( \15340 , \15339 );
xor \U$15095 ( \15341 , \15221 , \15340 );
not \U$15096 ( \15342 , \15341 );
xor \U$15097 ( \15343 , RIbe29380_53, RIbe2af28_112);
not \U$15098 ( \15344 , \15343 );
buf \U$15099 ( \15345 , \14423 );
not \U$15100 ( \15346 , \15345 );
or \U$15101 ( \15347 , \15344 , \15346 );
not \U$15102 ( \15348 , \14414 );
nand \U$15103 ( \15349 , \15348 , RIbe2af28_112);
nand \U$15104 ( \15350 , \15347 , \15349 );
xor \U$15105 ( \15351 , RIbe2b180_117, RIbe28048_12);
not \U$15106 ( \15352 , \15351 );
buf \U$15107 ( \15353 , \14851 );
not \U$15108 ( \15354 , \15353 );
or \U$15109 ( \15355 , \15352 , \15354 );
nand \U$15110 ( \15356 , \14966 , \14962 );
nand \U$15111 ( \15357 , \15355 , \15356 );
xor \U$15112 ( \15358 , \15350 , \15357 );
xor \U$15113 ( \15359 , RIbe285e8_24, RIbe29998_66);
not \U$15114 ( \15360 , \15359 );
not \U$15115 ( \15361 , \8267 );
or \U$15116 ( \15362 , \15360 , \15361 );
not \U$15117 ( \15363 , \14447 );
nand \U$15118 ( \15364 , \15363 , \8270 );
nand \U$15119 ( \15365 , \15362 , \15364 );
not \U$15120 ( \15366 , \15365 );
xor \U$15121 ( \15367 , RIbe2adc0_109, RIbe290b0_47);
not \U$15122 ( \15368 , \15367 );
not \U$15123 ( \15369 , \2730 );
or \U$15124 ( \15370 , \15368 , \15369 );
nand \U$15125 ( \15371 , \398 , \14616 );
nand \U$15126 ( \15372 , \15370 , \15371 );
not \U$15127 ( \15373 , \15372 );
or \U$15128 ( \15374 , \15366 , \15373 );
not \U$15129 ( \15375 , \15372 );
not \U$15130 ( \15376 , \15375 );
not \U$15131 ( \15377 , \15365 );
not \U$15132 ( \15378 , \15377 );
or \U$15133 ( \15379 , \15376 , \15378 );
xor \U$15134 ( \15380 , RIbe27ee0_9, RIbe2b180_117);
not \U$15135 ( \15381 , \15380 );
not \U$15136 ( \15382 , \14852 );
or \U$15137 ( \15383 , \15381 , \15382 );
nand \U$15138 ( \15384 , \14966 , \15351 );
nand \U$15139 ( \15385 , \15383 , \15384 );
nand \U$15140 ( \15386 , \15379 , \15385 );
nand \U$15141 ( \15387 , \15374 , \15386 );
and \U$15142 ( \15388 , \15358 , \15387 );
and \U$15143 ( \15389 , \15350 , \15357 );
or \U$15144 ( \15390 , \15388 , \15389 );
not \U$15145 ( \15391 , \15390 );
not \U$15146 ( \15392 , \15391 );
xor \U$15147 ( \15393 , RIbe2a910_99, RIbe293f8_54);
not \U$15148 ( \15394 , \15393 );
buf \U$15149 ( \15395 , \10987 );
not \U$15150 ( \15396 , \15395 );
or \U$15151 ( \15397 , \15394 , \15396 );
nand \U$15152 ( \15398 , \10401 , \14454 );
nand \U$15153 ( \15399 , \15397 , \15398 );
not \U$15154 ( \15400 , \15399 );
nand \U$15155 ( \15401 , RIbe27b98_2, RIbe2a730_95);
not \U$15156 ( \15402 , \15401 );
xor \U$15157 ( \15403 , RIbe29740_61, RIbe29e48_76);
not \U$15158 ( \15404 , \15403 );
not \U$15159 ( \15405 , \11039 );
or \U$15160 ( \15406 , \15404 , \15405 );
nand \U$15161 ( \15407 , \7368 , \14586 );
nand \U$15162 ( \15408 , \15406 , \15407 );
not \U$15163 ( \15409 , \15408 );
or \U$15164 ( \15410 , \15402 , \15409 );
or \U$15165 ( \15411 , \15408 , \15401 );
nand \U$15166 ( \15412 , \15410 , \15411 );
not \U$15167 ( \15413 , \15412 );
or \U$15168 ( \15414 , \15400 , \15413 );
not \U$15169 ( \15415 , \15401 );
nand \U$15170 ( \15416 , \15415 , \15408 );
nand \U$15171 ( \15417 , \15414 , \15416 );
not \U$15172 ( \15418 , \15417 );
xor \U$15173 ( \15419 , RIbe2a028_80, RIbe28138_14);
not \U$15174 ( \15420 , \15419 );
not \U$15175 ( \15421 , \8401 );
or \U$15176 ( \15422 , \15420 , \15421 );
nand \U$15177 ( \15423 , \8930 , \14511 );
nand \U$15178 ( \15424 , \15422 , \15423 );
xor \U$15179 ( \15425 , RIbe28de0_41, RIbe2ac58_106);
not \U$15180 ( \15426 , \15425 );
not \U$15181 ( \15427 , \923 );
or \U$15182 ( \15428 , \15426 , \15427 );
xor \U$15183 ( \15429 , RIbe28de0_41, RIbe2a640_93);
nand \U$15184 ( \15430 , \7472 , \15429 );
nand \U$15185 ( \15431 , \15428 , \15430 );
or \U$15186 ( \15432 , \15424 , \15431 );
xor \U$15187 ( \15433 , RIbe29470_55, RIbe2a2f8_86);
not \U$15188 ( \15434 , \15433 );
not \U$15189 ( \15435 , \10792 );
or \U$15190 ( \15436 , \15434 , \15435 );
nand \U$15191 ( \15437 , \11094 , \14403 );
nand \U$15192 ( \15438 , \15436 , \15437 );
nand \U$15193 ( \15439 , \15432 , \15438 );
nand \U$15194 ( \15440 , \15424 , \15431 );
nand \U$15195 ( \15441 , \15439 , \15440 );
xor \U$15196 ( \15442 , RIbe28228_16, RIbe2a898_98);
not \U$15197 ( \15443 , \15442 );
not \U$15198 ( \15444 , \14638 );
or \U$15199 ( \15445 , \15443 , \15444 );
nand \U$15200 ( \15446 , \885 , \14636 );
nand \U$15201 ( \15447 , \15445 , \15446 );
not \U$15202 ( \15448 , \15447 );
xor \U$15203 ( \15449 , RIbe27e68_8, RIbe27c88_4);
not \U$15204 ( \15450 , \15449 );
not \U$15205 ( \15451 , \2458 );
or \U$15206 ( \15452 , \15450 , \15451 );
nand \U$15207 ( \15453 , \2463 , \14528 );
nand \U$15208 ( \15454 , \15452 , \15453 );
not \U$15209 ( \15455 , \15454 );
or \U$15210 ( \15456 , \15448 , \15455 );
or \U$15211 ( \15457 , \15447 , \15454 );
xor \U$15212 ( \15458 , RIbe27c10_3, RIbe2a6b8_94);
not \U$15213 ( \15459 , \15458 );
not \U$15214 ( \15460 , \7440 );
or \U$15215 ( \15461 , \15459 , \15460 );
nand \U$15216 ( \15462 , \1498 , \14430 );
nand \U$15217 ( \15463 , \15461 , \15462 );
nand \U$15218 ( \15464 , \15457 , \15463 );
nand \U$15219 ( \15465 , \15456 , \15464 );
xor \U$15220 ( \15466 , \15441 , \15465 );
not \U$15221 ( \15467 , \15466 );
or \U$15222 ( \15468 , \15418 , \15467 );
nand \U$15223 ( \15469 , \15465 , \15441 );
nand \U$15224 ( \15470 , \15468 , \15469 );
not \U$15225 ( \15471 , \15470 );
or \U$15226 ( \15472 , \15392 , \15471 );
or \U$15227 ( \15473 , \15470 , \15391 );
nand \U$15228 ( \15474 , \15472 , \15473 );
not \U$15229 ( \15475 , \11544 );
not \U$15230 ( \15476 , \15475 );
xor \U$15231 ( \15477 , RIbe2a3e8_88, RIbe288b8_30);
not \U$15232 ( \15478 , \15477 );
or \U$15233 ( \15479 , \15476 , \15478 );
nand \U$15234 ( \15480 , \9268 , \14473 );
nand \U$15235 ( \15481 , \15479 , \15480 );
not \U$15236 ( \15482 , \15481 );
xor \U$15237 ( \15483 , RIbe2aa78_102, RIbe28930_31);
not \U$15238 ( \15484 , \15483 );
not \U$15239 ( \15485 , \965 );
or \U$15240 ( \15486 , \15484 , \15485 );
nand \U$15241 ( \15487 , \1199 , \14543 );
nand \U$15242 ( \15488 , \15486 , \15487 );
xor \U$15243 ( \15489 , RIbe2b360_121, RIbe296c8_60);
not \U$15244 ( \15490 , \15489 );
not \U$15245 ( \15491 , \8531 );
or \U$15246 ( \15492 , \15490 , \15491 );
nand \U$15247 ( \15493 , \1137 , \14629 );
nand \U$15248 ( \15494 , \15492 , \15493 );
and \U$15249 ( \15495 , \15488 , \15494 );
not \U$15250 ( \15496 , \15488 );
not \U$15251 ( \15497 , \15494 );
and \U$15252 ( \15498 , \15496 , \15497 );
nor \U$15253 ( \15499 , \15495 , \15498 );
not \U$15254 ( \15500 , \15499 );
or \U$15255 ( \15501 , \15482 , \15500 );
nand \U$15256 ( \15502 , \15488 , \15494 );
nand \U$15257 ( \15503 , \15501 , \15502 );
not \U$15258 ( \15504 , \15503 );
xor \U$15259 ( \15505 , RIbe2b108_116, RIbe28570_23);
not \U$15260 ( \15506 , \15505 );
not \U$15261 ( \15507 , \14297 );
or \U$15262 ( \15508 , \15506 , \15507 );
nand \U$15263 ( \15509 , \13534 , \14571 );
nand \U$15264 ( \15510 , \15508 , \15509 );
xor \U$15265 ( \15511 , RIbe2b540_125, RIbe27d78_6);
not \U$15266 ( \15512 , \15511 );
not \U$15267 ( \15513 , \2052 );
or \U$15268 ( \15514 , \15512 , \15513 );
nand \U$15269 ( \15515 , \314 , \14562 );
nand \U$15270 ( \15516 , \15514 , \15515 );
xor \U$15271 ( \15517 , \15510 , \15516 );
xor \U$15272 ( \15518 , RIbe28f48_44, RIbe29b00_69);
not \U$15273 ( \15519 , \15518 );
not \U$15274 ( \15520 , \8221 );
or \U$15275 ( \15521 , \15519 , \15520 );
nand \U$15276 ( \15522 , \3249 , \14600 );
nand \U$15277 ( \15523 , \15521 , \15522 );
and \U$15278 ( \15524 , \15517 , \15523 );
and \U$15279 ( \15525 , \15510 , \15516 );
or \U$15280 ( \15526 , \15524 , \15525 );
not \U$15281 ( \15527 , \15526 );
or \U$15282 ( \15528 , \15504 , \15527 );
xor \U$15283 ( \15529 , \15510 , \15516 );
and \U$15284 ( \15530 , \15529 , \15523 );
and \U$15285 ( \15531 , \15510 , \15516 );
or \U$15286 ( \15532 , \15530 , \15531 );
not \U$15287 ( \15533 , \15532 );
not \U$15288 ( \15534 , \15533 );
not \U$15289 ( \15535 , \15503 );
and \U$15290 ( \15536 , \15534 , \15535 );
and \U$15291 ( \15537 , \15503 , \15533 );
nor \U$15292 ( \15538 , \15536 , \15537 );
not \U$15293 ( \15539 , \10434 );
xor \U$15294 ( \15540 , RIbe2a550_91, RIbe28c00_37);
not \U$15295 ( \15541 , \15540 );
or \U$15296 ( \15542 , \15539 , \15541 );
not \U$15297 ( \15543 , \11228 );
not \U$15298 ( \15544 , \14608 );
or \U$15299 ( \15545 , \15543 , \15544 );
nand \U$15300 ( \15546 , \15542 , \15545 );
not \U$15301 ( \15547 , \15546 );
xor \U$15302 ( \15548 , RIbe29f38_78, RIbe28a20_33);
not \U$15303 ( \15549 , \15548 );
not \U$15304 ( \15550 , \2276 );
or \U$15305 ( \15551 , \15549 , \15550 );
nand \U$15306 ( \15552 , \2475 , \14488 );
nand \U$15307 ( \15553 , \15551 , \15552 );
not \U$15308 ( \15554 , \15553 );
xor \U$15309 ( \15555 , RIbe29b78_70, RIbe28390_19);
and \U$15310 ( \15556 , \2640 , \15555 );
and \U$15311 ( \15557 , \2648 , \14577 );
nor \U$15312 ( \15558 , \15556 , \15557 );
not \U$15313 ( \15559 , \15558 );
or \U$15314 ( \15560 , \15554 , \15559 );
or \U$15315 ( \15561 , \15553 , \15558 );
nand \U$15316 ( \15562 , \15560 , \15561 );
not \U$15317 ( \15563 , \15562 );
or \U$15318 ( \15564 , \15547 , \15563 );
not \U$15319 ( \15565 , \15558 );
nand \U$15320 ( \15566 , \15565 , \15553 );
nand \U$15321 ( \15567 , \15564 , \15566 );
not \U$15322 ( \15568 , \15567 );
or \U$15323 ( \15569 , \15538 , \15568 );
nand \U$15324 ( \15570 , \15528 , \15569 );
and \U$15325 ( \15571 , \15474 , \15570 );
and \U$15326 ( \15572 , \15470 , \15390 );
nor \U$15327 ( \15573 , \15571 , \15572 );
not \U$15328 ( \15574 , \15573 );
not \U$15329 ( \15575 , \15574 );
xor \U$15330 ( \15576 , \14946 , \14938 );
xnor \U$15331 ( \15577 , \15576 , \14955 );
not \U$15332 ( \15578 , \15577 );
not \U$15333 ( \15579 , \15012 );
not \U$15334 ( \15580 , \2730 );
or \U$15335 ( \15581 , \15579 , \15580 );
nand \U$15336 ( \15582 , \399 , \14354 );
nand \U$15337 ( \15583 , \15581 , \15582 );
not \U$15338 ( \15584 , \14980 );
or \U$15339 ( \15585 , \2700 , \15584 );
nand \U$15340 ( \15586 , \7549 , \14736 );
nand \U$15341 ( \15587 , \15585 , \15586 );
not \U$15342 ( \15588 , \15587 );
not \U$15343 ( \15589 , \14974 );
not \U$15344 ( \15590 , \14971 );
or \U$15345 ( \15591 , \15589 , \15590 );
nand \U$15346 ( \15592 , \4580 , \13572 );
nand \U$15347 ( \15593 , \15591 , \15592 );
not \U$15348 ( \15594 , \15593 );
not \U$15349 ( \15595 , \15594 );
or \U$15350 ( \15596 , \15588 , \15595 );
or \U$15351 ( \15597 , \15587 , \15594 );
nand \U$15352 ( \15598 , \15596 , \15597 );
xor \U$15353 ( \15599 , \15583 , \15598 );
xor \U$15354 ( \15600 , RIbe280c0_13, RIbe2aa00_101);
not \U$15355 ( \15601 , \15600 );
not \U$15356 ( \15602 , \858 );
or \U$15357 ( \15603 , \15601 , \15602 );
nand \U$15358 ( \15604 , \868 , \13624 );
nand \U$15359 ( \15605 , \15603 , \15604 );
not \U$15360 ( \15606 , \14289 );
not \U$15361 ( \15607 , \8804 );
or \U$15362 ( \15608 , \15606 , \15607 );
nand \U$15363 ( \15609 , \8793 , \13607 );
nand \U$15364 ( \15610 , \15608 , \15609 );
xor \U$15365 ( \15611 , \15605 , \15610 );
not \U$15366 ( \15612 , \15000 );
not \U$15367 ( \15613 , \2761 );
or \U$15368 ( \15614 , \15612 , \15613 );
nand \U$15369 ( \15615 , \8270 , \14756 );
nand \U$15370 ( \15616 , \15614 , \15615 );
xor \U$15371 ( \15617 , \15611 , \15616 );
and \U$15372 ( \15618 , \15599 , \15617 );
not \U$15373 ( \15619 , \15599 );
not \U$15374 ( \15620 , \15617 );
and \U$15375 ( \15621 , \15619 , \15620 );
nor \U$15376 ( \15622 , \15618 , \15621 );
not \U$15377 ( \15623 , \15622 );
or \U$15378 ( \15624 , \15578 , \15623 );
or \U$15379 ( \15625 , \15622 , \15577 );
nand \U$15380 ( \15626 , \15624 , \15625 );
xor \U$15381 ( \15627 , RIbe27fd0_11, RIbe29218_50);
not \U$15382 ( \15628 , \15627 );
not \U$15383 ( \15629 , \4893 );
or \U$15384 ( \15630 , \15628 , \15629 );
nand \U$15385 ( \15631 , \2707 , \14555 );
nand \U$15386 ( \15632 , \15630 , \15631 );
not \U$15387 ( \15633 , \15632 );
not \U$15388 ( \15634 , RIbe2a7a8_96);
and \U$15389 ( \15635 , RIbe27b98_2, \15634 );
not \U$15390 ( \15636 , RIbe27b98_2);
and \U$15391 ( \15637 , \15636 , RIbe2a7a8_96);
or \U$15392 ( \15638 , \15635 , \15637 );
not \U$15393 ( \15639 , \15638 );
not \U$15394 ( \15640 , \256 );
or \U$15395 ( \15641 , \15639 , \15640 );
nand \U$15396 ( \15642 , \7585 , \14520 );
nand \U$15397 ( \15643 , \15641 , \15642 );
not \U$15398 ( \15644 , \15643 );
or \U$15399 ( \15645 , \15633 , \15644 );
or \U$15400 ( \15646 , \15643 , \15632 );
xor \U$15401 ( \15647 , RIbe28cf0_39, RIbe28480_21);
not \U$15402 ( \15648 , \15647 );
not \U$15403 ( \15649 , \3483 );
or \U$15404 ( \15650 , \15648 , \15649 );
xor \U$15405 ( \15651 , RIbe298a8_64, RIbe28480_21);
nand \U$15406 ( \15652 , \11263 , \15651 );
nand \U$15407 ( \15653 , \15650 , \15652 );
nand \U$15408 ( \15654 , \15646 , \15653 );
nand \U$15409 ( \15655 , \15645 , \15654 );
not \U$15410 ( \15656 , \15655 );
xor \U$15411 ( \15657 , RIbe29c68_72, RIbe291a0_49);
not \U$15412 ( \15658 , \15657 );
not \U$15413 ( \15659 , \10720 );
or \U$15414 ( \15660 , \15658 , \15659 );
nand \U$15415 ( \15661 , \4580 , \14660 );
nand \U$15416 ( \15662 , \15660 , \15661 );
not \U$15417 ( \15663 , \15662 );
xor \U$15418 ( \15664 , RIbe28750_27, RIbe2a280_85);
not \U$15419 ( \15665 , \15664 );
not \U$15420 ( \15666 , \14942 );
or \U$15421 ( \15667 , \15665 , \15666 );
nand \U$15422 ( \15668 , \11348 , \14645 );
nand \U$15423 ( \15669 , \15667 , \15668 );
not \U$15424 ( \15670 , \15669 );
or \U$15425 ( \15671 , \15663 , \15670 );
or \U$15426 ( \15672 , \15669 , \15662 );
xor \U$15427 ( \15673 , RIbe2a4d8_90, RIbe29038_46);
not \U$15428 ( \15674 , \15673 );
not \U$15429 ( \15675 , \979 );
or \U$15430 ( \15676 , \15674 , \15675 );
nand \U$15431 ( \15677 , \1583 , \14461 );
nand \U$15432 ( \15678 , \15676 , \15677 );
nand \U$15433 ( \15679 , \15672 , \15678 );
nand \U$15434 ( \15680 , \15671 , \15679 );
not \U$15435 ( \15681 , \15680 );
nand \U$15436 ( \15682 , \15656 , \15681 );
not \U$15437 ( \15683 , \15682 );
not \U$15438 ( \15684 , RIbe28318_18);
not \U$15439 ( \15685 , RIbe2a190_83);
and \U$15440 ( \15686 , \15684 , \15685 );
and \U$15441 ( \15687 , RIbe28318_18, RIbe2a190_83);
nor \U$15442 ( \15688 , \15686 , \15687 );
not \U$15443 ( \15689 , \15688 );
not \U$15444 ( \15690 , \10689 );
not \U$15445 ( \15691 , \15690 );
or \U$15446 ( \15692 , \15689 , \15691 );
buf \U$15447 ( \15693 , \10695 );
nand \U$15448 ( \15694 , \15693 , \14675 );
nand \U$15449 ( \15695 , \15692 , \15694 );
not \U$15450 ( \15696 , \15695 );
xor \U$15451 ( \15697 , RIbe2a118_82, RIbe280c0_13);
not \U$15452 ( \15698 , \15697 );
not \U$15453 ( \15699 , \2379 );
or \U$15454 ( \15700 , \15698 , \15699 );
nand \U$15455 ( \15701 , \2369 , \14480 );
nand \U$15456 ( \15702 , \15700 , \15701 );
xor \U$15457 ( \15703 , RIbe29d58_74, RIbe28b88_36);
not \U$15458 ( \15704 , \15703 );
not \U$15459 ( \15705 , \2553 );
or \U$15460 ( \15706 , \15704 , \15705 );
nand \U$15461 ( \15707 , \7550 , \14668 );
nand \U$15462 ( \15708 , \15706 , \15707 );
xor \U$15463 ( \15709 , \15702 , \15708 );
not \U$15464 ( \15710 , \15709 );
or \U$15465 ( \15711 , \15696 , \15710 );
nand \U$15466 ( \15712 , \15708 , \15702 );
nand \U$15467 ( \15713 , \15711 , \15712 );
not \U$15468 ( \15714 , \15713 );
or \U$15469 ( \15715 , \15683 , \15714 );
nand \U$15470 ( \15716 , \15655 , \15680 );
nand \U$15471 ( \15717 , \15715 , \15716 );
not \U$15472 ( \15718 , \15717 );
not \U$15473 ( \15719 , \14604 );
not \U$15474 ( \15720 , \8221 );
or \U$15475 ( \15721 , \15719 , \15720 );
nand \U$15476 ( \15722 , \11201 , \14249 );
nand \U$15477 ( \15723 , \15721 , \15722 );
not \U$15478 ( \15724 , \14465 );
not \U$15479 ( \15725 , \281 );
or \U$15480 ( \15726 , \15724 , \15725 );
nand \U$15481 ( \15727 , \1583 , \14264 );
nand \U$15482 ( \15728 , \15726 , \15727 );
not \U$15483 ( \15729 , \14524 );
not \U$15484 ( \15730 , \256 );
or \U$15485 ( \15731 , \15729 , \15730 );
nand \U$15486 ( \15732 , \7585 , \15282 );
nand \U$15487 ( \15733 , \15731 , \15732 );
xor \U$15488 ( \15734 , \15728 , \15733 );
xor \U$15489 ( \15735 , \15723 , \15734 );
xor \U$15490 ( \15736 , \14312 , \14291 );
and \U$15491 ( \15737 , \15736 , \14302 );
not \U$15492 ( \15738 , \15736 );
and \U$15493 ( \15739 , \15738 , \14314 );
nor \U$15494 ( \15740 , \15737 , \15739 );
xnor \U$15495 ( \15741 , \15735 , \15740 );
not \U$15496 ( \15742 , \15741 );
or \U$15497 ( \15743 , \15718 , \15742 );
not \U$15498 ( \15744 , \15740 );
xor \U$15499 ( \15745 , \15723 , \15734 );
nand \U$15500 ( \15746 , \15744 , \15745 );
nand \U$15501 ( \15747 , \15743 , \15746 );
xor \U$15502 ( \15748 , \15626 , \15747 );
not \U$15503 ( \15749 , \15748 );
or \U$15504 ( \15750 , \15575 , \15749 );
nand \U$15505 ( \15751 , \15747 , \15626 );
nand \U$15506 ( \15752 , \15750 , \15751 );
xor \U$15507 ( \15753 , \14725 , \14791 );
xor \U$15508 ( \15754 , \15753 , \14876 );
xor \U$15509 ( \15755 , \15752 , \15754 );
xor \U$15510 ( \15756 , \14700 , \14401 );
and \U$15511 ( \15757 , \15755 , \15756 );
not \U$15512 ( \15758 , \15755 );
not \U$15513 ( \15759 , \15756 );
and \U$15514 ( \15760 , \15758 , \15759 );
nor \U$15515 ( \15761 , \15757 , \15760 );
not \U$15516 ( \15762 , \15761 );
not \U$15517 ( \15763 , \14679 );
not \U$15518 ( \15764 , \10689 );
not \U$15519 ( \15765 , \15764 );
or \U$15520 ( \15766 , \15763 , \15765 );
nand \U$15521 ( \15767 , \10834 , \14933 );
nand \U$15522 ( \15768 , \15766 , \15767 );
not \U$15523 ( \15769 , \15768 );
not \U$15524 ( \15770 , \14613 );
not \U$15525 ( \15771 , \11999 );
or \U$15526 ( \15772 , \15770 , \15771 );
nand \U$15527 ( \15773 , \11485 , \14258 );
nand \U$15528 ( \15774 , \15772 , \15773 );
not \U$15529 ( \15775 , \15774 );
or \U$15530 ( \15776 , \15769 , \15775 );
or \U$15531 ( \15777 , \15774 , \15768 );
not \U$15532 ( \15778 , \14582 );
not \U$15533 ( \15779 , \2639 );
or \U$15534 ( \15780 , \15778 , \15779 );
nand \U$15535 ( \15781 , \5831 , \14804 );
nand \U$15536 ( \15782 , \15780 , \15781 );
nand \U$15537 ( \15783 , \15777 , \15782 );
nand \U$15538 ( \15784 , \15776 , \15783 );
not \U$15539 ( \15785 , \15784 );
not \U$15540 ( \15786 , \14552 );
not \U$15541 ( \15787 , \4893 );
or \U$15542 ( \15788 , \15786 , \15787 );
nand \U$15543 ( \15789 , \7709 , \15269 );
nand \U$15544 ( \15790 , \15788 , \15789 );
not \U$15545 ( \15791 , \15790 );
not \U$15546 ( \15792 , \14654 );
buf \U$15547 ( \15793 , \13268 );
not \U$15548 ( \15794 , \15793 );
or \U$15549 ( \15795 , \15792 , \15794 );
nand \U$15550 ( \15796 , \11348 , \14940 );
nand \U$15551 ( \15797 , \15795 , \15796 );
not \U$15552 ( \15798 , \15797 );
or \U$15553 ( \15799 , \15791 , \15798 );
or \U$15554 ( \15800 , \15797 , \15790 );
not \U$15555 ( \15801 , \14458 );
not \U$15556 ( \15802 , \10987 );
or \U$15557 ( \15803 , \15801 , \15802 );
nand \U$15558 ( \15804 , \9726 , \14235 );
nand \U$15559 ( \15805 , \15803 , \15804 );
nand \U$15560 ( \15806 , \15800 , \15805 );
nand \U$15561 ( \15807 , \15799 , \15806 );
not \U$15562 ( \15808 , \15807 );
or \U$15563 ( \15809 , \15785 , \15808 );
not \U$15564 ( \15810 , \15807 );
not \U$15565 ( \15811 , \15784 );
nand \U$15566 ( \15812 , \15810 , \15811 );
not \U$15567 ( \15813 , \15723 );
not \U$15568 ( \15814 , \15734 );
or \U$15569 ( \15815 , \15813 , \15814 );
nand \U$15570 ( \15816 , \15728 , \15733 );
nand \U$15571 ( \15817 , \15815 , \15816 );
nand \U$15572 ( \15818 , \15812 , \15817 );
nand \U$15573 ( \15819 , \15809 , \15818 );
not \U$15574 ( \15820 , \15819 );
not \U$15575 ( \15821 , \15593 );
not \U$15576 ( \15822 , \15587 );
or \U$15577 ( \15823 , \15821 , \15822 );
or \U$15578 ( \15824 , \15587 , \15593 );
nand \U$15579 ( \15825 , \15824 , \15583 );
nand \U$15580 ( \15826 , \15823 , \15825 );
not \U$15581 ( \15827 , \14282 );
not \U$15582 ( \15828 , \14275 );
or \U$15583 ( \15829 , \15827 , \15828 );
nand \U$15584 ( \15830 , \14263 , \14270 );
nand \U$15585 ( \15831 , \15829 , \15830 );
not \U$15586 ( \15832 , \15831 );
xor \U$15587 ( \15833 , \15826 , \15832 );
not \U$15588 ( \15834 , \14797 );
not \U$15589 ( \15835 , \14815 );
or \U$15590 ( \15836 , \15834 , \15835 );
nand \U$15591 ( \15837 , \14803 , \14810 );
nand \U$15592 ( \15838 , \15836 , \15837 );
xor \U$15593 ( \15839 , \15833 , \15838 );
not \U$15594 ( \15840 , \15839 );
or \U$15595 ( \15841 , \15820 , \15840 );
or \U$15596 ( \15842 , \15839 , \15819 );
nand \U$15597 ( \15843 , \15841 , \15842 );
xor \U$15598 ( \15844 , \15267 , \15312 );
and \U$15599 ( \15845 , \15843 , \15844 );
not \U$15600 ( \15846 , \15843 );
not \U$15601 ( \15847 , \15844 );
and \U$15602 ( \15848 , \15846 , \15847 );
nor \U$15603 ( \15849 , \15845 , \15848 );
or \U$15604 ( \15850 , \14832 , \14839 );
nand \U$15605 ( \15851 , \15850 , \14834 );
not \U$15606 ( \15852 , \15851 );
not \U$15607 ( \15853 , \15616 );
not \U$15608 ( \15854 , \15611 );
or \U$15609 ( \15855 , \15853 , \15854 );
nand \U$15610 ( \15856 , \15610 , \15605 );
nand \U$15611 ( \15857 , \15855 , \15856 );
not \U$15612 ( \15858 , \15857 );
not \U$15613 ( \15859 , \15858 );
or \U$15614 ( \15860 , \15852 , \15859 );
or \U$15615 ( \15861 , \15858 , \15851 );
nand \U$15616 ( \15862 , \15860 , \15861 );
not \U$15617 ( \15863 , \14254 );
not \U$15618 ( \15864 , \14247 );
or \U$15619 ( \15865 , \15863 , \15864 );
nand \U$15620 ( \15866 , \14240 , \14246 );
nand \U$15621 ( \15867 , \15865 , \15866 );
and \U$15622 ( \15868 , \15862 , \15867 );
not \U$15623 ( \15869 , \15862 );
not \U$15624 ( \15870 , \15867 );
and \U$15625 ( \15871 , \15869 , \15870 );
nor \U$15626 ( \15872 , \15868 , \15871 );
xor \U$15627 ( \15873 , \15274 , \15288 );
not \U$15628 ( \15874 , \15873 );
not \U$15629 ( \15875 , \14492 );
not \U$15630 ( \15876 , \1780 );
or \U$15631 ( \15877 , \15875 , \15876 );
nand \U$15632 ( \15878 , \5055 , \14241 );
nand \U$15633 ( \15879 , \15877 , \15878 );
not \U$15634 ( \15880 , \15879 );
not \U$15635 ( \15881 , \14566 );
not \U$15636 ( \15882 , \8898 );
or \U$15637 ( \15883 , \15881 , \15882 );
nand \U$15638 ( \15884 , \10752 , \15276 );
nand \U$15639 ( \15885 , \15883 , \15884 );
not \U$15640 ( \15886 , \15885 );
or \U$15641 ( \15887 , \15880 , \15886 );
not \U$15642 ( \15888 , \15885 );
not \U$15643 ( \15889 , \15888 );
not \U$15644 ( \15890 , \15879 );
not \U$15645 ( \15891 , \15890 );
or \U$15646 ( \15892 , \15889 , \15891 );
not \U$15647 ( \15893 , \14484 );
not \U$15648 ( \15894 , \10542 );
or \U$15649 ( \15895 , \15893 , \15894 );
nand \U$15650 ( \15896 , \2369 , \15600 );
nand \U$15651 ( \15897 , \15895 , \15896 );
nand \U$15652 ( \15898 , \15892 , \15897 );
nand \U$15653 ( \15899 , \15887 , \15898 );
xor \U$15654 ( \15900 , \15299 , \15306 );
xnor \U$15655 ( \15901 , \15900 , \15297 );
xor \U$15656 ( \15902 , \15899 , \15901 );
not \U$15657 ( \15903 , \15902 );
or \U$15658 ( \15904 , \15874 , \15903 );
nand \U$15659 ( \15905 , \15901 , \15899 );
nand \U$15660 ( \15906 , \15904 , \15905 );
xor \U$15661 ( \15907 , \15872 , \15906 );
not \U$15662 ( \15908 , \15577 );
not \U$15663 ( \15909 , \15908 );
not \U$15664 ( \15910 , \15622 );
or \U$15665 ( \15911 , \15909 , \15910 );
nand \U$15666 ( \15912 , \15599 , \15617 );
nand \U$15667 ( \15913 , \15911 , \15912 );
xor \U$15668 ( \15914 , \15907 , \15913 );
xor \U$15669 ( \15915 , \15849 , \15914 );
xnor \U$15670 ( \15916 , \14870 , \14816 );
not \U$15671 ( \15917 , \15916 );
not \U$15672 ( \15918 , \15917 );
xnor \U$15673 ( \15919 , \15902 , \15873 );
not \U$15674 ( \15920 , \15919 );
not \U$15675 ( \15921 , \14255 );
not \U$15676 ( \15922 , \14320 );
or \U$15677 ( \15923 , \15921 , \15922 );
or \U$15678 ( \15924 , \14320 , \14255 );
nand \U$15679 ( \15925 , \15923 , \15924 );
not \U$15680 ( \15926 , \15925 );
or \U$15681 ( \15927 , \15920 , \15926 );
or \U$15682 ( \15928 , \15919 , \15925 );
nand \U$15683 ( \15929 , \15927 , \15928 );
not \U$15684 ( \15930 , \15929 );
or \U$15685 ( \15931 , \15918 , \15930 );
not \U$15686 ( \15932 , \15919 );
nand \U$15687 ( \15933 , \15932 , \15925 );
nand \U$15688 ( \15934 , \15931 , \15933 );
xor \U$15689 ( \15935 , \15915 , \15934 );
not \U$15690 ( \15936 , \15570 );
and \U$15691 ( \15937 , \15474 , \15936 );
not \U$15692 ( \15938 , \15474 );
and \U$15693 ( \15939 , \15938 , \15570 );
nor \U$15694 ( \15940 , \15937 , \15939 );
not \U$15695 ( \15941 , \15940 );
not \U$15696 ( \15942 , \15941 );
buf \U$15697 ( \15943 , \15741 );
xor \U$15698 ( \15944 , \15943 , \15717 );
xor \U$15699 ( \15945 , RIbe280c0_13, RIbe2a0a0_81);
not \U$15700 ( \15946 , \15945 );
not \U$15701 ( \15947 , \8551 );
or \U$15702 ( \15948 , \15946 , \15947 );
nand \U$15703 ( \15949 , \1263 , \15697 );
nand \U$15704 ( \15950 , \15948 , \15949 );
xor \U$15705 ( \15951 , RIbe2aaf0_103, RIbe2b630_127);
buf \U$15706 ( \15952 , \15951 );
buf \U$15707 ( \15953 , \15952 );
not \U$15708 ( \15954 , \15953 );
not \U$15709 ( \15955 , \15954 );
not \U$15710 ( \15956 , RIbe2b630_127);
not \U$15711 ( \15957 , \15956 );
not \U$15712 ( \15958 , RIbe2b018_114);
not \U$15713 ( \15959 , \15958 );
or \U$15714 ( \15960 , \15957 , \15959 );
and \U$15715 ( \15961 , RIbe2aaf0_103, RIbe2b018_114);
not \U$15716 ( \15962 , RIbe2aaf0_103);
and \U$15717 ( \15963 , \15962 , RIbe2b630_127);
nor \U$15718 ( \15964 , \15961 , \15963 );
nand \U$15719 ( \15965 , \15960 , \15964 );
buf \U$15720 ( \15966 , \15965 );
not \U$15721 ( \15967 , \15966 );
not \U$15722 ( \15968 , \15967 );
not \U$15723 ( \15969 , \15968 );
or \U$15724 ( \15970 , \15955 , \15969 );
nand \U$15725 ( \15971 , \15970 , RIbe2b018_114);
or \U$15726 ( \15972 , \15950 , \15971 );
xor \U$15727 ( \15973 , RIbe28a98_34, RIbe2a910_99);
not \U$15728 ( \15974 , \15973 );
not \U$15729 ( \15975 , \10987 );
or \U$15730 ( \15976 , \15974 , \15975 );
nand \U$15731 ( \15977 , \9726 , \15393 );
nand \U$15732 ( \15978 , \15976 , \15977 );
nand \U$15733 ( \15979 , \15972 , \15978 );
nand \U$15734 ( \15980 , \15971 , \15950 );
nand \U$15735 ( \15981 , \15979 , \15980 );
not \U$15736 ( \15982 , \10568 );
xor \U$15737 ( \15983 , RIbe2ad48_108, RIbe290b0_47);
not \U$15738 ( \15984 , \15983 );
or \U$15739 ( \15985 , \15982 , \15984 );
not \U$15740 ( \15986 , \15367 );
or \U$15741 ( \15987 , \3980 , \15986 );
nand \U$15742 ( \15988 , \15985 , \15987 );
xor \U$15743 ( \15989 , RIbe2a550_91, RIbe29308_52);
not \U$15744 ( \15990 , \15989 );
not \U$15745 ( \15991 , \10432 );
not \U$15746 ( \15992 , \15991 );
not \U$15747 ( \15993 , \15992 );
or \U$15748 ( \15994 , \15990 , \15993 );
not \U$15749 ( \15995 , \10439 );
nand \U$15750 ( \15996 , \15995 , \15540 );
nand \U$15751 ( \15997 , \15994 , \15996 );
nor \U$15752 ( \15998 , \15988 , \15997 );
xor \U$15753 ( \15999 , RIbe28f48_44, RIbe29a10_67);
not \U$15754 ( \16000 , \15999 );
not \U$15755 ( \16001 , \3256 );
or \U$15756 ( \16002 , \16000 , \16001 );
nand \U$15757 ( \16003 , \3249 , \15518 );
nand \U$15758 ( \16004 , \16002 , \16003 );
not \U$15759 ( \16005 , \16004 );
or \U$15760 ( \16006 , \15998 , \16005 );
nand \U$15761 ( \16007 , \15997 , \15988 );
nand \U$15762 ( \16008 , \16006 , \16007 );
xor \U$15763 ( \16009 , \15981 , \16008 );
not \U$15764 ( \16010 , \8270 );
not \U$15765 ( \16011 , \15359 );
or \U$15766 ( \16012 , \16010 , \16011 );
xnor \U$15767 ( \16013 , RIbe285e8_24, RIbe298a8_64);
or \U$15768 ( \16014 , \2762 , \16013 );
nand \U$15769 ( \16015 , \16012 , \16014 );
xor \U$15770 ( \16016 , RIbe29c68_72, RIbe29128_48);
not \U$15771 ( \16017 , \16016 );
not \U$15772 ( \16018 , \8595 );
or \U$15773 ( \16019 , \16017 , \16018 );
nand \U$15774 ( \16020 , \4580 , \15657 );
nand \U$15775 ( \16021 , \16019 , \16020 );
xor \U$15776 ( \16022 , \16015 , \16021 );
not \U$15777 ( \16023 , \15703 );
not \U$15778 ( \16024 , \2691 );
or \U$15779 ( \16025 , \16023 , \16024 );
xnor \U$15780 ( \16026 , RIbe28b88_36, RIbe29ec0_77);
or \U$15781 ( \16027 , \4541 , \16026 );
nand \U$15782 ( \16028 , \16025 , \16027 );
and \U$15783 ( \16029 , \16022 , \16028 );
and \U$15784 ( \16030 , \16015 , \16021 );
or \U$15785 ( \16031 , \16029 , \16030 );
and \U$15786 ( \16032 , \16009 , \16031 );
and \U$15787 ( \16033 , \15981 , \16008 );
or \U$15788 ( \16034 , \16032 , \16033 );
not \U$15789 ( \16035 , \16034 );
xnor \U$15790 ( \16036 , \14468 , \14452 );
not \U$15791 ( \16037 , \16036 );
xor \U$15792 ( \16038 , \15350 , \15357 );
xor \U$15793 ( \16039 , \16038 , \15387 );
not \U$15794 ( \16040 , \16039 );
or \U$15795 ( \16041 , \16037 , \16040 );
or \U$15796 ( \16042 , \16039 , \16036 );
nand \U$15797 ( \16043 , \16041 , \16042 );
not \U$15798 ( \16044 , \16043 );
or \U$15799 ( \16045 , \16035 , \16044 );
not \U$15800 ( \16046 , \16036 );
nand \U$15801 ( \16047 , \16046 , \16039 );
nand \U$15802 ( \16048 , \16045 , \16047 );
xor \U$15803 ( \16049 , \15944 , \16048 );
not \U$15804 ( \16050 , \16049 );
or \U$15805 ( \16051 , \15942 , \16050 );
nand \U$15806 ( \16052 , \16048 , \15944 );
nand \U$15807 ( \16053 , \16051 , \16052 );
not \U$15808 ( \16054 , \16053 );
not \U$15809 ( \16055 , \15916 );
not \U$15810 ( \16056 , \15929 );
or \U$15811 ( \16057 , \16055 , \16056 );
or \U$15812 ( \16058 , \15929 , \15916 );
nand \U$15813 ( \16059 , \16057 , \16058 );
not \U$15814 ( \16060 , \16059 );
not \U$15815 ( \16061 , \15573 );
not \U$15816 ( \16062 , \15748 );
or \U$15817 ( \16063 , \16061 , \16062 );
or \U$15818 ( \16064 , \15748 , \15573 );
nand \U$15819 ( \16065 , \16063 , \16064 );
not \U$15820 ( \16066 , \16065 );
not \U$15821 ( \16067 , \16066 );
or \U$15822 ( \16068 , \16060 , \16067 );
not \U$15823 ( \16069 , \16059 );
nand \U$15824 ( \16070 , \16069 , \16065 );
nand \U$15825 ( \16071 , \16068 , \16070 );
not \U$15826 ( \16072 , \16071 );
or \U$15827 ( \16073 , \16054 , \16072 );
nand \U$15828 ( \16074 , \16065 , \16059 );
nand \U$15829 ( \16075 , \16073 , \16074 );
and \U$15830 ( \16076 , \15935 , \16075 );
not \U$15831 ( \16077 , \15935 );
not \U$15832 ( \16078 , \16075 );
and \U$15833 ( \16079 , \16077 , \16078 );
nor \U$15834 ( \16080 , \16076 , \16079 );
not \U$15835 ( \16081 , \16080 );
or \U$15836 ( \16082 , \15762 , \16081 );
nand \U$15837 ( \16083 , \16075 , \15935 );
nand \U$15838 ( \16084 , \16082 , \16083 );
not \U$15839 ( \16085 , \16084 );
xor \U$15840 ( \16086 , \15774 , \15768 );
not \U$15841 ( \16087 , \15782 );
and \U$15842 ( \16088 , \16086 , \16087 );
not \U$15843 ( \16089 , \16086 );
and \U$15844 ( \16090 , \16089 , \15782 );
nor \U$15845 ( \16091 , \16088 , \16090 );
not \U$15846 ( \16092 , \15885 );
not \U$15847 ( \16093 , \15890 );
or \U$15848 ( \16094 , \16092 , \16093 );
nand \U$15849 ( \16095 , \15879 , \15888 );
nand \U$15850 ( \16096 , \16094 , \16095 );
and \U$15851 ( \16097 , \16096 , \15897 );
not \U$15852 ( \16098 , \16096 );
not \U$15853 ( \16099 , \15897 );
and \U$15854 ( \16100 , \16098 , \16099 );
nor \U$15855 ( \16101 , \16097 , \16100 );
xnor \U$15856 ( \16102 , \16091 , \16101 );
xor \U$15857 ( \16103 , \15797 , \15790 );
xor \U$15858 ( \16104 , \16103 , \15805 );
xor \U$15859 ( \16105 , \16102 , \16104 );
not \U$15860 ( \16106 , \16105 );
not \U$15861 ( \16107 , \15042 );
not \U$15862 ( \16108 , \15029 );
and \U$15863 ( \16109 , \16107 , \16108 );
and \U$15864 ( \16110 , \15042 , \15029 );
nor \U$15865 ( \16111 , \16109 , \16110 );
not \U$15866 ( \16112 , \16111 );
not \U$15867 ( \16113 , \15002 );
and \U$15868 ( \16114 , \15015 , \16113 );
not \U$15869 ( \16115 , \15015 );
and \U$15870 ( \16116 , \16115 , \15002 );
nor \U$15871 ( \16117 , \16114 , \16116 );
not \U$15872 ( \16118 , \16117 );
xor \U$15873 ( \16119 , \16112 , \16118 );
and \U$15874 ( \16120 , \3344 , \15651 );
nor \U$15875 ( \16121 , \2670 , \15049 );
nor \U$15876 ( \16122 , \16120 , \16121 );
not \U$15877 ( \16123 , \16122 );
not \U$15878 ( \16124 , \16123 );
not \U$15879 ( \16125 , \15429 );
not \U$15880 ( \16126 , \11321 );
or \U$15881 ( \16127 , \16125 , \16126 );
nand \U$15882 ( \16128 , \346 , \15076 );
nand \U$15883 ( \16129 , \16127 , \16128 );
nand \U$15884 ( \16130 , RIbe27b98_2, RIbe2a7a8_96);
and \U$15885 ( \16131 , \16129 , \16130 );
not \U$15886 ( \16132 , \16129 );
not \U$15887 ( \16133 , \16130 );
and \U$15888 ( \16134 , \16132 , \16133 );
or \U$15889 ( \16135 , \16131 , \16134 );
not \U$15890 ( \16136 , \16135 );
or \U$15891 ( \16137 , \16124 , \16136 );
nand \U$15892 ( \16138 , \16129 , \16133 );
nand \U$15893 ( \16139 , \16137 , \16138 );
xnor \U$15894 ( \16140 , \16119 , \16139 );
not \U$15895 ( \16141 , \16140 );
xor \U$15896 ( \16142 , \14968 , \14987 );
xor \U$15897 ( \16143 , \15063 , \15069 );
xnor \U$15898 ( \16144 , \16143 , \15054 );
xor \U$15899 ( \16145 , \16142 , \16144 );
xor \U$15900 ( \16146 , \15082 , \15094 );
buf \U$15901 ( \16147 , \16146 );
and \U$15902 ( \16148 , \16145 , \16147 );
not \U$15903 ( \16149 , \16145 );
not \U$15904 ( \16150 , \16147 );
and \U$15905 ( \16151 , \16149 , \16150 );
nor \U$15906 ( \16152 , \16148 , \16151 );
not \U$15907 ( \16153 , \16152 );
or \U$15908 ( \16154 , \16141 , \16153 );
or \U$15909 ( \16155 , \16152 , \16140 );
nand \U$15910 ( \16156 , \16154 , \16155 );
not \U$15911 ( \16157 , \16156 );
or \U$15912 ( \16158 , \16106 , \16157 );
not \U$15913 ( \16159 , \16140 );
nand \U$15914 ( \16160 , \16159 , \16152 );
nand \U$15915 ( \16161 , \16158 , \16160 );
not \U$15916 ( \16162 , \16161 );
not \U$15917 ( \16163 , \16146 );
not \U$15918 ( \16164 , \16144 );
or \U$15919 ( \16165 , \16163 , \16164 );
or \U$15920 ( \16166 , \16144 , \16146 );
nand \U$15921 ( \16167 , \16166 , \16142 );
nand \U$15922 ( \16168 , \16165 , \16167 );
not \U$15923 ( \16169 , \16112 );
not \U$15924 ( \16170 , \16118 );
or \U$15925 ( \16171 , \16169 , \16170 );
not \U$15926 ( \16172 , \16111 );
not \U$15927 ( \16173 , \16117 );
or \U$15928 ( \16174 , \16172 , \16173 );
nand \U$15929 ( \16175 , \16174 , \16139 );
nand \U$15930 ( \16176 , \16171 , \16175 );
xor \U$15931 ( \16177 , \16168 , \16176 );
not \U$15932 ( \16178 , \16104 );
not \U$15933 ( \16179 , \16102 );
or \U$15934 ( \16180 , \16178 , \16179 );
not \U$15935 ( \16181 , \16091 );
nand \U$15936 ( \16182 , \16181 , \16101 );
nand \U$15937 ( \16183 , \16180 , \16182 );
xor \U$15938 ( \16184 , \16177 , \16183 );
xor \U$15939 ( \16185 , \15807 , \15811 );
xnor \U$15940 ( \16186 , \16185 , \15817 );
buf \U$15941 ( \16187 , \15020 );
not \U$15942 ( \16188 , \14991 );
and \U$15943 ( \16189 , \16187 , \16188 );
not \U$15944 ( \16190 , \16187 );
and \U$15945 ( \16191 , \16190 , \14991 );
nor \U$15946 ( \16192 , \16189 , \16191 );
not \U$15947 ( \16193 , \16192 );
xor \U$15948 ( \16194 , \16186 , \16193 );
xor \U$15949 ( \16195 , \15098 , \15046 );
xor \U$15950 ( \16196 , \16195 , \15075 );
buf \U$15951 ( \16197 , \16196 );
xnor \U$15952 ( \16198 , \16194 , \16197 );
not \U$15953 ( \16199 , \16198 );
and \U$15954 ( \16200 , \16184 , \16199 );
not \U$15955 ( \16201 , \16184 );
and \U$15956 ( \16202 , \16201 , \16198 );
nor \U$15957 ( \16203 , \16200 , \16202 );
not \U$15958 ( \16204 , \16203 );
or \U$15959 ( \16205 , \16162 , \16204 );
nand \U$15960 ( \16206 , \16199 , \16184 );
nand \U$15961 ( \16207 , \16205 , \16206 );
not \U$15962 ( \16208 , \16207 );
not \U$15963 ( \16209 , \16186 );
not \U$15964 ( \16210 , \16196 );
not \U$15965 ( \16211 , \16192 );
or \U$15966 ( \16212 , \16210 , \16211 );
or \U$15967 ( \16213 , \16196 , \16192 );
nand \U$15968 ( \16214 , \16212 , \16213 );
not \U$15969 ( \16215 , \16214 );
or \U$15970 ( \16216 , \16209 , \16215 );
nand \U$15971 ( \16217 , \16197 , \16193 );
nand \U$15972 ( \16218 , \16216 , \16217 );
xor \U$15973 ( \16219 , \14961 , \15024 );
xor \U$15974 ( \16220 , \16219 , \15103 );
not \U$15975 ( \16221 , \16183 );
not \U$15976 ( \16222 , \16177 );
or \U$15977 ( \16223 , \16221 , \16222 );
nand \U$15978 ( \16224 , \16168 , \16176 );
nand \U$15979 ( \16225 , \16223 , \16224 );
and \U$15980 ( \16226 , \16220 , \16225 );
not \U$15981 ( \16227 , \16220 );
not \U$15982 ( \16228 , \16225 );
and \U$15983 ( \16229 , \16227 , \16228 );
nor \U$15984 ( \16230 , \16226 , \16229 );
xor \U$15985 ( \16231 , \16218 , \16230 );
xor \U$15986 ( \16232 , \14509 , \14696 );
not \U$15987 ( \16233 , \16232 );
xor \U$15988 ( \16234 , \14445 , \14505 );
not \U$15989 ( \16235 , \16234 );
not \U$15990 ( \16236 , \14541 );
not \U$15991 ( \16237 , \16236 );
not \U$15992 ( \16238 , \14595 );
and \U$15993 ( \16239 , \16237 , \16238 );
and \U$15994 ( \16240 , \14595 , \16236 );
nor \U$15995 ( \16241 , \16239 , \16240 );
not \U$15996 ( \16242 , \16241 );
xor \U$15997 ( \16243 , \14659 , \14689 );
xnor \U$15998 ( \16244 , \16243 , \14627 );
not \U$15999 ( \16245 , \16244 );
or \U$16000 ( \16246 , \16242 , \16245 );
or \U$16001 ( \16247 , \16244 , \16241 );
nand \U$16002 ( \16248 , \16246 , \16247 );
not \U$16003 ( \16249 , \16248 );
or \U$16004 ( \16250 , \16235 , \16249 );
not \U$16005 ( \16251 , \16241 );
nand \U$16006 ( \16252 , \16251 , \16244 );
nand \U$16007 ( \16253 , \16250 , \16252 );
buf \U$16008 ( \16254 , \14623 );
and \U$16009 ( \16255 , \16254 , \14606 );
not \U$16010 ( \16256 , \16254 );
not \U$16011 ( \16257 , \14606 );
and \U$16012 ( \16258 , \16256 , \16257 );
nor \U$16013 ( \16259 , \16255 , \16258 );
not \U$16014 ( \16260 , \16259 );
not \U$16015 ( \16261 , \14499 );
xor \U$16016 ( \16262 , \14478 , \16261 );
and \U$16017 ( \16263 , \14682 , \14666 );
not \U$16018 ( \16264 , \14682 );
not \U$16019 ( \16265 , \14666 );
and \U$16020 ( \16266 , \16264 , \16265 );
nor \U$16021 ( \16267 , \16263 , \16266 );
xnor \U$16022 ( \16268 , \16262 , \16267 );
not \U$16023 ( \16269 , \16268 );
or \U$16024 ( \16270 , \16260 , \16269 );
and \U$16025 ( \16271 , \14478 , \16261 );
not \U$16026 ( \16272 , \14478 );
and \U$16027 ( \16273 , \16272 , \14499 );
or \U$16028 ( \16274 , \16271 , \16273 );
nand \U$16029 ( \16275 , \16274 , \16267 );
nand \U$16030 ( \16276 , \16270 , \16275 );
not \U$16031 ( \16277 , \16122 );
not \U$16032 ( \16278 , \16135 );
or \U$16033 ( \16279 , \16277 , \16278 );
or \U$16034 ( \16280 , \16135 , \16122 );
nand \U$16035 ( \16281 , \16279 , \16280 );
not \U$16036 ( \16282 , \16281 );
xor \U$16037 ( \16283 , \14526 , \14535 );
xor \U$16038 ( \16284 , \16283 , \14518 );
not \U$16039 ( \16285 , \16284 );
or \U$16040 ( \16286 , \16282 , \16285 );
or \U$16041 ( \16287 , \16284 , \16281 );
nand \U$16042 ( \16288 , \16286 , \16287 );
not \U$16043 ( \16289 , \16288 );
xor \U$16044 ( \16290 , \14576 , \14591 );
xor \U$16045 ( \16291 , \16290 , \14584 );
not \U$16046 ( \16292 , \16291 );
or \U$16047 ( \16293 , \16289 , \16292 );
not \U$16048 ( \16294 , \16284 );
nand \U$16049 ( \16295 , \16294 , \16281 );
nand \U$16050 ( \16296 , \16293 , \16295 );
or \U$16051 ( \16297 , \16276 , \16296 );
xor \U$16052 ( \16298 , \14568 , \14558 );
xor \U$16053 ( \16299 , \14549 , \16298 );
not \U$16054 ( \16300 , \16299 );
xor \U$16055 ( \16301 , \14643 , \14635 );
xnor \U$16056 ( \16302 , \16301 , \14656 );
not \U$16057 ( \16303 , \16302 );
xnor \U$16058 ( \16304 , \14409 , \14440 );
not \U$16059 ( \16305 , \16304 );
or \U$16060 ( \16306 , \16303 , \16305 );
or \U$16061 ( \16307 , \16304 , \16302 );
nand \U$16062 ( \16308 , \16306 , \16307 );
not \U$16063 ( \16309 , \16308 );
or \U$16064 ( \16310 , \16300 , \16309 );
not \U$16065 ( \16311 , \16302 );
nand \U$16066 ( \16312 , \16311 , \16304 );
nand \U$16067 ( \16313 , \16310 , \16312 );
nand \U$16068 ( \16314 , \16297 , \16313 );
nand \U$16069 ( \16315 , \16296 , \16276 );
nand \U$16070 ( \16316 , \16314 , \16315 );
and \U$16071 ( \16317 , \16253 , \16316 );
not \U$16072 ( \16318 , \16253 );
not \U$16073 ( \16319 , \16316 );
and \U$16074 ( \16320 , \16318 , \16319 );
nor \U$16075 ( \16321 , \16317 , \16320 );
not \U$16076 ( \16322 , \16321 );
or \U$16077 ( \16323 , \16233 , \16322 );
nand \U$16078 ( \16324 , \16316 , \16253 );
nand \U$16079 ( \16325 , \16323 , \16324 );
and \U$16080 ( \16326 , \16231 , \16325 );
not \U$16081 ( \16327 , \16231 );
not \U$16082 ( \16328 , \16325 );
and \U$16083 ( \16329 , \16327 , \16328 );
nor \U$16084 ( \16330 , \16326 , \16329 );
not \U$16085 ( \16331 , \16330 );
or \U$16086 ( \16332 , \16208 , \16331 );
nand \U$16087 ( \16333 , \16325 , \16231 );
nand \U$16088 ( \16334 , \16332 , \16333 );
not \U$16089 ( \16335 , \16334 );
nor \U$16090 ( \16336 , \15857 , \15867 );
not \U$16091 ( \16337 , \15851 );
or \U$16092 ( \16338 , \16336 , \16337 );
nand \U$16093 ( \16339 , \15857 , \15867 );
nand \U$16094 ( \16340 , \16338 , \16339 );
not \U$16095 ( \16341 , \16340 );
not \U$16096 ( \16342 , \15826 );
nand \U$16097 ( \16343 , \16342 , \15832 );
not \U$16098 ( \16344 , \16343 );
not \U$16099 ( \16345 , \15838 );
or \U$16100 ( \16346 , \16344 , \16345 );
nand \U$16101 ( \16347 , \15831 , \15826 );
nand \U$16102 ( \16348 , \16346 , \16347 );
not \U$16103 ( \16349 , \16348 );
not \U$16104 ( \16350 , \16349 );
or \U$16105 ( \16351 , \16341 , \16350 );
not \U$16106 ( \16352 , \16340 );
nand \U$16107 ( \16353 , \16352 , \16348 );
nand \U$16108 ( \16354 , \16351 , \16353 );
not \U$16109 ( \16355 , \13579 );
and \U$16110 ( \16356 , \13638 , \16355 );
not \U$16111 ( \16357 , \13638 );
and \U$16112 ( \16358 , \16357 , \13579 );
nor \U$16113 ( \16359 , \16356 , \16358 );
not \U$16114 ( \16360 , \16359 );
and \U$16115 ( \16361 , \16354 , \16360 );
not \U$16116 ( \16362 , \16354 );
and \U$16117 ( \16363 , \16362 , \16359 );
nor \U$16118 ( \16364 , \16361 , \16363 );
xor \U$16119 ( \16365 , \15872 , \15906 );
and \U$16120 ( \16366 , \16365 , \15913 );
and \U$16121 ( \16367 , \15872 , \15906 );
or \U$16122 ( \16368 , \16366 , \16367 );
xor \U$16123 ( \16369 , \16364 , \16368 );
not \U$16124 ( \16370 , \15844 );
not \U$16125 ( \16371 , \15843 );
or \U$16126 ( \16372 , \16370 , \16371 );
not \U$16127 ( \16373 , \15839 );
nand \U$16128 ( \16374 , \16373 , \15819 );
nand \U$16129 ( \16375 , \16372 , \16374 );
xor \U$16130 ( \16376 , \16369 , \16375 );
not \U$16131 ( \16377 , \16376 );
not \U$16132 ( \16378 , \16218 );
not \U$16133 ( \16379 , \16230 );
or \U$16134 ( \16380 , \16378 , \16379 );
not \U$16135 ( \16381 , \16228 );
nand \U$16136 ( \16382 , \16381 , \16220 );
nand \U$16137 ( \16383 , \16380 , \16382 );
not \U$16138 ( \16384 , \16383 );
not \U$16139 ( \16385 , \16384 );
or \U$16140 ( \16386 , \16377 , \16385 );
or \U$16141 ( \16387 , \16384 , \16376 );
nand \U$16142 ( \16388 , \16386 , \16387 );
not \U$16143 ( \16389 , \16388 );
nand \U$16144 ( \16390 , \15934 , \15915 );
nand \U$16145 ( \16391 , \15914 , \15849 );
and \U$16146 ( \16392 , \16390 , \16391 );
not \U$16147 ( \16393 , \16392 );
and \U$16148 ( \16394 , \16389 , \16393 );
and \U$16149 ( \16395 , \16392 , \16388 );
nor \U$16150 ( \16396 , \16394 , \16395 );
not \U$16151 ( \16397 , \16396 );
or \U$16152 ( \16398 , \16335 , \16397 );
or \U$16153 ( \16399 , \16396 , \16334 );
nand \U$16154 ( \16400 , \16398 , \16399 );
not \U$16155 ( \16401 , \16400 );
or \U$16156 ( \16402 , \16085 , \16401 );
not \U$16157 ( \16403 , \16396 );
nand \U$16158 ( \16404 , \16403 , \16334 );
nand \U$16159 ( \16405 , \16402 , \16404 );
nand \U$16160 ( \16406 , \15342 , \16405 );
not \U$16161 ( \16407 , \16406 );
xor \U$16162 ( \16408 , \16364 , \16368 );
and \U$16163 ( \16409 , \16408 , \16375 );
and \U$16164 ( \16410 , \16364 , \16368 );
or \U$16165 ( \16411 , \16409 , \16410 );
xnor \U$16166 ( \16412 , \13642 , \13553 );
not \U$16167 ( \16413 , \16412 );
not \U$16168 ( \16414 , \16360 );
not \U$16169 ( \16415 , \16354 );
or \U$16170 ( \16416 , \16414 , \16415 );
nand \U$16171 ( \16417 , \16348 , \16340 );
nand \U$16172 ( \16418 , \16416 , \16417 );
not \U$16173 ( \16419 , \16418 );
or \U$16174 ( \16420 , \16413 , \16419 );
or \U$16175 ( \16421 , \16418 , \16412 );
nand \U$16176 ( \16422 , \16420 , \16421 );
not \U$16177 ( \16423 , \16422 );
not \U$16178 ( \16424 , \16423 );
not \U$16179 ( \16425 , \15167 );
not \U$16180 ( \16426 , \15178 );
or \U$16181 ( \16427 , \16425 , \16426 );
nand \U$16182 ( \16428 , \15172 , \15177 );
nand \U$16183 ( \16429 , \16427 , \16428 );
xor \U$16184 ( \16430 , \15145 , \15149 );
and \U$16185 ( \16431 , \16430 , \15156 );
and \U$16186 ( \16432 , \15145 , \15149 );
or \U$16187 ( \16433 , \16431 , \16432 );
not \U$16188 ( \16434 , \16433 );
not \U$16189 ( \16435 , \13476 );
not \U$16190 ( \16436 , \13413 );
not \U$16191 ( \16437 , \16436 );
and \U$16192 ( \16438 , \16435 , \16437 );
and \U$16193 ( \16439 , \13476 , \16436 );
nor \U$16194 ( \16440 , \16438 , \16439 );
not \U$16195 ( \16441 , \16440 );
or \U$16196 ( \16442 , \16434 , \16441 );
or \U$16197 ( \16443 , \16440 , \16433 );
nand \U$16198 ( \16444 , \16442 , \16443 );
xor \U$16199 ( \16445 , \16429 , \16444 );
not \U$16200 ( \16446 , \16445 );
or \U$16201 ( \16447 , \16424 , \16446 );
not \U$16202 ( \16448 , \16445 );
nand \U$16203 ( \16449 , \16448 , \16422 );
nand \U$16204 ( \16450 , \16447 , \16449 );
xor \U$16205 ( \16451 , \16411 , \16450 );
buf \U$16206 ( \16452 , \16451 );
and \U$16207 ( \16453 , \15254 , \15260 );
not \U$16208 ( \16454 , \15254 );
and \U$16209 ( \16455 , \16454 , \15259 );
nor \U$16210 ( \16456 , \16453 , \16455 );
xor \U$16211 ( \16457 , \16456 , \15316 );
xor \U$16212 ( \16458 , \15157 , \15162 );
xor \U$16213 ( \16459 , \16458 , \15179 );
xor \U$16214 ( \16460 , \16457 , \16459 );
xor \U$16215 ( \16461 , \15212 , \15200 );
and \U$16216 ( \16462 , \16460 , \16461 );
and \U$16217 ( \16463 , \16457 , \16459 );
or \U$16218 ( \16464 , \16462 , \16463 );
not \U$16219 ( \16465 , \16464 );
and \U$16220 ( \16466 , \16452 , \16465 );
not \U$16221 ( \16467 , \16452 );
and \U$16222 ( \16468 , \16467 , \16464 );
nor \U$16223 ( \16469 , \16466 , \16468 );
not \U$16224 ( \16470 , \16469 );
not \U$16225 ( \16471 , \16470 );
not \U$16226 ( \16472 , \16392 );
not \U$16227 ( \16473 , \16472 );
not \U$16228 ( \16474 , \16388 );
or \U$16229 ( \16475 , \16473 , \16474 );
not \U$16230 ( \16476 , \16384 );
nand \U$16231 ( \16477 , \16476 , \16376 );
nand \U$16232 ( \16478 , \16475 , \16477 );
not \U$16233 ( \16479 , \16478 );
not \U$16234 ( \16480 , \16479 );
or \U$16235 ( \16481 , \16471 , \16480 );
nand \U$16236 ( \16482 , \16478 , \16469 );
nand \U$16237 ( \16483 , \16481 , \16482 );
not \U$16238 ( \16484 , \14705 );
and \U$16239 ( \16485 , \15111 , \16484 );
not \U$16240 ( \16486 , \15111 );
and \U$16241 ( \16487 , \16486 , \14705 );
nor \U$16242 ( \16488 , \16485 , \16487 );
not \U$16243 ( \16489 , \16488 );
not \U$16244 ( \16490 , \16489 );
xor \U$16245 ( \16491 , \16457 , \16459 );
xor \U$16246 ( \16492 , \16491 , \16461 );
not \U$16247 ( \16493 , \15756 );
not \U$16248 ( \16494 , \15755 );
or \U$16249 ( \16495 , \16493 , \16494 );
nand \U$16250 ( \16496 , \15754 , \15752 );
nand \U$16251 ( \16497 , \16495 , \16496 );
xor \U$16252 ( \16498 , \16492 , \16497 );
not \U$16253 ( \16499 , \16498 );
or \U$16254 ( \16500 , \16490 , \16499 );
nand \U$16255 ( \16501 , \16497 , \16492 );
nand \U$16256 ( \16502 , \16500 , \16501 );
xnor \U$16257 ( \16503 , \16483 , \16502 );
not \U$16258 ( \16504 , \16503 );
not \U$16259 ( \16505 , \15341 );
not \U$16260 ( \16506 , \16405 );
or \U$16261 ( \16507 , \16505 , \16506 );
or \U$16262 ( \16508 , \15341 , \16405 );
nand \U$16263 ( \16509 , \16507 , \16508 );
nand \U$16264 ( \16510 , \16504 , \16509 );
not \U$16265 ( \16511 , \16510 );
or \U$16266 ( \16512 , \16407 , \16511 );
not \U$16267 ( \16513 , \15138 );
not \U$16268 ( \16514 , \15132 );
or \U$16269 ( \16515 , \16513 , \16514 );
nand \U$16270 ( \16516 , \15127 , \15121 );
nand \U$16271 ( \16517 , \16515 , \16516 );
xor \U$16272 ( \16518 , \13646 , \13669 );
xor \U$16273 ( \16519 , \16517 , \16518 );
not \U$16274 ( \16520 , \15328 );
nand \U$16275 ( \16521 , \15330 , \16520 );
not \U$16276 ( \16522 , \16521 );
not \U$16277 ( \16523 , \15320 );
or \U$16278 ( \16524 , \16522 , \16523 );
or \U$16279 ( \16525 , \15330 , \16520 );
nand \U$16280 ( \16526 , \16524 , \16525 );
xor \U$16281 ( \16527 , \16519 , \16526 );
not \U$16282 ( \16528 , \13107 );
and \U$16283 ( \16529 , \13169 , \16528 );
not \U$16284 ( \16530 , \13169 );
and \U$16285 ( \16531 , \16530 , \13107 );
nor \U$16286 ( \16532 , \16529 , \16531 );
buf \U$16287 ( \16533 , \13151 );
xor \U$16288 ( \16534 , \16532 , \16533 );
xor \U$16289 ( \16535 , \13230 , \13221 );
xor \U$16290 ( \16536 , \16535 , \13223 );
xor \U$16291 ( \16537 , \16534 , \16536 );
not \U$16292 ( \16538 , \16429 );
not \U$16293 ( \16539 , \16444 );
or \U$16294 ( \16540 , \16538 , \16539 );
not \U$16295 ( \16541 , \16440 );
nand \U$16296 ( \16542 , \16541 , \16433 );
nand \U$16297 ( \16543 , \16540 , \16542 );
not \U$16298 ( \16544 , \16543 );
xor \U$16299 ( \16545 , \16537 , \16544 );
xor \U$16300 ( \16546 , \16527 , \16545 );
not \U$16301 ( \16547 , \15248 );
not \U$16302 ( \16548 , \15335 );
not \U$16303 ( \16549 , \16548 );
or \U$16304 ( \16550 , \16547 , \16549 );
nand \U$16305 ( \16551 , \15247 , \15242 );
nand \U$16306 ( \16552 , \16550 , \16551 );
xor \U$16307 ( \16553 , \16546 , \16552 );
not \U$16308 ( \16554 , \16464 );
not \U$16309 ( \16555 , \16451 );
or \U$16310 ( \16556 , \16554 , \16555 );
nand \U$16311 ( \16557 , \16450 , \16411 );
nand \U$16312 ( \16558 , \16556 , \16557 );
not \U$16313 ( \16559 , \16558 );
not \U$16314 ( \16560 , \16422 );
not \U$16315 ( \16561 , \16445 );
or \U$16316 ( \16562 , \16560 , \16561 );
not \U$16317 ( \16563 , \16412 );
nand \U$16318 ( \16564 , \16563 , \16418 );
nand \U$16319 ( \16565 , \16562 , \16564 );
xor \U$16320 ( \16566 , \13322 , \13381 );
xor \U$16321 ( \16567 , \16566 , \13482 );
not \U$16322 ( \16568 , \16567 );
or \U$16323 ( \16569 , \15238 , \15227 );
nand \U$16324 ( \16570 , \16569 , \15240 );
not \U$16325 ( \16571 , \13189 );
not \U$16326 ( \16572 , \13186 );
or \U$16327 ( \16573 , \16571 , \16572 );
nand \U$16328 ( \16574 , \13185 , \13179 );
nand \U$16329 ( \16575 , \16573 , \16574 );
xor \U$16330 ( \16576 , \16575 , \13195 );
xor \U$16331 ( \16577 , \16570 , \16576 );
not \U$16332 ( \16578 , \16577 );
or \U$16333 ( \16579 , \16568 , \16578 );
or \U$16334 ( \16580 , \16567 , \16577 );
nand \U$16335 ( \16581 , \16579 , \16580 );
and \U$16336 ( \16582 , \16565 , \16581 );
not \U$16337 ( \16583 , \16565 );
not \U$16338 ( \16584 , \16581 );
and \U$16339 ( \16585 , \16583 , \16584 );
nor \U$16340 ( \16586 , \16582 , \16585 );
not \U$16341 ( \16587 , \15139 );
or \U$16342 ( \16588 , \15216 , \15182 );
not \U$16343 ( \16589 , \16588 );
or \U$16344 ( \16590 , \16587 , \16589 );
nand \U$16345 ( \16591 , \15216 , \15182 );
nand \U$16346 ( \16592 , \16590 , \16591 );
not \U$16347 ( \16593 , \16592 );
and \U$16348 ( \16594 , \16586 , \16593 );
not \U$16349 ( \16595 , \16586 );
and \U$16350 ( \16596 , \16595 , \16592 );
nor \U$16351 ( \16597 , \16594 , \16596 );
not \U$16352 ( \16598 , \16597 );
or \U$16353 ( \16599 , \16559 , \16598 );
or \U$16354 ( \16600 , \16597 , \16558 );
nand \U$16355 ( \16601 , \16599 , \16600 );
not \U$16356 ( \16602 , \15217 );
nand \U$16357 ( \16603 , \16602 , \15340 );
not \U$16358 ( \16604 , \15217 );
not \U$16359 ( \16605 , \15339 );
or \U$16360 ( \16606 , \16604 , \16605 );
nand \U$16361 ( \16607 , \16606 , \15116 );
nand \U$16362 ( \16608 , \16603 , \16607 );
not \U$16363 ( \16609 , \16608 );
and \U$16364 ( \16610 , \16601 , \16609 );
not \U$16365 ( \16611 , \16601 );
and \U$16366 ( \16612 , \16611 , \16608 );
nor \U$16367 ( \16613 , \16610 , \16612 );
xor \U$16368 ( \16614 , \16553 , \16613 );
not \U$16369 ( \16615 , \16479 );
not \U$16370 ( \16616 , \16469 );
and \U$16371 ( \16617 , \16615 , \16616 );
and \U$16372 ( \16618 , \16483 , \16502 );
nor \U$16373 ( \16619 , \16617 , \16618 );
xor \U$16374 ( \16620 , \16614 , \16619 );
not \U$16375 ( \16621 , \16620 );
nand \U$16376 ( \16622 , \16512 , \16621 );
not \U$16377 ( \16623 , \16622 );
not \U$16378 ( \16624 , \15940 );
not \U$16379 ( \16625 , \16049 );
or \U$16380 ( \16626 , \16624 , \16625 );
or \U$16381 ( \16627 , \16049 , \15940 );
nand \U$16382 ( \16628 , \16626 , \16627 );
not \U$16383 ( \16629 , \16628 );
xnor \U$16384 ( \16630 , \16156 , \16105 );
not \U$16385 ( \16631 , \16630 );
or \U$16386 ( \16632 , \16629 , \16631 );
or \U$16387 ( \16633 , \16628 , \16630 );
nand \U$16388 ( \16634 , \16632 , \16633 );
not \U$16389 ( \16635 , \16634 );
xor \U$16390 ( \16636 , RIbe296c8_60, RIbe2b2e8_120);
not \U$16391 ( \16637 , \16636 );
not \U$16392 ( \16638 , \8531 );
or \U$16393 ( \16639 , \16637 , \16638 );
nand \U$16394 ( \16640 , \907 , \15489 );
nand \U$16395 ( \16641 , \16639 , \16640 );
xor \U$16396 ( \16642 , RIbe286d8_26, RIbe2b180_117);
not \U$16397 ( \16643 , \16642 );
not \U$16398 ( \16644 , \14852 );
or \U$16399 ( \16645 , \16643 , \16644 );
buf \U$16400 ( \16646 , \14845 );
nand \U$16401 ( \16647 , \16646 , \15380 );
nand \U$16402 ( \16648 , \16645 , \16647 );
or \U$16403 ( \16649 , \16641 , \16648 );
xor \U$16404 ( \16650 , RIbe29e48_76, RIbe295d8_58);
not \U$16405 ( \16651 , \16650 );
not \U$16406 ( \16652 , \4841 );
not \U$16407 ( \16653 , \16652 );
or \U$16408 ( \16654 , \16651 , \16653 );
buf \U$16409 ( \16655 , \4849 );
nand \U$16410 ( \16656 , \16655 , \15403 );
nand \U$16411 ( \16657 , \16654 , \16656 );
nand \U$16412 ( \16658 , \16649 , \16657 );
nand \U$16413 ( \16659 , \16641 , \16648 );
and \U$16414 ( \16660 , \16658 , \16659 );
not \U$16415 ( \16661 , \16660 );
not \U$16416 ( \16662 , \16661 );
not \U$16417 ( \16663 , \15350 );
not \U$16418 ( \16664 , \16663 );
and \U$16419 ( \16665 , RIbe27b98_2, RIbe2b450_123);
xor \U$16420 ( \16666 , RIbe28de0_41, RIbe2abe0_105);
not \U$16421 ( \16667 , \16666 );
not \U$16422 ( \16668 , \11321 );
or \U$16423 ( \16669 , \16667 , \16668 );
nand \U$16424 ( \16670 , \7472 , \15425 );
nand \U$16425 ( \16671 , \16669 , \16670 );
xor \U$16426 ( \16672 , \16665 , \16671 );
xor \U$16427 ( \16673 , RIbe27b20_1, RIbe28480_21);
not \U$16428 ( \16674 , \16673 );
or \U$16429 ( \16675 , \15048 , \16674 );
buf \U$16430 ( \16676 , \2525 );
nand \U$16431 ( \16677 , \16676 , \15647 );
nand \U$16432 ( \16678 , \16675 , \16677 );
and \U$16433 ( \16679 , \16672 , \16678 );
and \U$16434 ( \16680 , \16665 , \16671 );
or \U$16435 ( \16681 , \16679 , \16680 );
not \U$16436 ( \16682 , \16681 );
not \U$16437 ( \16683 , \16682 );
or \U$16438 ( \16684 , \16664 , \16683 );
or \U$16439 ( \16685 , \16682 , \16663 );
nand \U$16440 ( \16686 , \16684 , \16685 );
not \U$16441 ( \16687 , \16686 );
or \U$16442 ( \16688 , \16662 , \16687 );
not \U$16443 ( \16689 , \16682 );
nand \U$16444 ( \16690 , \16689 , \16663 );
nand \U$16445 ( \16691 , \16688 , \16690 );
not \U$16446 ( \16692 , \15466 );
not \U$16447 ( \16693 , \15417 );
not \U$16448 ( \16694 , \16693 );
and \U$16449 ( \16695 , \16692 , \16694 );
and \U$16450 ( \16696 , \15466 , \16693 );
nor \U$16451 ( \16697 , \16695 , \16696 );
xor \U$16452 ( \16698 , \16691 , \16697 );
xor \U$16453 ( \16699 , RIbe28930_31, RIbe2aa00_101);
not \U$16454 ( \16700 , \16699 );
not \U$16455 ( \16701 , \1793 );
or \U$16456 ( \16702 , \16700 , \16701 );
nand \U$16457 ( \16703 , \1199 , \15483 );
nand \U$16458 ( \16704 , \16702 , \16703 );
xor \U$16459 ( \16705 , RIbe27c10_3, RIbe2a640_93);
not \U$16460 ( \16706 , \16705 );
not \U$16461 ( \16707 , \1103 );
or \U$16462 ( \16708 , \16706 , \16707 );
nand \U$16463 ( \16709 , \369 , \15458 );
nand \U$16464 ( \16710 , \16708 , \16709 );
or \U$16465 ( \16711 , \16704 , \16710 );
xor \U$16466 ( \16712 , RIbe2a2f8_86, RIbe282a0_17);
not \U$16467 ( \16713 , \16712 );
not \U$16468 ( \16714 , \8696 );
buf \U$16469 ( \16715 , \16714 );
not \U$16470 ( \16716 , \16715 );
or \U$16471 ( \16717 , \16713 , \16716 );
nand \U$16472 ( \16718 , \11094 , \15433 );
nand \U$16473 ( \16719 , \16717 , \16718 );
nand \U$16474 ( \16720 , \16711 , \16719 );
nand \U$16475 ( \16721 , \16704 , \16710 );
nand \U$16476 ( \16722 , \16720 , \16721 );
not \U$16477 ( \16723 , \16722 );
xor \U$16478 ( \16724 , RIbe28048_12, RIbe2af28_112);
not \U$16479 ( \16725 , \16724 );
not \U$16480 ( \16726 , \14423 );
or \U$16481 ( \16727 , \16725 , \16726 );
not \U$16482 ( \16728 , \14412 );
nand \U$16483 ( \16729 , \16728 , \15343 );
nand \U$16484 ( \16730 , \16727 , \16729 );
xor \U$16485 ( \16731 , RIbe27df0_7, RIbe27fd0_11);
not \U$16486 ( \16732 , \16731 );
not \U$16487 ( \16733 , \9825 );
or \U$16488 ( \16734 , \16732 , \16733 );
nand \U$16489 ( \16735 , \2707 , \15627 );
nand \U$16490 ( \16736 , \16734 , \16735 );
nor \U$16491 ( \16737 , \16730 , \16736 );
xor \U$16492 ( \16738 , RIbe27d78_6, RIbe2b4c8_124);
and \U$16493 ( \16739 , \5739 , \16738 );
and \U$16494 ( \16740 , \314 , \15511 );
nor \U$16495 ( \16741 , \16739 , \16740 );
or \U$16496 ( \16742 , \16737 , \16741 );
nand \U$16497 ( \16743 , \16730 , \16736 );
nand \U$16498 ( \16744 , \16742 , \16743 );
not \U$16499 ( \16745 , \16744 );
xor \U$16500 ( \16746 , RIbe27b98_2, RIbe2a730_95);
not \U$16501 ( \16747 , \16746 );
not \U$16502 ( \16748 , \9833 );
or \U$16503 ( \16749 , \16747 , \16748 );
nand \U$16504 ( \16750 , \7584 , \15638 );
nand \U$16505 ( \16751 , \16749 , \16750 );
xor \U$16506 ( \16752 , RIbe28d68_40, RIbe27e68_8);
not \U$16507 ( \16753 , \16752 );
not \U$16508 ( \16754 , \2457 );
or \U$16509 ( \16755 , \16753 , \16754 );
nand \U$16510 ( \16756 , \2463 , \15449 );
nand \U$16511 ( \16757 , \16755 , \16756 );
xor \U$16512 ( \16758 , \16751 , \16757 );
xor \U$16513 ( \16759 , RIbe297b8_62, RIbe2a028_80);
not \U$16514 ( \16760 , \16759 );
not \U$16515 ( \16761 , \8401 );
or \U$16516 ( \16762 , \16760 , \16761 );
nand \U$16517 ( \16763 , \8172 , \15419 );
nand \U$16518 ( \16764 , \16762 , \16763 );
nand \U$16519 ( \16765 , \16758 , \16764 );
nand \U$16520 ( \16766 , \16751 , \16757 );
nand \U$16521 ( \16767 , \16765 , \16766 );
not \U$16522 ( \16768 , \16767 );
not \U$16523 ( \16769 , \16768 );
or \U$16524 ( \16770 , \16745 , \16769 );
not \U$16525 ( \16771 , \16766 );
not \U$16526 ( \16772 , \16765 );
or \U$16527 ( \16773 , \16771 , \16772 );
not \U$16528 ( \16774 , \16744 );
nand \U$16529 ( \16775 , \16773 , \16774 );
nand \U$16530 ( \16776 , \16770 , \16775 );
not \U$16531 ( \16777 , \16776 );
or \U$16532 ( \16778 , \16723 , \16777 );
nand \U$16533 ( \16779 , \16767 , \16744 );
nand \U$16534 ( \16780 , \16778 , \16779 );
xnor \U$16535 ( \16781 , \16698 , \16780 );
xor \U$16536 ( \16782 , RIbe2a2f8_86, RIbe28138_14);
not \U$16537 ( \16783 , \16782 );
not \U$16538 ( \16784 , \10446 );
or \U$16539 ( \16785 , \16783 , \16784 );
nand \U$16540 ( \16786 , \8706 , \16712 );
nand \U$16541 ( \16787 , \16785 , \16786 );
not \U$16542 ( \16788 , \16787 );
xor \U$16543 ( \16789 , RIbe2a7a8_96, RIbe28de0_41);
not \U$16544 ( \16790 , \16789 );
not \U$16545 ( \16791 , \923 );
or \U$16546 ( \16792 , \16790 , \16791 );
nand \U$16547 ( \16793 , \346 , \16666 );
nand \U$16548 ( \16794 , \16792 , \16793 );
not \U$16549 ( \16795 , \16794 );
xor \U$16550 ( \16796 , RIbe29740_61, RIbe2a028_80);
not \U$16551 ( \16797 , \16796 );
not \U$16552 ( \16798 , \8400 );
or \U$16553 ( \16799 , \16797 , \16798 );
nand \U$16554 ( \16800 , \8930 , \16759 );
nand \U$16555 ( \16801 , \16799 , \16800 );
xnor \U$16556 ( \16802 , \16795 , \16801 );
not \U$16557 ( \16803 , \16802 );
or \U$16558 ( \16804 , \16788 , \16803 );
not \U$16559 ( \16805 , \16795 );
nand \U$16560 ( \16806 , \16805 , \16801 );
nand \U$16561 ( \16807 , \16804 , \16806 );
not \U$16562 ( \16808 , \16807 );
xor \U$16563 ( \16809 , RIbe2b018_114, RIbe29380_53);
not \U$16564 ( \16810 , \16809 );
not \U$16565 ( \16811 , \15965 );
buf \U$16566 ( \16812 , \16811 );
not \U$16567 ( \16813 , \16812 );
or \U$16568 ( \16814 , \16810 , \16813 );
nand \U$16569 ( \16815 , \15953 , RIbe2b018_114);
nand \U$16570 ( \16816 , \16814 , \16815 );
not \U$16571 ( \16817 , \16816 );
xor \U$16572 ( \16818 , RIbe27b98_2, RIbe2b450_123);
and \U$16573 ( \16819 , \16818 , \9833 );
and \U$16574 ( \16820 , \7584 , \16746 );
nor \U$16575 ( \16821 , \16819 , \16820 );
not \U$16576 ( \16822 , \16821 );
xor \U$16577 ( \16823 , RIbe2b540_125, RIbe290b0_47);
not \U$16578 ( \16824 , \16823 );
not \U$16579 ( \16825 , \2729 );
or \U$16580 ( \16826 , \16824 , \16825 );
nand \U$16581 ( \16827 , \398 , \15983 );
nand \U$16582 ( \16828 , \16826 , \16827 );
not \U$16583 ( \16829 , \16828 );
or \U$16584 ( \16830 , \16822 , \16829 );
or \U$16585 ( \16831 , \16821 , \16828 );
nand \U$16586 ( \16832 , \16830 , \16831 );
not \U$16587 ( \16833 , \16832 );
or \U$16588 ( \16834 , \16817 , \16833 );
not \U$16589 ( \16835 , \16821 );
nand \U$16590 ( \16836 , \16835 , \16828 );
nand \U$16591 ( \16837 , \16834 , \16836 );
not \U$16592 ( \16838 , \16837 );
xor \U$16593 ( \16839 , RIbe29b00_69, RIbe29c68_72);
not \U$16594 ( \16840 , \16839 );
not \U$16595 ( \16841 , \8259 );
or \U$16596 ( \16842 , \16840 , \16841 );
nand \U$16597 ( \16843 , \4580 , \16016 );
nand \U$16598 ( \16844 , \16842 , \16843 );
not \U$16599 ( \16845 , \16844 );
xor \U$16600 ( \16846 , RIbe29e48_76, RIbe291a0_49);
not \U$16601 ( \16847 , \16846 );
not \U$16602 ( \16848 , \14307 );
or \U$16603 ( \16849 , \16847 , \16848 );
nand \U$16604 ( \16850 , \4849 , \16650 );
nand \U$16605 ( \16851 , \16849 , \16850 );
xor \U$16606 ( \16852 , RIbe29038_46, RIbe2adc0_109);
not \U$16607 ( \16853 , \16852 );
buf \U$16608 ( \16854 , \280 );
not \U$16609 ( \16855 , \16854 );
or \U$16610 ( \16856 , \16853 , \16855 );
xor \U$16611 ( \16857 , RIbe29038_46, RIbe2a460_89);
nand \U$16612 ( \16858 , \286 , \16857 );
nand \U$16613 ( \16859 , \16856 , \16858 );
xor \U$16614 ( \16860 , \16851 , \16859 );
not \U$16615 ( \16861 , \16860 );
or \U$16616 ( \16862 , \16845 , \16861 );
nand \U$16617 ( \16863 , \16851 , \16859 );
nand \U$16618 ( \16864 , \16862 , \16863 );
not \U$16619 ( \16865 , \16864 );
not \U$16620 ( \16866 , \16865 );
or \U$16621 ( \16867 , \16838 , \16866 );
or \U$16622 ( \16868 , \16837 , \16865 );
nand \U$16623 ( \16869 , \16867 , \16868 );
not \U$16624 ( \16870 , \16869 );
or \U$16625 ( \16871 , \16808 , \16870 );
nand \U$16626 ( \16872 , \16864 , \16837 );
nand \U$16627 ( \16873 , \16871 , \16872 );
not \U$16628 ( \16874 , \16873 );
buf \U$16629 ( \16875 , \13533 );
not \U$16630 ( \16876 , \16875 );
not \U$16631 ( \16877 , \16876 );
not \U$16632 ( \16878 , \15505 );
not \U$16633 ( \16879 , \16878 );
and \U$16634 ( \16880 , \16877 , \16879 );
xor \U$16635 ( \16881 , RIbe28840_29, RIbe2b108_116);
and \U$16636 ( \16882 , \13543 , \16881 );
nor \U$16637 ( \16883 , \16880 , \16882 );
not \U$16638 ( \16884 , \16883 );
not \U$16639 ( \16885 , \16884 );
xor \U$16640 ( \16886 , RIbe29ce0_73, RIbe28390_19);
not \U$16641 ( \16887 , \16886 );
not \U$16642 ( \16888 , \2639 );
or \U$16643 ( \16889 , \16887 , \16888 );
nand \U$16644 ( \16890 , \2777 , \15555 );
nand \U$16645 ( \16891 , \16889 , \16890 );
not \U$16646 ( \16892 , \16891 );
xor \U$16647 ( \16893 , RIbe2b108_116, RIbe28750_27);
not \U$16648 ( \16894 , \16893 );
not \U$16649 ( \16895 , \14297 );
or \U$16650 ( \16896 , \16894 , \16895 );
not \U$16651 ( \16897 , \13533 );
not \U$16652 ( \16898 , \16897 );
nand \U$16653 ( \16899 , \16898 , \16881 );
nand \U$16654 ( \16900 , \16896 , \16899 );
not \U$16655 ( \16901 , \16900 );
not \U$16656 ( \16902 , \16901 );
or \U$16657 ( \16903 , \16892 , \16902 );
or \U$16658 ( \16904 , \16891 , \16901 );
nand \U$16659 ( \16905 , \16903 , \16904 );
not \U$16660 ( \16906 , \16905 );
or \U$16661 ( \16907 , \16885 , \16906 );
nand \U$16662 ( \16908 , \16891 , \16900 );
nand \U$16663 ( \16909 , \16907 , \16908 );
not \U$16664 ( \16910 , \16909 );
xor \U$16665 ( \16911 , RIbe27ee0_9, RIbe2af28_112);
not \U$16666 ( \16912 , \16911 );
buf \U$16667 ( \16913 , \14423 );
buf \U$16668 ( \16914 , \16913 );
not \U$16669 ( \16915 , \16914 );
or \U$16670 ( \16916 , \16912 , \16915 );
not \U$16671 ( \16917 , \14412 );
nand \U$16672 ( \16918 , \16917 , \16724 );
nand \U$16673 ( \16919 , \16916 , \16918 );
not \U$16674 ( \16920 , \16919 );
xor \U$16675 ( \16921 , RIbe2a550_91, RIbe293f8_54);
not \U$16676 ( \16922 , \16921 );
not \U$16677 ( \16923 , \12000 );
or \U$16678 ( \16924 , \16922 , \16923 );
nand \U$16679 ( \16925 , \11485 , \15989 );
nand \U$16680 ( \16926 , \16924 , \16925 );
not \U$16681 ( \16927 , \16926 );
xor \U$16682 ( \16928 , RIbe2a118_82, RIbe28228_16);
and \U$16683 ( \16929 , \879 , \16928 );
xor \U$16684 ( \16930 , RIbe28228_16, RIbe2a820_97);
and \U$16685 ( \16931 , \8680 , \16930 );
nor \U$16686 ( \16932 , \16929 , \16931 );
not \U$16687 ( \16933 , \16932 );
or \U$16688 ( \16934 , \16927 , \16933 );
or \U$16689 ( \16935 , \16926 , \16932 );
nand \U$16690 ( \16936 , \16934 , \16935 );
not \U$16691 ( \16937 , \16936 );
or \U$16692 ( \16938 , \16920 , \16937 );
not \U$16693 ( \16939 , \16932 );
nand \U$16694 ( \16940 , \16939 , \16926 );
nand \U$16695 ( \16941 , \16938 , \16940 );
not \U$16696 ( \16942 , \16941 );
xor \U$16697 ( \16943 , RIbe28390_19, RIbe29d58_74);
not \U$16698 ( \16944 , \16943 );
not \U$16699 ( \16945 , \14579 );
or \U$16700 ( \16946 , \16944 , \16945 );
nand \U$16701 ( \16947 , \8868 , \16886 );
nand \U$16702 ( \16948 , \16946 , \16947 );
not \U$16703 ( \16949 , \16948 );
xor \U$16704 ( \16950 , RIbe28480_21, RIbe29b78_70);
not \U$16705 ( \16951 , \16950 );
xor \U$16706 ( \16952 , RIbe28480_21, RIbe287c8_28);
and \U$16707 ( \16953 , \16952 , \2514 , \2516 );
not \U$16708 ( \16954 , \16953 );
or \U$16709 ( \16955 , \16951 , \16954 );
nand \U$16710 ( \16956 , \16676 , \16673 );
nand \U$16711 ( \16957 , \16955 , \16956 );
xor \U$16712 ( \16958 , RIbe28930_31, RIbe2a898_98);
not \U$16713 ( \16959 , \16958 );
not \U$16714 ( \16960 , \8887 );
or \U$16715 ( \16961 , \16959 , \16960 );
nand \U$16716 ( \16962 , \970 , \16699 );
nand \U$16717 ( \16963 , \16961 , \16962 );
xor \U$16718 ( \16964 , \16957 , \16963 );
not \U$16719 ( \16965 , \16964 );
or \U$16720 ( \16966 , \16949 , \16965 );
nand \U$16721 ( \16967 , \16963 , \16957 );
nand \U$16722 ( \16968 , \16966 , \16967 );
and \U$16723 ( \16969 , RIbe2b3d8_122, RIbe27b98_2);
xor \U$16724 ( \16970 , RIbe285e8_24, RIbe28cf0_39);
not \U$16725 ( \16971 , \16970 );
not \U$16726 ( \16972 , \11174 );
or \U$16727 ( \16973 , \16971 , \16972 );
not \U$16728 ( \16974 , \16013 );
nand \U$16729 ( \16975 , \16974 , \8270 );
nand \U$16730 ( \16976 , \16973 , \16975 );
xor \U$16731 ( \16977 , \16969 , \16976 );
xor \U$16732 ( \16978 , RIbe2ac58_106, RIbe27c10_3);
not \U$16733 ( \16979 , \16978 );
not \U$16734 ( \16980 , \1103 );
or \U$16735 ( \16981 , \16979 , \16980 );
nand \U$16736 ( \16982 , \1173 , \16705 );
nand \U$16737 ( \16983 , \16981 , \16982 );
and \U$16738 ( \16984 , \16977 , \16983 );
and \U$16739 ( \16985 , \16969 , \16976 );
or \U$16740 ( \16986 , \16984 , \16985 );
xor \U$16741 ( \16987 , \16968 , \16986 );
not \U$16742 ( \16988 , \16987 );
or \U$16743 ( \16989 , \16942 , \16988 );
nand \U$16744 ( \16990 , \16968 , \16986 );
nand \U$16745 ( \16991 , \16989 , \16990 );
not \U$16746 ( \16992 , \16991 );
not \U$16747 ( \16993 , \16992 );
or \U$16748 ( \16994 , \16910 , \16993 );
not \U$16749 ( \16995 , \16909 );
nand \U$16750 ( \16996 , \16995 , \16991 );
nand \U$16751 ( \16997 , \16994 , \16996 );
not \U$16752 ( \16998 , \16997 );
or \U$16753 ( \16999 , \16874 , \16998 );
nand \U$16754 ( \17000 , \16991 , \16909 );
nand \U$16755 ( \17001 , \16999 , \17000 );
xor \U$16756 ( \17002 , \16781 , \17001 );
xor \U$16757 ( \17003 , \15412 , \15399 );
xor \U$16758 ( \17004 , RIbe294e8_56, RIbe2a3e8_88);
not \U$16759 ( \17005 , \17004 );
not \U$16760 ( \17006 , \8806 );
or \U$16761 ( \17007 , \17005 , \17006 );
nand \U$16762 ( \17008 , \8794 , \15477 );
nand \U$16763 ( \17009 , \17007 , \17008 );
xor \U$16764 ( \17010 , RIbe28a20_33, RIbe2b6a8_128);
not \U$16765 ( \17011 , \17010 );
not \U$16766 ( \17012 , \1780 );
or \U$16767 ( \17013 , \17011 , \17012 );
nand \U$16768 ( \17014 , \5055 , \15548 );
nand \U$16769 ( \17015 , \17013 , \17014 );
nor \U$16770 ( \17016 , \17009 , \17015 );
buf \U$16771 ( \17017 , \17016 );
not \U$16772 ( \17018 , \16857 );
not \U$16773 ( \17019 , \979 );
or \U$16774 ( \17020 , \17018 , \17019 );
nand \U$16775 ( \17021 , \287 , \15673 );
nand \U$16776 ( \17022 , \17020 , \17021 );
not \U$16777 ( \17023 , \17022 );
or \U$16778 ( \17024 , \17017 , \17023 );
nand \U$16779 ( \17025 , \17015 , \17009 );
nand \U$16780 ( \17026 , \17024 , \17025 );
xor \U$16781 ( \17027 , RIbe28c78_38, RIbe2a190_83);
not \U$16782 ( \17028 , \17027 );
not \U$16783 ( \17029 , \11396 );
or \U$16784 ( \17030 , \17028 , \17029 );
nand \U$16785 ( \17031 , \15693 , \15688 );
nand \U$16786 ( \17032 , \17030 , \17031 );
not \U$16787 ( \17033 , \17032 );
xor \U$16788 ( \17034 , RIbe284f8_22, RIbe2a280_85);
not \U$16789 ( \17035 , \17034 );
not \U$16790 ( \17036 , \13268 );
or \U$16791 ( \17037 , \17035 , \17036 );
nand \U$16792 ( \17038 , \14649 , \15664 );
nand \U$16793 ( \17039 , \17037 , \17038 );
not \U$16794 ( \17040 , \16930 );
not \U$16795 ( \17041 , \14638 );
or \U$16796 ( \17042 , \17040 , \17041 );
nand \U$16797 ( \17043 , \885 , \15442 );
nand \U$16798 ( \17044 , \17042 , \17043 );
xor \U$16799 ( \17045 , \17039 , \17044 );
not \U$16800 ( \17046 , \17045 );
or \U$16801 ( \17047 , \17033 , \17046 );
nand \U$16802 ( \17048 , \17039 , \17044 );
nand \U$16803 ( \17049 , \17047 , \17048 );
and \U$16804 ( \17050 , \17026 , \17049 );
not \U$16805 ( \17051 , \17026 );
not \U$16806 ( \17052 , \17049 );
and \U$16807 ( \17053 , \17051 , \17052 );
nor \U$16808 ( \17054 , \17050 , \17053 );
xor \U$16809 ( \17055 , \17003 , \17054 );
xor \U$16810 ( \17056 , \15981 , \16008 );
xor \U$16811 ( \17057 , \17056 , \16031 );
xor \U$16812 ( \17058 , \17055 , \17057 );
not \U$16813 ( \17059 , \9262 );
not \U$16814 ( \17060 , \17059 );
xor \U$16815 ( \17061 , RIbe2a3e8_88, RIbe29470_55);
and \U$16816 ( \17062 , \17060 , \17061 );
and \U$16817 ( \17063 , \10476 , \17004 );
nor \U$16818 ( \17064 , \17062 , \17063 );
not \U$16819 ( \17065 , \17064 );
not \U$16820 ( \17066 , \17065 );
xor \U$16821 ( \17067 , RIbe296c8_60, RIbe2a4d8_90);
not \U$16822 ( \17068 , \17067 );
not \U$16823 ( \17069 , \10812 );
or \U$16824 ( \17070 , \17068 , \17069 );
nand \U$16825 ( \17071 , \8534 , \16636 );
nand \U$16826 ( \17072 , \17070 , \17071 );
not \U$16827 ( \17073 , \17072 );
not \U$16828 ( \17074 , \17073 );
xor \U$16829 ( \17075 , RIbe288b8_30, RIbe2a910_99);
not \U$16830 ( \17076 , \17075 );
not \U$16831 ( \17077 , \10987 );
or \U$16832 ( \17078 , \17076 , \17077 );
nand \U$16833 ( \17079 , \10400 , \15973 );
nand \U$16834 ( \17080 , \17078 , \17079 );
not \U$16835 ( \17081 , \17080 );
or \U$16836 ( \17082 , \17074 , \17081 );
or \U$16837 ( \17083 , \17080 , \17073 );
nand \U$16838 ( \17084 , \17082 , \17083 );
not \U$16839 ( \17085 , \17084 );
or \U$16840 ( \17086 , \17066 , \17085 );
nand \U$16841 ( \17087 , \17080 , \17072 );
nand \U$16842 ( \17088 , \17086 , \17087 );
not \U$16843 ( \17089 , \17088 );
xor \U$16844 ( \17090 , RIbe280c0_13, RIbe2b360_121);
not \U$16845 ( \17091 , \17090 );
not \U$16846 ( \17092 , \8624 );
or \U$16847 ( \17093 , \17091 , \17092 );
nand \U$16848 ( \17094 , \869 , \15945 );
nand \U$16849 ( \17095 , \17093 , \17094 );
xor \U$16850 ( \17096 , RIbe28c00_37, RIbe2a190_83);
not \U$16851 ( \17097 , \17096 );
not \U$16852 ( \17098 , \11396 );
or \U$16853 ( \17099 , \17097 , \17098 );
nand \U$16854 ( \17100 , \11400 , \17027 );
nand \U$16855 ( \17101 , \17099 , \17100 );
or \U$16856 ( \17102 , \17095 , \17101 );
xor \U$16857 ( \17103 , RIbe29f38_78, RIbe28b88_36);
not \U$16858 ( \17104 , \17103 );
not \U$16859 ( \17105 , \3401 );
or \U$16860 ( \17106 , \17104 , \17105 );
not \U$16861 ( \17107 , \16026 );
nand \U$16862 ( \17108 , \17107 , \7550 );
nand \U$16863 ( \17109 , \17106 , \17108 );
nand \U$16864 ( \17110 , \17102 , \17109 );
nand \U$16865 ( \17111 , \17095 , \17101 );
nand \U$16866 ( \17112 , \17110 , \17111 );
not \U$16867 ( \17113 , \17112 );
xor \U$16868 ( \17114 , RIbe27c88_4, RIbe27fd0_11);
not \U$16869 ( \17115 , \17114 );
not \U$16870 ( \17116 , \9825 );
or \U$16871 ( \17117 , \17115 , \17116 );
nand \U$16872 ( \17118 , \2707 , \16731 );
nand \U$16873 ( \17119 , \17117 , \17118 );
xor \U$16874 ( \17120 , RIbe28a20_33, RIbe2aa78_102);
not \U$16875 ( \17121 , \17120 );
not \U$16876 ( \17122 , \1780 );
or \U$16877 ( \17123 , \17121 , \17122 );
nand \U$16878 ( \17124 , \2475 , \17010 );
nand \U$16879 ( \17125 , \17123 , \17124 );
or \U$16880 ( \17126 , \17119 , \17125 );
xor \U$16881 ( \17127 , RIbe27d78_6, RIbe2a6b8_94);
not \U$16882 ( \17128 , \17127 );
not \U$16883 ( \17129 , \8768 );
or \U$16884 ( \17130 , \17128 , \17129 );
nand \U$16885 ( \17131 , \314 , \16738 );
nand \U$16886 ( \17132 , \17130 , \17131 );
nand \U$16887 ( \17133 , \17126 , \17132 );
nand \U$16888 ( \17134 , \17125 , \17119 );
nand \U$16889 ( \17135 , \17133 , \17134 );
not \U$16890 ( \17136 , \17135 );
not \U$16891 ( \17137 , \17136 );
or \U$16892 ( \17138 , \17113 , \17137 );
or \U$16893 ( \17139 , \17136 , \17112 );
nand \U$16894 ( \17140 , \17138 , \17139 );
not \U$16895 ( \17141 , \17140 );
or \U$16896 ( \17142 , \17089 , \17141 );
nand \U$16897 ( \17143 , \17135 , \17112 );
nand \U$16898 ( \17144 , \17142 , \17143 );
not \U$16899 ( \17145 , \17144 );
not \U$16900 ( \17146 , \17145 );
and \U$16901 ( \17147 , \17058 , \17146 );
and \U$16902 ( \17148 , \17055 , \17057 );
or \U$16903 ( \17149 , \17147 , \17148 );
not \U$16904 ( \17150 , \17149 );
not \U$16905 ( \17151 , \17150 );
and \U$16906 ( \17152 , \17002 , \17151 );
and \U$16907 ( \17153 , \16781 , \17001 );
or \U$16908 ( \17154 , \17152 , \17153 );
not \U$16909 ( \17155 , \17154 );
or \U$16910 ( \17156 , \16635 , \17155 );
not \U$16911 ( \17157 , \16630 );
nand \U$16912 ( \17158 , \17157 , \16628 );
nand \U$16913 ( \17159 , \17156 , \17158 );
not \U$16914 ( \17160 , \17159 );
not \U$16915 ( \17161 , \17160 );
xor \U$16916 ( \17162 , \16184 , \16161 );
xnor \U$16917 ( \17163 , \17162 , \16199 );
not \U$16918 ( \17164 , \17163 );
and \U$16919 ( \17165 , \16071 , \16053 );
not \U$16920 ( \17166 , \16071 );
not \U$16921 ( \17167 , \16053 );
and \U$16922 ( \17168 , \17166 , \17167 );
nor \U$16923 ( \17169 , \17165 , \17168 );
not \U$16924 ( \17170 , \17169 );
or \U$16925 ( \17171 , \17164 , \17170 );
or \U$16926 ( \17172 , \17169 , \17163 );
nand \U$16927 ( \17173 , \17171 , \17172 );
buf \U$16928 ( \17174 , \17173 );
not \U$16929 ( \17175 , \17174 );
or \U$16930 ( \17176 , \17161 , \17175 );
or \U$16931 ( \17177 , \17174 , \17160 );
nand \U$16932 ( \17178 , \17176 , \17177 );
not \U$16933 ( \17179 , \17178 );
buf \U$16934 ( \17180 , \16288 );
xor \U$16935 ( \17181 , \17180 , \16291 );
xor \U$16936 ( \17182 , \16268 , \16259 );
or \U$16937 ( \17183 , \17181 , \17182 );
xor \U$16938 ( \17184 , \16299 , \16302 );
xnor \U$16939 ( \17185 , \17184 , \16304 );
nand \U$16940 ( \17186 , \17183 , \17185 );
nand \U$16941 ( \17187 , \17181 , \17182 );
nand \U$16942 ( \17188 , \17186 , \17187 );
not \U$16943 ( \17189 , \16234 );
not \U$16944 ( \17190 , \17189 );
buf \U$16945 ( \17191 , \16248 );
not \U$16946 ( \17192 , \17191 );
or \U$16947 ( \17193 , \17190 , \17192 );
or \U$16948 ( \17194 , \17191 , \17189 );
nand \U$16949 ( \17195 , \17193 , \17194 );
xor \U$16950 ( \17196 , \17188 , \17195 );
not \U$16951 ( \17197 , \16313 );
not \U$16952 ( \17198 , \17197 );
xor \U$16953 ( \17199 , \16276 , \16296 );
not \U$16954 ( \17200 , \17199 );
or \U$16955 ( \17201 , \17198 , \17200 );
or \U$16956 ( \17202 , \17199 , \17197 );
nand \U$16957 ( \17203 , \17201 , \17202 );
and \U$16958 ( \17204 , \17196 , \17203 );
and \U$16959 ( \17205 , \17188 , \17195 );
or \U$16960 ( \17206 , \17204 , \17205 );
buf \U$16961 ( \17207 , \16321 );
buf \U$16962 ( \17208 , \16232 );
not \U$16963 ( \17209 , \17208 );
and \U$16964 ( \17210 , \17207 , \17209 );
not \U$16965 ( \17211 , \17207 );
and \U$16966 ( \17212 , \17211 , \17208 );
nor \U$16967 ( \17213 , \17210 , \17212 );
not \U$16968 ( \17214 , \17213 );
xor \U$16969 ( \17215 , \17206 , \17214 );
not \U$16970 ( \17216 , \16697 );
not \U$16971 ( \17217 , \17216 );
xor \U$16972 ( \17218 , \16691 , \16780 );
not \U$16973 ( \17219 , \17218 );
or \U$16974 ( \17220 , \17217 , \17219 );
nand \U$16975 ( \17221 , \16780 , \16691 );
nand \U$16976 ( \17222 , \17220 , \17221 );
not \U$16977 ( \17223 , \17222 );
xor \U$16978 ( \17224 , \15546 , \15562 );
not \U$16979 ( \17225 , \17224 );
xor \U$16980 ( \17226 , \15447 , \15463 );
xor \U$16981 ( \17227 , \17226 , \15454 );
not \U$16982 ( \17228 , \15695 );
and \U$16983 ( \17229 , \15709 , \17228 );
not \U$16984 ( \17230 , \15709 );
and \U$16985 ( \17231 , \17230 , \15695 );
or \U$16986 ( \17232 , \17229 , \17231 );
xor \U$16987 ( \17233 , \17227 , \17232 );
not \U$16988 ( \17234 , \17233 );
or \U$16989 ( \17235 , \17225 , \17234 );
nand \U$16990 ( \17236 , \17232 , \17227 );
nand \U$16991 ( \17237 , \17235 , \17236 );
not \U$16992 ( \17238 , \17237 );
not \U$16993 ( \17239 , \17003 );
not \U$16994 ( \17240 , \17054 );
or \U$16995 ( \17241 , \17239 , \17240 );
nand \U$16996 ( \17242 , \17049 , \17026 );
nand \U$16997 ( \17243 , \17241 , \17242 );
xor \U$16998 ( \17244 , \15431 , \15438 );
buf \U$16999 ( \17245 , \15424 );
xnor \U$17000 ( \17246 , \17244 , \17245 );
xor \U$17001 ( \17247 , \15365 , \15375 );
xor \U$17002 ( \17248 , \17247 , \15385 );
nand \U$17003 ( \17249 , \17246 , \17248 );
not \U$17004 ( \17250 , \17249 );
xor \U$17005 ( \17251 , \15669 , \15662 );
xor \U$17006 ( \17252 , \17251 , \15678 );
not \U$17007 ( \17253 , \17252 );
or \U$17008 ( \17254 , \17250 , \17253 );
not \U$17009 ( \17255 , \17248 );
not \U$17010 ( \17256 , \17246 );
nand \U$17011 ( \17257 , \17255 , \17256 );
nand \U$17012 ( \17258 , \17254 , \17257 );
xor \U$17013 ( \17259 , \17243 , \17258 );
not \U$17014 ( \17260 , \17259 );
or \U$17015 ( \17261 , \17238 , \17260 );
nand \U$17016 ( \17262 , \17243 , \17258 );
nand \U$17017 ( \17263 , \17261 , \17262 );
not \U$17018 ( \17264 , \17263 );
not \U$17019 ( \17265 , \17264 );
or \U$17020 ( \17266 , \17223 , \17265 );
or \U$17021 ( \17267 , \17264 , \17222 );
nand \U$17022 ( \17268 , \17266 , \17267 );
not \U$17023 ( \17269 , \17268 );
buf \U$17024 ( \17270 , \15538 );
xor \U$17025 ( \17271 , \17270 , \15567 );
not \U$17026 ( \17272 , \17271 );
xor \U$17027 ( \17273 , \15632 , \15643 );
xnor \U$17028 ( \17274 , \17273 , \15653 );
not \U$17029 ( \17275 , \17274 );
not \U$17030 ( \17276 , \15481 );
and \U$17031 ( \17277 , \15499 , \17276 );
not \U$17032 ( \17278 , \15499 );
and \U$17033 ( \17279 , \17278 , \15481 );
nor \U$17034 ( \17280 , \17277 , \17279 );
not \U$17035 ( \17281 , \17280 );
nand \U$17036 ( \17282 , \17275 , \17281 );
not \U$17037 ( \17283 , \17280 );
not \U$17038 ( \17284 , \17274 );
or \U$17039 ( \17285 , \17283 , \17284 );
xor \U$17040 ( \17286 , \15510 , \15516 );
xor \U$17041 ( \17287 , \17286 , \15523 );
nand \U$17042 ( \17288 , \17285 , \17287 );
nand \U$17043 ( \17289 , \17282 , \17288 );
not \U$17044 ( \17290 , \17289 );
and \U$17045 ( \17291 , \15655 , \15681 );
not \U$17046 ( \17292 , \15655 );
and \U$17047 ( \17293 , \17292 , \15680 );
nor \U$17048 ( \17294 , \17291 , \17293 );
xor \U$17049 ( \17295 , \17294 , \15713 );
not \U$17050 ( \17296 , \17295 );
or \U$17051 ( \17297 , \17290 , \17296 );
or \U$17052 ( \17298 , \17289 , \17295 );
nand \U$17053 ( \17299 , \17297 , \17298 );
nand \U$17054 ( \17300 , \17272 , \17299 );
not \U$17055 ( \17301 , \17295 );
nand \U$17056 ( \17302 , \17301 , \17289 );
and \U$17057 ( \17303 , \17300 , \17302 );
not \U$17058 ( \17304 , \17303 );
not \U$17059 ( \17305 , \17304 );
or \U$17060 ( \17306 , \17269 , \17305 );
nand \U$17061 ( \17307 , \17263 , \17222 );
nand \U$17062 ( \17308 , \17306 , \17307 );
not \U$17063 ( \17309 , \17308 );
xor \U$17064 ( \17310 , \17215 , \17309 );
xor \U$17065 ( \17311 , \17268 , \17303 );
not \U$17066 ( \17312 , \17311 );
not \U$17067 ( \17313 , \17312 );
not \U$17068 ( \17314 , \17299 );
not \U$17069 ( \17315 , \17271 );
and \U$17070 ( \17316 , \17314 , \17315 );
and \U$17071 ( \17317 , \17299 , \17271 );
nor \U$17072 ( \17318 , \17316 , \17317 );
not \U$17073 ( \17319 , \17318 );
xnor \U$17074 ( \17320 , \17259 , \17237 );
not \U$17075 ( \17321 , \17320 );
or \U$17076 ( \17322 , \17319 , \17321 );
not \U$17077 ( \17323 , \17252 );
and \U$17078 ( \17324 , \17248 , \17246 );
not \U$17079 ( \17325 , \17248 );
and \U$17080 ( \17326 , \17325 , \17256 );
nor \U$17081 ( \17327 , \17324 , \17326 );
not \U$17082 ( \17328 , \17327 );
not \U$17083 ( \17329 , \17328 );
or \U$17084 ( \17330 , \17323 , \17329 );
not \U$17085 ( \17331 , \17252 );
nand \U$17086 ( \17332 , \17331 , \17327 );
nand \U$17087 ( \17333 , \17330 , \17332 );
not \U$17088 ( \17334 , \17333 );
xor \U$17089 ( \17335 , \16665 , \16671 );
xor \U$17090 ( \17336 , \17335 , \16678 );
xor \U$17091 ( \17337 , \16758 , \16764 );
xor \U$17092 ( \17338 , \17336 , \17337 );
xor \U$17093 ( \17339 , RIbe29998_66, RIbe27e68_8);
not \U$17094 ( \17340 , \17339 );
not \U$17095 ( \17341 , \4443 );
or \U$17096 ( \17342 , \17340 , \17341 );
nand \U$17097 ( \17343 , \4447 , \16752 );
nand \U$17098 ( \17344 , \17342 , \17343 );
not \U$17099 ( \17345 , \17344 );
xor \U$17100 ( \17346 , RIbe28f48_44, RIbe29218_50);
not \U$17101 ( \17347 , \17346 );
not \U$17102 ( \17348 , \8221 );
or \U$17103 ( \17349 , \17347 , \17348 );
nand \U$17104 ( \17350 , \3249 , \15999 );
nand \U$17105 ( \17351 , \17349 , \17350 );
not \U$17106 ( \17352 , \17351 );
or \U$17107 ( \17353 , \17345 , \17352 );
or \U$17108 ( \17354 , \17344 , \17351 );
xor \U$17109 ( \17355 , RIbe28570_23, RIbe2b180_117);
not \U$17110 ( \17356 , \17355 );
not \U$17111 ( \17357 , \14852 );
or \U$17112 ( \17358 , \17356 , \17357 );
nand \U$17113 ( \17359 , \16646 , \16642 );
nand \U$17114 ( \17360 , \17358 , \17359 );
nand \U$17115 ( \17361 , \17354 , \17360 );
nand \U$17116 ( \17362 , \17353 , \17361 );
and \U$17117 ( \17363 , \17338 , \17362 );
and \U$17118 ( \17364 , \17336 , \17337 );
or \U$17119 ( \17365 , \17363 , \17364 );
not \U$17120 ( \17366 , \17365 );
xor \U$17121 ( \17367 , \16015 , \16021 );
xor \U$17122 ( \17368 , \17367 , \16028 );
not \U$17123 ( \17369 , \17368 );
not \U$17124 ( \17370 , \17016 );
nand \U$17125 ( \17371 , \17370 , \17025 );
xnor \U$17126 ( \17372 , \17371 , \17022 );
not \U$17127 ( \17373 , \17372 );
not \U$17128 ( \17374 , \17032 );
and \U$17129 ( \17375 , \17045 , \17374 );
not \U$17130 ( \17376 , \17045 );
and \U$17131 ( \17377 , \17376 , \17032 );
nor \U$17132 ( \17378 , \17375 , \17377 );
not \U$17133 ( \17379 , \17378 );
and \U$17134 ( \17380 , \17373 , \17379 );
and \U$17135 ( \17381 , \17372 , \17378 );
nor \U$17136 ( \17382 , \17380 , \17381 );
not \U$17137 ( \17383 , \17382 );
not \U$17138 ( \17384 , \17383 );
or \U$17139 ( \17385 , \17369 , \17384 );
not \U$17140 ( \17386 , \17378 );
nand \U$17141 ( \17387 , \17386 , \17372 );
nand \U$17142 ( \17388 , \17385 , \17387 );
xnor \U$17143 ( \17389 , \17366 , \17388 );
not \U$17144 ( \17390 , \17389 );
or \U$17145 ( \17391 , \17334 , \17390 );
nand \U$17146 ( \17392 , \17388 , \17365 );
nand \U$17147 ( \17393 , \17391 , \17392 );
nand \U$17148 ( \17394 , \17322 , \17393 );
not \U$17149 ( \17395 , \17320 );
not \U$17150 ( \17396 , \17318 );
nand \U$17151 ( \17397 , \17395 , \17396 );
nand \U$17152 ( \17398 , \17394 , \17397 );
xor \U$17153 ( \17399 , \15971 , \15978 );
xnor \U$17154 ( \17400 , \17399 , \15950 );
not \U$17155 ( \17401 , \15998 );
nand \U$17156 ( \17402 , \17401 , \16007 );
and \U$17157 ( \17403 , \17402 , \16004 );
not \U$17158 ( \17404 , \17402 );
and \U$17159 ( \17405 , \17404 , \16005 );
nor \U$17160 ( \17406 , \17403 , \17405 );
nand \U$17161 ( \17407 , \17400 , \17406 );
not \U$17162 ( \17408 , \17407 );
xnor \U$17163 ( \17409 , \16883 , \16905 );
not \U$17164 ( \17410 , \17409 );
or \U$17165 ( \17411 , \17408 , \17410 );
not \U$17166 ( \17412 , \17400 );
not \U$17167 ( \17413 , \17406 );
nand \U$17168 ( \17414 , \17412 , \17413 );
nand \U$17169 ( \17415 , \17411 , \17414 );
xnor \U$17170 ( \17416 , \17274 , \17287 );
and \U$17171 ( \17417 , \17416 , \17281 );
not \U$17172 ( \17418 , \17416 );
and \U$17173 ( \17419 , \17418 , \17280 );
nor \U$17174 ( \17420 , \17417 , \17419 );
xor \U$17175 ( \17421 , \17415 , \17420 );
xor \U$17176 ( \17422 , \17227 , \17232 );
xor \U$17177 ( \17423 , \17422 , \17224 );
and \U$17178 ( \17424 , \17421 , \17423 );
and \U$17179 ( \17425 , \17415 , \17420 );
or \U$17180 ( \17426 , \17424 , \17425 );
not \U$17181 ( \17427 , \17426 );
xor \U$17182 ( \17428 , \16704 , \16719 );
not \U$17183 ( \17429 , \16710 );
xor \U$17184 ( \17430 , \17428 , \17429 );
not \U$17185 ( \17431 , \17430 );
not \U$17186 ( \17432 , \17431 );
xor \U$17187 ( \17433 , \16730 , \16736 );
xnor \U$17188 ( \17434 , \17433 , \16741 );
not \U$17189 ( \17435 , \17434 );
xor \U$17190 ( \17436 , \16657 , \16641 );
xnor \U$17191 ( \17437 , \17436 , \16648 );
not \U$17192 ( \17438 , \17437 );
or \U$17193 ( \17439 , \17435 , \17438 );
or \U$17194 ( \17440 , \17437 , \17434 );
nand \U$17195 ( \17441 , \17439 , \17440 );
not \U$17196 ( \17442 , \17441 );
or \U$17197 ( \17443 , \17432 , \17442 );
not \U$17198 ( \17444 , \17437 );
nand \U$17199 ( \17445 , \17444 , \17434 );
nand \U$17200 ( \17446 , \17443 , \17445 );
not \U$17201 ( \17447 , \17446 );
xor \U$17202 ( \17448 , \16722 , \16776 );
not \U$17203 ( \17449 , \16686 );
not \U$17204 ( \17450 , \16660 );
and \U$17205 ( \17451 , \17449 , \17450 );
and \U$17206 ( \17452 , \16686 , \16660 );
nor \U$17207 ( \17453 , \17451 , \17452 );
xnor \U$17208 ( \17454 , \17448 , \17453 );
not \U$17209 ( \17455 , \17454 );
or \U$17210 ( \17456 , \17447 , \17455 );
not \U$17211 ( \17457 , \17453 );
xor \U$17212 ( \17458 , \16776 , \16722 );
nand \U$17213 ( \17459 , \17457 , \17458 );
nand \U$17214 ( \17460 , \17456 , \17459 );
not \U$17215 ( \17461 , \17460 );
xor \U$17216 ( \17462 , \16034 , \16043 );
not \U$17217 ( \17463 , \17462 );
and \U$17218 ( \17464 , \17461 , \17463 );
not \U$17219 ( \17465 , \17461 );
and \U$17220 ( \17466 , \17465 , \17462 );
nor \U$17221 ( \17467 , \17464 , \17466 );
not \U$17222 ( \17468 , \17467 );
or \U$17223 ( \17469 , \17427 , \17468 );
nand \U$17224 ( \17470 , \17460 , \17462 );
nand \U$17225 ( \17471 , \17469 , \17470 );
xor \U$17226 ( \17472 , \17398 , \17471 );
not \U$17227 ( \17473 , \17472 );
or \U$17228 ( \17474 , \17313 , \17473 );
nand \U$17229 ( \17475 , \17471 , \17398 );
nand \U$17230 ( \17476 , \17474 , \17475 );
xnor \U$17231 ( \17477 , \17310 , \17476 );
not \U$17232 ( \17478 , \17477 );
or \U$17233 ( \17479 , \17179 , \17478 );
not \U$17234 ( \17480 , \17310 );
nand \U$17235 ( \17481 , \17480 , \17476 );
nand \U$17236 ( \17482 , \17479 , \17481 );
not \U$17237 ( \17483 , \17159 );
not \U$17238 ( \17484 , \17173 );
or \U$17239 ( \17485 , \17483 , \17484 );
not \U$17240 ( \17486 , \17163 );
nand \U$17241 ( \17487 , \17486 , \17169 );
nand \U$17242 ( \17488 , \17485 , \17487 );
not \U$17243 ( \17489 , \15761 );
not \U$17244 ( \17490 , \16080 );
not \U$17245 ( \17491 , \17490 );
or \U$17246 ( \17492 , \17489 , \17491 );
not \U$17247 ( \17493 , \15761 );
nand \U$17248 ( \17494 , \17493 , \16080 );
nand \U$17249 ( \17495 , \17492 , \17494 );
xor \U$17250 ( \17496 , \17488 , \17495 );
xor \U$17251 ( \17497 , \16325 , \16231 );
xor \U$17252 ( \17498 , \17497 , \16207 );
not \U$17253 ( \17499 , \17206 );
not \U$17254 ( \17500 , \17214 );
or \U$17255 ( \17501 , \17499 , \17500 );
not \U$17256 ( \17502 , \17206 );
not \U$17257 ( \17503 , \17502 );
not \U$17258 ( \17504 , \17213 );
or \U$17259 ( \17505 , \17503 , \17504 );
nand \U$17260 ( \17506 , \17505 , \17308 );
nand \U$17261 ( \17507 , \17501 , \17506 );
and \U$17262 ( \17508 , \17498 , \17507 );
not \U$17263 ( \17509 , \17498 );
not \U$17264 ( \17510 , \17507 );
and \U$17265 ( \17511 , \17509 , \17510 );
nor \U$17266 ( \17512 , \17508 , \17511 );
xor \U$17267 ( \17513 , \17496 , \17512 );
xnor \U$17268 ( \17514 , \17482 , \17513 );
xor \U$17269 ( \17515 , \17178 , \17477 );
not \U$17270 ( \17516 , \17515 );
xor \U$17271 ( \17517 , \17415 , \17420 );
xor \U$17272 ( \17518 , \17517 , \17423 );
not \U$17273 ( \17519 , \17518 );
and \U$17274 ( \17520 , RIbe2aeb0_111, RIbe27b98_2);
xor \U$17275 ( \17521 , RIbe27d78_6, RIbe2a640_93);
not \U$17276 ( \17522 , \17521 );
not \U$17277 ( \17523 , \8898 );
or \U$17278 ( \17524 , \17522 , \17523 );
nand \U$17279 ( \17525 , \10752 , \17127 );
nand \U$17280 ( \17526 , \17524 , \17525 );
xor \U$17281 ( \17527 , \17520 , \17526 );
xor \U$17282 ( \17528 , RIbe2b108_116, RIbe284f8_22);
not \U$17283 ( \17529 , \17528 );
not \U$17284 ( \17530 , \13540 );
not \U$17285 ( \17531 , \17530 );
or \U$17286 ( \17532 , \17529 , \17531 );
nand \U$17287 ( \17533 , \16875 , \16893 );
nand \U$17288 ( \17534 , \17532 , \17533 );
xnor \U$17289 ( \17535 , \17527 , \17534 );
not \U$17290 ( \17536 , \17535 );
not \U$17291 ( \17537 , \17536 );
xor \U$17292 ( \17538 , RIbe27fd0_11, RIbe28d68_40);
not \U$17293 ( \17539 , \17538 );
not \U$17294 ( \17540 , \10466 );
or \U$17295 ( \17541 , \17539 , \17540 );
nand \U$17296 ( \17542 , \7709 , \17114 );
nand \U$17297 ( \17543 , \17541 , \17542 );
xor \U$17298 ( \17544 , RIbe28de0_41, RIbe2a730_95);
not \U$17299 ( \17545 , \17544 );
not \U$17300 ( \17546 , \331 );
or \U$17301 ( \17547 , \17545 , \17546 );
nand \U$17302 ( \17548 , \346 , \16789 );
nand \U$17303 ( \17549 , \17547 , \17548 );
xor \U$17304 ( \17550 , \17543 , \17549 );
xor \U$17305 ( \17551 , RIbe280c0_13, RIbe2b2e8_120);
not \U$17306 ( \17552 , \17551 );
not \U$17307 ( \17553 , \10542 );
or \U$17308 ( \17554 , \17552 , \17553 );
nand \U$17309 ( \17555 , \2369 , \17090 );
nand \U$17310 ( \17556 , \17554 , \17555 );
xor \U$17311 ( \17557 , \17550 , \17556 );
not \U$17312 ( \17558 , \17557 );
or \U$17313 ( \17559 , \17537 , \17558 );
or \U$17314 ( \17560 , \17557 , \17536 );
xor \U$17315 ( \17561 , RIbe29308_52, RIbe2a190_83);
not \U$17316 ( \17562 , \17561 );
not \U$17317 ( \17563 , \10689 );
not \U$17318 ( \17564 , \17563 );
or \U$17319 ( \17565 , \17562 , \17564 );
nand \U$17320 ( \17566 , \13278 , \17096 );
nand \U$17321 ( \17567 , \17565 , \17566 );
xor \U$17322 ( \17568 , RIbe28048_12, RIbe2b018_114);
not \U$17323 ( \17569 , \17568 );
not \U$17324 ( \17570 , \15965 );
buf \U$17325 ( \17571 , \17570 );
not \U$17326 ( \17572 , \17571 );
or \U$17327 ( \17573 , \17569 , \17572 );
nand \U$17328 ( \17574 , \15953 , \16809 );
nand \U$17329 ( \17575 , \17573 , \17574 );
xor \U$17330 ( \17576 , \17567 , \17575 );
xor \U$17331 ( \17577 , RIbe2a280_85, RIbe28c78_38);
not \U$17332 ( \17578 , \17577 );
not \U$17333 ( \17579 , \14383 );
or \U$17334 ( \17580 , \17578 , \17579 );
xor \U$17335 ( \17581 , RIbe2a280_85, RIbe28318_18);
nand \U$17336 ( \17582 , \11348 , \17581 );
nand \U$17337 ( \17583 , \17580 , \17582 );
xor \U$17338 ( \17584 , \17576 , \17583 );
nand \U$17339 ( \17585 , \17560 , \17584 );
nand \U$17340 ( \17586 , \17559 , \17585 );
not \U$17341 ( \17587 , \17586 );
not \U$17342 ( \17588 , \17587 );
xor \U$17343 ( \17589 , RIbe28840_29, RIbe2b180_117);
not \U$17344 ( \17590 , \17589 );
nand \U$17345 ( \17591 , \14848 , \14849 );
not \U$17346 ( \17592 , \17591 );
not \U$17347 ( \17593 , \17592 );
or \U$17348 ( \17594 , \17590 , \17593 );
nand \U$17349 ( \17595 , \16646 , \17355 );
nand \U$17350 ( \17596 , \17594 , \17595 );
xor \U$17351 ( \17597 , RIbe29a10_67, RIbe29c68_72);
not \U$17352 ( \17598 , \17597 );
not \U$17353 ( \17599 , \14971 );
or \U$17354 ( \17600 , \17598 , \17599 );
nand \U$17355 ( \17601 , \4580 , \16839 );
nand \U$17356 ( \17602 , \17600 , \17601 );
or \U$17357 ( \17603 , \17596 , \17602 );
xor \U$17358 ( \17604 , RIbe28480_21, RIbe29ce0_73);
not \U$17359 ( \17605 , \17604 );
not \U$17360 ( \17606 , \2518 );
or \U$17361 ( \17607 , \17605 , \17606 );
nand \U$17362 ( \17608 , \3074 , \16950 );
nand \U$17363 ( \17609 , \17607 , \17608 );
nand \U$17364 ( \17610 , \17603 , \17609 );
nand \U$17365 ( \17611 , \17596 , \17602 );
nand \U$17366 ( \17612 , \17610 , \17611 );
not \U$17367 ( \17613 , \17612 );
not \U$17368 ( \17614 , \17613 );
not \U$17369 ( \17615 , \17520 );
not \U$17370 ( \17616 , \17534 );
or \U$17371 ( \17617 , \17615 , \17616 );
or \U$17372 ( \17618 , \17534 , \17520 );
nand \U$17373 ( \17619 , \17618 , \17526 );
nand \U$17374 ( \17620 , \17617 , \17619 );
not \U$17375 ( \17621 , \17620 );
or \U$17376 ( \17622 , \17614 , \17621 );
or \U$17377 ( \17623 , \17620 , \17613 );
nand \U$17378 ( \17624 , \17622 , \17623 );
not \U$17379 ( \17625 , \17624 );
xor \U$17380 ( \17626 , \17567 , \17575 );
and \U$17381 ( \17627 , \17626 , \17583 );
and \U$17382 ( \17628 , \17567 , \17575 );
or \U$17383 ( \17629 , \17627 , \17628 );
not \U$17384 ( \17630 , \17629 );
not \U$17385 ( \17631 , \17630 );
and \U$17386 ( \17632 , \17625 , \17631 );
and \U$17387 ( \17633 , \17624 , \17630 );
nor \U$17388 ( \17634 , \17632 , \17633 );
not \U$17389 ( \17635 , \17634 );
or \U$17390 ( \17636 , \17588 , \17635 );
not \U$17391 ( \17637 , \13250 );
not \U$17392 ( \17638 , \17103 );
or \U$17393 ( \17639 , \17637 , \17638 );
not \U$17394 ( \17640 , \11938 );
xor \U$17395 ( \17641 , RIbe28b88_36, RIbe2b6a8_128);
nand \U$17396 ( \17642 , \17640 , \17641 );
nand \U$17397 ( \17643 , \17639 , \17642 );
xor \U$17398 ( \17644 , RIbe2a028_80, RIbe295d8_58);
not \U$17399 ( \17645 , \17644 );
not \U$17400 ( \17646 , \8401 );
or \U$17401 ( \17647 , \17645 , \17646 );
nand \U$17402 ( \17648 , \8930 , \16796 );
nand \U$17403 ( \17649 , \17647 , \17648 );
nor \U$17404 ( \17650 , \17643 , \17649 );
xor \U$17405 ( \17651 , RIbe29e48_76, RIbe29128_48);
not \U$17406 ( \17652 , \17651 );
not \U$17407 ( \17653 , \7372 );
or \U$17408 ( \17654 , \17652 , \17653 );
nand \U$17409 ( \17655 , \8245 , \16846 );
nand \U$17410 ( \17656 , \17654 , \17655 );
not \U$17411 ( \17657 , \17656 );
or \U$17412 ( \17658 , \17650 , \17657 );
nand \U$17413 ( \17659 , \17643 , \17649 );
nand \U$17414 ( \17660 , \17658 , \17659 );
not \U$17415 ( \17661 , \17660 );
not \U$17416 ( \17662 , \17661 );
xor \U$17417 ( \17663 , RIbe28f48_44, RIbe27df0_7);
not \U$17418 ( \17664 , \17663 );
not \U$17419 ( \17665 , \8221 );
or \U$17420 ( \17666 , \17664 , \17665 );
nand \U$17421 ( \17667 , \11201 , \17346 );
nand \U$17422 ( \17668 , \17666 , \17667 );
not \U$17423 ( \17669 , \17668 );
xor \U$17424 ( \17670 , RIbe296c8_60, RIbe2a460_89);
not \U$17425 ( \17671 , \17670 );
not \U$17426 ( \17672 , \10812 );
or \U$17427 ( \17673 , \17671 , \17672 );
nand \U$17428 ( \17674 , \907 , \17067 );
nand \U$17429 ( \17675 , \17673 , \17674 );
not \U$17430 ( \17676 , \17675 );
not \U$17431 ( \17677 , \17676 );
xor \U$17432 ( \17678 , RIbe2b4c8_124, RIbe290b0_47);
not \U$17433 ( \17679 , \17678 );
not \U$17434 ( \17680 , \2730 );
or \U$17435 ( \17681 , \17679 , \17680 );
nand \U$17436 ( \17682 , \399 , \16823 );
nand \U$17437 ( \17683 , \17681 , \17682 );
not \U$17438 ( \17684 , \17683 );
or \U$17439 ( \17685 , \17677 , \17684 );
or \U$17440 ( \17686 , \17676 , \17683 );
nand \U$17441 ( \17687 , \17685 , \17686 );
not \U$17442 ( \17688 , \17687 );
or \U$17443 ( \17689 , \17669 , \17688 );
nand \U$17444 ( \17690 , \17675 , \17683 );
nand \U$17445 ( \17691 , \17689 , \17690 );
xor \U$17446 ( \17692 , \17543 , \17549 );
and \U$17447 ( \17693 , \17692 , \17556 );
and \U$17448 ( \17694 , \17543 , \17549 );
or \U$17449 ( \17695 , \17693 , \17694 );
xor \U$17450 ( \17696 , \17691 , \17695 );
not \U$17451 ( \17697 , \17696 );
or \U$17452 ( \17698 , \17662 , \17697 );
or \U$17453 ( \17699 , \17661 , \17696 );
nand \U$17454 ( \17700 , \17698 , \17699 );
nand \U$17455 ( \17701 , \17636 , \17700 );
not \U$17456 ( \17702 , \17634 );
nand \U$17457 ( \17703 , \17702 , \17586 );
nand \U$17458 ( \17704 , \17701 , \17703 );
not \U$17459 ( \17705 , \17704 );
not \U$17460 ( \17706 , \17705 );
xor \U$17461 ( \17707 , RIbe293f8_54, RIbe2a190_83);
not \U$17462 ( \17708 , \17707 );
not \U$17463 ( \17709 , \14730 );
or \U$17464 ( \17710 , \17708 , \17709 );
nand \U$17465 ( \17711 , \10696 , \17561 );
nand \U$17466 ( \17712 , \17710 , \17711 );
not \U$17467 ( \17713 , \17712 );
not \U$17468 ( \17714 , \17713 );
xor \U$17469 ( \17715 , RIbe28138_14, RIbe2a3e8_88);
not \U$17470 ( \17716 , \17715 );
not \U$17471 ( \17717 , \8806 );
or \U$17472 ( \17718 , \17716 , \17717 );
xnor \U$17473 ( \17719 , RIbe282a0_17, RIbe2a3e8_88);
not \U$17474 ( \17720 , \17719 );
nand \U$17475 ( \17721 , \17720 , \9268 );
nand \U$17476 ( \17722 , \17718 , \17721 );
not \U$17477 ( \17723 , \17722 );
not \U$17478 ( \17724 , \17723 );
or \U$17479 ( \17725 , \17714 , \17724 );
xor \U$17480 ( \17726 , RIbe29740_61, RIbe2a2f8_86);
not \U$17481 ( \17727 , \17726 );
not \U$17482 ( \17728 , \10792 );
or \U$17483 ( \17729 , \17727 , \17728 );
xor \U$17484 ( \17730 , RIbe297b8_62, RIbe2a2f8_86);
nand \U$17485 ( \17731 , \8706 , \17730 );
nand \U$17486 ( \17732 , \17729 , \17731 );
nand \U$17487 ( \17733 , \17725 , \17732 );
not \U$17488 ( \17734 , \17723 );
nand \U$17489 ( \17735 , \17734 , \17712 );
nand \U$17490 ( \17736 , \17733 , \17735 );
xor \U$17491 ( \17737 , RIbe28930_31, RIbe2a118_82);
not \U$17492 ( \17738 , \17737 );
not \U$17493 ( \17739 , \3064 );
or \U$17494 ( \17740 , \17738 , \17739 );
xor \U$17495 ( \17741 , RIbe28930_31, RIbe2a820_97);
nand \U$17496 ( \17742 , \1199 , \17741 );
nand \U$17497 ( \17743 , \17740 , \17742 );
not \U$17498 ( \17744 , \17743 );
xor \U$17499 ( \17745 , RIbe27d78_6, RIbe2ac58_106);
not \U$17500 ( \17746 , \17745 );
not \U$17501 ( \17747 , \1043 );
or \U$17502 ( \17748 , \17746 , \17747 );
nand \U$17503 ( \17749 , \314 , \17521 );
nand \U$17504 ( \17750 , \17748 , \17749 );
not \U$17505 ( \17751 , \17750 );
not \U$17506 ( \17752 , \17751 );
xor \U$17507 ( \17753 , RIbe28cf0_39, RIbe27e68_8);
not \U$17508 ( \17754 , \17753 );
not \U$17509 ( \17755 , \2599 );
or \U$17510 ( \17756 , \17754 , \17755 );
xor \U$17511 ( \17757 , RIbe298a8_64, RIbe27e68_8);
nand \U$17512 ( \17758 , \2464 , \17757 );
nand \U$17513 ( \17759 , \17756 , \17758 );
not \U$17514 ( \17760 , \17759 );
or \U$17515 ( \17761 , \17752 , \17760 );
or \U$17516 ( \17762 , \17759 , \17751 );
nand \U$17517 ( \17763 , \17761 , \17762 );
not \U$17518 ( \17764 , \17763 );
or \U$17519 ( \17765 , \17744 , \17764 );
nand \U$17520 ( \17766 , \17759 , \17750 );
nand \U$17521 ( \17767 , \17765 , \17766 );
xor \U$17522 ( \17768 , \17736 , \17767 );
xor \U$17523 ( \17769 , RIbe29470_55, RIbe2a910_99);
not \U$17524 ( \17770 , \17769 );
not \U$17525 ( \17771 , \15395 );
or \U$17526 ( \17772 , \17770 , \17771 );
xor \U$17527 ( \17773 , RIbe294e8_56, RIbe2a910_99);
nand \U$17528 ( \17774 , \10401 , \17773 );
nand \U$17529 ( \17775 , \17772 , \17774 );
not \U$17530 ( \17776 , \17775 );
xor \U$17531 ( \17777 , RIbe2a4d8_90, RIbe280c0_13);
not \U$17532 ( \17778 , \17777 );
not \U$17533 ( \17779 , \2379 );
or \U$17534 ( \17780 , \17778 , \17779 );
nand \U$17535 ( \17781 , \869 , \17551 );
nand \U$17536 ( \17782 , \17780 , \17781 );
xor \U$17537 ( \17783 , RIbe2a898_98, RIbe28a20_33);
not \U$17538 ( \17784 , \17783 );
not \U$17539 ( \17785 , \1780 );
or \U$17540 ( \17786 , \17784 , \17785 );
xor \U$17541 ( \17787 , RIbe2aa00_101, RIbe28a20_33);
nand \U$17542 ( \17788 , \2475 , \17787 );
nand \U$17543 ( \17789 , \17786 , \17788 );
xor \U$17544 ( \17790 , \17782 , \17789 );
not \U$17545 ( \17791 , \17790 );
or \U$17546 ( \17792 , \17776 , \17791 );
nand \U$17547 ( \17793 , \17789 , \17782 );
nand \U$17548 ( \17794 , \17792 , \17793 );
and \U$17549 ( \17795 , \17768 , \17794 );
and \U$17550 ( \17796 , \17736 , \17767 );
or \U$17551 ( \17797 , \17795 , \17796 );
not \U$17552 ( \17798 , \17797 );
not \U$17553 ( \17799 , \17581 );
not \U$17554 ( \17800 , \14942 );
or \U$17555 ( \17801 , \17799 , \17800 );
nand \U$17556 ( \17802 , \11348 , \17034 );
nand \U$17557 ( \17803 , \17801 , \17802 );
xnor \U$17558 ( \17804 , \16900 , \17803 );
xor \U$17559 ( \17805 , RIbe286d8_26, RIbe2af28_112);
not \U$17560 ( \17806 , \17805 );
not \U$17561 ( \17807 , \15345 );
or \U$17562 ( \17808 , \17806 , \17807 );
not \U$17563 ( \17809 , \14412 );
buf \U$17564 ( \17810 , \17809 );
buf \U$17565 ( \17811 , \17810 );
nand \U$17566 ( \17812 , \17811 , \16911 );
nand \U$17567 ( \17813 , \17808 , \17812 );
not \U$17568 ( \17814 , \17813 );
xor \U$17569 ( \17815 , \17804 , \17814 );
not \U$17570 ( \17816 , \17815 );
xor \U$17571 ( \17817 , RIbe28b88_36, RIbe2aa78_102);
not \U$17572 ( \17818 , \17817 );
not \U$17573 ( \17819 , \8711 );
or \U$17574 ( \17820 , \17818 , \17819 );
nand \U$17575 ( \17821 , \13250 , \17641 );
nand \U$17576 ( \17822 , \17820 , \17821 );
not \U$17577 ( \17823 , \17822 );
xor \U$17578 ( \17824 , RIbe28570_23, RIbe2af28_112);
not \U$17579 ( \17825 , \17824 );
not \U$17580 ( \17826 , \16913 );
or \U$17581 ( \17827 , \17825 , \17826 );
nand \U$17582 ( \17828 , \17810 , \17805 );
nand \U$17583 ( \17829 , \17827 , \17828 );
not \U$17584 ( \17830 , \17829 );
or \U$17585 ( \17831 , \17823 , \17830 );
or \U$17586 ( \17832 , \17822 , \17829 );
xor \U$17587 ( \17833 , RIbe28f48_44, RIbe27c88_4);
not \U$17588 ( \17834 , \17833 );
not \U$17589 ( \17835 , \7609 );
or \U$17590 ( \17836 , \17834 , \17835 );
nand \U$17591 ( \17837 , \11201 , \17663 );
nand \U$17592 ( \17838 , \17836 , \17837 );
nand \U$17593 ( \17839 , \17832 , \17838 );
nand \U$17594 ( \17840 , \17831 , \17839 );
not \U$17595 ( \17841 , \17840 );
xor \U$17596 ( \17842 , RIbe29c68_72, RIbe29218_50);
not \U$17597 ( \17843 , \17842 );
not \U$17598 ( \17844 , \10720 );
or \U$17599 ( \17845 , \17843 , \17844 );
nand \U$17600 ( \17846 , \4580 , \17597 );
nand \U$17601 ( \17847 , \17845 , \17846 );
not \U$17602 ( \17848 , \17847 );
xor \U$17603 ( \17849 , RIbe2a280_85, RIbe28c00_37);
not \U$17604 ( \17850 , \17849 );
not \U$17605 ( \17851 , \11345 );
or \U$17606 ( \17852 , \17850 , \17851 );
nand \U$17607 ( \17853 , \14649 , \17577 );
nand \U$17608 ( \17854 , \17852 , \17853 );
not \U$17609 ( \17855 , \17854 );
or \U$17610 ( \17856 , \17848 , \17855 );
or \U$17611 ( \17857 , \17854 , \17847 );
xor \U$17612 ( \17858 , RIbe29f38_78, RIbe28390_19);
not \U$17613 ( \17859 , \17858 );
not \U$17614 ( \17860 , \14579 );
or \U$17615 ( \17861 , \17859 , \17860 );
xor \U$17616 ( \17862 , RIbe28390_19, RIbe29ec0_77);
nand \U$17617 ( \17863 , \5831 , \17862 );
nand \U$17618 ( \17864 , \17861 , \17863 );
nand \U$17619 ( \17865 , \17857 , \17864 );
nand \U$17620 ( \17866 , \17856 , \17865 );
not \U$17621 ( \17867 , \17866 );
or \U$17622 ( \17868 , \17841 , \17867 );
or \U$17623 ( \17869 , \17866 , \17840 );
xor \U$17624 ( \17870 , RIbe29d58_74, RIbe28480_21);
not \U$17625 ( \17871 , \17870 );
not \U$17626 ( \17872 , \2518 );
or \U$17627 ( \17873 , \17871 , \17872 );
nand \U$17628 ( \17874 , \16676 , \17604 );
nand \U$17629 ( \17875 , \17873 , \17874 );
not \U$17630 ( \17876 , \17875 );
nand \U$17631 ( \17877 , RIbe27b98_2, RIbe2ae38_110);
not \U$17632 ( \17878 , \17877 );
and \U$17633 ( \17879 , \17876 , \17878 );
and \U$17634 ( \17880 , \17875 , \17877 );
nor \U$17635 ( \17881 , \17879 , \17880 );
not \U$17636 ( \17882 , \17881 );
not \U$17637 ( \17883 , \17882 );
xor \U$17638 ( \17884 , RIbe2b450_123, RIbe28de0_41);
not \U$17639 ( \17885 , \17884 );
not \U$17640 ( \17886 , \332 );
or \U$17641 ( \17887 , \17885 , \17886 );
nand \U$17642 ( \17888 , \514 , \17544 );
nand \U$17643 ( \17889 , \17887 , \17888 );
not \U$17644 ( \17890 , \17889 );
or \U$17645 ( \17891 , \17883 , \17890 );
not \U$17646 ( \17892 , \17877 );
nand \U$17647 ( \17893 , \17892 , \17875 );
nand \U$17648 ( \17894 , \17891 , \17893 );
nand \U$17649 ( \17895 , \17869 , \17894 );
nand \U$17650 ( \17896 , \17868 , \17895 );
not \U$17651 ( \17897 , \17896 );
or \U$17652 ( \17898 , \17816 , \17897 );
or \U$17653 ( \17899 , \17896 , \17815 );
nand \U$17654 ( \17900 , \17898 , \17899 );
not \U$17655 ( \17901 , \17900 );
or \U$17656 ( \17902 , \17798 , \17901 );
not \U$17657 ( \17903 , \17815 );
nand \U$17658 ( \17904 , \17903 , \17896 );
nand \U$17659 ( \17905 , \17902 , \17904 );
not \U$17660 ( \17906 , \17905 );
not \U$17661 ( \17907 , \17906 );
or \U$17662 ( \17908 , \17706 , \17907 );
not \U$17663 ( \17909 , \17660 );
not \U$17664 ( \17910 , \17696 );
or \U$17665 ( \17911 , \17909 , \17910 );
nand \U$17666 ( \17912 , \17691 , \17695 );
nand \U$17667 ( \17913 , \17911 , \17912 );
not \U$17668 ( \17914 , \17913 );
not \U$17669 ( \17915 , \17914 );
not \U$17670 ( \17916 , \17813 );
not \U$17671 ( \17917 , \17804 );
or \U$17672 ( \17918 , \17916 , \17917 );
nand \U$17673 ( \17919 , \16901 , \17803 );
nand \U$17674 ( \17920 , \17918 , \17919 );
not \U$17675 ( \17921 , \17920 );
xor \U$17676 ( \17922 , RIbe2abe0_105, RIbe27c10_3);
not \U$17677 ( \17923 , \17922 );
not \U$17678 ( \17924 , \11907 );
or \U$17679 ( \17925 , \17923 , \17924 );
nand \U$17680 ( \17926 , \369 , \16978 );
nand \U$17681 ( \17927 , \17925 , \17926 );
not \U$17682 ( \17928 , \17757 );
not \U$17683 ( \17929 , \2599 );
or \U$17684 ( \17930 , \17928 , \17929 );
nand \U$17685 ( \17931 , \2463 , \17339 );
nand \U$17686 ( \17932 , \17930 , \17931 );
or \U$17687 ( \17933 , \17927 , \17932 );
xor \U$17688 ( \17934 , RIbe29038_46, RIbe2ad48_108);
not \U$17689 ( \17935 , \17934 );
not \U$17690 ( \17936 , \281 );
or \U$17691 ( \17937 , \17935 , \17936 );
nand \U$17692 ( \17938 , \1583 , \16852 );
nand \U$17693 ( \17939 , \17937 , \17938 );
nand \U$17694 ( \17940 , \17933 , \17939 );
nand \U$17695 ( \17941 , \17932 , \17927 );
nand \U$17696 ( \17942 , \17940 , \17941 );
not \U$17697 ( \17943 , \17942 );
not \U$17698 ( \17944 , \17943 );
not \U$17699 ( \17945 , \17741 );
not \U$17700 ( \17946 , \8887 );
or \U$17701 ( \17947 , \17945 , \17946 );
nand \U$17702 ( \17948 , \1797 , \16958 );
nand \U$17703 ( \17949 , \17947 , \17948 );
not \U$17704 ( \17950 , \17949 );
not \U$17705 ( \17951 , \17950 );
not \U$17706 ( \17952 , \17773 );
not \U$17707 ( \17953 , \9737 );
or \U$17708 ( \17954 , \17952 , \17953 );
nand \U$17709 ( \17955 , \9726 , \17075 );
nand \U$17710 ( \17956 , \17954 , \17955 );
not \U$17711 ( \17957 , \17956 );
or \U$17712 ( \17958 , \17951 , \17957 );
or \U$17713 ( \17959 , \17956 , \17950 );
nand \U$17714 ( \17960 , \17958 , \17959 );
xor \U$17715 ( \17961 , RIbe28a98_34, RIbe2a550_91);
not \U$17716 ( \17962 , \17961 );
not \U$17717 ( \17963 , \10434 );
or \U$17718 ( \17964 , \17962 , \17963 );
nand \U$17719 ( \17965 , \12004 , \16921 );
nand \U$17720 ( \17966 , \17964 , \17965 );
nand \U$17721 ( \17967 , \17960 , \17966 );
nand \U$17722 ( \17968 , \17956 , \17949 );
nand \U$17723 ( \17969 , \17967 , \17968 );
not \U$17724 ( \17970 , \17969 );
not \U$17725 ( \17971 , \17970 );
or \U$17726 ( \17972 , \17944 , \17971 );
xor \U$17727 ( \17973 , RIbe27b20_1, RIbe285e8_24);
not \U$17728 ( \17974 , \17973 );
not \U$17729 ( \17975 , \8813 );
or \U$17730 ( \17976 , \17974 , \17975 );
nand \U$17731 ( \17977 , \2625 , \16970 );
nand \U$17732 ( \17978 , \17976 , \17977 );
not \U$17733 ( \17979 , \17862 );
not \U$17734 ( \17980 , \14806 );
or \U$17735 ( \17981 , \17979 , \17980 );
nand \U$17736 ( \17982 , \2777 , \16943 );
nand \U$17737 ( \17983 , \17981 , \17982 );
nor \U$17738 ( \17984 , \17978 , \17983 );
xor \U$17739 ( \17985 , RIbe2a0a0_81, RIbe28228_16);
and \U$17740 ( \17986 , \879 , \17985 );
and \U$17741 ( \17987 , \885 , \16928 );
nor \U$17742 ( \17988 , \17986 , \17987 );
or \U$17743 ( \17989 , \17984 , \17988 );
nand \U$17744 ( \17990 , \17978 , \17983 );
nand \U$17745 ( \17991 , \17989 , \17990 );
nand \U$17746 ( \17992 , \17972 , \17991 );
nand \U$17747 ( \17993 , \17942 , \17969 );
nand \U$17748 ( \17994 , \17992 , \17993 );
not \U$17749 ( \17995 , \17994 );
not \U$17750 ( \17996 , \17995 );
or \U$17751 ( \17997 , \17921 , \17996 );
not \U$17752 ( \17998 , \17993 );
not \U$17753 ( \17999 , \17992 );
or \U$17754 ( \18000 , \17998 , \17999 );
not \U$17755 ( \18001 , \17920 );
nand \U$17756 ( \18002 , \18000 , \18001 );
nand \U$17757 ( \18003 , \17997 , \18002 );
not \U$17758 ( \18004 , \18003 );
or \U$17759 ( \18005 , \17915 , \18004 );
or \U$17760 ( \18006 , \18003 , \17914 );
nand \U$17761 ( \18007 , \18005 , \18006 );
nand \U$17762 ( \18008 , \17908 , \18007 );
nand \U$17763 ( \18009 , \17905 , \17704 );
nand \U$17764 ( \18010 , \18008 , \18009 );
not \U$17765 ( \18011 , \18010 );
not \U$17766 ( \18012 , \18011 );
or \U$17767 ( \18013 , \17519 , \18012 );
or \U$17768 ( \18014 , \18011 , \17518 );
nand \U$17769 ( \18015 , \18013 , \18014 );
not \U$17770 ( \18016 , \18015 );
xor \U$17771 ( \18017 , \17360 , \17344 );
xnor \U$17772 ( \18018 , \18017 , \17351 );
not \U$17773 ( \18019 , \18018 );
not \U$17774 ( \18020 , \18019 );
xor \U$17775 ( \18021 , \17064 , \17084 );
not \U$17776 ( \18022 , \18021 );
xor \U$17777 ( \18023 , \16802 , \16787 );
not \U$17778 ( \18024 , \18023 );
or \U$17779 ( \18025 , \18022 , \18024 );
or \U$17780 ( \18026 , \18023 , \18021 );
nand \U$17781 ( \18027 , \18025 , \18026 );
not \U$17782 ( \18028 , \18027 );
or \U$17783 ( \18029 , \18020 , \18028 );
not \U$17784 ( \18030 , \18021 );
nand \U$17785 ( \18031 , \18030 , \18023 );
nand \U$17786 ( \18032 , \18029 , \18031 );
not \U$17787 ( \18033 , \18032 );
xor \U$17788 ( \18034 , \16969 , \16976 );
xor \U$17789 ( \18035 , \18034 , \16983 );
or \U$17790 ( \18036 , \17095 , \17101 );
nand \U$17791 ( \18037 , \18036 , \17111 );
xnor \U$17792 ( \18038 , \18037 , \17109 );
xor \U$17793 ( \18039 , \18035 , \18038 );
xor \U$17794 ( \18040 , \16919 , \16936 );
and \U$17795 ( \18041 , \18039 , \18040 );
and \U$17796 ( \18042 , \18035 , \18038 );
or \U$17797 ( \18043 , \18041 , \18042 );
not \U$17798 ( \18044 , \18043 );
not \U$17799 ( \18045 , \16869 );
not \U$17800 ( \18046 , \16807 );
not \U$17801 ( \18047 , \18046 );
and \U$17802 ( \18048 , \18045 , \18047 );
and \U$17803 ( \18049 , \16869 , \18046 );
nor \U$17804 ( \18050 , \18048 , \18049 );
not \U$17805 ( \18051 , \18050 );
or \U$17806 ( \18052 , \18044 , \18051 );
or \U$17807 ( \18053 , \18050 , \18043 );
nand \U$17808 ( \18054 , \18052 , \18053 );
not \U$17809 ( \18055 , \18054 );
or \U$17810 ( \18056 , \18033 , \18055 );
not \U$17811 ( \18057 , \18050 );
nand \U$17812 ( \18058 , \18057 , \18043 );
nand \U$17813 ( \18059 , \18056 , \18058 );
not \U$17814 ( \18060 , \18059 );
not \U$17815 ( \18061 , \18060 );
not \U$17816 ( \18062 , \17913 );
not \U$17817 ( \18063 , \18003 );
or \U$17818 ( \18064 , \18062 , \18063 );
not \U$17819 ( \18065 , \17993 );
not \U$17820 ( \18066 , \17992 );
or \U$17821 ( \18067 , \18065 , \18066 );
nand \U$17822 ( \18068 , \18067 , \17920 );
nand \U$17823 ( \18069 , \18064 , \18068 );
not \U$17824 ( \18070 , \18069 );
not \U$17825 ( \18071 , \17629 );
not \U$17826 ( \18072 , \17624 );
or \U$17827 ( \18073 , \18071 , \18072 );
nand \U$17828 ( \18074 , \17620 , \17612 );
nand \U$17829 ( \18075 , \18073 , \18074 );
not \U$17830 ( \18076 , \18075 );
not \U$17831 ( \18077 , \18076 );
not \U$17832 ( \18078 , \16941 );
not \U$17833 ( \18079 , \18078 );
not \U$17834 ( \18080 , \16987 );
and \U$17835 ( \18081 , \18079 , \18080 );
and \U$17836 ( \18082 , \16987 , \18078 );
nor \U$17837 ( \18083 , \18081 , \18082 );
not \U$17838 ( \18084 , \18083 );
or \U$17839 ( \18085 , \18077 , \18084 );
xor \U$17840 ( \18086 , \17088 , \17140 );
nand \U$17841 ( \18087 , \18085 , \18086 );
not \U$17842 ( \18088 , \18076 );
not \U$17843 ( \18089 , \18083 );
nand \U$17844 ( \18090 , \18088 , \18089 );
nand \U$17845 ( \18091 , \18087 , \18090 );
not \U$17846 ( \18092 , \18091 );
and \U$17847 ( \18093 , \18070 , \18092 );
not \U$17848 ( \18094 , \18070 );
and \U$17849 ( \18095 , \18094 , \18091 );
nor \U$17850 ( \18096 , \18093 , \18095 );
not \U$17851 ( \18097 , \18096 );
or \U$17852 ( \18098 , \18061 , \18097 );
or \U$17853 ( \18099 , \18060 , \18096 );
nand \U$17854 ( \18100 , \18098 , \18099 );
not \U$17855 ( \18101 , \18100 );
or \U$17856 ( \18102 , \18016 , \18101 );
not \U$17857 ( \18103 , \18011 );
nand \U$17858 ( \18104 , \18103 , \17518 );
nand \U$17859 ( \18105 , \18102 , \18104 );
not \U$17860 ( \18106 , \18105 );
not \U$17861 ( \18107 , \17318 );
not \U$17862 ( \18108 , \17320 );
or \U$17863 ( \18109 , \18107 , \18108 );
nand \U$17864 ( \18110 , \18109 , \17397 );
and \U$17865 ( \18111 , \18110 , \17393 );
not \U$17866 ( \18112 , \18110 );
not \U$17867 ( \18113 , \17393 );
and \U$17868 ( \18114 , \18112 , \18113 );
nor \U$17869 ( \18115 , \18111 , \18114 );
not \U$17870 ( \18116 , \18115 );
not \U$17871 ( \18117 , \18116 );
or \U$17872 ( \18118 , \18106 , \18117 );
and \U$17873 ( \18119 , \18105 , \18115 );
not \U$17874 ( \18120 , \18105 );
and \U$17875 ( \18121 , \18120 , \18116 );
nor \U$17876 ( \18122 , \18119 , \18121 );
not \U$17877 ( \18123 , \18122 );
xor \U$17878 ( \18124 , \17182 , \17181 );
xor \U$17879 ( \18125 , \18124 , \17185 );
not \U$17880 ( \18126 , \18059 );
not \U$17881 ( \18127 , \18096 );
or \U$17882 ( \18128 , \18126 , \18127 );
not \U$17883 ( \18129 , \18070 );
nand \U$17884 ( \18130 , \18129 , \18091 );
nand \U$17885 ( \18131 , \18128 , \18130 );
not \U$17886 ( \18132 , \18131 );
xor \U$17887 ( \18133 , \18125 , \18132 );
xor \U$17888 ( \18134 , \17366 , \17333 );
xnor \U$17889 ( \18135 , \18134 , \17388 );
not \U$17890 ( \18136 , \18135 );
xnor \U$17891 ( \18137 , \17454 , \17446 );
not \U$17892 ( \18138 , \18137 );
xor \U$17893 ( \18139 , \17057 , \17145 );
xor \U$17894 ( \18140 , \18139 , \17055 );
not \U$17895 ( \18141 , \18140 );
xor \U$17896 ( \18142 , \18138 , \18141 );
not \U$17897 ( \18143 , \18142 );
or \U$17898 ( \18144 , \18136 , \18143 );
not \U$17899 ( \18145 , \18140 );
and \U$17900 ( \18146 , \18138 , \18145 );
not \U$17901 ( \18147 , \18146 );
nand \U$17902 ( \18148 , \18144 , \18147 );
xnor \U$17903 ( \18149 , \18133 , \18148 );
nand \U$17904 ( \18150 , \18123 , \18149 );
nand \U$17905 ( \18151 , \18118 , \18150 );
not \U$17906 ( \18152 , \18148 );
not \U$17907 ( \18153 , \18125 );
not \U$17908 ( \18154 , \18153 );
not \U$17909 ( \18155 , \18131 );
or \U$17910 ( \18156 , \18154 , \18155 );
or \U$17911 ( \18157 , \18131 , \18153 );
nand \U$17912 ( \18158 , \18156 , \18157 );
not \U$17913 ( \18159 , \18158 );
or \U$17914 ( \18160 , \18152 , \18159 );
nand \U$17915 ( \18161 , \18131 , \18125 );
nand \U$17916 ( \18162 , \18160 , \18161 );
not \U$17917 ( \18163 , \18162 );
not \U$17918 ( \18164 , \17311 );
not \U$17919 ( \18165 , \17472 );
or \U$17920 ( \18166 , \18164 , \18165 );
or \U$17921 ( \18167 , \17472 , \17311 );
nand \U$17922 ( \18168 , \18166 , \18167 );
not \U$17923 ( \18169 , \18168 );
nand \U$17924 ( \18170 , \18163 , \18169 );
and \U$17925 ( \18171 , \18151 , \18170 );
nand \U$17926 ( \18172 , \18168 , \18162 );
not \U$17927 ( \18173 , \18172 );
nor \U$17928 ( \18174 , \18171 , \18173 );
xor \U$17929 ( \18175 , \16634 , \17154 );
not \U$17930 ( \18176 , \18175 );
xor \U$17931 ( \18177 , \17188 , \17195 );
xor \U$17932 ( \18178 , \18177 , \17203 );
not \U$17933 ( \18179 , \18178 );
not \U$17934 ( \18180 , \18179 );
not \U$17935 ( \18181 , \9268 );
not \U$17936 ( \18182 , \17061 );
or \U$17937 ( \18183 , \18181 , \18182 );
not \U$17938 ( \18184 , \17719 );
nand \U$17939 ( \18185 , \18184 , \9096 );
nand \U$17940 ( \18186 , \18183 , \18185 );
not \U$17941 ( \18187 , \18186 );
not \U$17942 ( \18188 , \8380 );
xor \U$17943 ( \18189 , RIbe2b3d8_122, RIbe27b98_2);
not \U$17944 ( \18190 , \18189 );
or \U$17945 ( \18191 , \18188 , \18190 );
nand \U$17946 ( \18192 , \7585 , \16818 );
nand \U$17947 ( \18193 , \18191 , \18192 );
not \U$17948 ( \18194 , \18193 );
or \U$17949 ( \18195 , \18187 , \18194 );
or \U$17950 ( \18196 , \18193 , \18186 );
not \U$17951 ( \18197 , \17730 );
not \U$17952 ( \18198 , \9375 );
or \U$17953 ( \18199 , \18197 , \18198 );
nand \U$17954 ( \18200 , \8706 , \16782 );
nand \U$17955 ( \18201 , \18199 , \18200 );
nand \U$17956 ( \18202 , \18196 , \18201 );
nand \U$17957 ( \18203 , \18195 , \18202 );
and \U$17958 ( \18204 , \16832 , \16816 );
not \U$17959 ( \18205 , \16832 );
not \U$17960 ( \18206 , \16816 );
and \U$17961 ( \18207 , \18205 , \18206 );
nor \U$17962 ( \18208 , \18204 , \18207 );
xor \U$17963 ( \18209 , \18203 , \18208 );
and \U$17964 ( \18210 , \16860 , \16844 );
not \U$17965 ( \18211 , \16860 );
not \U$17966 ( \18212 , \16844 );
and \U$17967 ( \18213 , \18211 , \18212 );
nor \U$17968 ( \18214 , \18210 , \18213 );
and \U$17969 ( \18215 , \18209 , \18214 );
and \U$17970 ( \18216 , \18203 , \18208 );
or \U$17971 ( \18217 , \18215 , \18216 );
xor \U$17972 ( \18218 , \17336 , \17337 );
xor \U$17973 ( \18219 , \18218 , \17362 );
xor \U$17974 ( \18220 , \18217 , \18219 );
not \U$17975 ( \18221 , \17430 );
not \U$17976 ( \18222 , \17441 );
or \U$17977 ( \18223 , \18221 , \18222 );
or \U$17978 ( \18224 , \17441 , \17430 );
nand \U$17979 ( \18225 , \18223 , \18224 );
and \U$17980 ( \18226 , \18220 , \18225 );
and \U$17981 ( \18227 , \18217 , \18219 );
or \U$17982 ( \18228 , \18226 , \18227 );
not \U$17983 ( \18229 , \18228 );
xnor \U$17984 ( \18230 , \16997 , \16873 );
nand \U$17985 ( \18231 , \18229 , \18230 );
not \U$17986 ( \18232 , \18231 );
nand \U$17987 ( \18233 , \17407 , \17414 );
not \U$17988 ( \18234 , \17409 );
and \U$17989 ( \18235 , \18233 , \18234 );
not \U$17990 ( \18236 , \18233 );
and \U$17991 ( \18237 , \18236 , \17409 );
nor \U$17992 ( \18238 , \18235 , \18237 );
not \U$17993 ( \18239 , \18238 );
xor \U$17994 ( \18240 , \17368 , \17382 );
and \U$17995 ( \18241 , \16964 , \16948 );
not \U$17996 ( \18242 , \16964 );
not \U$17997 ( \18243 , \16948 );
and \U$17998 ( \18244 , \18242 , \18243 );
nor \U$17999 ( \18245 , \18241 , \18244 );
xor \U$18000 ( \18246 , \17132 , \17119 );
xor \U$18001 ( \18247 , \18246 , \17125 );
xor \U$18002 ( \18248 , \18245 , \18247 );
not \U$18003 ( \18249 , \17814 );
not \U$18004 ( \18250 , \17787 );
not \U$18005 ( \18251 , \7795 );
or \U$18006 ( \18252 , \18250 , \18251 );
nand \U$18007 ( \18253 , \2475 , \17120 );
nand \U$18008 ( \18254 , \18252 , \18253 );
and \U$18009 ( \18255 , \18254 , RIbe2aaf0_103);
not \U$18010 ( \18256 , \18254 );
not \U$18011 ( \18257 , RIbe2aaf0_103);
and \U$18012 ( \18258 , \18256 , \18257 );
or \U$18013 ( \18259 , \18255 , \18258 );
not \U$18014 ( \18260 , \18259 );
or \U$18015 ( \18261 , \18249 , \18260 );
nand \U$18016 ( \18262 , \18254 , \18257 );
nand \U$18017 ( \18263 , \18261 , \18262 );
and \U$18018 ( \18264 , \18248 , \18263 );
and \U$18019 ( \18265 , \18245 , \18247 );
or \U$18020 ( \18266 , \18264 , \18265 );
xnor \U$18021 ( \18267 , \18240 , \18266 );
not \U$18022 ( \18268 , \18267 );
or \U$18023 ( \18269 , \18239 , \18268 );
xor \U$18024 ( \18270 , \17368 , \17383 );
nand \U$18025 ( \18271 , \18270 , \18266 );
nand \U$18026 ( \18272 , \18269 , \18271 );
not \U$18027 ( \18273 , \18272 );
or \U$18028 ( \18274 , \18232 , \18273 );
not \U$18029 ( \18275 , \18230 );
nand \U$18030 ( \18276 , \18275 , \18228 );
nand \U$18031 ( \18277 , \18274 , \18276 );
xor \U$18032 ( \18278 , \17462 , \17461 );
xnor \U$18033 ( \18279 , \18278 , \17426 );
xor \U$18034 ( \18280 , \18277 , \18279 );
xor \U$18035 ( \18281 , \16781 , \17001 );
xnor \U$18036 ( \18282 , \18281 , \17150 );
and \U$18037 ( \18283 , \18280 , \18282 );
and \U$18038 ( \18284 , \18277 , \18279 );
or \U$18039 ( \18285 , \18283 , \18284 );
not \U$18040 ( \18286 , \18285 );
or \U$18041 ( \18287 , \18180 , \18286 );
or \U$18042 ( \18288 , \18285 , \18179 );
nand \U$18043 ( \18289 , \18287 , \18288 );
not \U$18044 ( \18290 , \18289 );
or \U$18045 ( \18291 , \18176 , \18290 );
nand \U$18046 ( \18292 , \18285 , \18178 );
nand \U$18047 ( \18293 , \18291 , \18292 );
not \U$18048 ( \18294 , \18293 );
and \U$18049 ( \18295 , \18174 , \18294 );
not \U$18050 ( \18296 , \18174 );
and \U$18051 ( \18297 , \18296 , \18293 );
nor \U$18052 ( \18298 , \18295 , \18297 );
not \U$18053 ( \18299 , \18298 );
or \U$18054 ( \18300 , \17516 , \18299 );
not \U$18055 ( \18301 , \18174 );
nand \U$18056 ( \18302 , \18301 , \18293 );
nand \U$18057 ( \18303 , \18300 , \18302 );
not \U$18058 ( \18304 , \18303 );
nor \U$18059 ( \18305 , \17514 , \18304 );
not \U$18060 ( \18306 , \18305 );
not \U$18061 ( \18307 , \16498 );
not \U$18062 ( \18308 , \16488 );
and \U$18063 ( \18309 , \18307 , \18308 );
and \U$18064 ( \18310 , \16498 , \16488 );
nor \U$18065 ( \18311 , \18309 , \18310 );
and \U$18066 ( \18312 , \16400 , \16084 );
not \U$18067 ( \18313 , \16400 );
not \U$18068 ( \18314 , \16084 );
and \U$18069 ( \18315 , \18313 , \18314 );
nor \U$18070 ( \18316 , \18312 , \18315 );
xor \U$18071 ( \18317 , \18311 , \18316 );
not \U$18072 ( \18318 , \17495 );
not \U$18073 ( \18319 , \17512 );
or \U$18074 ( \18320 , \18318 , \18319 );
not \U$18075 ( \18321 , \17510 );
nand \U$18076 ( \18322 , \18321 , \17498 );
nand \U$18077 ( \18323 , \18320 , \18322 );
xnor \U$18078 ( \18324 , \18317 , \18323 );
not \U$18079 ( \18325 , \18324 );
nand \U$18080 ( \18326 , \17513 , \17482 );
xor \U$18081 ( \18327 , \17512 , \17495 );
nand \U$18082 ( \18328 , \18327 , \17488 );
nand \U$18083 ( \18329 , \18325 , \18326 , \18328 );
not \U$18084 ( \18330 , \18329 );
or \U$18085 ( \18331 , \18306 , \18330 );
not \U$18086 ( \18332 , \16503 );
not \U$18087 ( \18333 , \16509 );
or \U$18088 ( \18334 , \18332 , \18333 );
or \U$18089 ( \18335 , \16509 , \16503 );
nand \U$18090 ( \18336 , \18334 , \18335 );
not \U$18091 ( \18337 , \18316 );
not \U$18092 ( \18338 , \18311 );
not \U$18093 ( \18339 , \18323 );
or \U$18094 ( \18340 , \18338 , \18339 );
or \U$18095 ( \18341 , \18323 , \18311 );
nand \U$18096 ( \18342 , \18340 , \18341 );
not \U$18097 ( \18343 , \18342 );
or \U$18098 ( \18344 , \18337 , \18343 );
not \U$18099 ( \18345 , \18311 );
nand \U$18100 ( \18346 , \18345 , \18323 );
nand \U$18101 ( \18347 , \18344 , \18346 );
nand \U$18102 ( \18348 , \18336 , \18347 );
not \U$18103 ( \18349 , \18328 );
not \U$18104 ( \18350 , \18326 );
or \U$18105 ( \18351 , \18349 , \18350 );
nand \U$18106 ( \18352 , \18351 , \18324 );
nand \U$18107 ( \18353 , \18348 , \18352 );
not \U$18108 ( \18354 , \18353 );
nand \U$18109 ( \18355 , \18331 , \18354 );
nor \U$18110 ( \18356 , \18347 , \18336 );
not \U$18111 ( \18357 , \18356 );
nand \U$18112 ( \18358 , \18355 , \18357 );
not \U$18113 ( \18359 , \18358 );
or \U$18114 ( \18360 , \16623 , \18359 );
not \U$18115 ( \18361 , \16608 );
not \U$18116 ( \18362 , \16601 );
or \U$18117 ( \18363 , \18361 , \18362 );
not \U$18118 ( \18364 , \16597 );
nand \U$18119 ( \18365 , \18364 , \16558 );
nand \U$18120 ( \18366 , \18363 , \18365 );
not \U$18121 ( \18367 , \16545 );
or \U$18122 ( \18368 , \18367 , \16552 );
nand \U$18123 ( \18369 , \18368 , \16527 );
nand \U$18124 ( \18370 , \16552 , \18367 );
nand \U$18125 ( \18371 , \18369 , \18370 );
nor \U$18126 ( \18372 , \18366 , \18371 );
not \U$18127 ( \18373 , \18372 );
not \U$18128 ( \18374 , \18371 );
not \U$18129 ( \18375 , \18374 );
nand \U$18130 ( \18376 , \18375 , \18366 );
nand \U$18131 ( \18377 , \18373 , \18376 );
not \U$18132 ( \18378 , \16567 );
not \U$18133 ( \18379 , \18378 );
not \U$18134 ( \18380 , \16577 );
or \U$18135 ( \18381 , \18379 , \18380 );
nand \U$18136 ( \18382 , \16570 , \16576 );
nand \U$18137 ( \18383 , \18381 , \18382 );
xor \U$18138 ( \18384 , \13197 , \13236 );
xor \U$18139 ( \18385 , \18384 , \13486 );
nor \U$18140 ( \18386 , \18383 , \18385 );
not \U$18141 ( \18387 , \18386 );
nand \U$18142 ( \18388 , \18383 , \18385 );
nand \U$18143 ( \18389 , \18387 , \18388 );
not \U$18144 ( \18390 , \18389 );
nand \U$18145 ( \18391 , \16536 , \16534 );
not \U$18146 ( \18392 , \18391 );
not \U$18147 ( \18393 , \16543 );
or \U$18148 ( \18394 , \18392 , \18393 );
or \U$18149 ( \18395 , \16536 , \16534 );
nand \U$18150 ( \18396 , \18394 , \18395 );
not \U$18151 ( \18397 , \18396 );
not \U$18152 ( \18398 , \18397 );
and \U$18153 ( \18399 , \18390 , \18398 );
and \U$18154 ( \18400 , \18389 , \18397 );
nor \U$18155 ( \18401 , \18399 , \18400 );
xor \U$18156 ( \18402 , \13094 , \13172 );
not \U$18157 ( \18403 , \18402 );
xor \U$18158 ( \18404 , \16517 , \16518 );
and \U$18159 ( \18405 , \18404 , \16526 );
and \U$18160 ( \18406 , \16517 , \16518 );
or \U$18161 ( \18407 , \18405 , \18406 );
not \U$18162 ( \18408 , \18407 );
not \U$18163 ( \18409 , \18408 );
or \U$18164 ( \18410 , \18403 , \18409 );
not \U$18165 ( \18411 , \18407 );
or \U$18166 ( \18412 , \18411 , \18402 );
nand \U$18167 ( \18413 , \18410 , \18412 );
not \U$18168 ( \18414 , \13507 );
not \U$18169 ( \18415 , \18414 );
buf \U$18170 ( \18416 , \13677 );
not \U$18171 ( \18417 , \18416 );
or \U$18172 ( \18418 , \18415 , \18417 );
or \U$18173 ( \18419 , \18416 , \18414 );
nand \U$18174 ( \18420 , \18418 , \18419 );
xor \U$18175 ( \18421 , \18413 , \18420 );
xor \U$18176 ( \18422 , \18401 , \18421 );
not \U$18177 ( \18423 , \16592 );
not \U$18178 ( \18424 , \16586 );
or \U$18179 ( \18425 , \18423 , \18424 );
not \U$18180 ( \18426 , \16584 );
nand \U$18181 ( \18427 , \18426 , \16565 );
nand \U$18182 ( \18428 , \18425 , \18427 );
xor \U$18183 ( \18429 , \18422 , \18428 );
not \U$18184 ( \18430 , \18429 );
and \U$18185 ( \18431 , \18377 , \18430 );
not \U$18186 ( \18432 , \18377 );
and \U$18187 ( \18433 , \18432 , \18429 );
nor \U$18188 ( \18434 , \18431 , \18433 );
not \U$18189 ( \18435 , \18434 );
xor \U$18190 ( \18436 , \16553 , \16613 );
and \U$18191 ( \18437 , \18436 , \16619 );
and \U$18192 ( \18438 , \16553 , \16613 );
or \U$18193 ( \18439 , \18437 , \18438 );
nand \U$18194 ( \18440 , \18435 , \18439 );
not \U$18195 ( \18441 , \18440 );
xor \U$18196 ( \18442 , \18401 , \18421 );
and \U$18197 ( \18443 , \18442 , \18428 );
and \U$18198 ( \18444 , \18401 , \18421 );
or \U$18199 ( \18445 , \18443 , \18444 );
not \U$18200 ( \18446 , \18445 );
xor \U$18201 ( \18447 , \13688 , \13505 );
not \U$18202 ( \18448 , \18447 );
not \U$18203 ( \18449 , \18420 );
not \U$18204 ( \18450 , \18413 );
or \U$18205 ( \18451 , \18449 , \18450 );
not \U$18206 ( \18452 , \18411 );
nand \U$18207 ( \18453 , \18452 , \18402 );
nand \U$18208 ( \18454 , \18451 , \18453 );
not \U$18209 ( \18455 , \18454 );
not \U$18210 ( \18456 , \18455 );
or \U$18211 ( \18457 , \18386 , \18397 );
nand \U$18212 ( \18458 , \18457 , \18388 );
not \U$18213 ( \18459 , \18458 );
not \U$18214 ( \18460 , \13495 );
nand \U$18215 ( \18461 , \18460 , \13497 );
and \U$18216 ( \18462 , \18461 , \13176 );
not \U$18217 ( \18463 , \18461 );
and \U$18218 ( \18464 , \18463 , \13177 );
nor \U$18219 ( \18465 , \18462 , \18464 );
not \U$18220 ( \18466 , \18465 );
or \U$18221 ( \18467 , \18459 , \18466 );
or \U$18222 ( \18468 , \18465 , \18458 );
nand \U$18223 ( \18469 , \18467 , \18468 );
not \U$18224 ( \18470 , \18469 );
not \U$18225 ( \18471 , \18470 );
or \U$18226 ( \18472 , \18456 , \18471 );
nand \U$18227 ( \18473 , \18469 , \18454 );
nand \U$18228 ( \18474 , \18472 , \18473 );
not \U$18229 ( \18475 , \18474 );
or \U$18230 ( \18476 , \18448 , \18475 );
or \U$18231 ( \18477 , \18447 , \18474 );
nand \U$18232 ( \18478 , \18476 , \18477 );
not \U$18233 ( \18479 , \18478 );
or \U$18234 ( \18480 , \18446 , \18479 );
or \U$18235 ( \18481 , \18445 , \18478 );
nand \U$18236 ( \18482 , \18480 , \18481 );
not \U$18237 ( \18483 , \18374 );
not \U$18238 ( \18484 , \18366 );
not \U$18239 ( \18485 , \18484 );
or \U$18240 ( \18486 , \18483 , \18485 );
nand \U$18241 ( \18487 , \18486 , \18429 );
buf \U$18242 ( \18488 , \18376 );
and \U$18243 ( \18489 , \18482 , \18487 , \18488 );
nor \U$18244 ( \18490 , \18441 , \18489 );
and \U$18245 ( \18491 , \16510 , \16620 , \16406 );
not \U$18246 ( \18492 , \18491 );
xnor \U$18247 ( \18493 , \12247 , \12196 );
buf \U$18248 ( \18494 , \12187 );
and \U$18249 ( \18495 , \18493 , \18494 );
not \U$18250 ( \18496 , \18493 );
not \U$18251 ( \18497 , \18494 );
and \U$18252 ( \18498 , \18496 , \18497 );
nor \U$18253 ( \18499 , \18495 , \18498 );
xor \U$18254 ( \18500 , \13498 , \13091 );
xor \U$18255 ( \18501 , \18500 , \13693 );
xor \U$18256 ( \18502 , \18499 , \18501 );
not \U$18257 ( \18503 , \18458 );
nand \U$18258 ( \18504 , \18503 , \18465 );
not \U$18259 ( \18505 , \18504 );
not \U$18260 ( \18506 , \18454 );
or \U$18261 ( \18507 , \18505 , \18506 );
not \U$18262 ( \18508 , \18465 );
nand \U$18263 ( \18509 , \18508 , \18458 );
nand \U$18264 ( \18510 , \18507 , \18509 );
not \U$18265 ( \18511 , \18510 );
xor \U$18266 ( \18512 , \18502 , \18511 );
not \U$18267 ( \18513 , \18447 );
not \U$18268 ( \18514 , \18513 );
not \U$18269 ( \18515 , \18474 );
or \U$18270 ( \18516 , \18514 , \18515 );
nand \U$18271 ( \18517 , \18516 , \18445 );
not \U$18272 ( \18518 , \18474 );
nand \U$18273 ( \18519 , \18518 , \18447 );
nand \U$18274 ( \18520 , \18517 , \18519 );
not \U$18275 ( \18521 , \18520 );
nand \U$18276 ( \18522 , \18512 , \18521 );
and \U$18277 ( \18523 , \13088 , \13698 );
not \U$18278 ( \18524 , \13088 );
and \U$18279 ( \18525 , \18524 , \13076 );
nor \U$18280 ( \18526 , \18523 , \18525 );
and \U$18281 ( \18527 , \18526 , \13695 );
not \U$18282 ( \18528 , \18526 );
not \U$18283 ( \18529 , \13694 );
nor \U$18284 ( \18530 , \13091 , \13502 );
nor \U$18285 ( \18531 , \18529 , \18530 );
and \U$18286 ( \18532 , \18528 , \18531 );
nor \U$18287 ( \18533 , \18527 , \18532 );
xor \U$18288 ( \18534 , \18499 , \18501 );
and \U$18289 ( \18535 , \18534 , \18511 );
and \U$18290 ( \18536 , \18499 , \18501 );
or \U$18291 ( \18537 , \18535 , \18536 );
nand \U$18292 ( \18538 , \18533 , \18537 );
and \U$18293 ( \18539 , \18522 , \18538 );
and \U$18294 ( \18540 , \18490 , \18492 , \18539 );
nand \U$18295 ( \18541 , \18360 , \18540 );
not \U$18296 ( \18542 , \18439 );
nand \U$18297 ( \18543 , \18434 , \18542 );
not \U$18298 ( \18544 , \18543 );
and \U$18299 ( \18545 , \18482 , \18487 , \18488 );
not \U$18300 ( \18546 , \18545 );
and \U$18301 ( \18547 , \18544 , \18546 );
and \U$18302 ( \18548 , \18487 , \18488 );
buf \U$18303 ( \18549 , \18482 );
nor \U$18304 ( \18550 , \18548 , \18549 );
nor \U$18305 ( \18551 , \18547 , \18550 );
not \U$18306 ( \18552 , \18512 );
nand \U$18307 ( \18553 , \18552 , \18520 );
nand \U$18308 ( \18554 , \18551 , \18553 );
and \U$18309 ( \18555 , \18554 , \18539 );
nor \U$18310 ( \18556 , \18533 , \18537 );
nor \U$18311 ( \18557 , \18555 , \18556 );
nand \U$18312 ( \18558 , \18541 , \18557 );
not \U$18313 ( \18559 , \13977 );
not \U$18314 ( \18560 , \13072 );
or \U$18315 ( \18561 , \13073 , \13700 );
nand \U$18316 ( \18562 , \18560 , \18561 );
nor \U$18317 ( \18563 , \18559 , \18562 );
and \U$18318 ( \18564 , \18563 , \10395 , \14154 );
and \U$18319 ( \18565 , \18564 , \14231 );
nand \U$18320 ( \18566 , \18558 , \18565 );
nand \U$18321 ( \18567 , \14234 , \18566 );
nand \U$18322 ( \18568 , \7202 , \18567 );
not \U$18323 ( \18569 , \18545 );
and \U$18324 ( \18570 , \18440 , \18569 , \18539 );
buf \U$18325 ( \18571 , \18329 );
nor \U$18326 ( \18572 , \18491 , \18356 );
not \U$18327 ( \18573 , \18303 );
nand \U$18328 ( \18574 , \18573 , \17514 );
and \U$18329 ( \18575 , \18570 , \18571 , \18572 , \18574 );
and \U$18330 ( \18576 , \18575 , \18565 );
xor \U$18331 ( \18577 , RIbe295d8_58, RIbe2a3e8_88);
not \U$18332 ( \18578 , \18577 );
not \U$18333 ( \18579 , \15475 );
or \U$18334 ( \18580 , \18578 , \18579 );
xor \U$18335 ( \18581 , RIbe29740_61, RIbe2a3e8_88);
nand \U$18336 ( \18582 , \11541 , \18581 );
nand \U$18337 ( \18583 , \18580 , \18582 );
not \U$18338 ( \18584 , \18583 );
xor \U$18339 ( \18585 , RIbe294e8_56, RIbe2a190_83);
not \U$18340 ( \18586 , \18585 );
not \U$18341 ( \18587 , \14730 );
or \U$18342 ( \18588 , \18586 , \18587 );
xor \U$18343 ( \18589 , RIbe288b8_30, RIbe2a190_83);
nand \U$18344 ( \18590 , \13278 , \18589 );
nand \U$18345 ( \18591 , \18588 , \18590 );
xor \U$18346 ( \18592 , RIbe28a20_33, RIbe2a0a0_81);
not \U$18347 ( \18593 , \18592 );
not \U$18348 ( \18594 , \7795 );
or \U$18349 ( \18595 , \18593 , \18594 );
xor \U$18350 ( \18596 , RIbe28a20_33, RIbe2a118_82);
nand \U$18351 ( \18597 , \2475 , \18596 );
nand \U$18352 ( \18598 , \18595 , \18597 );
xor \U$18353 ( \18599 , \18591 , \18598 );
not \U$18354 ( \18600 , \18599 );
or \U$18355 ( \18601 , \18584 , \18600 );
nand \U$18356 ( \18602 , \18598 , \18591 );
nand \U$18357 ( \18603 , \18601 , \18602 );
xor \U$18358 ( \18604 , RIbe296c8_60, RIbe2b4c8_124);
not \U$18359 ( \18605 , \18604 );
not \U$18360 ( \18606 , \900 );
or \U$18361 ( \18607 , \18605 , \18606 );
xor \U$18362 ( \18608 , RIbe2b540_125, RIbe296c8_60);
nand \U$18363 ( \18609 , \1939 , \18608 );
nand \U$18364 ( \18610 , \18607 , \18609 );
xor \U$18365 ( \18611 , RIbe28228_16, RIbe2a460_89);
not \U$18366 ( \18612 , \18611 );
not \U$18367 ( \18613 , \879 );
or \U$18368 ( \18614 , \18612 , \18613 );
xor \U$18369 ( \18615 , RIbe2a4d8_90, RIbe28228_16);
nand \U$18370 ( \18616 , \8680 , \18615 );
nand \U$18371 ( \18617 , \18614 , \18616 );
xor \U$18372 ( \18618 , \18610 , \18617 );
xor \U$18373 ( \18619 , RIbe28f48_44, RIbe298a8_64);
not \U$18374 ( \18620 , \18619 );
not \U$18375 ( \18621 , \8221 );
or \U$18376 ( \18622 , \18620 , \18621 );
xor \U$18377 ( \18623 , RIbe29998_66, RIbe28f48_44);
nand \U$18378 ( \18624 , \3249 , \18623 );
nand \U$18379 ( \18625 , \18622 , \18624 );
and \U$18380 ( \18626 , \18618 , \18625 );
and \U$18381 ( \18627 , \18610 , \18617 );
or \U$18382 ( \18628 , \18626 , \18627 );
nor \U$18383 ( \18629 , \18603 , \18628 );
not \U$18384 ( \18630 , \18629 );
nand \U$18385 ( \18631 , \18603 , \18628 );
nand \U$18386 ( \18632 , \18630 , \18631 );
xor \U$18387 ( \18633 , RIbe2a550_91, RIbe282a0_17);
not \U$18388 ( \18634 , \18633 );
buf \U$18389 ( \18635 , \10433 );
not \U$18390 ( \18636 , \18635 );
or \U$18391 ( \18637 , \18634 , \18636 );
xor \U$18392 ( \18638 , RIbe29470_55, RIbe2a550_91);
nand \U$18393 ( \18639 , \14612 , \18638 );
nand \U$18394 ( \18640 , \18637 , \18639 );
xor \U$18395 ( \18641 , RIbe29c68_72, RIbe28d68_40);
not \U$18396 ( \18642 , \18641 );
not \U$18397 ( \18643 , \4578 );
or \U$18398 ( \18644 , \18642 , \18643 );
xor \U$18399 ( \18645 , RIbe27c88_4, RIbe29c68_72);
nand \U$18400 ( \18646 , \4580 , \18645 );
nand \U$18401 ( \18647 , \18644 , \18646 );
xor \U$18402 ( \18648 , \18640 , \18647 );
not \U$18403 ( \18649 , \14424 );
xor \U$18404 ( \18650 , RIbe284f8_22, RIbe2af28_112);
and \U$18405 ( \18651 , \18649 , \18650 );
xor \U$18406 ( \18652 , RIbe2af28_112, RIbe28750_27);
and \U$18407 ( \18653 , \16917 , \18652 );
nor \U$18408 ( \18654 , \18651 , \18653 );
not \U$18409 ( \18655 , \18654 );
and \U$18410 ( \18656 , \18648 , \18655 );
and \U$18411 ( \18657 , \18647 , \18640 );
nor \U$18412 ( \18658 , \18656 , \18657 );
xnor \U$18413 ( \18659 , \18632 , \18658 );
not \U$18414 ( \18660 , \18659 );
not \U$18415 ( \18661 , \18660 );
xor \U$18416 ( \18662 , RIbe28a98_34, RIbe2a280_85);
not \U$18417 ( \18663 , \18662 );
not \U$18418 ( \18664 , \14382 );
or \U$18419 ( \18665 , \18663 , \18664 );
not \U$18420 ( \18666 , \10847 );
not \U$18421 ( \18667 , \18666 );
xor \U$18422 ( \18668 , RIbe2a280_85, RIbe293f8_54);
nand \U$18423 ( \18669 , \18667 , \18668 );
nand \U$18424 ( \18670 , \18665 , \18669 );
not \U$18425 ( \18671 , \18670 );
xor \U$18426 ( \18672 , RIbe2b108_116, RIbe29308_52);
not \U$18427 ( \18673 , \18672 );
not \U$18428 ( \18674 , \17530 );
or \U$18429 ( \18675 , \18673 , \18674 );
xor \U$18430 ( \18676 , RIbe2b108_116, RIbe28c00_37);
nand \U$18431 ( \18677 , \16898 , \18676 );
nand \U$18432 ( \18678 , \18675 , \18677 );
not \U$18433 ( \18679 , \18678 );
or \U$18434 ( \18680 , \18671 , \18679 );
or \U$18435 ( \18681 , \18678 , \18670 );
xor \U$18436 ( \18682 , RIbe27df0_7, RIbe29e48_76);
not \U$18437 ( \18683 , \18682 );
not \U$18438 ( \18684 , \7716 );
or \U$18439 ( \18685 , \18683 , \18684 );
xor \U$18440 ( \18686 , RIbe29e48_76, RIbe29218_50);
nand \U$18441 ( \18687 , \8245 , \18686 );
nand \U$18442 ( \18688 , \18685 , \18687 );
nand \U$18443 ( \18689 , \18681 , \18688 );
nand \U$18444 ( \18690 , \18680 , \18689 );
xor \U$18445 ( \18691 , RIbe29038_46, RIbe2a640_93);
not \U$18446 ( \18692 , \18691 );
not \U$18447 ( \18693 , \16854 );
or \U$18448 ( \18694 , \18692 , \18693 );
xor \U$18449 ( \18695 , RIbe29038_46, RIbe2a6b8_94);
nand \U$18450 ( \18696 , \286 , \18695 );
nand \U$18451 ( \18697 , \18694 , \18696 );
not \U$18452 ( \18698 , \18697 );
xor \U$18453 ( \18699 , RIbe27e68_8, RIbe29ce0_73);
not \U$18454 ( \18700 , \18699 );
not \U$18455 ( \18701 , \2600 );
or \U$18456 ( \18702 , \18700 , \18701 );
xor \U$18457 ( \18703 , RIbe27e68_8, RIbe29b78_70);
nand \U$18458 ( \18704 , \2603 , \18703 );
nand \U$18459 ( \18705 , \18702 , \18704 );
not \U$18460 ( \18706 , \18705 );
or \U$18461 ( \18707 , \18698 , \18706 );
or \U$18462 ( \18708 , \18697 , \18705 );
xor \U$18463 ( \18709 , RIbe28390_19, RIbe2aa00_101);
not \U$18464 ( \18710 , \18709 );
not \U$18465 ( \18711 , \14806 );
or \U$18466 ( \18712 , \18710 , \18711 );
xor \U$18467 ( \18713 , RIbe2aa78_102, RIbe28390_19);
nand \U$18468 ( \18714 , \3714 , \18713 );
nand \U$18469 ( \18715 , \18712 , \18714 );
nand \U$18470 ( \18716 , \18708 , \18715 );
nand \U$18471 ( \18717 , \18707 , \18716 );
xor \U$18472 ( \18718 , \18690 , \18717 );
xor \U$18473 ( \18719 , RIbe28930_31, RIbe2b2e8_120);
not \U$18474 ( \18720 , \18719 );
not \U$18475 ( \18721 , \965 );
or \U$18476 ( \18722 , \18720 , \18721 );
xor \U$18477 ( \18723 , RIbe28930_31, RIbe2b360_121);
nand \U$18478 ( \18724 , \970 , \18723 );
nand \U$18479 ( \18725 , \18722 , \18724 );
not \U$18480 ( \18726 , \18725 );
xor \U$18481 ( \18727 , RIbe2b180_117, RIbe28c78_38);
not \U$18482 ( \18728 , \18727 );
not \U$18483 ( \18729 , \14852 );
or \U$18484 ( \18730 , \18728 , \18729 );
xor \U$18485 ( \18731 , RIbe2b180_117, RIbe28318_18);
nand \U$18486 ( \18732 , \14966 , \18731 );
nand \U$18487 ( \18733 , \18730 , \18732 );
not \U$18488 ( \18734 , \18733 );
or \U$18489 ( \18735 , \18726 , \18734 );
or \U$18490 ( \18736 , \18733 , \18725 );
not \U$18491 ( \18737 , \16676 );
xor \U$18492 ( \18738 , RIbe29f38_78, RIbe28480_21);
not \U$18493 ( \18739 , \18738 );
or \U$18494 ( \18740 , \18737 , \18739 );
xnor \U$18495 ( \18741 , RIbe28480_21, RIbe2b6a8_128);
not \U$18496 ( \18742 , \18741 );
nand \U$18497 ( \18743 , \18742 , \2518 );
nand \U$18498 ( \18744 , \18740 , \18743 );
nand \U$18499 ( \18745 , \18736 , \18744 );
nand \U$18500 ( \18746 , \18735 , \18745 );
xor \U$18501 ( \18747 , \18718 , \18746 );
and \U$18502 ( \18748 , \18648 , \18655 );
not \U$18503 ( \18749 , \18648 );
and \U$18504 ( \18750 , \18749 , \18654 );
nor \U$18505 ( \18751 , \18748 , \18750 );
not \U$18506 ( \18752 , \18751 );
not \U$18507 ( \18753 , \18697 );
not \U$18508 ( \18754 , \18715 );
not \U$18509 ( \18755 , \18754 );
or \U$18510 ( \18756 , \18753 , \18755 );
or \U$18511 ( \18757 , \18697 , \18754 );
nand \U$18512 ( \18758 , \18756 , \18757 );
not \U$18513 ( \18759 , \18705 );
and \U$18514 ( \18760 , \18758 , \18759 );
not \U$18515 ( \18761 , \18758 );
and \U$18516 ( \18762 , \18761 , \18705 );
nor \U$18517 ( \18763 , \18760 , \18762 );
not \U$18518 ( \18764 , \18763 );
xor \U$18519 ( \18765 , RIbe28de0_41, RIbe2ae38_110);
not \U$18520 ( \18766 , \18765 );
not \U$18521 ( \18767 , \11321 );
or \U$18522 ( \18768 , \18766 , \18767 );
xor \U$18523 ( \18769 , RIbe28de0_41, RIbe2aeb0_111);
nand \U$18524 ( \18770 , \346 , \18769 );
nand \U$18525 ( \18771 , \18768 , \18770 );
not \U$18526 ( \18772 , \18771 );
xor \U$18527 ( \18773 , RIbe28840_29, RIbe2b018_114);
not \U$18528 ( \18774 , \18773 );
not \U$18529 ( \18775 , \17570 );
or \U$18530 ( \18776 , \18774 , \18775 );
buf \U$18531 ( \18777 , \15952 );
xor \U$18532 ( \18778 , RIbe28570_23, RIbe2b018_114);
nand \U$18533 ( \18779 , \18777 , \18778 );
nand \U$18534 ( \18780 , \18776 , \18779 );
not \U$18535 ( \18781 , \18780 );
not \U$18536 ( \18782 , \18781 );
or \U$18537 ( \18783 , \18772 , \18782 );
not \U$18538 ( \18784 , \18771 );
nand \U$18539 ( \18785 , \18780 , \18784 );
nand \U$18540 ( \18786 , \18783 , \18785 );
xor \U$18541 ( \18787 , RIbe290b0_47, RIbe2abe0_105);
not \U$18542 ( \18788 , \18787 );
not \U$18543 ( \18789 , \2730 );
or \U$18544 ( \18790 , \18788 , \18789 );
xor \U$18545 ( \18791 , RIbe290b0_47, RIbe2ac58_106);
nand \U$18546 ( \18792 , \398 , \18791 );
nand \U$18547 ( \18793 , \18790 , \18792 );
and \U$18548 ( \18794 , \18786 , \18793 );
not \U$18549 ( \18795 , \18786 );
not \U$18550 ( \18796 , \18793 );
and \U$18551 ( \18797 , \18795 , \18796 );
nor \U$18552 ( \18798 , \18794 , \18797 );
not \U$18553 ( \18799 , \18798 );
or \U$18554 ( \18800 , \18764 , \18799 );
or \U$18555 ( \18801 , \18798 , \18763 );
nand \U$18556 ( \18802 , \18800 , \18801 );
not \U$18557 ( \18803 , \18802 );
or \U$18558 ( \18804 , \18752 , \18803 );
not \U$18559 ( \18805 , \18763 );
nand \U$18560 ( \18806 , \18805 , \18798 );
nand \U$18561 ( \18807 , \18804 , \18806 );
xor \U$18562 ( \18808 , \18747 , \18807 );
not \U$18563 ( \18809 , \18808 );
or \U$18564 ( \18810 , \18661 , \18809 );
nand \U$18565 ( \18811 , \18807 , \18747 );
nand \U$18566 ( \18812 , \18810 , \18811 );
not \U$18567 ( \18813 , \18812 );
not \U$18568 ( \18814 , \18784 );
not \U$18569 ( \18815 , \18781 );
or \U$18570 ( \18816 , \18814 , \18815 );
nand \U$18571 ( \18817 , \18816 , \18793 );
nand \U$18572 ( \18818 , \18780 , \18771 );
nand \U$18573 ( \18819 , \18817 , \18818 );
xor \U$18574 ( \18820 , RIbe27b20_1, RIbe27fd0_11);
not \U$18575 ( \18821 , \18820 );
not \U$18576 ( \18822 , \10466 );
or \U$18577 ( \18823 , \18821 , \18822 );
xor \U$18578 ( \18824 , RIbe27fd0_11, RIbe28cf0_39);
nand \U$18579 ( \18825 , \2707 , \18824 );
nand \U$18580 ( \18826 , \18823 , \18825 );
not \U$18581 ( \18827 , \18826 );
xor \U$18582 ( \18828 , RIbe286d8_26, RIbe2aaf0_103);
not \U$18583 ( \18829 , \18828 );
not \U$18584 ( \18830 , RIbe2ab68_104);
nand \U$18585 ( \18831 , \18830 , RIbe2aaf0_103);
not \U$18586 ( \18832 , \18831 );
not \U$18587 ( \18833 , \18832 );
or \U$18588 ( \18834 , \18829 , \18833 );
xor \U$18589 ( \18835 , RIbe27ee0_9, RIbe2aaf0_103);
nand \U$18590 ( \18836 , \18835 , RIbe2ab68_104);
nand \U$18591 ( \18837 , \18834 , \18836 );
xor \U$18592 ( \18838 , RIbe29128_48, RIbe2a2f8_86);
not \U$18593 ( \18839 , \18838 );
not \U$18594 ( \18840 , \14826 );
or \U$18595 ( \18841 , \18839 , \18840 );
xor \U$18596 ( \18842 , RIbe291a0_49, RIbe2a2f8_86);
nand \U$18597 ( \18843 , \8705 , \18842 );
nand \U$18598 ( \18844 , \18841 , \18843 );
xor \U$18599 ( \18845 , \18837 , \18844 );
not \U$18600 ( \18846 , \18845 );
or \U$18601 ( \18847 , \18827 , \18846 );
nand \U$18602 ( \18848 , \18837 , \18844 );
nand \U$18603 ( \18849 , \18847 , \18848 );
xor \U$18604 ( \18850 , \18819 , \18849 );
xor \U$18605 ( \18851 , RIbe285e8_24, RIbe29ec0_77);
not \U$18606 ( \18852 , \18851 );
not \U$18607 ( \18853 , \8813 );
or \U$18608 ( \18854 , \18852 , \18853 );
xor \U$18609 ( \18855 , RIbe285e8_24, RIbe29d58_74);
nand \U$18610 ( \18856 , \2625 , \18855 );
nand \U$18611 ( \18857 , \18854 , \18856 );
xor \U$18612 ( \18858 , RIbe280c0_13, RIbe2ad48_108);
not \U$18613 ( \18859 , \18858 );
not \U$18614 ( \18860 , \10542 );
or \U$18615 ( \18861 , \18859 , \18860 );
xor \U$18616 ( \18862 , RIbe280c0_13, RIbe2adc0_109);
nand \U$18617 ( \18863 , \2369 , \18862 );
nand \U$18618 ( \18864 , \18861 , \18863 );
xor \U$18619 ( \18865 , \18857 , \18864 );
xor \U$18620 ( \18866 , RIbe2a028_80, RIbe29a10_67);
not \U$18621 ( \18867 , \18866 );
not \U$18622 ( \18868 , \8169 );
or \U$18623 ( \18869 , \18867 , \18868 );
xor \U$18624 ( \18870 , RIbe2a028_80, RIbe29b00_69);
nand \U$18625 ( \18871 , \8172 , \18870 );
nand \U$18626 ( \18872 , \18869 , \18871 );
and \U$18627 ( \18873 , \18865 , \18872 );
and \U$18628 ( \18874 , \18857 , \18864 );
or \U$18629 ( \18875 , \18873 , \18874 );
and \U$18630 ( \18876 , \18850 , \18875 );
and \U$18631 ( \18877 , \18819 , \18849 );
or \U$18632 ( \18878 , \18876 , \18877 );
xor \U$18633 ( \18879 , \18690 , \18717 );
and \U$18634 ( \18880 , \18879 , \18746 );
and \U$18635 ( \18881 , \18690 , \18717 );
or \U$18636 ( \18882 , \18880 , \18881 );
xor \U$18637 ( \18883 , \18878 , \18882 );
or \U$18638 ( \18884 , \18629 , \18658 );
nand \U$18639 ( \18885 , \18884 , \18631 );
xor \U$18640 ( \18886 , \18883 , \18885 );
not \U$18641 ( \18887 , \18886 );
xor \U$18642 ( \18888 , \18819 , \18849 );
xor \U$18643 ( \18889 , \18888 , \18875 );
not \U$18644 ( \18890 , \18889 );
not \U$18645 ( \18891 , \18826 );
and \U$18646 ( \18892 , \18845 , \18891 );
not \U$18647 ( \18893 , \18845 );
and \U$18648 ( \18894 , \18893 , \18826 );
nor \U$18649 ( \18895 , \18892 , \18894 );
not \U$18650 ( \18896 , \18895 );
xor \U$18651 ( \18897 , \18857 , \18864 );
xor \U$18652 ( \18898 , \18897 , \18872 );
not \U$18653 ( \18899 , \18898 );
or \U$18654 ( \18900 , \18896 , \18899 );
or \U$18655 ( \18901 , \18898 , \18895 );
nand \U$18656 ( \18902 , \18900 , \18901 );
not \U$18657 ( \18903 , \18902 );
xor \U$18658 ( \18904 , \18599 , \18583 );
not \U$18659 ( \18905 , \18904 );
or \U$18660 ( \18906 , \18903 , \18905 );
not \U$18661 ( \18907 , \18895 );
nand \U$18662 ( \18908 , \18907 , \18898 );
nand \U$18663 ( \18909 , \18906 , \18908 );
not \U$18664 ( \18910 , \18909 );
or \U$18665 ( \18911 , \18890 , \18910 );
or \U$18666 ( \18912 , \18909 , \18889 );
xor \U$18667 ( \18913 , \18744 , \18725 );
xnor \U$18668 ( \18914 , \18913 , \18733 );
not \U$18669 ( \18915 , \18914 );
not \U$18670 ( \18916 , \18915 );
xor \U$18671 ( \18917 , RIbe2af28_112, RIbe28318_18);
not \U$18672 ( \18918 , \18917 );
not \U$18673 ( \18919 , \16913 );
or \U$18674 ( \18920 , \18918 , \18919 );
nand \U$18675 ( \18921 , \16728 , \18650 );
nand \U$18676 ( \18922 , \18920 , \18921 );
not \U$18677 ( \18923 , \18922 );
xor \U$18678 ( \18924 , RIbe27fd0_11, RIbe29b78_70);
not \U$18679 ( \18925 , \18924 );
not \U$18680 ( \18926 , \9082 );
or \U$18681 ( \18927 , \18925 , \18926 );
nand \U$18682 ( \18928 , \2707 , \18820 );
nand \U$18683 ( \18929 , \18927 , \18928 );
not \U$18684 ( \18930 , \18929 );
or \U$18685 ( \18931 , \18923 , \18930 );
or \U$18686 ( \18932 , \18922 , \18929 );
xor \U$18687 ( \18933 , RIbe280c0_13, RIbe2b540_125);
not \U$18688 ( \18934 , \18933 );
not \U$18689 ( \18935 , \1053 );
or \U$18690 ( \18936 , \18934 , \18935 );
nand \U$18691 ( \18937 , \1263 , \18858 );
nand \U$18692 ( \18938 , \18936 , \18937 );
nand \U$18693 ( \18939 , \18932 , \18938 );
nand \U$18694 ( \18940 , \18931 , \18939 );
not \U$18695 ( \18941 , \18940 );
xor \U$18696 ( \18942 , RIbe285e8_24, RIbe29f38_78);
not \U$18697 ( \18943 , \18942 );
not \U$18698 ( \18944 , \7618 );
or \U$18699 ( \18945 , \18943 , \18944 );
nand \U$18700 ( \18946 , \8270 , \18851 );
nand \U$18701 ( \18947 , \18945 , \18946 );
not \U$18702 ( \18948 , \18947 );
xor \U$18703 ( \18949 , RIbe28570_23, RIbe2aaf0_103);
not \U$18704 ( \18950 , \18949 );
not \U$18705 ( \18951 , \18832 );
or \U$18706 ( \18952 , \18950 , \18951 );
nand \U$18707 ( \18953 , \18828 , RIbe2ab68_104);
nand \U$18708 ( \18954 , \18952 , \18953 );
xor \U$18709 ( \18955 , RIbe29b00_69, RIbe2a2f8_86);
not \U$18710 ( \18956 , \18955 );
not \U$18711 ( \18957 , \14826 );
or \U$18712 ( \18958 , \18956 , \18957 );
not \U$18713 ( \18959 , RIbe2a370_87);
not \U$18714 ( \18960 , RIbe2a3e8_88);
and \U$18715 ( \18961 , \18959 , \18960 );
and \U$18716 ( \18962 , RIbe2a370_87, RIbe2a3e8_88);
nor \U$18717 ( \18963 , \18961 , \18962 );
nand \U$18718 ( \18964 , \18963 , \18838 );
nand \U$18719 ( \18965 , \18958 , \18964 );
xor \U$18720 ( \18966 , \18954 , \18965 );
not \U$18721 ( \18967 , \18966 );
or \U$18722 ( \18968 , \18948 , \18967 );
nand \U$18723 ( \18969 , \18965 , \18954 );
nand \U$18724 ( \18970 , \18968 , \18969 );
not \U$18725 ( \18971 , \18970 );
not \U$18726 ( \18972 , \18971 );
or \U$18727 ( \18973 , \18941 , \18972 );
or \U$18728 ( \18974 , \18940 , \18971 );
nand \U$18729 ( \18975 , \18973 , \18974 );
not \U$18730 ( \18976 , \18975 );
or \U$18731 ( \18977 , \18916 , \18976 );
nand \U$18732 ( \18978 , \18970 , \18940 );
nand \U$18733 ( \18979 , \18977 , \18978 );
nand \U$18734 ( \18980 , \18912 , \18979 );
nand \U$18735 ( \18981 , \18911 , \18980 );
not \U$18736 ( \18982 , \18981 );
nand \U$18737 ( \18983 , \18887 , \18982 );
not \U$18738 ( \18984 , \18983 );
or \U$18739 ( \18985 , \18813 , \18984 );
nand \U$18740 ( \18986 , \18981 , \18886 );
nand \U$18741 ( \18987 , \18985 , \18986 );
not \U$18742 ( \18988 , \18987 );
xor \U$18743 ( \18989 , RIbe27c10_3, RIbe2aeb0_111);
not \U$18744 ( \18990 , \18989 );
not \U$18745 ( \18991 , \7440 );
or \U$18746 ( \18992 , \18990 , \18991 );
xor \U$18747 ( \18993 , RIbe27c10_3, RIbe2b3d8_122);
nand \U$18748 ( \18994 , \1173 , \18993 );
nand \U$18749 ( \18995 , \18992 , \18994 );
xor \U$18750 ( \18996 , RIbe29470_55, RIbe2a190_83);
not \U$18751 ( \18997 , \18996 );
not \U$18752 ( \18998 , \15764 );
or \U$18753 ( \18999 , \18997 , \18998 );
nand \U$18754 ( \19000 , \11400 , \18585 );
nand \U$18755 ( \19001 , \18999 , \19000 );
xor \U$18756 ( \19002 , \18995 , \19001 );
not \U$18757 ( \19003 , \19002 );
xor \U$18758 ( \19004 , RIbe2a3e8_88, RIbe291a0_49);
and \U$18759 ( \19005 , \9264 , \19004 );
and \U$18760 ( \19006 , \10476 , \18577 );
nor \U$18761 ( \19007 , \19005 , \19006 );
not \U$18762 ( \19008 , \19007 );
not \U$18763 ( \19009 , \19008 );
or \U$18764 ( \19010 , \19003 , \19009 );
nand \U$18765 ( \19011 , \19001 , \18995 );
nand \U$18766 ( \19012 , \19010 , \19011 );
not \U$18767 ( \19013 , \19012 );
xor \U$18768 ( \19014 , RIbe290b0_47, RIbe2a7a8_96);
not \U$18769 ( \19015 , \19014 );
not \U$18770 ( \19016 , \2729 );
or \U$18771 ( \19017 , \19015 , \19016 );
nand \U$18772 ( \19018 , \398 , \18787 );
nand \U$18773 ( \19019 , \19017 , \19018 );
xor \U$18774 ( \19020 , RIbe29740_61, RIbe2a910_99);
not \U$18775 ( \19021 , \19020 );
not \U$18776 ( \19022 , \9736 );
or \U$18777 ( \19023 , \19021 , \19022 );
xor \U$18778 ( \19024 , RIbe297b8_62, RIbe2a910_99);
nand \U$18779 ( \19025 , \9726 , \19024 );
nand \U$18780 ( \19026 , \19023 , \19025 );
xor \U$18781 ( \19027 , \19019 , \19026 );
xor \U$18782 ( \19028 , RIbe28cf0_39, RIbe28f48_44);
not \U$18783 ( \19029 , \19028 );
not \U$18784 ( \19030 , \12721 );
or \U$18785 ( \19031 , \19029 , \19030 );
nand \U$18786 ( \19032 , \11201 , \18619 );
nand \U$18787 ( \19033 , \19031 , \19032 );
and \U$18788 ( \19034 , \19027 , \19033 );
and \U$18789 ( \19035 , \19019 , \19026 );
or \U$18790 ( \19036 , \19034 , \19035 );
xor \U$18791 ( \19037 , RIbe2ac58_106, RIbe29038_46);
not \U$18792 ( \19038 , \19037 );
not \U$18793 ( \19039 , \281 );
or \U$18794 ( \19040 , \19038 , \19039 );
nand \U$18795 ( \19041 , \1583 , \18691 );
nand \U$18796 ( \19042 , \19040 , \19041 );
xor \U$18797 ( \19043 , RIbe28b88_36, RIbe2a118_82);
not \U$18798 ( \19044 , \19043 );
not \U$18799 ( \19045 , \2701 );
or \U$18800 ( \19046 , \19044 , \19045 );
xor \U$18801 ( \19047 , RIbe28b88_36, RIbe2a820_97);
nand \U$18802 ( \19048 , \13250 , \19047 );
nand \U$18803 ( \19049 , \19046 , \19048 );
xor \U$18804 ( \19050 , \19042 , \19049 );
xor \U$18805 ( \19051 , RIbe29998_66, RIbe29c68_72);
not \U$18806 ( \19052 , \19051 );
not \U$18807 ( \19053 , \8595 );
or \U$18808 ( \19054 , \19052 , \19053 );
nand \U$18809 ( \19055 , \4580 , \18641 );
nand \U$18810 ( \19056 , \19054 , \19055 );
and \U$18811 ( \19057 , \19050 , \19056 );
and \U$18812 ( \19058 , \19042 , \19049 );
or \U$18813 ( \19059 , \19057 , \19058 );
xor \U$18814 ( \19060 , \19036 , \19059 );
not \U$18815 ( \19061 , \19060 );
or \U$18816 ( \19062 , \19013 , \19061 );
nand \U$18817 ( \19063 , \19059 , \19036 );
nand \U$18818 ( \19064 , \19062 , \19063 );
not \U$18819 ( \19065 , \19064 );
not \U$18820 ( \19066 , RIbe28e58_42);
nand \U$18821 ( \19067 , \19066 , \363 );
and \U$18822 ( \19068 , \19067 , RIbe2ae38_110);
nand \U$18823 ( \19069 , RIbe27c10_3, RIbe28e58_42);
nand \U$18824 ( \19070 , \19069 , RIbe28de0_41);
nor \U$18825 ( \19071 , \19068 , \19070 );
not \U$18826 ( \19072 , \18993 );
not \U$18827 ( \19073 , \7440 );
or \U$18828 ( \19074 , \19072 , \19073 );
xor \U$18829 ( \19075 , RIbe27c10_3, RIbe2b450_123);
nand \U$18830 ( \19076 , \369 , \19075 );
nand \U$18831 ( \19077 , \19074 , \19076 );
xor \U$18832 ( \19078 , \19071 , \19077 );
nand \U$18833 ( \19079 , \7472 , RIbe2ae38_110);
not \U$18834 ( \19080 , \19079 );
not \U$18835 ( \19081 , \19080 );
xor \U$18836 ( \19082 , RIbe29d58_74, RIbe27e68_8);
not \U$18837 ( \19083 , \19082 );
not \U$18838 ( \19084 , \2458 );
or \U$18839 ( \19085 , \19083 , \19084 );
nand \U$18840 ( \19086 , \2464 , \18699 );
nand \U$18841 ( \19087 , \19085 , \19086 );
not \U$18842 ( \19088 , \19087 );
or \U$18843 ( \19089 , \19081 , \19088 );
or \U$18844 ( \19090 , \19087 , \19080 );
xor \U$18845 ( \19091 , RIbe27d78_6, RIbe2b450_123);
not \U$18846 ( \19092 , \19091 );
not \U$18847 ( \19093 , \8898 );
or \U$18848 ( \19094 , \19092 , \19093 );
xor \U$18849 ( \19095 , RIbe27d78_6, RIbe2a730_95);
nand \U$18850 ( \19096 , \10752 , \19095 );
nand \U$18851 ( \19097 , \19094 , \19096 );
nand \U$18852 ( \19098 , \19090 , \19097 );
nand \U$18853 ( \19099 , \19089 , \19098 );
xor \U$18854 ( \19100 , \19078 , \19099 );
xor \U$18855 ( \19101 , RIbe2a028_80, RIbe29218_50);
not \U$18856 ( \19102 , \19101 );
not \U$18857 ( \19103 , \8400 );
or \U$18858 ( \19104 , \19102 , \19103 );
nand \U$18859 ( \19105 , \8930 , \18866 );
nand \U$18860 ( \19106 , \19104 , \19105 );
xor \U$18861 ( \19107 , RIbe293f8_54, RIbe2b108_116);
not \U$18862 ( \19108 , \19107 );
not \U$18863 ( \19109 , \13529 );
or \U$18864 ( \19110 , \19108 , \19109 );
nand \U$18865 ( \19111 , \13533 , \18672 );
nand \U$18866 ( \19112 , \19110 , \19111 );
or \U$18867 ( \19113 , \19106 , \19112 );
xor \U$18868 ( \19114 , RIbe28480_21, RIbe2aa78_102);
not \U$18869 ( \19115 , \19114 );
not \U$18870 ( \19116 , \3483 );
or \U$18871 ( \19117 , \19115 , \19116 );
not \U$18872 ( \19118 , \18741 );
nand \U$18873 ( \19119 , \19118 , \2527 );
nand \U$18874 ( \19120 , \19117 , \19119 );
nand \U$18875 ( \19121 , \19113 , \19120 );
nand \U$18876 ( \19122 , \19106 , \19112 );
nand \U$18877 ( \19123 , \19121 , \19122 );
and \U$18878 ( \19124 , \19100 , \19123 );
and \U$18879 ( \19125 , \19078 , \19099 );
or \U$18880 ( \19126 , \19124 , \19125 );
xor \U$18881 ( \19127 , RIbe28c00_37, RIbe2b180_117);
not \U$18882 ( \19128 , \19127 );
not \U$18883 ( \19129 , \17592 );
or \U$18884 ( \19130 , \19128 , \19129 );
nand \U$18885 ( \19131 , \16646 , \18727 );
nand \U$18886 ( \19132 , \19130 , \19131 );
not \U$18887 ( \19133 , \19132 );
xor \U$18888 ( \19134 , RIbe28a20_33, RIbe2b360_121);
not \U$18889 ( \19135 , \19134 );
not \U$18890 ( \19136 , \1779 );
or \U$18891 ( \19137 , \19135 , \19136 );
nand \U$18892 ( \19138 , \18592 , \1767 );
nand \U$18893 ( \19139 , \19137 , \19138 );
not \U$18894 ( \19140 , \19139 );
nand \U$18895 ( \19141 , \19133 , \19140 );
xor \U$18896 ( \19142 , RIbe28228_16, RIbe2adc0_109);
not \U$18897 ( \19143 , \19142 );
not \U$18898 ( \19144 , \15059 );
or \U$18899 ( \19145 , \19143 , \19144 );
nand \U$18900 ( \19146 , \8679 , \18611 );
nand \U$18901 ( \19147 , \19145 , \19146 );
and \U$18902 ( \19148 , \19141 , \19147 );
not \U$18903 ( \19149 , \19140 );
and \U$18904 ( \19150 , \19132 , \19149 );
nor \U$18905 ( \19151 , \19148 , \19150 );
not \U$18906 ( \19152 , \19151 );
xor \U$18907 ( \19153 , RIbe28930_31, RIbe2a4d8_90);
not \U$18908 ( \19154 , \19153 );
not \U$18909 ( \19155 , \965 );
or \U$18910 ( \19156 , \19154 , \19155 );
nand \U$18911 ( \19157 , \1797 , \18719 );
nand \U$18912 ( \19158 , \19156 , \19157 );
not \U$18913 ( \19159 , \19158 );
xor \U$18914 ( \19160 , RIbe28390_19, RIbe2a898_98);
not \U$18915 ( \19161 , \19160 );
nand \U$18916 ( \19162 , \2645 , \2636 );
not \U$18917 ( \19163 , \19162 );
not \U$18918 ( \19164 , \19163 );
or \U$18919 ( \19165 , \19161 , \19164 );
nand \U$18920 ( \19166 , \2776 , \18709 );
nand \U$18921 ( \19167 , \19165 , \19166 );
xor \U$18922 ( \19168 , RIbe2a550_91, RIbe28138_14);
not \U$18923 ( \19169 , \19168 );
not \U$18924 ( \19170 , \10432 );
or \U$18925 ( \19171 , \19169 , \19170 );
nand \U$18926 ( \19172 , \11484 , \18633 );
nand \U$18927 ( \19173 , \19171 , \19172 );
xor \U$18928 ( \19174 , \19167 , \19173 );
not \U$18929 ( \19175 , \19174 );
or \U$18930 ( \19176 , \19159 , \19175 );
nand \U$18931 ( \19177 , \19173 , \19167 );
nand \U$18932 ( \19178 , \19176 , \19177 );
not \U$18933 ( \19179 , \19178 );
not \U$18934 ( \19180 , \19179 );
or \U$18935 ( \19181 , \19152 , \19180 );
xor \U$18936 ( \19182 , RIbe288b8_30, RIbe2a280_85);
not \U$18937 ( \19183 , \19182 );
not \U$18938 ( \19184 , \10845 );
or \U$18939 ( \19185 , \19183 , \19184 );
nand \U$18940 ( \19186 , \11348 , \18662 );
nand \U$18941 ( \19187 , \19185 , \19186 );
not \U$18942 ( \19188 , \19187 );
not \U$18943 ( \19189 , \19188 );
xor \U$18944 ( \19190 , RIbe296c8_60, RIbe2a6b8_94);
not \U$18945 ( \19191 , \19190 );
not \U$18946 ( \19192 , \9793 );
or \U$18947 ( \19193 , \19191 , \19192 );
nand \U$18948 ( \19194 , \1937 , \18604 );
nand \U$18949 ( \19195 , \19193 , \19194 );
not \U$18950 ( \19196 , \19195 );
not \U$18951 ( \19197 , \19196 );
or \U$18952 ( \19198 , \19189 , \19197 );
xor \U$18953 ( \19199 , RIbe27c88_4, RIbe29e48_76);
not \U$18954 ( \19200 , \19199 );
not \U$18955 ( \19201 , \14307 );
or \U$18956 ( \19202 , \19200 , \19201 );
nand \U$18957 ( \19203 , \4849 , \18682 );
nand \U$18958 ( \19204 , \19202 , \19203 );
nand \U$18959 ( \19205 , \19198 , \19204 );
nand \U$18960 ( \19206 , \19187 , \19195 );
nand \U$18961 ( \19207 , \19205 , \19206 );
nand \U$18962 ( \19208 , \19181 , \19207 );
not \U$18963 ( \19209 , \19179 );
not \U$18964 ( \19210 , \19132 );
not \U$18965 ( \19211 , \19147 );
not \U$18966 ( \19212 , \19140 );
or \U$18967 ( \19213 , \19211 , \19212 );
or \U$18968 ( \19214 , \19140 , \19147 );
nand \U$18969 ( \19215 , \19213 , \19214 );
not \U$18970 ( \19216 , \19215 );
or \U$18971 ( \19217 , \19210 , \19216 );
nand \U$18972 ( \19218 , \19149 , \19147 );
nand \U$18973 ( \19219 , \19217 , \19218 );
nand \U$18974 ( \19220 , \19209 , \19219 );
nand \U$18975 ( \19221 , \19208 , \19220 );
xor \U$18976 ( \19222 , \19126 , \19221 );
not \U$18977 ( \19223 , \19222 );
or \U$18978 ( \19224 , \19065 , \19223 );
nand \U$18979 ( \19225 , \19221 , \19126 );
nand \U$18980 ( \19226 , \19224 , \19225 );
not \U$18981 ( \19227 , \19226 );
and \U$18982 ( \19228 , \19071 , \19077 );
not \U$18983 ( \19229 , \19228 );
not \U$18984 ( \19230 , \19229 );
not \U$18985 ( \19231 , \18731 );
not \U$18986 ( \19232 , \15353 );
or \U$18987 ( \19233 , \19231 , \19232 );
xor \U$18988 ( \19234 , RIbe284f8_22, RIbe2b180_117);
nand \U$18989 ( \19235 , \14966 , \19234 );
nand \U$18990 ( \19236 , \19233 , \19235 );
not \U$18991 ( \19237 , \2518 );
not \U$18992 ( \19238 , \18738 );
or \U$18993 ( \19239 , \19237 , \19238 );
xnor \U$18994 ( \19240 , RIbe29ec0_77, RIbe28480_21);
or \U$18995 ( \19241 , \2670 , \19240 );
nand \U$18996 ( \19242 , \19239 , \19241 );
xor \U$18997 ( \19243 , \19236 , \19242 );
not \U$18998 ( \19244 , \19243 );
and \U$18999 ( \19245 , \19230 , \19244 );
and \U$19000 ( \19246 , \19243 , \19229 );
nor \U$19001 ( \19247 , \19245 , \19246 );
not \U$19002 ( \19248 , \19247 );
not \U$19003 ( \19249 , \19248 );
not \U$19004 ( \19250 , \18668 );
not \U$19005 ( \19251 , \11345 );
or \U$19006 ( \19252 , \19250 , \19251 );
xor \U$19007 ( \19253 , RIbe2a280_85, RIbe29308_52);
nand \U$19008 ( \19254 , \10849 , \19253 );
nand \U$19009 ( \19255 , \19252 , \19254 );
not \U$19010 ( \19256 , \18676 );
not \U$19011 ( \19257 , \17530 );
or \U$19012 ( \19258 , \19256 , \19257 );
xor \U$19013 ( \19259 , RIbe28c78_38, RIbe2b108_116);
nand \U$19014 ( \19260 , \13534 , \19259 );
nand \U$19015 ( \19261 , \19258 , \19260 );
xor \U$19016 ( \19262 , \19255 , \19261 );
not \U$19017 ( \19263 , \18723 );
not \U$19018 ( \19264 , \965 );
or \U$19019 ( \19265 , \19263 , \19264 );
xor \U$19020 ( \19266 , RIbe28930_31, RIbe2a0a0_81);
nand \U$19021 ( \19267 , \1199 , \19266 );
nand \U$19022 ( \19268 , \19265 , \19267 );
xnor \U$19023 ( \19269 , \19262 , \19268 );
not \U$19024 ( \19270 , \19269 );
not \U$19025 ( \19271 , \19270 );
not \U$19026 ( \19272 , \18842 );
not \U$19027 ( \19273 , \8989 );
or \U$19028 ( \19274 , \19272 , \19273 );
xor \U$19029 ( \19275 , RIbe295d8_58, RIbe2a2f8_86);
nand \U$19030 ( \19276 , \11094 , \19275 );
nand \U$19031 ( \19277 , \19274 , \19276 );
not \U$19032 ( \19278 , \18769 );
not \U$19033 ( \19279 , \11321 );
or \U$19034 ( \19280 , \19278 , \19279 );
xor \U$19035 ( \19281 , RIbe28de0_41, RIbe2b3d8_122);
nand \U$19036 ( \19282 , \7472 , \19281 );
nand \U$19037 ( \19283 , \19280 , \19282 );
not \U$19038 ( \19284 , \19283 );
not \U$19039 ( \19285 , \18824 );
not \U$19040 ( \19286 , \10466 );
or \U$19041 ( \19287 , \19285 , \19286 );
xor \U$19042 ( \19288 , RIbe27fd0_11, RIbe298a8_64);
nand \U$19043 ( \19289 , \7709 , \19288 );
nand \U$19044 ( \19290 , \19287 , \19289 );
not \U$19045 ( \19291 , \19290 );
not \U$19046 ( \19292 , \19291 );
or \U$19047 ( \19293 , \19284 , \19292 );
or \U$19048 ( \19294 , \19291 , \19283 );
nand \U$19049 ( \19295 , \19293 , \19294 );
xor \U$19050 ( \19296 , \19277 , \19295 );
not \U$19051 ( \19297 , \19296 );
not \U$19052 ( \19298 , \19297 );
or \U$19053 ( \19299 , \19271 , \19298 );
nand \U$19054 ( \19300 , \19296 , \19269 );
nand \U$19055 ( \19301 , \19299 , \19300 );
not \U$19056 ( \19302 , \19301 );
or \U$19057 ( \19303 , \19249 , \19302 );
nand \U$19058 ( \19304 , \19296 , \19270 );
nand \U$19059 ( \19305 , \19303 , \19304 );
not \U$19060 ( \19306 , \19305 );
not \U$19061 ( \19307 , \19306 );
xor \U$19062 ( \19308 , RIbe28390_19, RIbe2b6a8_128);
not \U$19063 ( \19309 , \19308 );
not \U$19064 ( \19310 , \3712 );
or \U$19065 ( \19311 , \19309 , \19310 );
nand \U$19066 ( \19312 , \3714 , \17858 );
nand \U$19067 ( \19313 , \19311 , \19312 );
not \U$19068 ( \19314 , \19313 );
not \U$19069 ( \19315 , \19281 );
not \U$19070 ( \19316 , \331 );
or \U$19071 ( \19317 , \19315 , \19316 );
nand \U$19072 ( \19318 , \346 , \17884 );
nand \U$19073 ( \19319 , \19317 , \19318 );
not \U$19074 ( \19320 , \19319 );
or \U$19075 ( \19321 , RIbe28de0_41, RIbe29920_65);
nand \U$19076 ( \19322 , \19321 , RIbe2ae38_110);
nand \U$19077 ( \19323 , RIbe28de0_41, RIbe29920_65);
nand \U$19078 ( \19324 , \19322 , \19323 , RIbe27b98_2);
not \U$19079 ( \19325 , \19324 );
and \U$19080 ( \19326 , \19320 , \19325 );
and \U$19081 ( \19327 , \19319 , \19324 );
nor \U$19082 ( \19328 , \19326 , \19327 );
not \U$19083 ( \19329 , \19328 );
or \U$19084 ( \19330 , \19314 , \19329 );
or \U$19085 ( \19331 , \19313 , \19328 );
nand \U$19086 ( \19332 , \19330 , \19331 );
not \U$19087 ( \19333 , \18855 );
not \U$19088 ( \19334 , \2618 );
or \U$19089 ( \19335 , \19333 , \19334 );
xor \U$19090 ( \19336 , RIbe29ce0_73, RIbe285e8_24);
nand \U$19091 ( \19337 , \2626 , \19336 );
nand \U$19092 ( \19338 , \19335 , \19337 );
not \U$19093 ( \19339 , \19338 );
not \U$19094 ( \19340 , \19075 );
not \U$19095 ( \19341 , \1103 );
or \U$19096 ( \19342 , \19340 , \19341 );
xor \U$19097 ( \19343 , RIbe27c10_3, RIbe2a730_95);
nand \U$19098 ( \19344 , \1498 , \19343 );
nand \U$19099 ( \19345 , \19342 , \19344 );
nand \U$19100 ( \19346 , \1734 , RIbe2ae38_110);
not \U$19101 ( \19347 , \19346 );
and \U$19102 ( \19348 , \19345 , \19347 );
not \U$19103 ( \19349 , \19345 );
and \U$19104 ( \19350 , \19349 , \19346 );
nor \U$19105 ( \19351 , \19348 , \19350 );
not \U$19106 ( \19352 , \19351 );
or \U$19107 ( \19353 , \19339 , \19352 );
nand \U$19108 ( \19354 , \19345 , \19347 );
nand \U$19109 ( \19355 , \19353 , \19354 );
not \U$19110 ( \19356 , \19355 );
and \U$19111 ( \19357 , \19332 , \19356 );
not \U$19112 ( \19358 , \19332 );
and \U$19113 ( \19359 , \19358 , \19355 );
nor \U$19114 ( \19360 , \19357 , \19359 );
not \U$19115 ( \19361 , \19360 );
not \U$19116 ( \19362 , \19228 );
not \U$19117 ( \19363 , \19243 );
or \U$19118 ( \19364 , \19362 , \19363 );
nand \U$19119 ( \19365 , \19236 , \19242 );
nand \U$19120 ( \19366 , \19364 , \19365 );
xor \U$19121 ( \19367 , RIbe286d8_26, RIbe2b018_114);
not \U$19122 ( \19368 , \19367 );
not \U$19123 ( \19369 , \15967 );
or \U$19124 ( \19370 , \19368 , \19369 );
buf \U$19125 ( \19371 , \15952 );
xor \U$19126 ( \19372 , RIbe27ee0_9, RIbe2b018_114);
nand \U$19127 ( \19373 , \19371 , \19372 );
nand \U$19128 ( \19374 , \19370 , \19373 );
xor \U$19129 ( \19375 , RIbe297b8_62, RIbe2a3e8_88);
not \U$19130 ( \19376 , \19375 );
not \U$19131 ( \19377 , \9263 );
or \U$19132 ( \19378 , \19376 , \19377 );
nand \U$19133 ( \19379 , \9268 , \17715 );
nand \U$19134 ( \19380 , \19378 , \19379 );
xor \U$19135 ( \19381 , \19374 , \19380 );
xor \U$19136 ( \19382 , RIbe2b4c8_124, RIbe29038_46);
not \U$19137 ( \19383 , \19382 );
not \U$19138 ( \19384 , \979 );
or \U$19139 ( \19385 , \19383 , \19384 );
xor \U$19140 ( \19386 , RIbe29038_46, RIbe2b540_125);
nand \U$19141 ( \19387 , \1805 , \19386 );
nand \U$19142 ( \19388 , \19385 , \19387 );
and \U$19143 ( \19389 , \19381 , \19388 );
not \U$19144 ( \19390 , \19381 );
not \U$19145 ( \19391 , \19388 );
and \U$19146 ( \19392 , \19390 , \19391 );
nor \U$19147 ( \19393 , \19389 , \19392 );
xor \U$19148 ( \19394 , \19366 , \19393 );
not \U$19149 ( \19395 , \19394 );
or \U$19150 ( \19396 , \19361 , \19395 );
or \U$19151 ( \19397 , \19394 , \19360 );
nand \U$19152 ( \19398 , \19396 , \19397 );
not \U$19153 ( \19399 , \19398 );
or \U$19154 ( \19400 , \19307 , \19399 );
or \U$19155 ( \19401 , \19398 , \19306 );
nand \U$19156 ( \19402 , \19400 , \19401 );
not \U$19157 ( \19403 , \19402 );
or \U$19158 ( \19404 , \19227 , \19403 );
not \U$19159 ( \19405 , \19306 );
nand \U$19160 ( \19406 , \19405 , \19398 );
nand \U$19161 ( \19407 , \19404 , \19406 );
not \U$19162 ( \19408 , \19407 );
xor \U$19163 ( \19409 , \17847 , \17854 );
and \U$19164 ( \19410 , \19409 , \17864 );
not \U$19165 ( \19411 , \19409 );
not \U$19166 ( \19412 , \17864 );
and \U$19167 ( \19413 , \19411 , \19412 );
nor \U$19168 ( \19414 , \19410 , \19413 );
xor \U$19169 ( \19415 , RIbe29380_53, RIbe2aaf0_103);
not \U$19170 ( \19416 , \19415 );
not \U$19171 ( \19417 , \18832 );
or \U$19172 ( \19418 , \19416 , \19417 );
nand \U$19173 ( \19419 , RIbe2aaf0_103, RIbe2ab68_104);
nand \U$19174 ( \19420 , \19418 , \19419 );
xor \U$19175 ( \19421 , RIbe2aeb0_111, RIbe27b98_2);
not \U$19176 ( \19422 , \19421 );
not \U$19177 ( \19423 , \4827 );
or \U$19178 ( \19424 , \19422 , \19423 );
nand \U$19179 ( \19425 , \267 , \18189 );
nand \U$19180 ( \19426 , \19424 , \19425 );
xor \U$19181 ( \19427 , \19420 , \19426 );
xor \U$19182 ( \19428 , RIbe2a028_80, RIbe291a0_49);
not \U$19183 ( \19429 , \19428 );
not \U$19184 ( \19430 , \9530 );
or \U$19185 ( \19431 , \19429 , \19430 );
nand \U$19186 ( \19432 , \8930 , \17644 );
nand \U$19187 ( \19433 , \19431 , \19432 );
and \U$19188 ( \19434 , \19427 , \19433 );
not \U$19189 ( \19435 , \19427 );
not \U$19190 ( \19436 , \19433 );
and \U$19191 ( \19437 , \19435 , \19436 );
nor \U$19192 ( \19438 , \19434 , \19437 );
xor \U$19193 ( \19439 , \19414 , \19438 );
xor \U$19194 ( \19440 , RIbe285e8_24, RIbe29b78_70);
not \U$19195 ( \19441 , \19440 );
not \U$19196 ( \19442 , \11174 );
or \U$19197 ( \19443 , \19441 , \19442 );
nand \U$19198 ( \19444 , \8270 , \17973 );
nand \U$19199 ( \19445 , \19443 , \19444 );
xor \U$19200 ( \19446 , RIbe288b8_30, RIbe2a550_91);
not \U$19201 ( \19447 , \19446 );
not \U$19202 ( \19448 , \10433 );
or \U$19203 ( \19449 , \19447 , \19448 );
nand \U$19204 ( \19450 , \11485 , \17961 );
nand \U$19205 ( \19451 , \19449 , \19450 );
xor \U$19206 ( \19452 , \19445 , \19451 );
xor \U$19207 ( \19453 , RIbe290b0_47, RIbe2a6b8_94);
not \U$19208 ( \19454 , \19453 );
not \U$19209 ( \19455 , \9114 );
or \U$19210 ( \19456 , \19454 , \19455 );
nand \U$19211 ( \19457 , \399 , \17678 );
nand \U$19212 ( \19458 , \19456 , \19457 );
xor \U$19213 ( \19459 , \19452 , \19458 );
xor \U$19214 ( \19460 , \19439 , \19459 );
xor \U$19215 ( \19461 , RIbe29e48_76, RIbe29b00_69);
not \U$19216 ( \19462 , \19461 );
not \U$19217 ( \19463 , \7716 );
or \U$19218 ( \19464 , \19462 , \19463 );
nand \U$19219 ( \19465 , \4850 , \17651 );
nand \U$19220 ( \19466 , \19464 , \19465 );
xor \U$19221 ( \19467 , RIbe28750_27, RIbe2b180_117);
not \U$19222 ( \19468 , \19467 );
not \U$19223 ( \19469 , \14852 );
or \U$19224 ( \19470 , \19468 , \19469 );
nand \U$19225 ( \19471 , \16646 , \17589 );
nand \U$19226 ( \19472 , \19470 , \19471 );
xor \U$19227 ( \19473 , \19466 , \19472 );
xor \U$19228 ( \19474 , RIbe2adc0_109, RIbe296c8_60);
not \U$19229 ( \19475 , \19474 );
not \U$19230 ( \19476 , \1130 );
or \U$19231 ( \19477 , \19475 , \19476 );
nand \U$19232 ( \19478 , \908 , \17670 );
nand \U$19233 ( \19479 , \19477 , \19478 );
xor \U$19234 ( \19480 , \19473 , \19479 );
xor \U$19235 ( \19481 , RIbe27fd0_11, RIbe29998_66);
not \U$19236 ( \19482 , \19481 );
not \U$19237 ( \19483 , \11366 );
or \U$19238 ( \19484 , \19482 , \19483 );
nand \U$19239 ( \19485 , \2707 , \17538 );
nand \U$19240 ( \19486 , \19484 , \19485 );
xor \U$19241 ( \19487 , RIbe28318_18, RIbe2b108_116);
not \U$19242 ( \19488 , \19487 );
not \U$19243 ( \19489 , \17530 );
or \U$19244 ( \19490 , \19488 , \19489 );
nand \U$19245 ( \19491 , \16875 , \17528 );
nand \U$19246 ( \19492 , \19490 , \19491 );
xor \U$19247 ( \19493 , \19486 , \19492 );
xor \U$19248 ( \19494 , RIbe2b360_121, RIbe28228_16);
not \U$19249 ( \19495 , \19494 );
not \U$19250 ( \19496 , \879 );
or \U$19251 ( \19497 , \19495 , \19496 );
nand \U$19252 ( \19498 , \8680 , \17985 );
nand \U$19253 ( \19499 , \19497 , \19498 );
and \U$19254 ( \19500 , \19493 , \19499 );
not \U$19255 ( \19501 , \19493 );
not \U$19256 ( \19502 , \19499 );
and \U$19257 ( \19503 , \19501 , \19502 );
nor \U$19258 ( \19504 , \19500 , \19503 );
and \U$19259 ( \19505 , \19480 , \19504 );
not \U$19260 ( \19506 , \19480 );
not \U$19261 ( \19507 , \19504 );
and \U$19262 ( \19508 , \19506 , \19507 );
nor \U$19263 ( \19509 , \19505 , \19508 );
xor \U$19264 ( \19510 , \17763 , \17743 );
and \U$19265 ( \19511 , \19509 , \19510 );
not \U$19266 ( \19512 , \19509 );
not \U$19267 ( \19513 , \19510 );
and \U$19268 ( \19514 , \19512 , \19513 );
nor \U$19269 ( \19515 , \19511 , \19514 );
xor \U$19270 ( \19516 , \19460 , \19515 );
not \U$19271 ( \19517 , \19372 );
not \U$19272 ( \19518 , \16811 );
or \U$19273 ( \19519 , \19517 , \19518 );
nand \U$19274 ( \19520 , \15953 , \17568 );
nand \U$19275 ( \19521 , \19519 , \19520 );
not \U$19276 ( \19522 , \19386 );
not \U$19277 ( \19523 , \281 );
or \U$19278 ( \19524 , \19522 , \19523 );
nand \U$19279 ( \19525 , \1583 , \17934 );
nand \U$19280 ( \19526 , \19524 , \19525 );
not \U$19281 ( \19527 , \19526 );
xor \U$19282 ( \19528 , \19521 , \19527 );
xor \U$19283 ( \19529 , RIbe2a7a8_96, RIbe27c10_3);
not \U$19284 ( \19530 , \19529 );
not \U$19285 ( \19531 , \1493 );
or \U$19286 ( \19532 , \19530 , \19531 );
nand \U$19287 ( \19533 , \1174 , \17922 );
nand \U$19288 ( \19534 , \19532 , \19533 );
xor \U$19289 ( \19535 , \19528 , \19534 );
not \U$19290 ( \19536 , \19535 );
not \U$19291 ( \19537 , \17732 );
not \U$19292 ( \19538 , \17723 );
or \U$19293 ( \19539 , \19537 , \19538 );
or \U$19294 ( \19540 , \17732 , \17723 );
nand \U$19295 ( \19541 , \19539 , \19540 );
xor \U$19296 ( \19542 , \17713 , \19541 );
not \U$19297 ( \19543 , \19542 );
xor \U$19298 ( \19544 , \19536 , \19543 );
xor \U$19299 ( \19545 , \17790 , \17775 );
xor \U$19300 ( \19546 , \19544 , \19545 );
xor \U$19301 ( \19547 , \19516 , \19546 );
not \U$19302 ( \19548 , \19547 );
nand \U$19303 ( \19549 , \19408 , \19548 );
not \U$19304 ( \19550 , \19549 );
or \U$19305 ( \19551 , \18988 , \19550 );
nand \U$19306 ( \19552 , \19407 , \19547 );
nand \U$19307 ( \19553 , \19551 , \19552 );
not \U$19308 ( \19554 , \19553 );
not \U$19309 ( \19555 , \19536 );
not \U$19310 ( \19556 , \19543 );
or \U$19311 ( \19557 , \19555 , \19556 );
not \U$19312 ( \19558 , \19535 );
not \U$19313 ( \19559 , \19542 );
or \U$19314 ( \19560 , \19558 , \19559 );
nand \U$19315 ( \19561 , \19560 , \19545 );
nand \U$19316 ( \19562 , \19557 , \19561 );
not \U$19317 ( \19563 , \19438 );
not \U$19318 ( \19564 , \19459 );
or \U$19319 ( \19565 , \19563 , \19564 );
or \U$19320 ( \19566 , \19459 , \19438 );
nand \U$19321 ( \19567 , \19566 , \19414 );
nand \U$19322 ( \19568 , \19565 , \19567 );
xor \U$19323 ( \19569 , \19562 , \19568 );
xor \U$19324 ( \19570 , RIbe27b20_1, RIbe27e68_8);
not \U$19325 ( \19571 , \19570 );
not \U$19326 ( \19572 , \2458 );
or \U$19327 ( \19573 , \19571 , \19572 );
nand \U$19328 ( \19574 , \13306 , \17753 );
nand \U$19329 ( \19575 , \19573 , \19574 );
xor \U$19330 ( \19576 , RIbe2aaf0_103, RIbe28048_12);
not \U$19331 ( \19577 , \19576 );
not \U$19332 ( \19578 , RIbe2ab68_104);
nand \U$19333 ( \19579 , \19578 , RIbe2aaf0_103);
buf \U$19334 ( \19580 , \19579 );
not \U$19335 ( \19581 , \19580 );
not \U$19336 ( \19582 , \19581 );
or \U$19337 ( \19583 , \19577 , \19582 );
nand \U$19338 ( \19584 , \19415 , RIbe2ab68_104);
nand \U$19339 ( \19585 , \19583 , \19584 );
or \U$19340 ( \19586 , \19575 , \19585 );
xor \U$19341 ( \19587 , RIbe27d78_6, RIbe2abe0_105);
not \U$19342 ( \19588 , \19587 );
not \U$19343 ( \19589 , \1043 );
or \U$19344 ( \19590 , \19588 , \19589 );
nand \U$19345 ( \19591 , \314 , \17745 );
nand \U$19346 ( \19592 , \19590 , \19591 );
nand \U$19347 ( \19593 , \19586 , \19592 );
nand \U$19348 ( \19594 , \19575 , \19585 );
nand \U$19349 ( \19595 , \19593 , \19594 );
xnor \U$19350 ( \19596 , \17881 , \17889 );
xor \U$19351 ( \19597 , \19595 , \19596 );
xor \U$19352 ( \19598 , RIbe280c0_13, RIbe2a460_89);
not \U$19353 ( \19599 , \19598 );
not \U$19354 ( \19600 , \861 );
or \U$19355 ( \19601 , \19599 , \19600 );
nand \U$19356 ( \19602 , \1265 , \17777 );
nand \U$19357 ( \19603 , \19601 , \19602 );
not \U$19358 ( \19604 , \19603 );
xor \U$19359 ( \19605 , RIbe294e8_56, RIbe2a550_91);
not \U$19360 ( \19606 , \19605 );
buf \U$19361 ( \19607 , \10433 );
not \U$19362 ( \19608 , \19607 );
or \U$19363 ( \19609 , \19606 , \19608 );
nand \U$19364 ( \19610 , \12004 , \19446 );
nand \U$19365 ( \19611 , \19609 , \19610 );
not \U$19366 ( \19612 , \19611 );
or \U$19367 ( \19613 , \19604 , \19612 );
or \U$19368 ( \19614 , \19611 , \19603 );
xor \U$19369 ( \19615 , RIbe290b0_47, RIbe2a640_93);
not \U$19370 ( \19616 , \19615 );
not \U$19371 ( \19617 , \2731 );
or \U$19372 ( \19618 , \19616 , \19617 );
nand \U$19373 ( \19619 , \2071 , \19453 );
nand \U$19374 ( \19620 , \19618 , \19619 );
nand \U$19375 ( \19621 , \19614 , \19620 );
nand \U$19376 ( \19622 , \19613 , \19621 );
and \U$19377 ( \19623 , \19597 , \19622 );
and \U$19378 ( \19624 , \19595 , \19596 );
or \U$19379 ( \19625 , \19623 , \19624 );
xor \U$19380 ( \19626 , \19569 , \19625 );
xor \U$19381 ( \19627 , \17866 , \17840 );
buf \U$19382 ( \19628 , \17894 );
xnor \U$19383 ( \19629 , \19627 , \19628 );
not \U$19384 ( \19630 , \19504 );
not \U$19385 ( \19631 , \19510 );
or \U$19386 ( \19632 , \19630 , \19631 );
or \U$19387 ( \19633 , \19504 , \19510 );
nand \U$19388 ( \19634 , \19633 , \19480 );
nand \U$19389 ( \19635 , \19632 , \19634 );
xor \U$19390 ( \19636 , \19629 , \19635 );
or \U$19391 ( \19637 , \19492 , \19486 );
nand \U$19392 ( \19638 , \19637 , \19499 );
nand \U$19393 ( \19639 , \19492 , \19486 );
nand \U$19394 ( \19640 , \19638 , \19639 );
buf \U$19395 ( \19641 , \19640 );
not \U$19396 ( \19642 , \19641 );
and \U$19397 ( \19643 , \19427 , \19433 );
and \U$19398 ( \19644 , \19426 , \19420 );
nor \U$19399 ( \19645 , \19643 , \19644 );
not \U$19400 ( \19646 , \19645 );
or \U$19401 ( \19647 , \19642 , \19646 );
not \U$19402 ( \19648 , \19645 );
not \U$19403 ( \19649 , \19640 );
nand \U$19404 ( \19650 , \19648 , \19649 );
nand \U$19405 ( \19651 , \19647 , \19650 );
not \U$19406 ( \19652 , \19479 );
not \U$19407 ( \19653 , \19473 );
or \U$19408 ( \19654 , \19652 , \19653 );
nand \U$19409 ( \19655 , \19466 , \19472 );
nand \U$19410 ( \19656 , \19654 , \19655 );
buf \U$19411 ( \19657 , \19656 );
not \U$19412 ( \19658 , \19657 );
and \U$19413 ( \19659 , \19651 , \19658 );
not \U$19414 ( \19660 , \19651 );
and \U$19415 ( \19661 , \19660 , \19657 );
nor \U$19416 ( \19662 , \19659 , \19661 );
buf \U$19417 ( \19663 , \19662 );
xor \U$19418 ( \19664 , \19636 , \19663 );
xor \U$19419 ( \19665 , \19626 , \19664 );
xor \U$19420 ( \19666 , \19460 , \19515 );
and \U$19421 ( \19667 , \19666 , \19546 );
and \U$19422 ( \19668 , \19460 , \19515 );
or \U$19423 ( \19669 , \19667 , \19668 );
xor \U$19424 ( \19670 , \19665 , \19669 );
not \U$19425 ( \19671 , \19670 );
not \U$19426 ( \19672 , \19671 );
or \U$19427 ( \19673 , \19554 , \19672 );
or \U$19428 ( \19674 , \19553 , \19671 );
nand \U$19429 ( \19675 , \19673 , \19674 );
not \U$19430 ( \19676 , \19675 );
xor \U$19431 ( \19677 , \18878 , \18882 );
and \U$19432 ( \19678 , \19677 , \18885 );
and \U$19433 ( \19679 , \18878 , \18882 );
or \U$19434 ( \19680 , \19678 , \19679 );
not \U$19435 ( \19681 , \19680 );
not \U$19436 ( \19682 , \19360 );
not \U$19437 ( \19683 , \19682 );
not \U$19438 ( \19684 , \19394 );
or \U$19439 ( \19685 , \19683 , \19684 );
nand \U$19440 ( \19686 , \19366 , \19393 );
nand \U$19441 ( \19687 , \19685 , \19686 );
not \U$19442 ( \19688 , \19687 );
nand \U$19443 ( \19689 , \19681 , \19688 );
not \U$19444 ( \19690 , \19689 );
not \U$19445 ( \19691 , \18638 );
not \U$19446 ( \19692 , \10433 );
or \U$19447 ( \19693 , \19691 , \19692 );
nand \U$19448 ( \19694 , \11227 , \19605 );
nand \U$19449 ( \19695 , \19693 , \19694 );
not \U$19450 ( \19696 , \18623 );
not \U$19451 ( \19697 , \9618 );
or \U$19452 ( \19698 , \19696 , \19697 );
xor \U$19453 ( \19699 , RIbe28f48_44, RIbe28d68_40);
nand \U$19454 ( \19700 , \3249 , \19699 );
nand \U$19455 ( \19701 , \19698 , \19700 );
xor \U$19456 ( \19702 , \19695 , \19701 );
not \U$19457 ( \19703 , \18615 );
not \U$19458 ( \19704 , \1061 );
or \U$19459 ( \19705 , \19703 , \19704 );
xor \U$19460 ( \19706 , RIbe2b2e8_120, RIbe28228_16);
nand \U$19461 ( \19707 , \8680 , \19706 );
nand \U$19462 ( \19708 , \19705 , \19707 );
and \U$19463 ( \19709 , \19702 , \19708 );
and \U$19464 ( \19710 , \19695 , \19701 );
or \U$19465 ( \19711 , \19709 , \19710 );
not \U$19466 ( \19712 , \18645 );
not \U$19467 ( \19713 , \8594 );
or \U$19468 ( \19714 , \19712 , \19713 );
xor \U$19469 ( \19715 , RIbe27df0_7, RIbe29c68_72);
nand \U$19470 ( \19716 , \4580 , \19715 );
nand \U$19471 ( \19717 , \19714 , \19716 );
not \U$19472 ( \19718 , \18652 );
not \U$19473 ( \19719 , \15345 );
or \U$19474 ( \19720 , \19718 , \19719 );
buf \U$19475 ( \19721 , \16728 );
xor \U$19476 ( \19722 , RIbe28840_29, RIbe2af28_112);
nand \U$19477 ( \19723 , \19721 , \19722 );
nand \U$19478 ( \19724 , \19720 , \19723 );
xor \U$19479 ( \19725 , \19717 , \19724 );
not \U$19480 ( \19726 , \18695 );
not \U$19481 ( \19727 , \979 );
or \U$19482 ( \19728 , \19726 , \19727 );
nand \U$19483 ( \19729 , \287 , \19382 );
nand \U$19484 ( \19730 , \19728 , \19729 );
and \U$19485 ( \19731 , \19725 , \19730 );
and \U$19486 ( \19732 , \19717 , \19724 );
or \U$19487 ( \19733 , \19731 , \19732 );
xor \U$19488 ( \19734 , \19711 , \19733 );
not \U$19489 ( \19735 , \1131 );
not \U$19490 ( \19736 , \18608 );
not \U$19491 ( \19737 , \19736 );
and \U$19492 ( \19738 , \19735 , \19737 );
xor \U$19493 ( \19739 , RIbe2ad48_108, RIbe296c8_60);
and \U$19494 ( \19740 , \1137 , \19739 );
nor \U$19495 ( \19741 , \19738 , \19740 );
not \U$19496 ( \19742 , \19741 );
not \U$19497 ( \19743 , \19742 );
xor \U$19498 ( \19744 , RIbe28138_14, RIbe2a910_99);
not \U$19499 ( \19745 , \19744 );
not \U$19500 ( \19746 , \11453 );
or \U$19501 ( \19747 , \19745 , \19746 );
xor \U$19502 ( \19748 , RIbe2a910_99, RIbe282a0_17);
nand \U$19503 ( \19749 , \10401 , \19748 );
nand \U$19504 ( \19750 , \19747 , \19749 );
not \U$19505 ( \19751 , \19750 );
xor \U$19506 ( \19752 , RIbe28b88_36, RIbe2a898_98);
not \U$19507 ( \19753 , \19752 );
not \U$19508 ( \19754 , \2701 );
or \U$19509 ( \19755 , \19753 , \19754 );
xor \U$19510 ( \19756 , RIbe28b88_36, RIbe2aa00_101);
nand \U$19511 ( \19757 , \13250 , \19756 );
nand \U$19512 ( \19758 , \19755 , \19757 );
not \U$19513 ( \19759 , \19758 );
not \U$19514 ( \19760 , \19759 );
or \U$19515 ( \19761 , \19751 , \19760 );
or \U$19516 ( \19762 , \19750 , \19759 );
nand \U$19517 ( \19763 , \19761 , \19762 );
not \U$19518 ( \19764 , \19763 );
or \U$19519 ( \19765 , \19743 , \19764 );
not \U$19520 ( \19766 , \19759 );
nand \U$19521 ( \19767 , \19766 , \19750 );
nand \U$19522 ( \19768 , \19765 , \19767 );
xor \U$19523 ( \19769 , \19734 , \19768 );
not \U$19524 ( \19770 , \19769 );
not \U$19525 ( \19771 , \19261 );
not \U$19526 ( \19772 , \19255 );
or \U$19527 ( \19773 , \19771 , \19772 );
or \U$19528 ( \19774 , \19261 , \19255 );
nand \U$19529 ( \19775 , \19774 , \19268 );
nand \U$19530 ( \19776 , \19773 , \19775 );
not \U$19531 ( \19777 , \19776 );
not \U$19532 ( \19778 , \18581 );
not \U$19533 ( \19779 , \9262 );
or \U$19534 ( \19780 , \19778 , \19779 );
nand \U$19535 ( \19781 , \9089 , \19375 );
nand \U$19536 ( \19782 , \19780 , \19781 );
not \U$19537 ( \19783 , \19782 );
not \U$19538 ( \19784 , \18596 );
not \U$19539 ( \19785 , \9192 );
or \U$19540 ( \19786 , \19784 , \19785 );
xor \U$19541 ( \19787 , RIbe28a20_33, RIbe2a820_97);
nand \U$19542 ( \19788 , \5055 , \19787 );
nand \U$19543 ( \19789 , \19786 , \19788 );
not \U$19544 ( \19790 , \19789 );
or \U$19545 ( \19791 , \19783 , \19790 );
not \U$19546 ( \19792 , \19789 );
not \U$19547 ( \19793 , \19792 );
not \U$19548 ( \19794 , \19782 );
not \U$19549 ( \19795 , \19794 );
or \U$19550 ( \19796 , \19793 , \19795 );
xor \U$19551 ( \19797 , RIbe27d78_6, RIbe2a7a8_96);
not \U$19552 ( \19798 , \19797 );
not \U$19553 ( \19799 , \1043 );
or \U$19554 ( \19800 , \19798 , \19799 );
nand \U$19555 ( \19801 , \314 , \19587 );
nand \U$19556 ( \19802 , \19800 , \19801 );
nand \U$19557 ( \19803 , \19796 , \19802 );
nand \U$19558 ( \19804 , \19791 , \19803 );
not \U$19559 ( \19805 , \19804 );
not \U$19560 ( \19806 , \19805 );
or \U$19561 ( \19807 , \19777 , \19806 );
not \U$19562 ( \19808 , \19776 );
nand \U$19563 ( \19809 , \19808 , \19804 );
nand \U$19564 ( \19810 , \19807 , \19809 );
not \U$19565 ( \19811 , \18686 );
not \U$19566 ( \19812 , \10938 );
or \U$19567 ( \19813 , \19811 , \19812 );
xor \U$19568 ( \19814 , RIbe29a10_67, RIbe29e48_76);
nand \U$19569 ( \19815 , \7368 , \19814 );
nand \U$19570 ( \19816 , \19813 , \19815 );
not \U$19571 ( \19817 , \19816 );
not \U$19572 ( \19818 , \18713 );
not \U$19573 ( \19819 , \14806 );
or \U$19574 ( \19820 , \19818 , \19819 );
nand \U$19575 ( \19821 , \2777 , \19308 );
nand \U$19576 ( \19822 , \19820 , \19821 );
not \U$19577 ( \19823 , \19822 );
not \U$19578 ( \19824 , \19823 );
not \U$19579 ( \19825 , \18703 );
not \U$19580 ( \19826 , \2458 );
or \U$19581 ( \19827 , \19825 , \19826 );
nand \U$19582 ( \19828 , \13306 , \19570 );
nand \U$19583 ( \19829 , \19827 , \19828 );
not \U$19584 ( \19830 , \19829 );
or \U$19585 ( \19831 , \19824 , \19830 );
or \U$19586 ( \19832 , \19829 , \19823 );
nand \U$19587 ( \19833 , \19831 , \19832 );
not \U$19588 ( \19834 , \19833 );
or \U$19589 ( \19835 , \19817 , \19834 );
nand \U$19590 ( \19836 , \19829 , \19822 );
nand \U$19591 ( \19837 , \19835 , \19836 );
not \U$19592 ( \19838 , \19837 );
and \U$19593 ( \19839 , \19810 , \19838 );
not \U$19594 ( \19840 , \19810 );
and \U$19595 ( \19841 , \19840 , \19837 );
nor \U$19596 ( \19842 , \19839 , \19841 );
not \U$19597 ( \19843 , \19842 );
not \U$19598 ( \19844 , \19843 );
not \U$19599 ( \19845 , \19816 );
not \U$19600 ( \19846 , \19833 );
not \U$19601 ( \19847 , \19846 );
or \U$19602 ( \19848 , \19845 , \19847 );
not \U$19603 ( \19849 , \19816 );
nand \U$19604 ( \19850 , \19849 , \19833 );
nand \U$19605 ( \19851 , \19848 , \19850 );
not \U$19606 ( \19852 , \18778 );
or \U$19607 ( \19853 , RIbe2b018_114, RIbe2b630_127);
nand \U$19608 ( \19854 , \19853 , \15964 );
not \U$19609 ( \19855 , \19854 );
not \U$19610 ( \19856 , \19855 );
or \U$19611 ( \19857 , \19852 , \19856 );
nand \U$19612 ( \19858 , \15952 , \19367 );
nand \U$19613 ( \19859 , \19857 , \19858 );
not \U$19614 ( \19860 , \18589 );
not \U$19615 ( \19861 , \10831 );
or \U$19616 ( \19862 , \19860 , \19861 );
xor \U$19617 ( \19863 , RIbe28a98_34, RIbe2a190_83);
nand \U$19618 ( \19864 , \11399 , \19863 );
nand \U$19619 ( \19865 , \19862 , \19864 );
xor \U$19620 ( \19866 , \19859 , \19865 );
not \U$19621 ( \19867 , \18791 );
not \U$19622 ( \19868 , \10567 );
or \U$19623 ( \19869 , \19867 , \19868 );
nand \U$19624 ( \19870 , \398 , \19615 );
nand \U$19625 ( \19871 , \19869 , \19870 );
and \U$19626 ( \19872 , \19866 , \19871 );
not \U$19627 ( \19873 , \19866 );
not \U$19628 ( \19874 , \19871 );
and \U$19629 ( \19875 , \19873 , \19874 );
nor \U$19630 ( \19876 , \19872 , \19875 );
xor \U$19631 ( \19877 , \19851 , \19876 );
not \U$19632 ( \19878 , \18835 );
not \U$19633 ( \19879 , \18832 );
or \U$19634 ( \19880 , \19878 , \19879 );
nand \U$19635 ( \19881 , \19576 , RIbe2ab68_104);
nand \U$19636 ( \19882 , \19880 , \19881 );
not \U$19637 ( \19883 , \18862 );
not \U$19638 ( \19884 , \1053 );
or \U$19639 ( \19885 , \19883 , \19884 );
nand \U$19640 ( \19886 , \1263 , \19598 );
nand \U$19641 ( \19887 , \19885 , \19886 );
xor \U$19642 ( \19888 , \19882 , \19887 );
not \U$19643 ( \19889 , \18870 );
not \U$19644 ( \19890 , \8400 );
or \U$19645 ( \19891 , \19889 , \19890 );
xor \U$19646 ( \19892 , RIbe2a028_80, RIbe29128_48);
nand \U$19647 ( \19893 , \8172 , \19892 );
nand \U$19648 ( \19894 , \19891 , \19893 );
xnor \U$19649 ( \19895 , \19888 , \19894 );
not \U$19650 ( \19896 , \19895 );
and \U$19651 ( \19897 , \19877 , \19896 );
and \U$19652 ( \19898 , \19851 , \19876 );
or \U$19653 ( \19899 , \19897 , \19898 );
not \U$19654 ( \19900 , \19899 );
not \U$19655 ( \19901 , \19900 );
or \U$19656 ( \19902 , \19844 , \19901 );
or \U$19657 ( \19903 , \19900 , \19843 );
nand \U$19658 ( \19904 , \19902 , \19903 );
not \U$19659 ( \19905 , \19904 );
or \U$19660 ( \19906 , \19770 , \19905 );
nand \U$19661 ( \19907 , \19899 , \19843 );
nand \U$19662 ( \19908 , \19906 , \19907 );
not \U$19663 ( \19909 , \19908 );
or \U$19664 ( \19910 , \19690 , \19909 );
not \U$19665 ( \19911 , \19688 );
nand \U$19666 ( \19912 , \19911 , \19680 );
nand \U$19667 ( \19913 , \19910 , \19912 );
xor \U$19668 ( \19914 , \17535 , \17557 );
xnor \U$19669 ( \19915 , \19914 , \17584 );
xor \U$19670 ( \19916 , \17596 , \17602 );
xor \U$19671 ( \19917 , \19916 , \17609 );
not \U$19672 ( \19918 , \17960 );
xnor \U$19673 ( \19919 , \17966 , \19918 );
xor \U$19674 ( \19920 , \19917 , \19919 );
not \U$19675 ( \19921 , \17650 );
nand \U$19676 ( \19922 , \19921 , \17659 );
and \U$19677 ( \19923 , \19922 , \17656 );
not \U$19678 ( \19924 , \19922 );
and \U$19679 ( \19925 , \19924 , \17657 );
nor \U$19680 ( \19926 , \19923 , \19925 );
xnor \U$19681 ( \19927 , \19920 , \19926 );
xor \U$19682 ( \19928 , \19915 , \19927 );
xor \U$19683 ( \19929 , \18201 , \18193 );
xor \U$19684 ( \19930 , \19929 , \18186 );
xor \U$19685 ( \19931 , \17927 , \17932 );
xnor \U$19686 ( \19932 , \19931 , \17939 );
xor \U$19687 ( \19933 , \17988 , \17983 );
xnor \U$19688 ( \19934 , \19933 , \17978 );
xnor \U$19689 ( \19935 , \19932 , \19934 );
xor \U$19690 ( \19936 , \19930 , \19935 );
xor \U$19691 ( \19937 , \19928 , \19936 );
and \U$19692 ( \19938 , \19913 , \19937 );
not \U$19693 ( \19939 , \19913 );
not \U$19694 ( \19940 , \19937 );
and \U$19695 ( \19941 , \19939 , \19940 );
nor \U$19696 ( \19942 , \19938 , \19941 );
xor \U$19697 ( \19943 , \17829 , \17822 );
xor \U$19698 ( \19944 , \19943 , \17838 );
not \U$19699 ( \19945 , \19355 );
not \U$19700 ( \19946 , \19332 );
or \U$19701 ( \19947 , \19945 , \19946 );
not \U$19702 ( \19948 , \19328 );
nand \U$19703 ( \19949 , \19948 , \19313 );
nand \U$19704 ( \19950 , \19947 , \19949 );
xor \U$19705 ( \19951 , \19944 , \19950 );
xor \U$19706 ( \19952 , \19711 , \19733 );
and \U$19707 ( \19953 , \19952 , \19768 );
and \U$19708 ( \19954 , \19711 , \19733 );
or \U$19709 ( \19955 , \19953 , \19954 );
and \U$19710 ( \19956 , \19951 , \19955 );
not \U$19711 ( \19957 , \19951 );
not \U$19712 ( \19958 , \19955 );
and \U$19713 ( \19959 , \19957 , \19958 );
nor \U$19714 ( \19960 , \19956 , \19959 );
not \U$19715 ( \19961 , \19960 );
not \U$19716 ( \19962 , \19324 );
nand \U$19717 ( \19963 , \19962 , \19319 );
not \U$19718 ( \19964 , \19963 );
not \U$19719 ( \19965 , \19259 );
or \U$19720 ( \19966 , \13540 , \19965 );
not \U$19721 ( \19967 , \13533 );
not \U$19722 ( \19968 , \19487 );
or \U$19723 ( \19969 , \19967 , \19968 );
nand \U$19724 ( \19970 , \19966 , \19969 );
not \U$19725 ( \19971 , \19234 );
not \U$19726 ( \19972 , \17592 );
or \U$19727 ( \19973 , \19971 , \19972 );
nand \U$19728 ( \19974 , \14966 , \19467 );
nand \U$19729 ( \19975 , \19973 , \19974 );
or \U$19730 ( \19976 , \19970 , \19975 );
not \U$19731 ( \19977 , \19814 );
not \U$19732 ( \19978 , \4841 );
not \U$19733 ( \19979 , \19978 );
or \U$19734 ( \19980 , \19977 , \19979 );
nand \U$19735 ( \19981 , \16655 , \19461 );
nand \U$19736 ( \19982 , \19980 , \19981 );
nand \U$19737 ( \19983 , \19976 , \19982 );
nand \U$19738 ( \19984 , \19970 , \19975 );
nand \U$19739 ( \19985 , \19983 , \19984 );
not \U$19740 ( \19986 , \19985 );
or \U$19741 ( \19987 , \19964 , \19986 );
or \U$19742 ( \19988 , \19963 , \19985 );
nand \U$19743 ( \19989 , \19987 , \19988 );
buf \U$19744 ( \19990 , \19989 );
not \U$19745 ( \19991 , \19706 );
not \U$19746 ( \19992 , \879 );
or \U$19747 ( \19993 , \19991 , \19992 );
nand \U$19748 ( \19994 , \885 , \19494 );
nand \U$19749 ( \19995 , \19993 , \19994 );
not \U$19750 ( \19996 , \19288 );
not \U$19751 ( \19997 , \4893 );
or \U$19752 ( \19998 , \19996 , \19997 );
nand \U$19753 ( \19999 , \2707 , \19481 );
nand \U$19754 ( \20000 , \19998 , \19999 );
nor \U$19755 ( \20001 , \19995 , \20000 );
not \U$19756 ( \20002 , \2670 );
not \U$19757 ( \20003 , \17870 );
not \U$19758 ( \20004 , \20003 );
and \U$19759 ( \20005 , \20002 , \20004 );
not \U$19760 ( \20006 , \19240 );
and \U$19761 ( \20007 , \3485 , \20006 );
nor \U$19762 ( \20008 , \20005 , \20007 );
or \U$19763 ( \20009 , \20001 , \20008 );
nand \U$19764 ( \20010 , \19995 , \20000 );
nand \U$19765 ( \20011 , \20009 , \20010 );
buf \U$19766 ( \20012 , \20011 );
not \U$19767 ( \20013 , \20012 );
and \U$19768 ( \20014 , \19990 , \20013 );
not \U$19769 ( \20015 , \19990 );
and \U$19770 ( \20016 , \20015 , \20012 );
nor \U$19771 ( \20017 , \20014 , \20016 );
not \U$19772 ( \20018 , \20017 );
or \U$19773 ( \20019 , \19894 , \19882 );
nand \U$19774 ( \20020 , \20019 , \19887 );
nand \U$19775 ( \20021 , \19894 , \19882 );
nand \U$19776 ( \20022 , \20020 , \20021 );
or \U$19777 ( \20023 , \19865 , \19859 );
nand \U$19778 ( \20024 , \20023 , \19871 );
nand \U$19779 ( \20025 , \19865 , \19859 );
and \U$19780 ( \20026 , \20024 , \20025 );
xnor \U$19781 ( \20027 , \20022 , \20026 );
not \U$19782 ( \20028 , \20027 );
not \U$19783 ( \20029 , \19277 );
not \U$19784 ( \20030 , \19295 );
or \U$19785 ( \20031 , \20029 , \20030 );
nand \U$19786 ( \20032 , \19290 , \19283 );
nand \U$19787 ( \20033 , \20031 , \20032 );
not \U$19788 ( \20034 , \20033 );
or \U$19789 ( \20035 , \20028 , \20034 );
not \U$19790 ( \20036 , \20026 );
nand \U$19791 ( \20037 , \20036 , \20022 );
nand \U$19792 ( \20038 , \20035 , \20037 );
not \U$19793 ( \20039 , \19808 );
not \U$19794 ( \20040 , \19805 );
or \U$19795 ( \20041 , \20039 , \20040 );
nand \U$19796 ( \20042 , \20041 , \19837 );
nand \U$19797 ( \20043 , \19804 , \19776 );
nand \U$19798 ( \20044 , \20042 , \20043 );
xor \U$19799 ( \20045 , \20038 , \20044 );
not \U$19800 ( \20046 , \20045 );
or \U$19801 ( \20047 , \20018 , \20046 );
or \U$19802 ( \20048 , \20045 , \20017 );
nand \U$19803 ( \20049 , \20047 , \20048 );
not \U$19804 ( \20050 , \20049 );
xor \U$19805 ( \20051 , \19717 , \19724 );
xor \U$19806 ( \20052 , \20051 , \19730 );
xor \U$19807 ( \20053 , \19695 , \19701 );
xor \U$19808 ( \20054 , \20053 , \19708 );
xor \U$19809 ( \20055 , \20052 , \20054 );
not \U$19810 ( \20056 , \19763 );
not \U$19811 ( \20057 , \19741 );
or \U$19812 ( \20058 , \20056 , \20057 );
or \U$19813 ( \20059 , \19763 , \19741 );
nand \U$19814 ( \20060 , \20058 , \20059 );
and \U$19815 ( \20061 , \20055 , \20060 );
and \U$19816 ( \20062 , \20052 , \20054 );
or \U$19817 ( \20063 , \20061 , \20062 );
not \U$19818 ( \20064 , \20063 );
not \U$19819 ( \20065 , \19782 );
not \U$19820 ( \20066 , \19792 );
or \U$19821 ( \20067 , \20065 , \20066 );
nand \U$19822 ( \20068 , \19794 , \19789 );
nand \U$19823 ( \20069 , \20067 , \20068 );
not \U$19824 ( \20070 , \19802 );
and \U$19825 ( \20071 , \20069 , \20070 );
not \U$19826 ( \20072 , \20069 );
and \U$19827 ( \20073 , \20072 , \19802 );
nor \U$19828 ( \20074 , \20071 , \20073 );
not \U$19829 ( \20075 , \20074 );
not \U$19830 ( \20076 , \19095 );
not \U$19831 ( \20077 , \1043 );
or \U$19832 ( \20078 , \20076 , \20077 );
nand \U$19833 ( \20079 , \314 , \19797 );
nand \U$19834 ( \20080 , \20078 , \20079 );
not \U$19835 ( \20081 , \20080 );
not \U$19836 ( \20082 , \19047 );
not \U$19837 ( \20083 , \9052 );
or \U$19838 ( \20084 , \20082 , \20083 );
nand \U$19839 ( \20085 , \2559 , \19752 );
nand \U$19840 ( \20086 , \20084 , \20085 );
not \U$19841 ( \20087 , \20086 );
or \U$19842 ( \20088 , \20081 , \20087 );
or \U$19843 ( \20089 , \20086 , \20080 );
not \U$19844 ( \20090 , \19024 );
not \U$19845 ( \20091 , \11453 );
or \U$19846 ( \20092 , \20090 , \20091 );
nand \U$19847 ( \20093 , \10401 , \19744 );
nand \U$19848 ( \20094 , \20092 , \20093 );
nand \U$19849 ( \20095 , \20089 , \20094 );
nand \U$19850 ( \20096 , \20088 , \20095 );
or \U$19851 ( \20097 , \20075 , \20096 );
xor \U$19852 ( \20098 , \19338 , \19351 );
nand \U$19853 ( \20099 , \20097 , \20098 );
nand \U$19854 ( \20100 , \20075 , \20096 );
nand \U$19855 ( \20101 , \20099 , \20100 );
not \U$19856 ( \20102 , \20101 );
xnor \U$19857 ( \20103 , \20027 , \20033 );
nand \U$19858 ( \20104 , \20102 , \20103 );
not \U$19859 ( \20105 , \20104 );
or \U$19860 ( \20106 , \20064 , \20105 );
not \U$19861 ( \20107 , \20103 );
buf \U$19862 ( \20108 , \20101 );
nand \U$19863 ( \20109 , \20107 , \20108 );
nand \U$19864 ( \20110 , \20106 , \20109 );
not \U$19865 ( \20111 , \20110 );
not \U$19866 ( \20112 , \20111 );
or \U$19867 ( \20113 , \20050 , \20112 );
or \U$19868 ( \20114 , \20049 , \20111 );
nand \U$19869 ( \20115 , \20113 , \20114 );
not \U$19870 ( \20116 , \20115 );
or \U$19871 ( \20117 , \19961 , \20116 );
not \U$19872 ( \20118 , \20111 );
buf \U$19873 ( \20119 , \20049 );
nand \U$19874 ( \20120 , \20118 , \20119 );
nand \U$19875 ( \20121 , \20117 , \20120 );
buf \U$19876 ( \20122 , \20121 );
xor \U$19877 ( \20123 , \19942 , \20122 );
not \U$19878 ( \20124 , \20123 );
and \U$19879 ( \20125 , \19676 , \20124 );
and \U$19880 ( \20126 , \19675 , \20123 );
nor \U$19881 ( \20127 , \20125 , \20126 );
not \U$19882 ( \20128 , \19863 );
not \U$19883 ( \20129 , \15764 );
or \U$19884 ( \20130 , \20128 , \20129 );
nand \U$19885 ( \20131 , \11400 , \17707 );
nand \U$19886 ( \20132 , \20130 , \20131 );
not \U$19887 ( \20133 , \19266 );
not \U$19888 ( \20134 , \965 );
or \U$19889 ( \20135 , \20133 , \20134 );
nand \U$19890 ( \20136 , \1199 , \17737 );
nand \U$19891 ( \20137 , \20135 , \20136 );
xor \U$19892 ( \20138 , \20132 , \20137 );
not \U$19893 ( \20139 , \19275 );
not \U$19894 ( \20140 , \16715 );
or \U$19895 ( \20141 , \20139 , \20140 );
nand \U$19896 ( \20142 , \11094 , \17726 );
nand \U$19897 ( \20143 , \20141 , \20142 );
xor \U$19898 ( \20144 , \20138 , \20143 );
not \U$19899 ( \20145 , \19343 );
not \U$19900 ( \20146 , \1103 );
or \U$19901 ( \20147 , \20145 , \20146 );
nand \U$19902 ( \20148 , \369 , \19529 );
nand \U$19903 ( \20149 , \20147 , \20148 );
not \U$19904 ( \20150 , \19787 );
not \U$19905 ( \20151 , \9194 );
or \U$19906 ( \20152 , \20150 , \20151 );
nand \U$19907 ( \20153 , \1769 , \17783 );
nand \U$19908 ( \20154 , \20152 , \20153 );
xor \U$19909 ( \20155 , \20149 , \20154 );
not \U$19910 ( \20156 , \19748 );
not \U$19911 ( \20157 , \10987 );
or \U$19912 ( \20158 , \20156 , \20157 );
nand \U$19913 ( \20159 , \9726 , \17769 );
nand \U$19914 ( \20160 , \20158 , \20159 );
xor \U$19915 ( \20161 , \20155 , \20160 );
xor \U$19916 ( \20162 , \20144 , \20161 );
xor \U$19917 ( \20163 , \19611 , \19603 );
and \U$19918 ( \20164 , \20163 , \19620 );
not \U$19919 ( \20165 , \20163 );
not \U$19920 ( \20166 , \19620 );
and \U$19921 ( \20167 , \20165 , \20166 );
nor \U$19922 ( \20168 , \20164 , \20167 );
xor \U$19923 ( \20169 , \20162 , \20168 );
not \U$19924 ( \20170 , \20169 );
not \U$19925 ( \20171 , \19892 );
not \U$19926 ( \20172 , \10674 );
or \U$19927 ( \20173 , \20171 , \20172 );
nand \U$19928 ( \20174 , \8930 , \19428 );
nand \U$19929 ( \20175 , \20173 , \20174 );
xor \U$19930 ( \20176 , RIbe27b98_2, RIbe2ae38_110);
not \U$19931 ( \20177 , \20176 );
not \U$19932 ( \20178 , \256 );
or \U$19933 ( \20179 , \20177 , \20178 );
nand \U$19934 ( \20180 , \267 , \19421 );
nand \U$19935 ( \20181 , \20179 , \20180 );
not \U$19936 ( \20182 , \20181 );
xor \U$19937 ( \20183 , \20175 , \20182 );
not \U$19938 ( \20184 , \19739 );
not \U$19939 ( \20185 , \1452 );
or \U$19940 ( \20186 , \20184 , \20185 );
nand \U$19941 ( \20187 , \907 , \19474 );
nand \U$19942 ( \20188 , \20186 , \20187 );
and \U$19943 ( \20189 , \20183 , \20188 );
not \U$19944 ( \20190 , \20183 );
not \U$19945 ( \20191 , \20188 );
and \U$19946 ( \20192 , \20190 , \20191 );
nor \U$19947 ( \20193 , \20189 , \20192 );
not \U$19948 ( \20194 , \20193 );
xor \U$19949 ( \20195 , \19585 , \19592 );
xnor \U$19950 ( \20196 , \20195 , \19575 );
not \U$19951 ( \20197 , \20196 );
nand \U$19952 ( \20198 , \20194 , \20197 );
nand \U$19953 ( \20199 , \20193 , \20196 );
nand \U$19954 ( \20200 , \20198 , \20199 );
not \U$19955 ( \20201 , \19756 );
not \U$19956 ( \20202 , \3402 );
or \U$19957 ( \20203 , \20201 , \20202 );
nand \U$19958 ( \20204 , \2691 , \17817 );
nand \U$19959 ( \20205 , \20203 , \20204 );
not \U$19960 ( \20206 , \19336 );
not \U$19961 ( \20207 , \2890 );
or \U$19962 ( \20208 , \20206 , \20207 );
nand \U$19963 ( \20209 , \8270 , \19440 );
nand \U$19964 ( \20210 , \20208 , \20209 );
not \U$19965 ( \20211 , \20210 );
not \U$19966 ( \20212 , \20211 );
not \U$19967 ( \20213 , \19699 );
not \U$19968 ( \20214 , \12721 );
or \U$19969 ( \20215 , \20213 , \20214 );
nand \U$19970 ( \20216 , \9524 , \17833 );
nand \U$19971 ( \20217 , \20215 , \20216 );
not \U$19972 ( \20218 , \20217 );
or \U$19973 ( \20219 , \20212 , \20218 );
or \U$19974 ( \20220 , \20217 , \20211 );
nand \U$19975 ( \20221 , \20219 , \20220 );
xor \U$19976 ( \20222 , \20205 , \20221 );
and \U$19977 ( \20223 , \20200 , \20222 );
not \U$19978 ( \20224 , \20200 );
not \U$19979 ( \20225 , \20222 );
and \U$19980 ( \20226 , \20224 , \20225 );
nor \U$19981 ( \20227 , \20223 , \20226 );
not \U$19982 ( \20228 , \20227 );
or \U$19983 ( \20229 , \20170 , \20228 );
or \U$19984 ( \20230 , \20227 , \20169 );
nand \U$19985 ( \20231 , \20229 , \20230 );
not \U$19986 ( \20232 , \20001 );
nand \U$19987 ( \20233 , \20232 , \20010 );
xor \U$19988 ( \20234 , \20233 , \20008 );
not \U$19989 ( \20235 , \20234 );
not \U$19990 ( \20236 , \19253 );
not \U$19991 ( \20237 , \11344 );
not \U$19992 ( \20238 , \20237 );
or \U$19993 ( \20239 , \20236 , \20238 );
nand \U$19994 ( \20240 , \11348 , \17849 );
nand \U$19995 ( \20241 , \20239 , \20240 );
not \U$19996 ( \20242 , \19722 );
not \U$19997 ( \20243 , \15345 );
or \U$19998 ( \20244 , \20242 , \20243 );
nand \U$19999 ( \20245 , \19721 , \17824 );
nand \U$20000 ( \20246 , \20244 , \20245 );
xor \U$20001 ( \20247 , \20241 , \20246 );
not \U$20002 ( \20248 , \19715 );
not \U$20003 ( \20249 , \8595 );
or \U$20004 ( \20250 , \20248 , \20249 );
nand \U$20005 ( \20251 , \7642 , \17842 );
nand \U$20006 ( \20252 , \20250 , \20251 );
not \U$20007 ( \20253 , \20252 );
and \U$20008 ( \20254 , \20247 , \20253 );
not \U$20009 ( \20255 , \20247 );
and \U$20010 ( \20256 , \20255 , \20252 );
nor \U$20011 ( \20257 , \20254 , \20256 );
not \U$20012 ( \20258 , \19970 );
xor \U$20013 ( \20259 , \20258 , \19982 );
and \U$20014 ( \20260 , \20259 , \19975 );
not \U$20015 ( \20261 , \20259 );
not \U$20016 ( \20262 , \19975 );
and \U$20017 ( \20263 , \20261 , \20262 );
nor \U$20018 ( \20264 , \20260 , \20263 );
nand \U$20019 ( \20265 , \20257 , \20264 );
or \U$20020 ( \20266 , \20257 , \20264 );
nand \U$20021 ( \20267 , \20265 , \20266 );
not \U$20022 ( \20268 , \20267 );
or \U$20023 ( \20269 , \20235 , \20268 );
or \U$20024 ( \20270 , \20267 , \20234 );
nand \U$20025 ( \20271 , \20269 , \20270 );
and \U$20026 ( \20272 , \20231 , \20271 );
not \U$20027 ( \20273 , \20231 );
not \U$20028 ( \20274 , \20271 );
and \U$20029 ( \20275 , \20273 , \20274 );
nor \U$20030 ( \20276 , \20272 , \20275 );
xor \U$20031 ( \20277 , \19226 , \19402 );
xor \U$20032 ( \20278 , \20276 , \20277 );
xor \U$20033 ( \20279 , RIbe280c0_13, RIbe2b4c8_124);
not \U$20034 ( \20280 , \20279 );
not \U$20035 ( \20281 , \8551 );
or \U$20036 ( \20282 , \20280 , \20281 );
nand \U$20037 ( \20283 , \869 , \18933 );
nand \U$20038 ( \20284 , \20282 , \20283 );
xor \U$20039 ( \20285 , RIbe2af28_112, RIbe28c78_38);
not \U$20040 ( \20286 , \20285 );
not \U$20041 ( \20287 , \14423 );
or \U$20042 ( \20288 , \20286 , \20287 );
nand \U$20043 ( \20289 , \17810 , \18917 );
nand \U$20044 ( \20290 , \20288 , \20289 );
xor \U$20045 ( \20291 , \20284 , \20290 );
xor \U$20046 ( \20292 , RIbe28390_19, RIbe2a820_97);
not \U$20047 ( \20293 , \20292 );
not \U$20048 ( \20294 , \14579 );
or \U$20049 ( \20295 , \20293 , \20294 );
nand \U$20050 ( \20296 , \3714 , \19160 );
nand \U$20051 ( \20297 , \20295 , \20296 );
and \U$20052 ( \20298 , \20291 , \20297 );
and \U$20053 ( \20299 , \20284 , \20290 );
or \U$20054 ( \20300 , \20298 , \20299 );
not \U$20055 ( \20301 , \20300 );
xor \U$20056 ( \20302 , RIbe296c8_60, RIbe2a640_93);
not \U$20057 ( \20303 , \20302 );
not \U$20058 ( \20304 , \9793 );
or \U$20059 ( \20305 , \20303 , \20304 );
nand \U$20060 ( \20306 , \1937 , \19190 );
nand \U$20061 ( \20307 , \20305 , \20306 );
not \U$20062 ( \20308 , \20307 );
xor \U$20063 ( \20309 , RIbe2a028_80, RIbe27df0_7);
not \U$20064 ( \20310 , \20309 );
not \U$20065 ( \20311 , \8168 );
or \U$20066 ( \20312 , \20310 , \20311 );
nand \U$20067 ( \20313 , \8171 , \19101 );
nand \U$20068 ( \20314 , \20312 , \20313 );
not \U$20069 ( \20315 , \20314 );
or \U$20070 ( \20316 , \20308 , \20315 );
or \U$20071 ( \20317 , \20314 , \20307 );
xor \U$20072 ( \20318 , RIbe28480_21, RIbe2aa00_101);
not \U$20073 ( \20319 , \20318 );
not \U$20074 ( \20320 , \2518 );
or \U$20075 ( \20321 , \20319 , \20320 );
nand \U$20076 ( \20322 , \7483 , \19114 );
nand \U$20077 ( \20323 , \20321 , \20322 );
nand \U$20078 ( \20324 , \20317 , \20323 );
nand \U$20079 ( \20325 , \20316 , \20324 );
xor \U$20080 ( \20326 , RIbe295d8_58, RIbe2a910_99);
not \U$20081 ( \20327 , \20326 );
not \U$20082 ( \20328 , \9737 );
or \U$20083 ( \20329 , \20327 , \20328 );
nand \U$20084 ( \20330 , \9726 , \19020 );
nand \U$20085 ( \20331 , \20329 , \20330 );
xor \U$20086 ( \20332 , RIbe297b8_62, RIbe2a550_91);
not \U$20087 ( \20333 , \20332 );
not \U$20088 ( \20334 , \10433 );
or \U$20089 ( \20335 , \20333 , \20334 );
not \U$20090 ( \20336 , \10439 );
nand \U$20091 ( \20337 , \20336 , \19168 );
nand \U$20092 ( \20338 , \20335 , \20337 );
or \U$20093 ( \20339 , \20331 , \20338 );
xor \U$20094 ( \20340 , RIbe28930_31, RIbe2a460_89);
not \U$20095 ( \20341 , \20340 );
not \U$20096 ( \20342 , \965 );
or \U$20097 ( \20343 , \20341 , \20342 );
nand \U$20098 ( \20344 , \1199 , \19153 );
nand \U$20099 ( \20345 , \20343 , \20344 );
nand \U$20100 ( \20346 , \20339 , \20345 );
nand \U$20101 ( \20347 , \20331 , \20338 );
nand \U$20102 ( \20348 , \20346 , \20347 );
xor \U$20103 ( \20349 , \20325 , \20348 );
not \U$20104 ( \20350 , \20349 );
or \U$20105 ( \20351 , \20301 , \20350 );
nand \U$20106 ( \20352 , \20348 , \20325 );
nand \U$20107 ( \20353 , \20351 , \20352 );
not \U$20108 ( \20354 , \20353 );
xor \U$20109 ( \20355 , RIbe28a20_33, RIbe2b2e8_120);
not \U$20110 ( \20356 , \20355 );
not \U$20111 ( \20357 , \1780 );
or \U$20112 ( \20358 , \20356 , \20357 );
nand \U$20113 ( \20359 , \2475 , \19134 );
nand \U$20114 ( \20360 , \20358 , \20359 );
not \U$20115 ( \20361 , \20360 );
xor \U$20116 ( \20362 , RIbe2b108_116, RIbe28a98_34);
not \U$20117 ( \20363 , \20362 );
not \U$20118 ( \20364 , \14297 );
or \U$20119 ( \20365 , \20363 , \20364 );
nand \U$20120 ( \20366 , \13533 , \19107 );
nand \U$20121 ( \20367 , \20365 , \20366 );
not \U$20122 ( \20368 , \20367 );
or \U$20123 ( \20369 , \20361 , \20368 );
or \U$20124 ( \20370 , \20367 , \20360 );
xor \U$20125 ( \20371 , RIbe2ad48_108, RIbe28228_16);
not \U$20126 ( \20372 , \20371 );
not \U$20127 ( \20373 , \3056 );
or \U$20128 ( \20374 , \20372 , \20373 );
nand \U$20129 ( \20375 , \8680 , \19142 );
nand \U$20130 ( \20376 , \20374 , \20375 );
nand \U$20131 ( \20377 , \20370 , \20376 );
nand \U$20132 ( \20378 , \20369 , \20377 );
not \U$20133 ( \20379 , \20378 );
xor \U$20134 ( \20380 , RIbe27d78_6, RIbe2b3d8_122);
not \U$20135 ( \20381 , \20380 );
not \U$20136 ( \20382 , \8898 );
or \U$20137 ( \20383 , \20381 , \20382 );
nand \U$20138 ( \20384 , \10752 , \19091 );
nand \U$20139 ( \20385 , \20383 , \20384 );
not \U$20140 ( \20386 , \20385 );
or \U$20141 ( \20387 , RIbe27d00_5, RIbe27d78_6);
nand \U$20142 ( \20388 , \20387 , RIbe2ae38_110);
nand \U$20143 ( \20389 , RIbe27d00_5, RIbe27d78_6);
nand \U$20144 ( \20390 , \20388 , \20389 , RIbe27c10_3);
nor \U$20145 ( \20391 , \20386 , \20390 );
not \U$20146 ( \20392 , \20391 );
xor \U$20147 ( \20393 , RIbe2b018_114, RIbe28750_27);
not \U$20148 ( \20394 , \20393 );
not \U$20149 ( \20395 , \15966 );
buf \U$20150 ( \20396 , \20395 );
not \U$20151 ( \20397 , \20396 );
or \U$20152 ( \20398 , \20394 , \20397 );
nand \U$20153 ( \20399 , \19371 , \18773 );
nand \U$20154 ( \20400 , \20398 , \20399 );
not \U$20155 ( \20401 , \20400 );
not \U$20156 ( \20402 , \20401 );
or \U$20157 ( \20403 , \20392 , \20402 );
or \U$20158 ( \20404 , \20391 , \20401 );
nand \U$20159 ( \20405 , \20403 , \20404 );
not \U$20160 ( \20406 , \20405 );
or \U$20161 ( \20407 , \20379 , \20406 );
not \U$20162 ( \20408 , \20401 );
nand \U$20163 ( \20409 , \20408 , \20391 );
nand \U$20164 ( \20410 , \20407 , \20409 );
xor \U$20165 ( \20411 , RIbe29ec0_77, RIbe27e68_8);
not \U$20166 ( \20412 , \20411 );
not \U$20167 ( \20413 , \2599 );
or \U$20168 ( \20414 , \20412 , \20413 );
nand \U$20169 ( \20415 , \2603 , \19082 );
nand \U$20170 ( \20416 , \20414 , \20415 );
not \U$20171 ( \20417 , \20416 );
xor \U$20172 ( \20418 , RIbe282a0_17, RIbe2a190_83);
not \U$20173 ( \20419 , \20418 );
not \U$20174 ( \20420 , \10831 );
or \U$20175 ( \20421 , \20419 , \20420 );
nand \U$20176 ( \20422 , \11399 , \18996 );
nand \U$20177 ( \20423 , \20421 , \20422 );
not \U$20178 ( \20424 , \20423 );
not \U$20179 ( \20425 , \20424 );
and \U$20180 ( \20426 , RIbe2a3e8_88, \5592 );
not \U$20181 ( \20427 , RIbe2a3e8_88);
and \U$20182 ( \20428 , \20427 , RIbe29128_48);
or \U$20183 ( \20429 , \20426 , \20428 );
not \U$20184 ( \20430 , \20429 );
not \U$20185 ( \20431 , \8805 );
or \U$20186 ( \20432 , \20430 , \20431 );
nand \U$20187 ( \20433 , \9089 , \19004 );
nand \U$20188 ( \20434 , \20432 , \20433 );
not \U$20189 ( \20435 , \20434 );
or \U$20190 ( \20436 , \20425 , \20435 );
or \U$20191 ( \20437 , \20424 , \20434 );
nand \U$20192 ( \20438 , \20436 , \20437 );
not \U$20193 ( \20439 , \20438 );
or \U$20194 ( \20440 , \20417 , \20439 );
nand \U$20195 ( \20441 , \20423 , \20434 );
nand \U$20196 ( \20442 , \20440 , \20441 );
not \U$20197 ( \20443 , \20442 );
xor \U$20198 ( \20444 , RIbe27c10_3, RIbe2ae38_110);
not \U$20199 ( \20445 , \20444 );
not \U$20200 ( \20446 , \11907 );
or \U$20201 ( \20447 , \20445 , \20446 );
nand \U$20202 ( \20448 , \1173 , \18989 );
nand \U$20203 ( \20449 , \20447 , \20448 );
xor \U$20204 ( \20450 , RIbe298a8_64, RIbe29c68_72);
not \U$20205 ( \20451 , \20450 );
not \U$20206 ( \20452 , \14971 );
or \U$20207 ( \20453 , \20451 , \20452 );
nand \U$20208 ( \20454 , \4580 , \19051 );
nand \U$20209 ( \20455 , \20453 , \20454 );
or \U$20210 ( \20456 , \20449 , \20455 );
xor \U$20211 ( \20457 , RIbe29038_46, RIbe2abe0_105);
not \U$20212 ( \20458 , \20457 );
not \U$20213 ( \20459 , \281 );
or \U$20214 ( \20460 , \20458 , \20459 );
nand \U$20215 ( \20461 , \287 , \19037 );
nand \U$20216 ( \20462 , \20460 , \20461 );
nand \U$20217 ( \20463 , \20456 , \20462 );
nand \U$20218 ( \20464 , \20449 , \20455 );
nand \U$20219 ( \20465 , \20443 , \20463 , \20464 );
xor \U$20220 ( \20466 , RIbe290b0_47, RIbe2a730_95);
not \U$20221 ( \20467 , \20466 );
not \U$20222 ( \20468 , \2729 );
or \U$20223 ( \20469 , \20467 , \20468 );
nand \U$20224 ( \20470 , \398 , \19014 );
nand \U$20225 ( \20471 , \20469 , \20470 );
xor \U$20226 ( \20472 , RIbe27b20_1, RIbe28f48_44);
not \U$20227 ( \20473 , \20472 );
not \U$20228 ( \20474 , \12721 );
or \U$20229 ( \20475 , \20473 , \20474 );
nand \U$20230 ( \20476 , \11201 , \19028 );
nand \U$20231 ( \20477 , \20475 , \20476 );
xor \U$20232 ( \20478 , \20471 , \20477 );
xor \U$20233 ( \20479 , RIbe28b88_36, RIbe2a0a0_81);
not \U$20234 ( \20480 , \20479 );
not \U$20235 ( \20481 , \9052 );
or \U$20236 ( \20482 , \20480 , \20481 );
nand \U$20237 ( \20483 , \2559 , \19043 );
nand \U$20238 ( \20484 , \20482 , \20483 );
and \U$20239 ( \20485 , \20478 , \20484 );
and \U$20240 ( \20486 , \20471 , \20477 );
or \U$20241 ( \20487 , \20485 , \20486 );
nand \U$20242 ( \20488 , \20465 , \20487 );
nand \U$20243 ( \20489 , \20463 , \20464 );
buf \U$20244 ( \20490 , \20442 );
nand \U$20245 ( \20491 , \20489 , \20490 );
nand \U$20246 ( \20492 , \20488 , \20491 );
and \U$20247 ( \20493 , \20410 , \20492 );
not \U$20248 ( \20494 , \20410 );
and \U$20249 ( \20495 , \20491 , \20488 );
and \U$20250 ( \20496 , \20494 , \20495 );
nor \U$20251 ( \20497 , \20493 , \20496 );
not \U$20252 ( \20498 , \20497 );
or \U$20253 ( \20499 , \20354 , \20498 );
nand \U$20254 ( \20500 , \20492 , \20410 );
nand \U$20255 ( \20501 , \20499 , \20500 );
not \U$20256 ( \20502 , \20501 );
xor \U$20257 ( \20503 , \20052 , \20054 );
xor \U$20258 ( \20504 , \20503 , \20060 );
not \U$20259 ( \20505 , \19301 );
not \U$20260 ( \20506 , \19247 );
and \U$20261 ( \20507 , \20505 , \20506 );
and \U$20262 ( \20508 , \19301 , \19247 );
nor \U$20263 ( \20509 , \20507 , \20508 );
not \U$20264 ( \20510 , \20509 );
xor \U$20265 ( \20511 , \20504 , \20510 );
not \U$20266 ( \20512 , \20511 );
or \U$20267 ( \20513 , \20502 , \20512 );
not \U$20268 ( \20514 , \20509 );
and \U$20269 ( \20515 , \20504 , \20514 );
not \U$20270 ( \20516 , \20515 );
nand \U$20271 ( \20517 , \20513 , \20516 );
xor \U$20272 ( \20518 , \20278 , \20517 );
not \U$20273 ( \20519 , \20518 );
not \U$20274 ( \20520 , \20108 );
not \U$20275 ( \20521 , \20103 );
and \U$20276 ( \20522 , \20520 , \20521 );
and \U$20277 ( \20523 , \20103 , \20108 );
nor \U$20278 ( \20524 , \20522 , \20523 );
xnor \U$20279 ( \20525 , \20063 , \20524 );
and \U$20280 ( \20526 , \20096 , \20074 );
not \U$20281 ( \20527 , \20096 );
and \U$20282 ( \20528 , \20527 , \20075 );
or \U$20283 ( \20529 , \20526 , \20528 );
and \U$20284 ( \20530 , \20529 , \20098 );
not \U$20285 ( \20531 , \20529 );
not \U$20286 ( \20532 , \20098 );
and \U$20287 ( \20533 , \20531 , \20532 );
nor \U$20288 ( \20534 , \20530 , \20533 );
not \U$20289 ( \20535 , \20534 );
xor \U$20290 ( \20536 , \18610 , \18617 );
xor \U$20291 ( \20537 , \20536 , \18625 );
not \U$20292 ( \20538 , \20537 );
xor \U$20293 ( \20539 , \20080 , \20086 );
xnor \U$20294 ( \20540 , \20539 , \20094 );
not \U$20295 ( \20541 , \20540 );
not \U$20296 ( \20542 , \20541 );
or \U$20297 ( \20543 , \20538 , \20542 );
or \U$20298 ( \20544 , \20541 , \20537 );
xor \U$20299 ( \20545 , \18678 , \18670 );
not \U$20300 ( \20546 , \18688 );
and \U$20301 ( \20547 , \20545 , \20546 );
not \U$20302 ( \20548 , \20545 );
and \U$20303 ( \20549 , \20548 , \18688 );
nor \U$20304 ( \20550 , \20547 , \20549 );
not \U$20305 ( \20551 , \20550 );
nand \U$20306 ( \20552 , \20544 , \20551 );
nand \U$20307 ( \20553 , \20543 , \20552 );
xor \U$20308 ( \20554 , \19876 , \19895 );
xnor \U$20309 ( \20555 , \20554 , \19851 );
and \U$20310 ( \20556 , \20553 , \20555 );
not \U$20311 ( \20557 , \20553 );
not \U$20312 ( \20558 , \20555 );
and \U$20313 ( \20559 , \20557 , \20558 );
nor \U$20314 ( \20560 , \20556 , \20559 );
not \U$20315 ( \20561 , \20560 );
or \U$20316 ( \20562 , \20535 , \20561 );
not \U$20317 ( \20563 , \20558 );
nand \U$20318 ( \20564 , \20563 , \20553 );
nand \U$20319 ( \20565 , \20562 , \20564 );
not \U$20320 ( \20566 , \20565 );
xor \U$20321 ( \20567 , \20525 , \20566 );
xor \U$20322 ( \20568 , \19842 , \19769 );
xnor \U$20323 ( \20569 , \20568 , \19900 );
xnor \U$20324 ( \20570 , \20567 , \20569 );
not \U$20325 ( \20571 , \20570 );
xor \U$20326 ( \20572 , RIbe2aaf0_103, RIbe28840_29);
not \U$20327 ( \20573 , \20572 );
not \U$20328 ( \20574 , \19580 );
not \U$20329 ( \20575 , \20574 );
or \U$20330 ( \20576 , \20573 , \20575 );
nand \U$20331 ( \20577 , \18949 , RIbe2ab68_104);
nand \U$20332 ( \20578 , \20576 , \20577 );
xor \U$20333 ( \20579 , RIbe284f8_22, RIbe2b018_114);
not \U$20334 ( \20580 , \20579 );
not \U$20335 ( \20581 , \17571 );
or \U$20336 ( \20582 , \20580 , \20581 );
buf \U$20337 ( \20583 , \18777 );
nand \U$20338 ( \20584 , \20393 , \20583 );
nand \U$20339 ( \20585 , \20582 , \20584 );
xor \U$20340 ( \20586 , \20578 , \20585 );
not \U$20341 ( \20587 , \20390 );
not \U$20342 ( \20588 , \20385 );
or \U$20343 ( \20589 , \20587 , \20588 );
or \U$20344 ( \20590 , \20385 , \20390 );
nand \U$20345 ( \20591 , \20589 , \20590 );
and \U$20346 ( \20592 , \20586 , \20591 );
and \U$20347 ( \20593 , \20578 , \20585 );
or \U$20348 ( \20594 , \20592 , \20593 );
xor \U$20349 ( \20595 , \20405 , \20378 );
xor \U$20350 ( \20596 , \20594 , \20595 );
xor \U$20351 ( \20597 , RIbe296c8_60, RIbe2ac58_106);
not \U$20352 ( \20598 , \20597 );
not \U$20353 ( \20599 , \2875 );
or \U$20354 ( \20600 , \20598 , \20599 );
nand \U$20355 ( \20601 , \907 , \20302 );
nand \U$20356 ( \20602 , \20600 , \20601 );
xor \U$20357 ( \20603 , RIbe27d78_6, RIbe2aeb0_111);
not \U$20358 ( \20604 , \20603 );
not \U$20359 ( \20605 , \1043 );
or \U$20360 ( \20606 , \20604 , \20605 );
nand \U$20361 ( \20607 , \314 , \20380 );
nand \U$20362 ( \20608 , \20606 , \20607 );
or \U$20363 ( \20609 , \20602 , \20608 );
xor \U$20364 ( \20610 , RIbe29e48_76, RIbe29998_66);
not \U$20365 ( \20611 , \20610 );
not \U$20366 ( \20612 , \9252 );
or \U$20367 ( \20613 , \20611 , \20612 );
xor \U$20368 ( \20614 , RIbe28d68_40, RIbe29e48_76);
nand \U$20369 ( \20615 , \7368 , \20614 );
nand \U$20370 ( \20616 , \20613 , \20615 );
nand \U$20371 ( \20617 , \20609 , \20616 );
nand \U$20372 ( \20618 , \20608 , \20602 );
nand \U$20373 ( \20619 , \20617 , \20618 );
not \U$20374 ( \20620 , \20619 );
xor \U$20375 ( \20621 , RIbe29d58_74, RIbe27fd0_11);
not \U$20376 ( \20622 , \20621 );
not \U$20377 ( \20623 , \12808 );
or \U$20378 ( \20624 , \20622 , \20623 );
xor \U$20379 ( \20625 , RIbe27fd0_11, RIbe29ce0_73);
nand \U$20380 ( \20626 , \2707 , \20625 );
nand \U$20381 ( \20627 , \20624 , \20626 );
not \U$20382 ( \20628 , \20627 );
and \U$20383 ( \20629 , \369 , RIbe2ae38_110);
xor \U$20384 ( \20630 , RIbe2b450_123, RIbe290b0_47);
not \U$20385 ( \20631 , \20630 );
not \U$20386 ( \20632 , \523 );
or \U$20387 ( \20633 , \20631 , \20632 );
nand \U$20388 ( \20634 , \399 , \20466 );
nand \U$20389 ( \20635 , \20633 , \20634 );
xor \U$20390 ( \20636 , \20629 , \20635 );
not \U$20391 ( \20637 , \20636 );
or \U$20392 ( \20638 , \20628 , \20637 );
nand \U$20393 ( \20639 , \20635 , \20629 );
nand \U$20394 ( \20640 , \20638 , \20639 );
not \U$20395 ( \20641 , \20640 );
or \U$20396 ( \20642 , \20620 , \20641 );
or \U$20397 ( \20643 , \20640 , \20619 );
xor \U$20398 ( \20644 , RIbe29f38_78, RIbe27e68_8);
not \U$20399 ( \20645 , \20644 );
not \U$20400 ( \20646 , \4443 );
or \U$20401 ( \20647 , \20645 , \20646 );
nand \U$20402 ( \20648 , \4447 , \20411 );
nand \U$20403 ( \20649 , \20647 , \20648 );
not \U$20404 ( \20650 , \20649 );
xor \U$20405 ( \20651 , RIbe29470_55, RIbe2a280_85);
not \U$20406 ( \20652 , \20651 );
not \U$20407 ( \20653 , \11345 );
or \U$20408 ( \20654 , \20652 , \20653 );
xor \U$20409 ( \20655 , RIbe294e8_56, RIbe2a280_85);
nand \U$20410 ( \20656 , \18667 , \20655 );
nand \U$20411 ( \20657 , \20654 , \20656 );
xor \U$20412 ( \20658 , RIbe29b00_69, RIbe2a3e8_88);
not \U$20413 ( \20659 , \20658 );
not \U$20414 ( \20660 , \8806 );
or \U$20415 ( \20661 , \20659 , \20660 );
nand \U$20416 ( \20662 , \10476 , \20429 );
nand \U$20417 ( \20663 , \20661 , \20662 );
and \U$20418 ( \20664 , \20657 , \20663 );
not \U$20419 ( \20665 , \20657 );
not \U$20420 ( \20666 , \20663 );
and \U$20421 ( \20667 , \20665 , \20666 );
nor \U$20422 ( \20668 , \20664 , \20667 );
not \U$20423 ( \20669 , \20668 );
or \U$20424 ( \20670 , \20650 , \20669 );
nand \U$20425 ( \20671 , \20657 , \20663 );
nand \U$20426 ( \20672 , \20670 , \20671 );
nand \U$20427 ( \20673 , \20643 , \20672 );
nand \U$20428 ( \20674 , \20642 , \20673 );
and \U$20429 ( \20675 , \20596 , \20674 );
and \U$20430 ( \20676 , \20594 , \20595 );
or \U$20431 ( \20677 , \20675 , \20676 );
not \U$20432 ( \20678 , \20677 );
xor \U$20433 ( \20679 , \18802 , \18751 );
not \U$20434 ( \20680 , \20679 );
not \U$20435 ( \20681 , \20680 );
not \U$20436 ( \20682 , \20551 );
not \U$20437 ( \20683 , \20541 );
or \U$20438 ( \20684 , \20682 , \20683 );
nand \U$20439 ( \20685 , \20540 , \20550 );
nand \U$20440 ( \20686 , \20684 , \20685 );
and \U$20441 ( \20687 , \20686 , \20537 );
not \U$20442 ( \20688 , \20686 );
not \U$20443 ( \20689 , \20537 );
and \U$20444 ( \20690 , \20688 , \20689 );
nor \U$20445 ( \20691 , \20687 , \20690 );
not \U$20446 ( \20692 , \20691 );
not \U$20447 ( \20693 , \20692 );
or \U$20448 ( \20694 , \20681 , \20693 );
nand \U$20449 ( \20695 , \20691 , \20679 );
nand \U$20450 ( \20696 , \20694 , \20695 );
not \U$20451 ( \20697 , \20696 );
or \U$20452 ( \20698 , \20678 , \20697 );
nand \U$20453 ( \20699 , \20692 , \20679 );
nand \U$20454 ( \20700 , \20698 , \20699 );
not \U$20455 ( \20701 , \20700 );
xor \U$20456 ( \20702 , \20534 , \20553 );
xor \U$20457 ( \20703 , \20702 , \20558 );
not \U$20458 ( \20704 , \20703 );
xor \U$20459 ( \20705 , \20504 , \20509 );
xnor \U$20460 ( \20706 , \20705 , \20501 );
not \U$20461 ( \20707 , \20706 );
or \U$20462 ( \20708 , \20704 , \20707 );
or \U$20463 ( \20709 , \20706 , \20703 );
nand \U$20464 ( \20710 , \20708 , \20709 );
not \U$20465 ( \20711 , \20710 );
or \U$20466 ( \20712 , \20701 , \20711 );
not \U$20467 ( \20713 , \20703 );
buf \U$20468 ( \20714 , \20706 );
nand \U$20469 ( \20715 , \20713 , \20714 );
nand \U$20470 ( \20716 , \20712 , \20715 );
not \U$20471 ( \20717 , \20716 );
or \U$20472 ( \20718 , \20571 , \20717 );
or \U$20473 ( \20719 , \20716 , \20570 );
nand \U$20474 ( \20720 , \20718 , \20719 );
not \U$20475 ( \20721 , \20720 );
or \U$20476 ( \20722 , \20519 , \20721 );
not \U$20477 ( \20723 , \20570 );
nand \U$20478 ( \20724 , \20723 , \20716 );
nand \U$20479 ( \20725 , \20722 , \20724 );
not \U$20480 ( \20726 , \20725 );
xor \U$20481 ( \20727 , \18886 , \18982 );
xnor \U$20482 ( \20728 , \20727 , \18812 );
not \U$20483 ( \20729 , \20728 );
not \U$20484 ( \20730 , \19012 );
and \U$20485 ( \20731 , \19060 , \20730 );
not \U$20486 ( \20732 , \19060 );
and \U$20487 ( \20733 , \20732 , \19012 );
nor \U$20488 ( \20734 , \20731 , \20733 );
not \U$20489 ( \20735 , \20734 );
not \U$20490 ( \20736 , \20735 );
not \U$20491 ( \20737 , \18975 );
not \U$20492 ( \20738 , \18914 );
and \U$20493 ( \20739 , \20737 , \20738 );
and \U$20494 ( \20740 , \18975 , \18914 );
nor \U$20495 ( \20741 , \20739 , \20740 );
not \U$20496 ( \20742 , \20741 );
and \U$20497 ( \20743 , \19207 , \19178 );
not \U$20498 ( \20744 , \19207 );
and \U$20499 ( \20745 , \20744 , \19179 );
or \U$20500 ( \20746 , \20743 , \20745 );
not \U$20501 ( \20747 , \19219 );
xor \U$20502 ( \20748 , \20746 , \20747 );
not \U$20503 ( \20749 , \20748 );
or \U$20504 ( \20750 , \20742 , \20749 );
or \U$20505 ( \20751 , \20741 , \20748 );
nand \U$20506 ( \20752 , \20750 , \20751 );
not \U$20507 ( \20753 , \20752 );
or \U$20508 ( \20754 , \20736 , \20753 );
not \U$20509 ( \20755 , \20741 );
nand \U$20510 ( \20756 , \20755 , \20748 );
nand \U$20511 ( \20757 , \20754 , \20756 );
not \U$20512 ( \20758 , \20757 );
xor \U$20513 ( \20759 , \19215 , \19132 );
xor \U$20514 ( \20760 , \19019 , \19026 );
xor \U$20515 ( \20761 , \20760 , \19033 );
or \U$20516 ( \20762 , \20759 , \20761 );
xor \U$20517 ( \20763 , \19106 , \19112 );
xor \U$20518 ( \20764 , \20763 , \19120 );
nand \U$20519 ( \20765 , \20762 , \20764 );
nand \U$20520 ( \20766 , \20761 , \20759 );
nand \U$20521 ( \20767 , \20765 , \20766 );
xor \U$20522 ( \20768 , \19078 , \19099 );
xor \U$20523 ( \20769 , \20768 , \19123 );
nor \U$20524 ( \20770 , \20767 , \20769 );
buf \U$20525 ( \20771 , \20770 );
xor \U$20526 ( \20772 , \18966 , \18947 );
not \U$20527 ( \20773 , \20772 );
not \U$20528 ( \20774 , \20773 );
xor \U$20529 ( \20775 , \19097 , \19079 );
xor \U$20530 ( \20776 , \20775 , \19087 );
not \U$20531 ( \20777 , \20776 );
or \U$20532 ( \20778 , \20774 , \20777 );
xor \U$20533 ( \20779 , \19042 , \19049 );
xor \U$20534 ( \20780 , \20779 , \19056 );
nand \U$20535 ( \20781 , \20778 , \20780 );
not \U$20536 ( \20782 , \20776 );
nand \U$20537 ( \20783 , \20782 , \20772 );
nand \U$20538 ( \20784 , \20781 , \20783 );
not \U$20539 ( \20785 , \20784 );
or \U$20540 ( \20786 , \20771 , \20785 );
nand \U$20541 ( \20787 , \20767 , \20769 );
nand \U$20542 ( \20788 , \20786 , \20787 );
not \U$20543 ( \20789 , \20788 );
not \U$20544 ( \20790 , \20789 );
xor \U$20545 ( \20791 , \19064 , \19222 );
not \U$20546 ( \20792 , \20791 );
or \U$20547 ( \20793 , \20790 , \20792 );
or \U$20548 ( \20794 , \20791 , \20789 );
nand \U$20549 ( \20795 , \20793 , \20794 );
not \U$20550 ( \20796 , \20795 );
or \U$20551 ( \20797 , \20758 , \20796 );
nand \U$20552 ( \20798 , \20791 , \20788 );
nand \U$20553 ( \20799 , \20797 , \20798 );
not \U$20554 ( \20800 , \20799 );
xor \U$20555 ( \20801 , \18889 , \18979 );
xnor \U$20556 ( \20802 , \20801 , \18909 );
not \U$20557 ( \20803 , \20802 );
not \U$20558 ( \20804 , \20625 );
not \U$20559 ( \20805 , \9082 );
or \U$20560 ( \20806 , \20804 , \20805 );
nand \U$20561 ( \20807 , \2707 , \18924 );
nand \U$20562 ( \20808 , \20806 , \20807 );
not \U$20563 ( \20809 , \20808 );
not \U$20564 ( \20810 , \20655 );
not \U$20565 ( \20811 , \10845 );
or \U$20566 ( \20812 , \20810 , \20811 );
nand \U$20567 ( \20813 , \18667 , \19182 );
nand \U$20568 ( \20814 , \20812 , \20813 );
not \U$20569 ( \20815 , \20814 );
or \U$20570 ( \20816 , \20809 , \20815 );
or \U$20571 ( \20817 , \20814 , \20808 );
not \U$20572 ( \20818 , \20614 );
not \U$20573 ( \20819 , \16652 );
or \U$20574 ( \20820 , \20818 , \20819 );
nand \U$20575 ( \20821 , \4849 , \19199 );
nand \U$20576 ( \20822 , \20820 , \20821 );
nand \U$20577 ( \20823 , \20817 , \20822 );
nand \U$20578 ( \20824 , \20816 , \20823 );
xor \U$20579 ( \20825 , RIbe285e8_24, RIbe2b6a8_128);
not \U$20580 ( \20826 , \20825 );
not \U$20581 ( \20827 , \10863 );
or \U$20582 ( \20828 , \20826 , \20827 );
nand \U$20583 ( \20829 , \2758 , \18942 );
nand \U$20584 ( \20830 , \20828 , \20829 );
xor \U$20585 ( \20831 , RIbe29a10_67, RIbe2a2f8_86);
not \U$20586 ( \20832 , \20831 );
not \U$20587 ( \20833 , \16714 );
or \U$20588 ( \20834 , \20832 , \20833 );
nand \U$20589 ( \20835 , \8705 , \18955 );
nand \U$20590 ( \20836 , \20834 , \20835 );
xor \U$20591 ( \20837 , \20830 , \20836 );
xor \U$20592 ( \20838 , RIbe29308_52, RIbe2b180_117);
not \U$20593 ( \20839 , \20838 );
not \U$20594 ( \20840 , \15353 );
or \U$20595 ( \20841 , \20839 , \20840 );
nand \U$20596 ( \20842 , \14966 , \19127 );
nand \U$20597 ( \20843 , \20841 , \20842 );
and \U$20598 ( \20844 , \20837 , \20843 );
and \U$20599 ( \20845 , \20830 , \20836 );
or \U$20600 ( \20846 , \20844 , \20845 );
xor \U$20601 ( \20847 , \20824 , \20846 );
not \U$20602 ( \20848 , \20847 );
not \U$20603 ( \20849 , \19007 );
not \U$20604 ( \20850 , \19002 );
or \U$20605 ( \20851 , \20849 , \20850 );
or \U$20606 ( \20852 , \19002 , \19007 );
nand \U$20607 ( \20853 , \20851 , \20852 );
not \U$20608 ( \20854 , \20853 );
or \U$20609 ( \20855 , \20848 , \20854 );
nand \U$20610 ( \20856 , \20846 , \20824 );
nand \U$20611 ( \20857 , \20855 , \20856 );
not \U$20612 ( \20858 , \20857 );
xor \U$20613 ( \20859 , \18895 , \18898 );
xnor \U$20614 ( \20860 , \20859 , \18904 );
not \U$20615 ( \20861 , \20860 );
or \U$20616 ( \20862 , \20858 , \20861 );
or \U$20617 ( \20863 , \20860 , \20857 );
xor \U$20618 ( \20864 , \18929 , \18938 );
xnor \U$20619 ( \20865 , \20864 , \18922 );
not \U$20620 ( \20866 , \20865 );
not \U$20621 ( \20867 , \20866 );
not \U$20622 ( \20868 , \19158 );
not \U$20623 ( \20869 , \20868 );
not \U$20624 ( \20870 , \19174 );
or \U$20625 ( \20871 , \20869 , \20870 );
or \U$20626 ( \20872 , \19174 , \20868 );
nand \U$20627 ( \20873 , \20871 , \20872 );
not \U$20628 ( \20874 , \20873 );
not \U$20629 ( \20875 , \20874 );
not \U$20630 ( \20876 , \19204 );
not \U$20631 ( \20877 , \19188 );
or \U$20632 ( \20878 , \20876 , \20877 );
not \U$20633 ( \20879 , \19204 );
nand \U$20634 ( \20880 , \20879 , \19187 );
nand \U$20635 ( \20881 , \20878 , \20880 );
and \U$20636 ( \20882 , \20881 , \19196 );
not \U$20637 ( \20883 , \20881 );
and \U$20638 ( \20884 , \20883 , \19195 );
nor \U$20639 ( \20885 , \20882 , \20884 );
not \U$20640 ( \20886 , \20885 );
not \U$20641 ( \20887 , \20886 );
or \U$20642 ( \20888 , \20875 , \20887 );
nand \U$20643 ( \20889 , \20873 , \20885 );
nand \U$20644 ( \20890 , \20888 , \20889 );
not \U$20645 ( \20891 , \20890 );
or \U$20646 ( \20892 , \20867 , \20891 );
nand \U$20647 ( \20893 , \20873 , \20886 );
nand \U$20648 ( \20894 , \20892 , \20893 );
nand \U$20649 ( \20895 , \20863 , \20894 );
nand \U$20650 ( \20896 , \20862 , \20895 );
not \U$20651 ( \20897 , \20896 );
not \U$20652 ( \20898 , \20897 );
or \U$20653 ( \20899 , \20803 , \20898 );
not \U$20654 ( \20900 , \18659 );
not \U$20655 ( \20901 , \18808 );
or \U$20656 ( \20902 , \20900 , \20901 );
or \U$20657 ( \20903 , \18808 , \18659 );
nand \U$20658 ( \20904 , \20902 , \20903 );
nand \U$20659 ( \20905 , \20899 , \20904 );
not \U$20660 ( \20906 , \20802 );
nand \U$20661 ( \20907 , \20906 , \20896 );
and \U$20662 ( \20908 , \20905 , \20907 );
not \U$20663 ( \20909 , \20908 );
or \U$20664 ( \20910 , \20800 , \20909 );
or \U$20665 ( \20911 , \20908 , \20799 );
nand \U$20666 ( \20912 , \20910 , \20911 );
not \U$20667 ( \20913 , \20912 );
or \U$20668 ( \20914 , \20729 , \20913 );
not \U$20669 ( \20915 , \20908 );
nand \U$20670 ( \20916 , \20915 , \20799 );
nand \U$20671 ( \20917 , \20914 , \20916 );
not \U$20672 ( \20918 , \20917 );
not \U$20673 ( \20919 , \19688 );
not \U$20674 ( \20920 , \19680 );
or \U$20675 ( \20921 , \20919 , \20920 );
or \U$20676 ( \20922 , \19680 , \19688 );
nand \U$20677 ( \20923 , \20921 , \20922 );
or \U$20678 ( \20924 , \20923 , \19908 );
nand \U$20679 ( \20925 , \19908 , \20923 );
nand \U$20680 ( \20926 , \20924 , \20925 );
xor \U$20681 ( \20927 , \20110 , \19960 );
xnor \U$20682 ( \20928 , \20927 , \20119 );
xor \U$20683 ( \20929 , \20926 , \20928 );
not \U$20684 ( \20930 , \20929 );
not \U$20685 ( \20931 , \20525 );
not \U$20686 ( \20932 , \20565 );
not \U$20687 ( \20933 , \20569 );
or \U$20688 ( \20934 , \20932 , \20933 );
or \U$20689 ( \20935 , \20565 , \20569 );
nand \U$20690 ( \20936 , \20934 , \20935 );
not \U$20691 ( \20937 , \20936 );
or \U$20692 ( \20938 , \20931 , \20937 );
not \U$20693 ( \20939 , \20569 );
nand \U$20694 ( \20940 , \20939 , \20565 );
nand \U$20695 ( \20941 , \20938 , \20940 );
not \U$20696 ( \20942 , \20941 );
not \U$20697 ( \20943 , \20942 );
and \U$20698 ( \20944 , \20930 , \20943 );
and \U$20699 ( \20945 , \20942 , \20929 );
nor \U$20700 ( \20946 , \20944 , \20945 );
not \U$20701 ( \20947 , \20946 );
or \U$20702 ( \20948 , \20918 , \20947 );
or \U$20703 ( \20949 , \20917 , \20946 );
nand \U$20704 ( \20950 , \20948 , \20949 );
not \U$20705 ( \20951 , \20950 );
or \U$20706 ( \20952 , \20726 , \20951 );
not \U$20707 ( \20953 , \20946 );
nand \U$20708 ( \20954 , \20953 , \20917 );
nand \U$20709 ( \20955 , \20952 , \20954 );
xor \U$20710 ( \20956 , \20127 , \20955 );
not \U$20711 ( \20957 , \20271 );
not \U$20712 ( \20958 , \20231 );
or \U$20713 ( \20959 , \20957 , \20958 );
not \U$20714 ( \20960 , \20227 );
nand \U$20715 ( \20961 , \20960 , \20169 );
nand \U$20716 ( \20962 , \20959 , \20961 );
not \U$20717 ( \20963 , \20962 );
not \U$20718 ( \20964 , \19374 );
not \U$20719 ( \20965 , \19380 );
or \U$20720 ( \20966 , \20964 , \20965 );
or \U$20721 ( \20967 , \19380 , \19374 );
nand \U$20722 ( \20968 , \20967 , \19388 );
nand \U$20723 ( \20969 , \20966 , \20968 );
not \U$20724 ( \20970 , \20181 );
not \U$20725 ( \20971 , \20175 );
or \U$20726 ( \20972 , \20970 , \20971 );
or \U$20727 ( \20973 , \20175 , \20181 );
nand \U$20728 ( \20974 , \20973 , \20188 );
nand \U$20729 ( \20975 , \20972 , \20974 );
xor \U$20730 ( \20976 , \20969 , \20975 );
not \U$20731 ( \20977 , \20143 );
not \U$20732 ( \20978 , \20138 );
or \U$20733 ( \20979 , \20977 , \20978 );
nand \U$20734 ( \20980 , \20137 , \20132 );
nand \U$20735 ( \20981 , \20979 , \20980 );
xor \U$20736 ( \20982 , \20976 , \20981 );
xor \U$20737 ( \20983 , \19595 , \19596 );
xor \U$20738 ( \20984 , \20983 , \19622 );
xor \U$20739 ( \20985 , \20982 , \20984 );
xor \U$20740 ( \20986 , \20149 , \20154 );
and \U$20741 ( \20987 , \20986 , \20160 );
and \U$20742 ( \20988 , \20149 , \20154 );
or \U$20743 ( \20989 , \20987 , \20988 );
not \U$20744 ( \20990 , \20246 );
not \U$20745 ( \20991 , \20241 );
or \U$20746 ( \20992 , \20990 , \20991 );
or \U$20747 ( \20993 , \20241 , \20246 );
nand \U$20748 ( \20994 , \20993 , \20252 );
nand \U$20749 ( \20995 , \20992 , \20994 );
xor \U$20750 ( \20996 , \20989 , \20995 );
not \U$20751 ( \20997 , \20205 );
not \U$20752 ( \20998 , \20221 );
or \U$20753 ( \20999 , \20997 , \20998 );
nand \U$20754 ( \21000 , \20217 , \20210 );
nand \U$20755 ( \21001 , \20999 , \21000 );
xor \U$20756 ( \21002 , \20996 , \21001 );
xnor \U$20757 ( \21003 , \20985 , \21002 );
not \U$20758 ( \21004 , \20234 );
not \U$20759 ( \21005 , \20265 );
or \U$20760 ( \21006 , \21004 , \21005 );
nand \U$20761 ( \21007 , \21006 , \20266 );
not \U$20762 ( \21008 , \21007 );
not \U$20763 ( \21009 , \20199 );
not \U$20764 ( \21010 , \20222 );
or \U$20765 ( \21011 , \21009 , \21010 );
nand \U$20766 ( \21012 , \21011 , \20198 );
not \U$20767 ( \21013 , \21012 );
not \U$20768 ( \21014 , \21013 );
or \U$20769 ( \21015 , \21008 , \21014 );
not \U$20770 ( \21016 , \21007 );
nand \U$20771 ( \21017 , \21016 , \21012 );
nand \U$20772 ( \21018 , \21015 , \21017 );
xor \U$20773 ( \21019 , \20144 , \20161 );
and \U$20774 ( \21020 , \21019 , \20168 );
and \U$20775 ( \21021 , \20144 , \20161 );
or \U$20776 ( \21022 , \21020 , \21021 );
not \U$20777 ( \21023 , \21022 );
and \U$20778 ( \21024 , \21018 , \21023 );
not \U$20779 ( \21025 , \21018 );
and \U$20780 ( \21026 , \21025 , \21022 );
nor \U$20781 ( \21027 , \21024 , \21026 );
nand \U$20782 ( \21028 , \21003 , \21027 );
not \U$20783 ( \21029 , \21028 );
or \U$20784 ( \21030 , \20963 , \21029 );
not \U$20785 ( \21031 , \21003 );
not \U$20786 ( \21032 , \21027 );
nand \U$20787 ( \21033 , \21031 , \21032 );
nand \U$20788 ( \21034 , \21030 , \21033 );
not \U$20789 ( \21035 , \21034 );
not \U$20790 ( \21036 , \21035 );
not \U$20791 ( \21037 , \19955 );
not \U$20792 ( \21038 , \19951 );
or \U$20793 ( \21039 , \21037 , \21038 );
nand \U$20794 ( \21040 , \19950 , \19944 );
nand \U$20795 ( \21041 , \21039 , \21040 );
not \U$20796 ( \21042 , \21001 );
not \U$20797 ( \21043 , \20996 );
or \U$20798 ( \21044 , \21042 , \21043 );
nand \U$20799 ( \21045 , \20989 , \20995 );
nand \U$20800 ( \21046 , \21044 , \21045 );
not \U$20801 ( \21047 , \21046 );
not \U$20802 ( \21048 , \21047 );
and \U$20803 ( \21049 , \18259 , \17813 );
not \U$20804 ( \21050 , \18259 );
and \U$20805 ( \21051 , \21050 , \17814 );
nor \U$20806 ( \21052 , \21049 , \21051 );
not \U$20807 ( \21053 , \21052 );
not \U$20808 ( \21054 , \20011 );
not \U$20809 ( \21055 , \19989 );
or \U$20810 ( \21056 , \21054 , \21055 );
not \U$20811 ( \21057 , \19963 );
nand \U$20812 ( \21058 , \21057 , \19985 );
nand \U$20813 ( \21059 , \21056 , \21058 );
not \U$20814 ( \21060 , \21059 );
or \U$20815 ( \21061 , \21053 , \21060 );
or \U$20816 ( \21062 , \21059 , \21052 );
nand \U$20817 ( \21063 , \21061 , \21062 );
buf \U$20818 ( \21064 , \21063 );
not \U$20819 ( \21065 , \21064 );
or \U$20820 ( \21066 , \21048 , \21065 );
or \U$20821 ( \21067 , \21064 , \21047 );
nand \U$20822 ( \21068 , \21066 , \21067 );
xor \U$20823 ( \21069 , \21041 , \21068 );
not \U$20824 ( \21070 , \20017 );
not \U$20825 ( \21071 , \21070 );
not \U$20826 ( \21072 , \20045 );
or \U$20827 ( \21073 , \21071 , \21072 );
nand \U$20828 ( \21074 , \20044 , \20038 );
nand \U$20829 ( \21075 , \21073 , \21074 );
xor \U$20830 ( \21076 , \21069 , \21075 );
not \U$20831 ( \21077 , \21076 );
not \U$20832 ( \21078 , \21077 );
or \U$20833 ( \21079 , \21036 , \21078 );
nand \U$20834 ( \21080 , \21034 , \21076 );
nand \U$20835 ( \21081 , \21079 , \21080 );
not \U$20836 ( \21082 , \21012 );
not \U$20837 ( \21083 , \21022 );
or \U$20838 ( \21084 , \21082 , \21083 );
or \U$20839 ( \21085 , \21022 , \21012 );
nand \U$20840 ( \21086 , \21085 , \21007 );
nand \U$20841 ( \21087 , \21084 , \21086 );
not \U$20842 ( \21088 , \20982 );
not \U$20843 ( \21089 , \20984 );
or \U$20844 ( \21090 , \21088 , \21089 );
or \U$20845 ( \21091 , \20984 , \20982 );
nand \U$20846 ( \21092 , \21091 , \21002 );
nand \U$20847 ( \21093 , \21090 , \21092 );
xor \U$20848 ( \21094 , \21087 , \21093 );
xor \U$20849 ( \21095 , \20969 , \20975 );
and \U$20850 ( \21096 , \21095 , \20981 );
and \U$20851 ( \21097 , \20969 , \20975 );
or \U$20852 ( \21098 , \21096 , \21097 );
xor \U$20853 ( \21099 , \17687 , \17668 );
xor \U$20854 ( \21100 , \19445 , \19451 );
and \U$20855 ( \21101 , \21100 , \19458 );
and \U$20856 ( \21102 , \19445 , \19451 );
or \U$20857 ( \21103 , \21101 , \21102 );
not \U$20858 ( \21104 , \19521 );
not \U$20859 ( \21105 , \19526 );
or \U$20860 ( \21106 , \21104 , \21105 );
not \U$20861 ( \21107 , \19521 );
not \U$20862 ( \21108 , \21107 );
not \U$20863 ( \21109 , \19527 );
or \U$20864 ( \21110 , \21108 , \21109 );
nand \U$20865 ( \21111 , \21110 , \19534 );
nand \U$20866 ( \21112 , \21106 , \21111 );
xor \U$20867 ( \21113 , \21103 , \21112 );
xor \U$20868 ( \21114 , \21099 , \21113 );
xor \U$20869 ( \21115 , \21098 , \21114 );
xor \U$20870 ( \21116 , \17736 , \17767 );
xor \U$20871 ( \21117 , \21116 , \17794 );
xor \U$20872 ( \21118 , \21115 , \21117 );
and \U$20873 ( \21119 , \21094 , \21118 );
not \U$20874 ( \21120 , \21094 );
not \U$20875 ( \21121 , \21118 );
and \U$20876 ( \21122 , \21120 , \21121 );
nor \U$20877 ( \21123 , \21119 , \21122 );
and \U$20878 ( \21124 , \21081 , \21123 );
not \U$20879 ( \21125 , \21081 );
not \U$20880 ( \21126 , \21123 );
and \U$20881 ( \21127 , \21125 , \21126 );
nor \U$20882 ( \21128 , \21124 , \21127 );
not \U$20883 ( \21129 , \21128 );
buf \U$20884 ( \21130 , \20926 );
not \U$20885 ( \21131 , \21130 );
not \U$20886 ( \21132 , \20928 );
nand \U$20887 ( \21133 , \21131 , \21132 );
not \U$20888 ( \21134 , \21133 );
nor \U$20889 ( \21135 , \21134 , \20941 );
and \U$20890 ( \21136 , \20926 , \20928 );
nor \U$20891 ( \21137 , \21135 , \21136 );
not \U$20892 ( \21138 , \21137 );
or \U$20893 ( \21139 , \21129 , \21138 );
not \U$20894 ( \21140 , \21136 );
not \U$20895 ( \21141 , \21140 );
nand \U$20896 ( \21142 , \20942 , \21133 );
not \U$20897 ( \21143 , \21142 );
or \U$20898 ( \21144 , \21141 , \21143 );
not \U$20899 ( \21145 , \21128 );
nand \U$20900 ( \21146 , \21144 , \21145 );
nand \U$20901 ( \21147 , \21139 , \21146 );
nand \U$20902 ( \21148 , \21033 , \21028 );
not \U$20903 ( \21149 , \20962 );
and \U$20904 ( \21150 , \21148 , \21149 );
not \U$20905 ( \21151 , \21148 );
and \U$20906 ( \21152 , \21151 , \20962 );
nor \U$20907 ( \21153 , \21150 , \21152 );
xor \U$20908 ( \21154 , \19407 , \19547 );
xor \U$20909 ( \21155 , \21154 , \18987 );
xor \U$20910 ( \21156 , \21153 , \21155 );
not \U$20911 ( \21157 , \20517 );
xnor \U$20912 ( \21158 , \20231 , \20271 );
not \U$20913 ( \21159 , \21158 );
not \U$20914 ( \21160 , \20277 );
or \U$20915 ( \21161 , \21159 , \21160 );
or \U$20916 ( \21162 , \20277 , \21158 );
nand \U$20917 ( \21163 , \21161 , \21162 );
not \U$20918 ( \21164 , \21163 );
or \U$20919 ( \21165 , \21157 , \21164 );
not \U$20920 ( \21166 , \21158 );
nand \U$20921 ( \21167 , \21166 , \20277 );
nand \U$20922 ( \21168 , \21165 , \21167 );
and \U$20923 ( \21169 , \21156 , \21168 );
and \U$20924 ( \21170 , \21153 , \21155 );
or \U$20925 ( \21171 , \21169 , \21170 );
not \U$20926 ( \21172 , \21171 );
and \U$20927 ( \21173 , \21147 , \21172 );
not \U$20928 ( \21174 , \21147 );
and \U$20929 ( \21175 , \21174 , \21171 );
nor \U$20930 ( \21176 , \21173 , \21175 );
xnor \U$20931 ( \21177 , \20956 , \21176 );
not \U$20932 ( \21178 , \21177 );
xnor \U$20933 ( \21179 , \20912 , \20728 );
not \U$20934 ( \21180 , \21179 );
xor \U$20935 ( \21181 , \20795 , \20757 );
not \U$20936 ( \21182 , \21181 );
xnor \U$20937 ( \21183 , \20752 , \20734 );
not \U$20938 ( \21184 , \20338 );
and \U$20939 ( \21185 , \20331 , \21184 );
not \U$20940 ( \21186 , \20331 );
and \U$20941 ( \21187 , \21186 , \20338 );
nor \U$20942 ( \21188 , \21185 , \21187 );
not \U$20943 ( \21189 , \20345 );
and \U$20944 ( \21190 , \21188 , \21189 );
not \U$20945 ( \21191 , \21188 );
and \U$20946 ( \21192 , \21191 , \20345 );
nor \U$20947 ( \21193 , \21190 , \21192 );
not \U$20948 ( \21194 , \21193 );
not \U$20949 ( \21195 , \8270 );
not \U$20950 ( \21196 , \20825 );
or \U$20951 ( \21197 , \21195 , \21196 );
xor \U$20952 ( \21198 , RIbe285e8_24, RIbe2aa78_102);
not \U$20953 ( \21199 , \21198 );
or \U$20954 ( \21200 , \2762 , \21199 );
nand \U$20955 ( \21201 , \21197 , \21200 );
not \U$20956 ( \21202 , \11094 );
not \U$20957 ( \21203 , \20831 );
or \U$20958 ( \21204 , \21202 , \21203 );
xnor \U$20959 ( \21205 , RIbe2a2f8_86, RIbe29218_50);
or \U$20960 ( \21206 , \8988 , \21205 );
nand \U$20961 ( \21207 , \21204 , \21206 );
nor \U$20962 ( \21208 , \21201 , \21207 );
xor \U$20963 ( \21209 , RIbe280c0_13, RIbe2a6b8_94);
and \U$20964 ( \21210 , \2379 , \21209 );
and \U$20965 ( \21211 , \2369 , \20279 );
nor \U$20966 ( \21212 , \21210 , \21211 );
or \U$20967 ( \21213 , \21208 , \21212 );
nand \U$20968 ( \21214 , \21207 , \21201 );
nand \U$20969 ( \21215 , \21213 , \21214 );
not \U$20970 ( \21216 , \20416 );
and \U$20971 ( \21217 , \20438 , \21216 );
not \U$20972 ( \21218 , \20438 );
and \U$20973 ( \21219 , \21218 , \20416 );
nor \U$20974 ( \21220 , \21217 , \21219 );
and \U$20975 ( \21221 , \21215 , \21220 );
not \U$20976 ( \21222 , \21215 );
not \U$20977 ( \21223 , \21220 );
and \U$20978 ( \21224 , \21222 , \21223 );
or \U$20979 ( \21225 , \21221 , \21224 );
not \U$20980 ( \21226 , \21225 );
or \U$20981 ( \21227 , \21194 , \21226 );
nand \U$20982 ( \21228 , \21215 , \21223 );
nand \U$20983 ( \21229 , \21227 , \21228 );
not \U$20984 ( \21230 , \21229 );
xor \U$20985 ( \21231 , \20865 , \20890 );
xor \U$20986 ( \21232 , \20471 , \20477 );
xor \U$20987 ( \21233 , \21232 , \20484 );
xor \U$20988 ( \21234 , \20830 , \20836 );
xor \U$20989 ( \21235 , \21234 , \20843 );
or \U$20990 ( \21236 , \21233 , \21235 );
xor \U$20991 ( \21237 , \20449 , \20455 );
xor \U$20992 ( \21238 , \21237 , \20462 );
nand \U$20993 ( \21239 , \21236 , \21238 );
nand \U$20994 ( \21240 , \21233 , \21235 );
nand \U$20995 ( \21241 , \21239 , \21240 );
xnor \U$20996 ( \21242 , \21231 , \21241 );
not \U$20997 ( \21243 , \21242 );
or \U$20998 ( \21244 , \21230 , \21243 );
nand \U$20999 ( \21245 , \20890 , \20865 );
not \U$21000 ( \21246 , \21245 );
not \U$21001 ( \21247 , \20890 );
nand \U$21002 ( \21248 , \21247 , \20866 );
not \U$21003 ( \21249 , \21248 );
or \U$21004 ( \21250 , \21246 , \21249 );
nand \U$21005 ( \21251 , \21250 , \21241 );
nand \U$21006 ( \21252 , \21244 , \21251 );
or \U$21007 ( \21253 , \21183 , \21252 );
not \U$21008 ( \21254 , \20770 );
nand \U$21009 ( \21255 , \21254 , \20787 );
and \U$21010 ( \21256 , \21255 , \20784 );
not \U$21011 ( \21257 , \21255 );
and \U$21012 ( \21258 , \21257 , \20785 );
nor \U$21013 ( \21259 , \21256 , \21258 );
not \U$21014 ( \21260 , \21259 );
nand \U$21015 ( \21261 , \21253 , \21260 );
nand \U$21016 ( \21262 , \21183 , \21252 );
nand \U$21017 ( \21263 , \21261 , \21262 );
not \U$21018 ( \21264 , \21263 );
xor \U$21019 ( \21265 , \20284 , \20290 );
xor \U$21020 ( \21266 , \21265 , \20297 );
xor \U$21021 ( \21267 , \20314 , \20307 );
xnor \U$21022 ( \21268 , \21267 , \20323 );
not \U$21023 ( \21269 , \21268 );
or \U$21024 ( \21270 , \21266 , \21269 );
xor \U$21025 ( \21271 , \20814 , \20808 );
xor \U$21026 ( \21272 , \21271 , \20822 );
nand \U$21027 ( \21273 , \21270 , \21272 );
nand \U$21028 ( \21274 , \21266 , \21269 );
nand \U$21029 ( \21275 , \21273 , \21274 );
xor \U$21030 ( \21276 , \20489 , \20487 );
xor \U$21031 ( \21277 , \21276 , \20490 );
xor \U$21032 ( \21278 , \21275 , \21277 );
xor \U$21033 ( \21279 , \20847 , \20853 );
and \U$21034 ( \21280 , \21278 , \21279 );
and \U$21035 ( \21281 , \21275 , \21277 );
or \U$21036 ( \21282 , \21280 , \21281 );
not \U$21037 ( \21283 , \21282 );
xor \U$21038 ( \21284 , RIbe28228_16, RIbe2b540_125);
not \U$21039 ( \21285 , \21284 );
not \U$21040 ( \21286 , \3056 );
or \U$21041 ( \21287 , \21285 , \21286 );
nand \U$21042 ( \21288 , \885 , \20371 );
nand \U$21043 ( \21289 , \21287 , \21288 );
not \U$21044 ( \21290 , \21289 );
xor \U$21045 ( \21291 , RIbe288b8_30, RIbe2b108_116);
not \U$21046 ( \21292 , \21291 );
not \U$21047 ( \21293 , \13541 );
or \U$21048 ( \21294 , \21292 , \21293 );
nand \U$21049 ( \21295 , \16875 , \20362 );
nand \U$21050 ( \21296 , \21294 , \21295 );
not \U$21051 ( \21297 , \21296 );
or \U$21052 ( \21298 , \21290 , \21297 );
or \U$21053 ( \21299 , \21296 , \21289 );
xor \U$21054 ( \21300 , RIbe28930_31, RIbe2adc0_109);
not \U$21055 ( \21301 , \21300 );
not \U$21056 ( \21302 , \965 );
or \U$21057 ( \21303 , \21301 , \21302 );
nand \U$21058 ( \21304 , \1199 , \20340 );
nand \U$21059 ( \21305 , \21303 , \21304 );
nand \U$21060 ( \21306 , \21299 , \21305 );
nand \U$21061 ( \21307 , \21298 , \21306 );
not \U$21062 ( \21308 , \21307 );
xor \U$21063 ( \21309 , RIbe2af28_112, RIbe28c00_37);
not \U$21064 ( \21310 , \21309 );
not \U$21065 ( \21311 , \14423 );
or \U$21066 ( \21312 , \21310 , \21311 );
nand \U$21067 ( \21313 , \14413 , \20285 );
nand \U$21068 ( \21314 , \21312 , \21313 );
not \U$21069 ( \21315 , \21314 );
xor \U$21070 ( \21316 , RIbe28b88_36, RIbe2b360_121);
not \U$21071 ( \21317 , \21316 );
not \U$21072 ( \21318 , \9052 );
or \U$21073 ( \21319 , \21317 , \21318 );
nand \U$21074 ( \21320 , \2559 , \20479 );
nand \U$21075 ( \21321 , \21319 , \21320 );
not \U$21076 ( \21322 , \21321 );
nand \U$21077 ( \21323 , \21315 , \21322 );
not \U$21078 ( \21324 , \21323 );
xor \U$21079 ( \21325 , RIbe2b180_117, RIbe293f8_54);
not \U$21080 ( \21326 , \21325 );
not \U$21081 ( \21327 , \15353 );
or \U$21082 ( \21328 , \21326 , \21327 );
nand \U$21083 ( \21329 , \14966 , \20838 );
nand \U$21084 ( \21330 , \21328 , \21329 );
not \U$21085 ( \21331 , \21330 );
or \U$21086 ( \21332 , \21324 , \21331 );
nand \U$21087 ( \21333 , \21314 , \21321 );
nand \U$21088 ( \21334 , \21332 , \21333 );
not \U$21089 ( \21335 , \21334 );
nand \U$21090 ( \21336 , \21308 , \21335 );
not \U$21091 ( \21337 , \21336 );
xor \U$21092 ( \21338 , RIbe28cf0_39, RIbe29c68_72);
not \U$21093 ( \21339 , \21338 );
not \U$21094 ( \21340 , \4578 );
or \U$21095 ( \21341 , \21339 , \21340 );
nand \U$21096 ( \21342 , \7237 , \20450 );
nand \U$21097 ( \21343 , \21341 , \21342 );
not \U$21098 ( \21344 , \21343 );
not \U$21099 ( \21345 , \19580 );
xor \U$21100 ( \21346 , RIbe28750_27, RIbe2aaf0_103);
not \U$21101 ( \21347 , \21346 );
not \U$21102 ( \21348 , \21347 );
and \U$21103 ( \21349 , \21345 , \21348 );
and \U$21104 ( \21350 , \20572 , RIbe2ab68_104);
nor \U$21105 ( \21351 , \21349 , \21350 );
not \U$21106 ( \21352 , \21351 );
xor \U$21107 ( \21353 , RIbe291a0_49, RIbe2a910_99);
not \U$21108 ( \21354 , \21353 );
not \U$21109 ( \21355 , \9737 );
or \U$21110 ( \21356 , \21354 , \21355 );
nand \U$21111 ( \21357 , \11456 , \20326 );
nand \U$21112 ( \21358 , \21356 , \21357 );
not \U$21113 ( \21359 , \21358 );
or \U$21114 ( \21360 , \21352 , \21359 );
or \U$21115 ( \21361 , \21358 , \21351 );
nand \U$21116 ( \21362 , \21360 , \21361 );
not \U$21117 ( \21363 , \21362 );
or \U$21118 ( \21364 , \21344 , \21363 );
not \U$21119 ( \21365 , \21351 );
nand \U$21120 ( \21366 , \21365 , \21358 );
nand \U$21121 ( \21367 , \21364 , \21366 );
not \U$21122 ( \21368 , \21367 );
or \U$21123 ( \21369 , \21337 , \21368 );
nand \U$21124 ( \21370 , \21334 , \21307 );
nand \U$21125 ( \21371 , \21369 , \21370 );
not \U$21126 ( \21372 , \21371 );
not \U$21127 ( \21373 , \20349 );
not \U$21128 ( \21374 , \20300 );
not \U$21129 ( \21375 , \21374 );
and \U$21130 ( \21376 , \21373 , \21375 );
and \U$21131 ( \21377 , \20349 , \21374 );
nor \U$21132 ( \21378 , \21376 , \21377 );
nand \U$21133 ( \21379 , \21372 , \21378 );
not \U$21134 ( \21380 , \21379 );
xor \U$21135 ( \21381 , RIbe2a190_83, RIbe28138_14);
not \U$21136 ( \21382 , \21381 );
or \U$21137 ( \21383 , \11973 , \21382 );
not \U$21138 ( \21384 , \20418 );
or \U$21139 ( \21385 , \11971 , \21384 );
nand \U$21140 ( \21386 , \21383 , \21385 );
not \U$21141 ( \21387 , \21386 );
not \U$21142 ( \21388 , \9524 );
not \U$21143 ( \21389 , \20472 );
or \U$21144 ( \21390 , \21388 , \21389 );
xnor \U$21145 ( \21391 , RIbe28f48_44, RIbe29b78_70);
not \U$21146 ( \21392 , \21391 );
nand \U$21147 ( \21393 , \21392 , \11461 );
nand \U$21148 ( \21394 , \21390 , \21393 );
not \U$21149 ( \21395 , \21394 );
xor \U$21150 ( \21396 , RIbe28a20_33, RIbe2a4d8_90);
not \U$21151 ( \21397 , \21396 );
not \U$21152 ( \21398 , \1781 );
or \U$21153 ( \21399 , \21397 , \21398 );
nand \U$21154 ( \21400 , \2475 , \20355 );
nand \U$21155 ( \21401 , \21399 , \21400 );
not \U$21156 ( \21402 , \21401 );
not \U$21157 ( \21403 , \21402 );
or \U$21158 ( \21404 , \21395 , \21403 );
or \U$21159 ( \21405 , \21394 , \21402 );
nand \U$21160 ( \21406 , \21404 , \21405 );
not \U$21161 ( \21407 , \21406 );
or \U$21162 ( \21408 , \21387 , \21407 );
nand \U$21163 ( \21409 , \21401 , \21394 );
nand \U$21164 ( \21410 , \21408 , \21409 );
not \U$21165 ( \21411 , \21410 );
xor \U$21166 ( \21412 , RIbe29740_61, RIbe2a550_91);
not \U$21167 ( \21413 , \21412 );
not \U$21168 ( \21414 , \10433 );
or \U$21169 ( \21415 , \21413 , \21414 );
nand \U$21170 ( \21416 , \11485 , \20332 );
nand \U$21171 ( \21417 , \21415 , \21416 );
not \U$21172 ( \21418 , \21417 );
xor \U$21173 ( \21419 , RIbe29038_46, RIbe2a7a8_96);
not \U$21174 ( \21420 , \21419 );
not \U$21175 ( \21421 , \281 );
or \U$21176 ( \21422 , \21420 , \21421 );
nand \U$21177 ( \21423 , \1583 , \20457 );
nand \U$21178 ( \21424 , \21422 , \21423 );
not \U$21179 ( \21425 , \21424 );
or \U$21180 ( \21426 , \21418 , \21425 );
or \U$21181 ( \21427 , \21424 , \21417 );
xor \U$21182 ( \21428 , RIbe28390_19, RIbe2a118_82);
not \U$21183 ( \21429 , \21428 );
not \U$21184 ( \21430 , \14806 );
or \U$21185 ( \21431 , \21429 , \21430 );
nand \U$21186 ( \21432 , \2777 , \20292 );
nand \U$21187 ( \21433 , \21431 , \21432 );
nand \U$21188 ( \21434 , \21427 , \21433 );
nand \U$21189 ( \21435 , \21426 , \21434 );
not \U$21190 ( \21436 , \21435 );
not \U$21191 ( \21437 , \21436 );
xor \U$21192 ( \21438 , RIbe28318_18, RIbe2b018_114);
not \U$21193 ( \21439 , \21438 );
not \U$21194 ( \21440 , \16811 );
or \U$21195 ( \21441 , \21439 , \21440 );
buf \U$21196 ( \21442 , \15952 );
nand \U$21197 ( \21443 , \21442 , \20579 );
nand \U$21198 ( \21444 , \21441 , \21443 );
buf \U$21199 ( \21445 , \21444 );
not \U$21200 ( \21446 , \21445 );
xor \U$21201 ( \21447 , RIbe2a028_80, RIbe27c88_4);
not \U$21202 ( \21448 , \21447 );
not \U$21203 ( \21449 , \8400 );
or \U$21204 ( \21450 , \21448 , \21449 );
nand \U$21205 ( \21451 , \8930 , \20309 );
nand \U$21206 ( \21452 , \21450 , \21451 );
not \U$21207 ( \21453 , \21452 );
or \U$21208 ( \21454 , \21446 , \21453 );
or \U$21209 ( \21455 , \21445 , \21452 );
xor \U$21210 ( \21456 , RIbe2a898_98, RIbe28480_21);
not \U$21211 ( \21457 , \21456 );
not \U$21212 ( \21458 , \3344 );
or \U$21213 ( \21459 , \21457 , \21458 );
nand \U$21214 ( \21460 , \3074 , \20318 );
nand \U$21215 ( \21461 , \21459 , \21460 );
nand \U$21216 ( \21462 , \21455 , \21461 );
nand \U$21217 ( \21463 , \21454 , \21462 );
not \U$21218 ( \21464 , \21463 );
or \U$21219 ( \21465 , \21437 , \21464 );
or \U$21220 ( \21466 , \21463 , \21436 );
nand \U$21221 ( \21467 , \21465 , \21466 );
not \U$21222 ( \21468 , \21467 );
or \U$21223 ( \21469 , \21411 , \21468 );
nand \U$21224 ( \21470 , \21463 , \21435 );
nand \U$21225 ( \21471 , \21469 , \21470 );
not \U$21226 ( \21472 , \21471 );
or \U$21227 ( \21473 , \21380 , \21472 );
not \U$21228 ( \21474 , \21378 );
nand \U$21229 ( \21475 , \21474 , \21371 );
nand \U$21230 ( \21476 , \21473 , \21475 );
not \U$21231 ( \21477 , \20353 );
not \U$21232 ( \21478 , \21477 );
not \U$21233 ( \21479 , \20497 );
or \U$21234 ( \21480 , \21478 , \21479 );
or \U$21235 ( \21481 , \20497 , \21477 );
nand \U$21236 ( \21482 , \21480 , \21481 );
xor \U$21237 ( \21483 , \21476 , \21482 );
not \U$21238 ( \21484 , \21483 );
or \U$21239 ( \21485 , \21283 , \21484 );
nand \U$21240 ( \21486 , \21482 , \21476 );
nand \U$21241 ( \21487 , \21485 , \21486 );
and \U$21242 ( \21488 , \21264 , \21487 );
not \U$21243 ( \21489 , \21264 );
not \U$21244 ( \21490 , \21487 );
and \U$21245 ( \21491 , \21489 , \21490 );
nor \U$21246 ( \21492 , \21488 , \21491 );
not \U$21247 ( \21493 , \21492 );
not \U$21248 ( \21494 , \21493 );
or \U$21249 ( \21495 , \21182 , \21494 );
not \U$21250 ( \21496 , \21264 );
nand \U$21251 ( \21497 , \21496 , \21487 );
nand \U$21252 ( \21498 , \21495 , \21497 );
not \U$21253 ( \21499 , \21498 );
not \U$21254 ( \21500 , \21499 );
or \U$21255 ( \21501 , \21180 , \21500 );
not \U$21256 ( \21502 , \20703 );
xor \U$21257 ( \21503 , \20700 , \21502 );
xnor \U$21258 ( \21504 , \21503 , \20714 );
not \U$21259 ( \21505 , \21504 );
not \U$21260 ( \21506 , \21505 );
not \U$21261 ( \21507 , \20677 );
not \U$21262 ( \21508 , \21507 );
not \U$21263 ( \21509 , \20696 );
or \U$21264 ( \21510 , \21508 , \21509 );
or \U$21265 ( \21511 , \20696 , \21507 );
nand \U$21266 ( \21512 , \21510 , \21511 );
not \U$21267 ( \21513 , \21512 );
xor \U$21268 ( \21514 , \20367 , \20360 );
not \U$21269 ( \21515 , \20376 );
and \U$21270 ( \21516 , \21514 , \21515 );
not \U$21271 ( \21517 , \21514 );
and \U$21272 ( \21518 , \21517 , \20376 );
nor \U$21273 ( \21519 , \21516 , \21518 );
xor \U$21274 ( \21520 , \20578 , \20585 );
xor \U$21275 ( \21521 , \21520 , \20591 );
xnor \U$21276 ( \21522 , \21519 , \21521 );
not \U$21277 ( \21523 , \21522 );
xor \U$21278 ( \21524 , RIbe2ae38_110, RIbe27d78_6);
not \U$21279 ( \21525 , \21524 );
not \U$21280 ( \21526 , \8768 );
or \U$21281 ( \21527 , \21525 , \21526 );
nand \U$21282 ( \21528 , \314 , \20603 );
nand \U$21283 ( \21529 , \21527 , \21528 );
xor \U$21284 ( \21530 , RIbe29ec0_77, RIbe27fd0_11);
not \U$21285 ( \21531 , \21530 );
not \U$21286 ( \21532 , \3378 );
or \U$21287 ( \21533 , \21531 , \21532 );
nand \U$21288 ( \21534 , \2707 , \20621 );
nand \U$21289 ( \21535 , \21533 , \21534 );
xor \U$21290 ( \21536 , \21529 , \21535 );
xor \U$21291 ( \21537 , RIbe298a8_64, RIbe29e48_76);
not \U$21292 ( \21538 , \21537 );
not \U$21293 ( \21539 , \4843 );
or \U$21294 ( \21540 , \21538 , \21539 );
nand \U$21295 ( \21541 , \8245 , \20610 );
nand \U$21296 ( \21542 , \21540 , \21541 );
and \U$21297 ( \21543 , \21536 , \21542 );
and \U$21298 ( \21544 , \21529 , \21535 );
or \U$21299 ( \21545 , \21543 , \21544 );
not \U$21300 ( \21546 , \21545 );
xor \U$21301 ( \21547 , RIbe290b0_47, RIbe2b3d8_122);
not \U$21302 ( \21548 , \21547 );
not \U$21303 ( \21549 , \9114 );
or \U$21304 ( \21550 , \21548 , \21549 );
nand \U$21305 ( \21551 , \399 , \20630 );
nand \U$21306 ( \21552 , \21550 , \21551 );
not \U$21307 ( \21553 , RIbe29a88_68);
nand \U$21308 ( \21554 , \21553 , \387 );
and \U$21309 ( \21555 , \21554 , RIbe2ae38_110);
nand \U$21310 ( \21556 , RIbe290b0_47, RIbe29a88_68);
nand \U$21311 ( \21557 , \21556 , RIbe27d78_6);
nor \U$21312 ( \21558 , \21555 , \21557 );
nand \U$21313 ( \21559 , \21552 , \21558 );
not \U$21314 ( \21560 , \21559 );
xor \U$21315 ( \21561 , RIbe2abe0_105, RIbe296c8_60);
not \U$21316 ( \21562 , \21561 );
not \U$21317 ( \21563 , \1129 );
or \U$21318 ( \21564 , \21562 , \21563 );
nand \U$21319 ( \21565 , \1939 , \20597 );
nand \U$21320 ( \21566 , \21564 , \21565 );
not \U$21321 ( \21567 , \21566 );
xor \U$21322 ( \21568 , RIbe29038_46, RIbe2a730_95);
not \U$21323 ( \21569 , \21568 );
not \U$21324 ( \21570 , \281 );
or \U$21325 ( \21571 , \21569 , \21570 );
nand \U$21326 ( \21572 , \1583 , \21419 );
nand \U$21327 ( \21573 , \21571 , \21572 );
not \U$21328 ( \21574 , \21573 );
or \U$21329 ( \21575 , \21567 , \21574 );
or \U$21330 ( \21576 , \21573 , \21566 );
xor \U$21331 ( \21577 , RIbe2a0a0_81, RIbe28390_19);
not \U$21332 ( \21578 , \21577 );
not \U$21333 ( \21579 , \14579 );
or \U$21334 ( \21580 , \21578 , \21579 );
nand \U$21335 ( \21581 , \2777 , \21428 );
nand \U$21336 ( \21582 , \21580 , \21581 );
nand \U$21337 ( \21583 , \21576 , \21582 );
nand \U$21338 ( \21584 , \21575 , \21583 );
not \U$21339 ( \21585 , \21584 );
or \U$21340 ( \21586 , \21560 , \21585 );
or \U$21341 ( \21587 , \21584 , \21559 );
nand \U$21342 ( \21588 , \21586 , \21587 );
not \U$21343 ( \21589 , \21588 );
or \U$21344 ( \21590 , \21546 , \21589 );
not \U$21345 ( \21591 , \21559 );
nand \U$21346 ( \21592 , \21591 , \21584 );
nand \U$21347 ( \21593 , \21590 , \21592 );
not \U$21348 ( \21594 , \21593 );
or \U$21349 ( \21595 , \21523 , \21594 );
not \U$21350 ( \21596 , \21519 );
nand \U$21351 ( \21597 , \21596 , \21521 );
nand \U$21352 ( \21598 , \21595 , \21597 );
not \U$21353 ( \21599 , \21598 );
not \U$21354 ( \21600 , \20773 );
not \U$21355 ( \21601 , \20776 );
not \U$21356 ( \21602 , \21601 );
or \U$21357 ( \21603 , \21600 , \21602 );
nand \U$21358 ( \21604 , \20776 , \20772 );
nand \U$21359 ( \21605 , \21603 , \21604 );
not \U$21360 ( \21606 , \20780 );
and \U$21361 ( \21607 , \21605 , \21606 );
not \U$21362 ( \21608 , \21605 );
and \U$21363 ( \21609 , \21608 , \20780 );
nor \U$21364 ( \21610 , \21607 , \21609 );
not \U$21365 ( \21611 , \21610 );
xor \U$21366 ( \21612 , \20759 , \20761 );
xor \U$21367 ( \21613 , \21612 , \20764 );
not \U$21368 ( \21614 , \21613 );
or \U$21369 ( \21615 , \21611 , \21614 );
or \U$21370 ( \21616 , \21613 , \21610 );
nand \U$21371 ( \21617 , \21615 , \21616 );
not \U$21372 ( \21618 , \21617 );
or \U$21373 ( \21619 , \21599 , \21618 );
not \U$21374 ( \21620 , \21610 );
nand \U$21375 ( \21621 , \21620 , \21613 );
nand \U$21376 ( \21622 , \21619 , \21621 );
xor \U$21377 ( \21623 , \20857 , \20894 );
xnor \U$21378 ( \21624 , \21623 , \20860 );
and \U$21379 ( \21625 , \21622 , \21624 );
not \U$21380 ( \21626 , \21622 );
not \U$21381 ( \21627 , \21624 );
and \U$21382 ( \21628 , \21626 , \21627 );
or \U$21383 ( \21629 , \21625 , \21628 );
not \U$21384 ( \21630 , \21629 );
or \U$21385 ( \21631 , \21513 , \21630 );
nand \U$21386 ( \21632 , \21627 , \21622 );
nand \U$21387 ( \21633 , \21631 , \21632 );
and \U$21388 ( \21634 , \20896 , \20802 );
not \U$21389 ( \21635 , \20896 );
and \U$21390 ( \21636 , \21635 , \20906 );
nor \U$21391 ( \21637 , \21634 , \21636 );
not \U$21392 ( \21638 , \20904 );
and \U$21393 ( \21639 , \21637 , \21638 );
not \U$21394 ( \21640 , \21637 );
and \U$21395 ( \21641 , \21640 , \20904 );
nor \U$21396 ( \21642 , \21639 , \21641 );
and \U$21397 ( \21643 , \21633 , \21642 );
not \U$21398 ( \21644 , \21633 );
not \U$21399 ( \21645 , \21642 );
and \U$21400 ( \21646 , \21644 , \21645 );
nor \U$21401 ( \21647 , \21643 , \21646 );
not \U$21402 ( \21648 , \21647 );
or \U$21403 ( \21649 , \21506 , \21648 );
not \U$21404 ( \21650 , \21645 );
nand \U$21405 ( \21651 , \21650 , \21633 );
nand \U$21406 ( \21652 , \21649 , \21651 );
nand \U$21407 ( \21653 , \21501 , \21652 );
not \U$21408 ( \21654 , \21179 );
nand \U$21409 ( \21655 , \21654 , \21498 );
nand \U$21410 ( \21656 , \21653 , \21655 );
xor \U$21411 ( \21657 , \21153 , \21155 );
xor \U$21412 ( \21658 , \21657 , \21168 );
not \U$21413 ( \21659 , \21658 );
and \U$21414 ( \21660 , \21656 , \21659 );
not \U$21415 ( \21661 , \21656 );
and \U$21416 ( \21662 , \21661 , \21658 );
or \U$21417 ( \21663 , \21660 , \21662 );
not \U$21418 ( \21664 , \21663 );
buf \U$21419 ( \21665 , \20950 );
buf \U$21420 ( \21666 , \20725 );
not \U$21421 ( \21667 , \21666 );
and \U$21422 ( \21668 , \21665 , \21667 );
not \U$21423 ( \21669 , \21665 );
and \U$21424 ( \21670 , \21669 , \21666 );
nor \U$21425 ( \21671 , \21668 , \21670 );
not \U$21426 ( \21672 , \21671 );
not \U$21427 ( \21673 , \21672 );
or \U$21428 ( \21674 , \21664 , \21673 );
not \U$21429 ( \21675 , \21655 );
not \U$21430 ( \21676 , \21653 );
or \U$21431 ( \21677 , \21675 , \21676 );
nand \U$21432 ( \21678 , \21677 , \21658 );
nand \U$21433 ( \21679 , \21674 , \21678 );
not \U$21434 ( \21680 , \21679 );
nand \U$21435 ( \21681 , \21178 , \21680 );
buf \U$21436 ( \21682 , \21681 );
not \U$21437 ( \21683 , \21671 );
not \U$21438 ( \21684 , \21663 );
or \U$21439 ( \21685 , \21683 , \21684 );
or \U$21440 ( \21686 , \21663 , \21671 );
nand \U$21441 ( \21687 , \21685 , \21686 );
xor \U$21442 ( \21688 , \20594 , \20595 );
xor \U$21443 ( \21689 , \21688 , \20674 );
xor \U$21444 ( \21690 , \21275 , \21277 );
xor \U$21445 ( \21691 , \21690 , \21279 );
xor \U$21446 ( \21692 , \21689 , \21691 );
xor \U$21447 ( \21693 , \21229 , \21242 );
and \U$21448 ( \21694 , \21692 , \21693 );
and \U$21449 ( \21695 , \21689 , \21691 );
or \U$21450 ( \21696 , \21694 , \21695 );
xor \U$21451 ( \21697 , \21282 , \21483 );
xor \U$21452 ( \21698 , \21696 , \21697 );
xor \U$21453 ( \21699 , \21433 , \21424 );
and \U$21454 ( \21700 , \21699 , \21417 );
not \U$21455 ( \21701 , \21699 );
not \U$21456 ( \21702 , \21417 );
and \U$21457 ( \21703 , \21701 , \21702 );
nor \U$21458 ( \21704 , \21700 , \21703 );
and \U$21459 ( \21705 , \20668 , \20649 );
not \U$21460 ( \21706 , \20668 );
not \U$21461 ( \21707 , \20649 );
and \U$21462 ( \21708 , \21706 , \21707 );
nor \U$21463 ( \21709 , \21705 , \21708 );
xor \U$21464 ( \21710 , \21704 , \21709 );
xor \U$21465 ( \21711 , \20627 , \20636 );
and \U$21466 ( \21712 , \21710 , \21711 );
and \U$21467 ( \21713 , \21704 , \21709 );
or \U$21468 ( \21714 , \21712 , \21713 );
not \U$21469 ( \21715 , \21714 );
not \U$21470 ( \21716 , \21410 );
not \U$21471 ( \21717 , \21716 );
not \U$21472 ( \21718 , \21467 );
or \U$21473 ( \21719 , \21717 , \21718 );
or \U$21474 ( \21720 , \21467 , \21716 );
nand \U$21475 ( \21721 , \21719 , \21720 );
not \U$21476 ( \21722 , \21721 );
xor \U$21477 ( \21723 , \20619 , \20672 );
xnor \U$21478 ( \21724 , \21723 , \20640 );
not \U$21479 ( \21725 , \21724 );
or \U$21480 ( \21726 , \21722 , \21725 );
or \U$21481 ( \21727 , \21724 , \21721 );
nand \U$21482 ( \21728 , \21726 , \21727 );
not \U$21483 ( \21729 , \21728 );
or \U$21484 ( \21730 , \21715 , \21729 );
not \U$21485 ( \21731 , \21724 );
nand \U$21486 ( \21732 , \21731 , \21721 );
nand \U$21487 ( \21733 , \21730 , \21732 );
not \U$21488 ( \21734 , \21733 );
xor \U$21489 ( \21735 , \21371 , \21378 );
xor \U$21490 ( \21736 , \21735 , \21471 );
not \U$21491 ( \21737 , \21736 );
xor \U$21492 ( \21738 , RIbe285e8_24, RIbe2aa00_101);
not \U$21493 ( \21739 , \21738 );
not \U$21494 ( \21740 , \8813 );
or \U$21495 ( \21741 , \21739 , \21740 );
not \U$21496 ( \21742 , \21199 );
nand \U$21497 ( \21743 , \21742 , \8270 );
nand \U$21498 ( \21744 , \21741 , \21743 );
not \U$21499 ( \21745 , \21744 );
xor \U$21500 ( \21746 , RIbe2b2e8_120, RIbe28b88_36);
not \U$21501 ( \21747 , \21746 );
not \U$21502 ( \21748 , \2701 );
or \U$21503 ( \21749 , \21747 , \21748 );
nand \U$21504 ( \21750 , \7550 , \21316 );
nand \U$21505 ( \21751 , \21749 , \21750 );
not \U$21506 ( \21752 , \21751 );
or \U$21507 ( \21753 , \21745 , \21752 );
or \U$21508 ( \21754 , \21751 , \21744 );
xor \U$21509 ( \21755 , RIbe2b180_117, RIbe28a98_34);
not \U$21510 ( \21756 , \21755 );
not \U$21511 ( \21757 , \14852 );
or \U$21512 ( \21758 , \21756 , \21757 );
not \U$21513 ( \21759 , \14846 );
nand \U$21514 ( \21760 , \21759 , \21325 );
nand \U$21515 ( \21761 , \21758 , \21760 );
nand \U$21516 ( \21762 , \21754 , \21761 );
nand \U$21517 ( \21763 , \21753 , \21762 );
xor \U$21518 ( \21764 , RIbe29a10_67, RIbe2a3e8_88);
not \U$21519 ( \21765 , \21764 );
not \U$21520 ( \21766 , \9262 );
or \U$21521 ( \21767 , \21765 , \21766 );
nand \U$21522 ( \21768 , \8794 , \20658 );
nand \U$21523 ( \21769 , \21767 , \21768 );
xor \U$21524 ( \21770 , RIbe29308_52, RIbe2af28_112);
not \U$21525 ( \21771 , \21770 );
not \U$21526 ( \21772 , \16913 );
or \U$21527 ( \21773 , \21771 , \21772 );
nand \U$21528 ( \21774 , \16917 , \21309 );
nand \U$21529 ( \21775 , \21773 , \21774 );
xor \U$21530 ( \21776 , \21769 , \21775 );
xor \U$21531 ( \21777 , RIbe282a0_17, RIbe2a280_85);
not \U$21532 ( \21778 , \21777 );
not \U$21533 ( \21779 , \15793 );
or \U$21534 ( \21780 , \21778 , \21779 );
nand \U$21535 ( \21781 , \14649 , \20651 );
nand \U$21536 ( \21782 , \21780 , \21781 );
and \U$21537 ( \21783 , \21776 , \21782 );
and \U$21538 ( \21784 , \21769 , \21775 );
or \U$21539 ( \21785 , \21783 , \21784 );
xor \U$21540 ( \21786 , \21763 , \21785 );
xor \U$21541 ( \21787 , RIbe27df0_7, RIbe2a2f8_86);
not \U$21542 ( \21788 , \21787 );
not \U$21543 ( \21789 , \8989 );
or \U$21544 ( \21790 , \21788 , \21789 );
not \U$21545 ( \21791 , \21205 );
nand \U$21546 ( \21792 , \21791 , \8706 );
nand \U$21547 ( \21793 , \21790 , \21792 );
not \U$21548 ( \21794 , \21793 );
xor \U$21549 ( \21795 , RIbe2ad48_108, RIbe28930_31);
not \U$21550 ( \21796 , \21795 );
not \U$21551 ( \21797 , \965 );
or \U$21552 ( \21798 , \21796 , \21797 );
nand \U$21553 ( \21799 , \1199 , \21300 );
nand \U$21554 ( \21800 , \21798 , \21799 );
xor \U$21555 ( \21801 , RIbe2a640_93, RIbe280c0_13);
not \U$21556 ( \21802 , \21801 );
not \U$21557 ( \21803 , \2379 );
or \U$21558 ( \21804 , \21802 , \21803 );
nand \U$21559 ( \21805 , \2369 , \21209 );
nand \U$21560 ( \21806 , \21804 , \21805 );
xor \U$21561 ( \21807 , \21800 , \21806 );
not \U$21562 ( \21808 , \21807 );
or \U$21563 ( \21809 , \21794 , \21808 );
nand \U$21564 ( \21810 , \21806 , \21800 );
nand \U$21565 ( \21811 , \21809 , \21810 );
and \U$21566 ( \21812 , \21786 , \21811 );
and \U$21567 ( \21813 , \21763 , \21785 );
or \U$21568 ( \21814 , \21812 , \21813 );
xor \U$21569 ( \21815 , \21307 , \21335 );
xnor \U$21570 ( \21816 , \21815 , \21367 );
xor \U$21571 ( \21817 , \21814 , \21816 );
xor \U$21572 ( \21818 , RIbe28a20_33, RIbe2a460_89);
not \U$21573 ( \21819 , \21818 );
not \U$21574 ( \21820 , \7795 );
or \U$21575 ( \21821 , \21819 , \21820 );
nand \U$21576 ( \21822 , \5055 , \21396 );
nand \U$21577 ( \21823 , \21821 , \21822 );
not \U$21578 ( \21824 , \21823 );
xor \U$21579 ( \21825 , RIbe295d8_58, RIbe2a550_91);
not \U$21580 ( \21826 , \21825 );
not \U$21581 ( \21827 , \10433 );
or \U$21582 ( \21828 , \21826 , \21827 );
nand \U$21583 ( \21829 , \20336 , \21412 );
nand \U$21584 ( \21830 , \21828 , \21829 );
not \U$21585 ( \21831 , \21830 );
or \U$21586 ( \21832 , \21824 , \21831 );
not \U$21587 ( \21833 , \21830 );
not \U$21588 ( \21834 , \21833 );
not \U$21589 ( \21835 , \21823 );
not \U$21590 ( \21836 , \21835 );
or \U$21591 ( \21837 , \21834 , \21836 );
not \U$21592 ( \21838 , \9524 );
not \U$21593 ( \21839 , \21838 );
not \U$21594 ( \21840 , \21391 );
and \U$21595 ( \21841 , \21839 , \21840 );
not \U$21596 ( \21842 , \7609 );
xnor \U$21597 ( \21843 , RIbe28f48_44, RIbe29ce0_73);
nor \U$21598 ( \21844 , \21842 , \21843 );
nor \U$21599 ( \21845 , \21841 , \21844 );
not \U$21600 ( \21846 , \21845 );
nand \U$21601 ( \21847 , \21837 , \21846 );
nand \U$21602 ( \21848 , \21832 , \21847 );
not \U$21603 ( \21849 , \21848 );
xor \U$21604 ( \21850 , RIbe2b108_116, RIbe294e8_56);
not \U$21605 ( \21851 , \21850 );
buf \U$21606 ( \21852 , \14296 );
not \U$21607 ( \21853 , \21852 );
or \U$21608 ( \21854 , \21851 , \21853 );
nand \U$21609 ( \21855 , \13534 , \21291 );
nand \U$21610 ( \21856 , \21854 , \21855 );
not \U$21611 ( \21857 , \21856 );
xor \U$21612 ( \21858 , RIbe28228_16, RIbe2b4c8_124);
not \U$21613 ( \21859 , \21858 );
not \U$21614 ( \21860 , \14638 );
or \U$21615 ( \21861 , \21859 , \21860 );
nand \U$21616 ( \21862 , \885 , \21284 );
nand \U$21617 ( \21863 , \21861 , \21862 );
xor \U$21618 ( \21864 , RIbe28c78_38, RIbe2b018_114);
not \U$21619 ( \21865 , \21864 );
not \U$21620 ( \21866 , \17570 );
or \U$21621 ( \21867 , \21865 , \21866 );
nand \U$21622 ( \21868 , \18777 , \21438 );
nand \U$21623 ( \21869 , \21867 , \21868 );
and \U$21624 ( \21870 , \21863 , \21869 );
not \U$21625 ( \21871 , \21863 );
not \U$21626 ( \21872 , \21869 );
and \U$21627 ( \21873 , \21871 , \21872 );
nor \U$21628 ( \21874 , \21870 , \21873 );
not \U$21629 ( \21875 , \21874 );
or \U$21630 ( \21876 , \21857 , \21875 );
not \U$21631 ( \21877 , \21872 );
nand \U$21632 ( \21878 , \21877 , \21863 );
nand \U$21633 ( \21879 , \21876 , \21878 );
xor \U$21634 ( \21880 , RIbe2a028_80, RIbe28d68_40);
not \U$21635 ( \21881 , \21880 );
not \U$21636 ( \21882 , \8401 );
or \U$21637 ( \21883 , \21881 , \21882 );
nand \U$21638 ( \21884 , \8172 , \21447 );
nand \U$21639 ( \21885 , \21883 , \21884 );
not \U$21640 ( \21886 , \21885 );
xor \U$21641 ( \21887 , RIbe2a190_83, RIbe297b8_62);
not \U$21642 ( \21888 , \21887 );
not \U$21643 ( \21889 , \15690 );
or \U$21644 ( \21890 , \21888 , \21889 );
nand \U$21645 ( \21891 , \15693 , \21381 );
nand \U$21646 ( \21892 , \21890 , \21891 );
not \U$21647 ( \21893 , \21892 );
or \U$21648 ( \21894 , \21886 , \21893 );
or \U$21649 ( \21895 , \21892 , \21885 );
xor \U$21650 ( \21896 , RIbe2a820_97, RIbe28480_21);
not \U$21651 ( \21897 , \21896 );
not \U$21652 ( \21898 , \3344 );
or \U$21653 ( \21899 , \21897 , \21898 );
nand \U$21654 ( \21900 , \2527 , \21456 );
nand \U$21655 ( \21901 , \21899 , \21900 );
nand \U$21656 ( \21902 , \21895 , \21901 );
nand \U$21657 ( \21903 , \21894 , \21902 );
xor \U$21658 ( \21904 , \21879 , \21903 );
not \U$21659 ( \21905 , \21904 );
or \U$21660 ( \21906 , \21849 , \21905 );
nand \U$21661 ( \21907 , \21879 , \21903 );
nand \U$21662 ( \21908 , \21906 , \21907 );
and \U$21663 ( \21909 , \21817 , \21908 );
and \U$21664 ( \21910 , \21814 , \21816 );
or \U$21665 ( \21911 , \21909 , \21910 );
not \U$21666 ( \21912 , \21911 );
or \U$21667 ( \21913 , \21737 , \21912 );
or \U$21668 ( \21914 , \21736 , \21911 );
nand \U$21669 ( \21915 , \21913 , \21914 );
not \U$21670 ( \21916 , \21915 );
or \U$21671 ( \21917 , \21734 , \21916 );
not \U$21672 ( \21918 , \21736 );
nand \U$21673 ( \21919 , \21918 , \21911 );
nand \U$21674 ( \21920 , \21917 , \21919 );
and \U$21675 ( \21921 , \21698 , \21920 );
and \U$21676 ( \21922 , \21696 , \21697 );
or \U$21677 ( \21923 , \21921 , \21922 );
not \U$21678 ( \21924 , \21923 );
not \U$21679 ( \21925 , \21181 );
not \U$21680 ( \21926 , \21925 );
not \U$21681 ( \21927 , \21493 );
or \U$21682 ( \21928 , \21926 , \21927 );
nand \U$21683 ( \21929 , \21492 , \21181 );
nand \U$21684 ( \21930 , \21928 , \21929 );
not \U$21685 ( \21931 , \21930 );
not \U$21686 ( \21932 , \21931 );
not \U$21687 ( \21933 , \21932 );
or \U$21688 ( \21934 , \21924 , \21933 );
not \U$21689 ( \21935 , \21923 );
not \U$21690 ( \21936 , \21935 );
not \U$21691 ( \21937 , \21931 );
or \U$21692 ( \21938 , \21936 , \21937 );
not \U$21693 ( \21939 , \21183 );
and \U$21694 ( \21940 , \21252 , \21259 );
not \U$21695 ( \21941 , \21252 );
and \U$21696 ( \21942 , \21941 , \21260 );
nor \U$21697 ( \21943 , \21940 , \21942 );
not \U$21698 ( \21944 , \21943 );
or \U$21699 ( \21945 , \21939 , \21944 );
or \U$21700 ( \21946 , \21943 , \21183 );
nand \U$21701 ( \21947 , \21945 , \21946 );
xor \U$21702 ( \21948 , \21512 , \21629 );
xor \U$21703 ( \21949 , \21947 , \21948 );
not \U$21704 ( \21950 , \21193 );
and \U$21705 ( \21951 , \21225 , \21950 );
not \U$21706 ( \21952 , \21225 );
and \U$21707 ( \21953 , \21952 , \21193 );
nor \U$21708 ( \21954 , \21951 , \21953 );
not \U$21709 ( \21955 , \21954 );
xor \U$21710 ( \21956 , \21272 , \21268 );
xnor \U$21711 ( \21957 , \21956 , \21266 );
not \U$21712 ( \21958 , \21957 );
and \U$21713 ( \21959 , \21955 , \21958 );
and \U$21714 ( \21960 , \21954 , \21957 );
nor \U$21715 ( \21961 , \21959 , \21960 );
not \U$21716 ( \21962 , \21961 );
not \U$21717 ( \21963 , \21962 );
xor \U$21718 ( \21964 , \21444 , \21452 );
xnor \U$21719 ( \21965 , \21964 , \21461 );
not \U$21720 ( \21966 , \21965 );
not \U$21721 ( \21967 , \21296 );
xor \U$21722 ( \21968 , \21305 , \21967 );
xnor \U$21723 ( \21969 , \21968 , \21289 );
not \U$21724 ( \21970 , \21969 );
or \U$21725 ( \21971 , \21966 , \21970 );
or \U$21726 ( \21972 , \21969 , \21965 );
nand \U$21727 ( \21973 , \21971 , \21972 );
not \U$21728 ( \21974 , \21973 );
xor \U$21729 ( \21975 , RIbe29f38_78, RIbe27fd0_11);
not \U$21730 ( \21976 , \21975 );
not \U$21731 ( \21977 , \12808 );
or \U$21732 ( \21978 , \21976 , \21977 );
nand \U$21733 ( \21979 , \2707 , \21530 );
nand \U$21734 ( \21980 , \21978 , \21979 );
not \U$21735 ( \21981 , \21980 );
xor \U$21736 ( \21982 , RIbe29e48_76, RIbe28cf0_39);
and \U$21737 ( \21983 , \21982 , \11039 );
and \U$21738 ( \21984 , \4849 , \21537 );
nor \U$21739 ( \21985 , \21983 , \21984 );
not \U$21740 ( \21986 , \21985 );
xor \U$21741 ( \21987 , RIbe29b00_69, RIbe2a910_99);
not \U$21742 ( \21988 , \21987 );
not \U$21743 ( \21989 , \9737 );
or \U$21744 ( \21990 , \21988 , \21989 );
xor \U$21745 ( \21991 , RIbe29128_48, RIbe2a910_99);
nand \U$21746 ( \21992 , \11456 , \21991 );
nand \U$21747 ( \21993 , \21990 , \21992 );
not \U$21748 ( \21994 , \21993 );
or \U$21749 ( \21995 , \21986 , \21994 );
or \U$21750 ( \21996 , \21985 , \21993 );
nand \U$21751 ( \21997 , \21995 , \21996 );
not \U$21752 ( \21998 , \21997 );
or \U$21753 ( \21999 , \21981 , \21998 );
not \U$21754 ( \22000 , \21985 );
nand \U$21755 ( \22001 , \22000 , \21993 );
nand \U$21756 ( \22002 , \21999 , \22001 );
not \U$21757 ( \22003 , \22002 );
xor \U$21758 ( \22004 , RIbe29218_50, RIbe2a3e8_88);
not \U$21759 ( \22005 , \22004 );
not \U$21760 ( \22006 , \9262 );
or \U$21761 ( \22007 , \22005 , \22006 );
nand \U$21762 ( \22008 , \8794 , \21764 );
nand \U$21763 ( \22009 , \22007 , \22008 );
xor \U$21764 ( \22010 , RIbe2aa78_102, RIbe27e68_8);
not \U$21765 ( \22011 , \22010 );
not \U$21766 ( \22012 , \2458 );
or \U$21767 ( \22013 , \22011 , \22012 );
xor \U$21768 ( \22014 , RIbe27e68_8, RIbe2b6a8_128);
nand \U$21769 ( \22015 , \2464 , \22014 );
nand \U$21770 ( \22016 , \22013 , \22015 );
nor \U$21771 ( \22017 , \22009 , \22016 );
xor \U$21772 ( \22018 , RIbe28228_16, RIbe2a6b8_94);
not \U$21773 ( \22019 , \22018 );
not \U$21774 ( \22020 , \3056 );
or \U$21775 ( \22021 , \22019 , \22020 );
nand \U$21776 ( \22022 , \8679 , \21858 );
nand \U$21777 ( \22023 , \22021 , \22022 );
not \U$21778 ( \22024 , \22023 );
or \U$21779 ( \22025 , \22017 , \22024 );
nand \U$21780 ( \22026 , \22016 , \22009 );
nand \U$21781 ( \22027 , \22025 , \22026 );
xor \U$21782 ( \22028 , RIbe28a20_33, RIbe2adc0_109);
not \U$21783 ( \22029 , \22028 );
not \U$21784 ( \22030 , \1780 );
or \U$21785 ( \22031 , \22029 , \22030 );
nand \U$21786 ( \22032 , \2475 , \21818 );
nand \U$21787 ( \22033 , \22031 , \22032 );
xor \U$21788 ( \22034 , RIbe288b8_30, RIbe2b180_117);
not \U$21789 ( \22035 , \22034 );
not \U$21790 ( \22036 , \15353 );
or \U$21791 ( \22037 , \22035 , \22036 );
nand \U$21792 ( \22038 , \16646 , \21755 );
nand \U$21793 ( \22039 , \22037 , \22038 );
or \U$21794 ( \22040 , \22033 , \22039 );
xor \U$21795 ( \22041 , RIbe28930_31, RIbe2b540_125);
not \U$21796 ( \22042 , \22041 );
not \U$21797 ( \22043 , \11374 );
or \U$21798 ( \22044 , \22042 , \22043 );
nand \U$21799 ( \22045 , \1797 , \21795 );
nand \U$21800 ( \22046 , \22044 , \22045 );
nand \U$21801 ( \22047 , \22040 , \22046 );
nand \U$21802 ( \22048 , \22033 , \22039 );
nand \U$21803 ( \22049 , \22047 , \22048 );
xor \U$21804 ( \22050 , \22027 , \22049 );
not \U$21805 ( \22051 , \22050 );
or \U$21806 ( \22052 , \22003 , \22051 );
nand \U$21807 ( \22053 , \22049 , \22027 );
nand \U$21808 ( \22054 , \22052 , \22053 );
not \U$21809 ( \22055 , \22054 );
or \U$21810 ( \22056 , \21974 , \22055 );
not \U$21811 ( \22057 , \21965 );
nand \U$21812 ( \22058 , \22057 , \21969 );
nand \U$21813 ( \22059 , \22056 , \22058 );
not \U$21814 ( \22060 , \22059 );
or \U$21815 ( \22061 , \21963 , \22060 );
not \U$21816 ( \22062 , \21954 );
nand \U$21817 ( \22063 , \22062 , \21957 );
nand \U$21818 ( \22064 , \22061 , \22063 );
not \U$21819 ( \22065 , \22064 );
xnor \U$21820 ( \22066 , \21617 , \21598 );
not \U$21821 ( \22067 , \22066 );
xor \U$21822 ( \22068 , \21235 , \21238 );
xor \U$21823 ( \22069 , \22068 , \21233 );
and \U$21824 ( \22070 , \21314 , \21322 );
not \U$21825 ( \22071 , \21314 );
and \U$21826 ( \22072 , \22071 , \21321 );
or \U$21827 ( \22073 , \22070 , \22072 );
and \U$21828 ( \22074 , \22073 , \21330 );
not \U$21829 ( \22075 , \22073 );
not \U$21830 ( \22076 , \21330 );
and \U$21831 ( \22077 , \22075 , \22076 );
nor \U$21832 ( \22078 , \22074 , \22077 );
not \U$21833 ( \22079 , \22078 );
xor \U$21834 ( \22080 , \21386 , \21406 );
not \U$21835 ( \22081 , \22080 );
or \U$21836 ( \22082 , \22079 , \22081 );
or \U$21837 ( \22083 , \22080 , \22078 );
not \U$21838 ( \22084 , \21214 );
nor \U$21839 ( \22085 , \22084 , \21208 );
xor \U$21840 ( \22086 , \22085 , \21212 );
not \U$21841 ( \22087 , \22086 );
nand \U$21842 ( \22088 , \22083 , \22087 );
nand \U$21843 ( \22089 , \22082 , \22088 );
xor \U$21844 ( \22090 , \22069 , \22089 );
xor \U$21845 ( \22091 , \20608 , \20616 );
xor \U$21846 ( \22092 , \22091 , \20602 );
not \U$21847 ( \22093 , \22092 );
not \U$21848 ( \22094 , \21991 );
not \U$21849 ( \22095 , \13325 );
or \U$21850 ( \22096 , \22094 , \22095 );
nand \U$21851 ( \22097 , \10401 , \21353 );
nand \U$21852 ( \22098 , \22096 , \22097 );
not \U$21853 ( \22099 , \22098 );
xor \U$21854 ( \22100 , RIbe27b20_1, RIbe29c68_72);
not \U$21855 ( \22101 , \22100 );
not \U$21856 ( \22102 , \7513 );
or \U$21857 ( \22103 , \22101 , \22102 );
nand \U$21858 ( \22104 , \4580 , \21338 );
nand \U$21859 ( \22105 , \22103 , \22104 );
not \U$21860 ( \22106 , \22105 );
not \U$21861 ( \22107 , \22106 );
not \U$21862 ( \22108 , \22014 );
not \U$21863 ( \22109 , \2458 );
or \U$21864 ( \22110 , \22108 , \22109 );
nand \U$21865 ( \22111 , \2603 , \20644 );
nand \U$21866 ( \22112 , \22110 , \22111 );
not \U$21867 ( \22113 , \22112 );
or \U$21868 ( \22114 , \22107 , \22113 );
or \U$21869 ( \22115 , \22112 , \22106 );
nand \U$21870 ( \22116 , \22114 , \22115 );
not \U$21871 ( \22117 , \22116 );
or \U$21872 ( \22118 , \22099 , \22117 );
nand \U$21873 ( \22119 , \22112 , \22105 );
nand \U$21874 ( \22120 , \22118 , \22119 );
not \U$21875 ( \22121 , \21343 );
not \U$21876 ( \22122 , \21362 );
not \U$21877 ( \22123 , \22122 );
or \U$21878 ( \22124 , \22121 , \22123 );
not \U$21879 ( \22125 , \21343 );
nand \U$21880 ( \22126 , \22125 , \21362 );
nand \U$21881 ( \22127 , \22124 , \22126 );
xor \U$21882 ( \22128 , \22120 , \22127 );
not \U$21883 ( \22129 , \22128 );
or \U$21884 ( \22130 , \22093 , \22129 );
nand \U$21885 ( \22131 , \22120 , \22127 );
nand \U$21886 ( \22132 , \22130 , \22131 );
and \U$21887 ( \22133 , \22090 , \22132 );
and \U$21888 ( \22134 , \22069 , \22089 );
or \U$21889 ( \22135 , \22133 , \22134 );
not \U$21890 ( \22136 , \22135 );
or \U$21891 ( \22137 , \22067 , \22136 );
or \U$21892 ( \22138 , \22135 , \22066 );
nand \U$21893 ( \22139 , \22137 , \22138 );
not \U$21894 ( \22140 , \22139 );
or \U$21895 ( \22141 , \22065 , \22140 );
not \U$21896 ( \22142 , \22066 );
nand \U$21897 ( \22143 , \22142 , \22135 );
nand \U$21898 ( \22144 , \22141 , \22143 );
and \U$21899 ( \22145 , \21949 , \22144 );
and \U$21900 ( \22146 , \21947 , \21948 );
or \U$21901 ( \22147 , \22145 , \22146 );
nand \U$21902 ( \22148 , \21938 , \22147 );
nand \U$21903 ( \22149 , \21934 , \22148 );
buf \U$21904 ( \22150 , \22149 );
xor \U$21905 ( \22151 , \20518 , \20720 );
nor \U$21906 ( \22152 , \22150 , \22151 );
xor \U$21907 ( \22153 , \21499 , \21179 );
not \U$21908 ( \22154 , \21652 );
xor \U$21909 ( \22155 , \22153 , \22154 );
or \U$21910 ( \22156 , \22152 , \22155 );
nand \U$21911 ( \22157 , \22150 , \22151 );
nand \U$21912 ( \22158 , \22156 , \22157 );
or \U$21913 ( \22159 , \21687 , \22158 );
and \U$21914 ( \22160 , \21682 , \22159 );
not \U$21915 ( \22161 , \20123 );
not \U$21916 ( \22162 , \22161 );
not \U$21917 ( \22163 , \19675 );
or \U$21918 ( \22164 , \22162 , \22163 );
not \U$21919 ( \22165 , \19553 );
nand \U$21920 ( \22166 , \22165 , \19671 );
nand \U$21921 ( \22167 , \22164 , \22166 );
not \U$21922 ( \22168 , \21046 );
not \U$21923 ( \22169 , \21063 );
or \U$21924 ( \22170 , \22168 , \22169 );
not \U$21925 ( \22171 , \21052 );
nand \U$21926 ( \22172 , \22171 , \21059 );
nand \U$21927 ( \22173 , \22170 , \22172 );
xor \U$21928 ( \22174 , \17797 , \17900 );
xor \U$21929 ( \22175 , \22173 , \22174 );
xor \U$21930 ( \22176 , \21098 , \21114 );
and \U$21931 ( \22177 , \22176 , \21117 );
and \U$21932 ( \22178 , \21098 , \21114 );
or \U$21933 ( \22179 , \22177 , \22178 );
xor \U$21934 ( \22180 , \22175 , \22179 );
not \U$21935 ( \22181 , \22180 );
not \U$21936 ( \22182 , \22181 );
not \U$21937 ( \22183 , \19930 );
not \U$21938 ( \22184 , \19935 );
or \U$21939 ( \22185 , \22183 , \22184 );
not \U$21940 ( \22186 , \19932 );
nand \U$21941 ( \22187 , \22186 , \19934 );
nand \U$21942 ( \22188 , \22185 , \22187 );
not \U$21943 ( \22189 , \22188 );
not \U$21944 ( \22190 , \22189 );
not \U$21945 ( \22191 , \19648 );
not \U$21946 ( \22192 , \19641 );
or \U$21947 ( \22193 , \22191 , \22192 );
not \U$21948 ( \22194 , \19649 );
not \U$21949 ( \22195 , \19645 );
or \U$21950 ( \22196 , \22194 , \22195 );
nand \U$21951 ( \22197 , \22196 , \19656 );
nand \U$21952 ( \22198 , \22193 , \22197 );
not \U$21953 ( \22199 , \22198 );
not \U$21954 ( \22200 , \22199 );
not \U$21955 ( \22201 , \17942 );
not \U$21956 ( \22202 , \17991 );
not \U$21957 ( \22203 , \22202 );
or \U$21958 ( \22204 , \22201 , \22203 );
nand \U$21959 ( \22205 , \17943 , \17991 );
nand \U$21960 ( \22206 , \22204 , \22205 );
and \U$21961 ( \22207 , \22206 , \17969 );
not \U$21962 ( \22208 , \22206 );
and \U$21963 ( \22209 , \22208 , \17970 );
nor \U$21964 ( \22210 , \22207 , \22209 );
not \U$21965 ( \22211 , \22210 );
or \U$21966 ( \22212 , \22200 , \22211 );
or \U$21967 ( \22213 , \22210 , \22199 );
nand \U$21968 ( \22214 , \22212 , \22213 );
buf \U$21969 ( \22215 , \22214 );
not \U$21970 ( \22216 , \22215 );
or \U$21971 ( \22217 , \22190 , \22216 );
or \U$21972 ( \22218 , \22215 , \22189 );
nand \U$21973 ( \22219 , \22217 , \22218 );
not \U$21974 ( \22220 , \22219 );
not \U$21975 ( \22221 , \19562 );
not \U$21976 ( \22222 , \19568 );
or \U$21977 ( \22223 , \22221 , \22222 );
or \U$21978 ( \22224 , \19562 , \19568 );
nand \U$21979 ( \22225 , \22224 , \19625 );
nand \U$21980 ( \22226 , \22223 , \22225 );
not \U$21981 ( \22227 , \22226 );
not \U$21982 ( \22228 , \22227 );
not \U$21983 ( \22229 , \19629 );
not \U$21984 ( \22230 , \19662 );
or \U$21985 ( \22231 , \22229 , \22230 );
nand \U$21986 ( \22232 , \22231 , \19635 );
not \U$21987 ( \22233 , \19662 );
not \U$21988 ( \22234 , \19629 );
nand \U$21989 ( \22235 , \22233 , \22234 );
nand \U$21990 ( \22236 , \22232 , \22235 );
not \U$21991 ( \22237 , \22236 );
or \U$21992 ( \22238 , \22228 , \22237 );
or \U$21993 ( \22239 , \22227 , \22236 );
nand \U$21994 ( \22240 , \22238 , \22239 );
not \U$21995 ( \22241 , \22240 );
not \U$21996 ( \22242 , \22241 );
or \U$21997 ( \22243 , \22220 , \22242 );
not \U$21998 ( \22244 , \22219 );
nand \U$21999 ( \22245 , \22244 , \22240 );
nand \U$22000 ( \22246 , \22243 , \22245 );
not \U$22001 ( \22247 , \21093 );
not \U$22002 ( \22248 , \21118 );
or \U$22003 ( \22249 , \22247 , \22248 );
or \U$22004 ( \22250 , \21118 , \21093 );
nand \U$22005 ( \22251 , \22250 , \21087 );
nand \U$22006 ( \22252 , \22249 , \22251 );
and \U$22007 ( \22253 , \22246 , \22252 );
not \U$22008 ( \22254 , \22246 );
not \U$22009 ( \22255 , \22252 );
and \U$22010 ( \22256 , \22254 , \22255 );
nor \U$22011 ( \22257 , \22253 , \22256 );
not \U$22012 ( \22258 , \22257 );
or \U$22013 ( \22259 , \22182 , \22258 );
not \U$22014 ( \22260 , \22257 );
nand \U$22015 ( \22261 , \22260 , \22180 );
nand \U$22016 ( \22262 , \22259 , \22261 );
xor \U$22017 ( \22263 , \18203 , \18208 );
xor \U$22018 ( \22264 , \22263 , \18214 );
xor \U$22019 ( \22265 , \18245 , \18247 );
xor \U$22020 ( \22266 , \22265 , \18263 );
xor \U$22021 ( \22267 , \22264 , \22266 );
not \U$22022 ( \22268 , \18018 );
not \U$22023 ( \22269 , \18027 );
or \U$22024 ( \22270 , \22268 , \22269 );
or \U$22025 ( \22271 , \18027 , \18018 );
nand \U$22026 ( \22272 , \22270 , \22271 );
xor \U$22027 ( \22273 , \22267 , \22272 );
not \U$22028 ( \22274 , \22273 );
xor \U$22029 ( \22275 , \21041 , \21068 );
and \U$22030 ( \22276 , \22275 , \21075 );
and \U$22031 ( \22277 , \21041 , \21068 );
or \U$22032 ( \22278 , \22276 , \22277 );
not \U$22033 ( \22279 , \22278 );
not \U$22034 ( \22280 , \22279 );
or \U$22035 ( \22281 , \22274 , \22280 );
not \U$22036 ( \22282 , \22273 );
nand \U$22037 ( \22283 , \22282 , \22278 );
nand \U$22038 ( \22284 , \22281 , \22283 );
xor \U$22039 ( \22285 , \19626 , \19664 );
and \U$22040 ( \22286 , \22285 , \19669 );
and \U$22041 ( \22287 , \19626 , \19664 );
or \U$22042 ( \22288 , \22286 , \22287 );
and \U$22043 ( \22289 , \22284 , \22288 );
not \U$22044 ( \22290 , \22284 );
not \U$22045 ( \22291 , \22288 );
and \U$22046 ( \22292 , \22290 , \22291 );
nor \U$22047 ( \22293 , \22289 , \22292 );
xor \U$22048 ( \22294 , \22262 , \22293 );
not \U$22049 ( \22295 , \22294 );
nand \U$22050 ( \22296 , \17634 , \17587 );
nand \U$22051 ( \22297 , \17703 , \22296 );
buf \U$22052 ( \22298 , \17700 );
and \U$22053 ( \22299 , \22297 , \22298 );
not \U$22054 ( \22300 , \22297 );
not \U$22055 ( \22301 , \22298 );
and \U$22056 ( \22302 , \22300 , \22301 );
nor \U$22057 ( \22303 , \22299 , \22302 );
not \U$22058 ( \22304 , \22303 );
xor \U$22059 ( \22305 , \19915 , \19927 );
and \U$22060 ( \22306 , \22305 , \19936 );
and \U$22061 ( \22307 , \19915 , \19927 );
or \U$22062 ( \22308 , \22306 , \22307 );
not \U$22063 ( \22309 , \22308 );
or \U$22064 ( \22310 , \22304 , \22309 );
or \U$22065 ( \22311 , \22308 , \22303 );
nand \U$22066 ( \22312 , \22310 , \22311 );
not \U$22067 ( \22313 , \19919 );
nand \U$22068 ( \22314 , \19926 , \22313 );
and \U$22069 ( \22315 , \22314 , \19917 );
nor \U$22070 ( \22316 , \22313 , \19926 );
nor \U$22071 ( \22317 , \22315 , \22316 );
not \U$22072 ( \22318 , \21099 );
not \U$22073 ( \22319 , \21113 );
or \U$22074 ( \22320 , \22318 , \22319 );
nand \U$22075 ( \22321 , \21103 , \21112 );
nand \U$22076 ( \22322 , \22320 , \22321 );
not \U$22077 ( \22323 , \22322 );
xnor \U$22078 ( \22324 , \22317 , \22323 );
xor \U$22079 ( \22325 , \18035 , \18038 );
xor \U$22080 ( \22326 , \22325 , \18040 );
not \U$22081 ( \22327 , \22326 );
and \U$22082 ( \22328 , \22324 , \22327 );
not \U$22083 ( \22329 , \22324 );
and \U$22084 ( \22330 , \22329 , \22326 );
nor \U$22085 ( \22331 , \22328 , \22330 );
xor \U$22086 ( \22332 , \22312 , \22331 );
not \U$22087 ( \22333 , \22332 );
or \U$22088 ( \22334 , \20121 , \19937 );
nand \U$22089 ( \22335 , \22334 , \19913 );
nand \U$22090 ( \22336 , \20121 , \19937 );
nand \U$22091 ( \22337 , \22335 , \22336 );
not \U$22092 ( \22338 , \22337 );
not \U$22093 ( \22339 , \22338 );
or \U$22094 ( \22340 , \22333 , \22339 );
not \U$22095 ( \22341 , \22335 );
not \U$22096 ( \22342 , \22336 );
or \U$22097 ( \22343 , \22341 , \22342 );
not \U$22098 ( \22344 , \22332 );
nand \U$22099 ( \22345 , \22343 , \22344 );
nand \U$22100 ( \22346 , \22340 , \22345 );
not \U$22101 ( \22347 , \21035 );
not \U$22102 ( \22348 , \21077 );
or \U$22103 ( \22349 , \22347 , \22348 );
nand \U$22104 ( \22350 , \22349 , \21123 );
nand \U$22105 ( \22351 , \22350 , \21080 );
and \U$22106 ( \22352 , \22346 , \22351 );
not \U$22107 ( \22353 , \22346 );
not \U$22108 ( \22354 , \22351 );
and \U$22109 ( \22355 , \22353 , \22354 );
nor \U$22110 ( \22356 , \22352 , \22355 );
not \U$22111 ( \22357 , \22356 );
and \U$22112 ( \22358 , \22295 , \22357 );
and \U$22113 ( \22359 , \22294 , \22356 );
nor \U$22114 ( \22360 , \22358 , \22359 );
xor \U$22115 ( \22361 , \22167 , \22360 );
nand \U$22116 ( \22362 , \21147 , \21172 );
not \U$22117 ( \22363 , \21140 );
not \U$22118 ( \22364 , \21142 );
or \U$22119 ( \22365 , \22363 , \22364 );
nand \U$22120 ( \22366 , \22365 , \21128 );
nand \U$22121 ( \22367 , \22362 , \22366 );
xnor \U$22122 ( \22368 , \22361 , \22367 );
xnor \U$22123 ( \22369 , \21147 , \21171 );
not \U$22124 ( \22370 , \22369 );
not \U$22125 ( \22371 , \20955 );
not \U$22126 ( \22372 , \20127 );
not \U$22127 ( \22373 , \22372 );
or \U$22128 ( \22374 , \22371 , \22373 );
or \U$22129 ( \22375 , \20955 , \22372 );
nand \U$22130 ( \22376 , \22374 , \22375 );
not \U$22131 ( \22377 , \22376 );
or \U$22132 ( \22378 , \22370 , \22377 );
not \U$22133 ( \22379 , \20955 );
nand \U$22134 ( \22380 , \22379 , \22372 );
nand \U$22135 ( \22381 , \22378 , \22380 );
nand \U$22136 ( \22382 , \22368 , \22381 );
nand \U$22137 ( \22383 , \22367 , \22167 );
not \U$22138 ( \22384 , \22383 );
not \U$22139 ( \22385 , \22167 );
nand \U$22140 ( \22386 , \22385 , \22367 );
not \U$22141 ( \22387 , \22386 );
nand \U$22142 ( \22388 , \22362 , \22366 , \22167 );
not \U$22143 ( \22389 , \22388 );
or \U$22144 ( \22390 , \22387 , \22389 );
not \U$22145 ( \22391 , \22360 );
nand \U$22146 ( \22392 , \22390 , \22391 );
not \U$22147 ( \22393 , \22392 );
or \U$22148 ( \22394 , \22384 , \22393 );
not \U$22149 ( \22395 , \22252 );
not \U$22150 ( \22396 , \22246 );
or \U$22151 ( \22397 , \22395 , \22396 );
or \U$22152 ( \22398 , \22246 , \22252 );
nand \U$22153 ( \22399 , \22398 , \22180 );
nand \U$22154 ( \22400 , \22397 , \22399 );
not \U$22155 ( \22401 , \22188 );
not \U$22156 ( \22402 , \22214 );
or \U$22157 ( \22403 , \22401 , \22402 );
nand \U$22158 ( \22404 , \22210 , \22198 );
nand \U$22159 ( \22405 , \22403 , \22404 );
xor \U$22160 ( \22406 , \22264 , \22266 );
and \U$22161 ( \22407 , \22406 , \22272 );
and \U$22162 ( \22408 , \22264 , \22266 );
or \U$22163 ( \22409 , \22407 , \22408 );
xor \U$22164 ( \22410 , \22405 , \22409 );
not \U$22165 ( \22411 , \18032 );
not \U$22166 ( \22412 , \22411 );
not \U$22167 ( \22413 , \18054 );
or \U$22168 ( \22414 , \22412 , \22413 );
or \U$22169 ( \22415 , \18054 , \22411 );
nand \U$22170 ( \22416 , \22414 , \22415 );
xor \U$22171 ( \22417 , \22410 , \22416 );
xor \U$22172 ( \22418 , \22400 , \22417 );
not \U$22173 ( \22419 , \22331 );
not \U$22174 ( \22420 , \22312 );
or \U$22175 ( \22421 , \22419 , \22420 );
not \U$22176 ( \22422 , \22303 );
nand \U$22177 ( \22423 , \22422 , \22308 );
nand \U$22178 ( \22424 , \22421 , \22423 );
xor \U$22179 ( \22425 , \18267 , \18238 );
not \U$22180 ( \22426 , \22425 );
nand \U$22181 ( \22427 , \22175 , \22179 );
not \U$22182 ( \22428 , \22427 );
and \U$22183 ( \22429 , \22173 , \22174 );
nor \U$22184 ( \22430 , \22428 , \22429 );
not \U$22185 ( \22431 , \22430 );
or \U$22186 ( \22432 , \22426 , \22431 );
not \U$22187 ( \22433 , \22429 );
not \U$22188 ( \22434 , \22433 );
not \U$22189 ( \22435 , \22427 );
or \U$22190 ( \22436 , \22434 , \22435 );
not \U$22191 ( \22437 , \22425 );
nand \U$22192 ( \22438 , \22436 , \22437 );
nand \U$22193 ( \22439 , \22432 , \22438 );
xor \U$22194 ( \22440 , \22424 , \22439 );
xnor \U$22195 ( \22441 , \22418 , \22440 );
or \U$22196 ( \22442 , \22293 , \22262 );
and \U$22197 ( \22443 , \22442 , \22356 );
and \U$22198 ( \22444 , \22262 , \22293 );
nor \U$22199 ( \22445 , \22443 , \22444 );
xor \U$22200 ( \22446 , \22441 , \22445 );
not \U$22201 ( \22447 , \22317 );
not \U$22202 ( \22448 , \22447 );
not \U$22203 ( \22449 , \22322 );
or \U$22204 ( \22450 , \22448 , \22449 );
not \U$22205 ( \22451 , \22323 );
not \U$22206 ( \22452 , \22317 );
or \U$22207 ( \22453 , \22451 , \22452 );
nand \U$22208 ( \22454 , \22453 , \22326 );
nand \U$22209 ( \22455 , \22450 , \22454 );
xor \U$22210 ( \22456 , \18217 , \18219 );
xor \U$22211 ( \22457 , \22456 , \18225 );
xor \U$22212 ( \22458 , \22455 , \22457 );
not \U$22213 ( \22459 , \18083 );
not \U$22214 ( \22460 , \22459 );
not \U$22215 ( \22461 , \18076 );
not \U$22216 ( \22462 , \18086 );
or \U$22217 ( \22463 , \22461 , \22462 );
or \U$22218 ( \22464 , \18086 , \18076 );
nand \U$22219 ( \22465 , \22463 , \22464 );
not \U$22220 ( \22466 , \22465 );
or \U$22221 ( \22467 , \22460 , \22466 );
or \U$22222 ( \22468 , \22465 , \22459 );
nand \U$22223 ( \22469 , \22467 , \22468 );
buf \U$22224 ( \22470 , \22469 );
xor \U$22225 ( \22471 , \22458 , \22470 );
not \U$22226 ( \22472 , \22471 );
not \U$22227 ( \22473 , \17704 );
not \U$22228 ( \22474 , \17906 );
or \U$22229 ( \22475 , \22473 , \22474 );
or \U$22230 ( \22476 , \17906 , \17704 );
nand \U$22231 ( \22477 , \22475 , \22476 );
and \U$22232 ( \22478 , \22477 , \18007 );
not \U$22233 ( \22479 , \22477 );
not \U$22234 ( \22480 , \18007 );
and \U$22235 ( \22481 , \22479 , \22480 );
nor \U$22236 ( \22482 , \22478 , \22481 );
not \U$22237 ( \22483 , \22219 );
not \U$22238 ( \22484 , \22240 );
or \U$22239 ( \22485 , \22483 , \22484 );
not \U$22240 ( \22486 , \22227 );
nand \U$22241 ( \22487 , \22486 , \22236 );
nand \U$22242 ( \22488 , \22485 , \22487 );
xor \U$22243 ( \22489 , \22482 , \22488 );
not \U$22244 ( \22490 , \22489 );
or \U$22245 ( \22491 , \22472 , \22490 );
or \U$22246 ( \22492 , \22489 , \22471 );
nand \U$22247 ( \22493 , \22491 , \22492 );
not \U$22248 ( \22494 , \22288 );
not \U$22249 ( \22495 , \22284 );
or \U$22250 ( \22496 , \22494 , \22495 );
nand \U$22251 ( \22497 , \22278 , \22273 );
nand \U$22252 ( \22498 , \22496 , \22497 );
nor \U$22253 ( \22499 , \22493 , \22498 );
not \U$22254 ( \22500 , \22499 );
nand \U$22255 ( \22501 , \22493 , \22498 );
nand \U$22256 ( \22502 , \22500 , \22501 );
not \U$22257 ( \22503 , \22351 );
not \U$22258 ( \22504 , \22346 );
or \U$22259 ( \22505 , \22503 , \22504 );
not \U$22260 ( \22506 , \22336 );
not \U$22261 ( \22507 , \22335 );
or \U$22262 ( \22508 , \22506 , \22507 );
nand \U$22263 ( \22509 , \22508 , \22332 );
nand \U$22264 ( \22510 , \22505 , \22509 );
xor \U$22265 ( \22511 , \22502 , \22510 );
xor \U$22266 ( \22512 , \22446 , \22511 );
nand \U$22267 ( \22513 , \22394 , \22512 );
and \U$22268 ( \22514 , \22382 , \22513 );
xor \U$22269 ( \22515 , \18178 , \18175 );
xnor \U$22270 ( \22516 , \22515 , \18285 );
xor \U$22271 ( \22517 , \18277 , \18279 );
xor \U$22272 ( \22518 , \22517 , \18282 );
not \U$22273 ( \22519 , \22518 );
not \U$22274 ( \22520 , \22519 );
buf \U$22275 ( \22521 , \18228 );
xor \U$22276 ( \22522 , \18230 , \22521 );
buf \U$22277 ( \22523 , \18272 );
xnor \U$22278 ( \22524 , \22522 , \22523 );
not \U$22279 ( \22525 , \22524 );
not \U$22280 ( \22526 , \22525 );
xor \U$22281 ( \22527 , \18100 , \18015 );
not \U$22282 ( \22528 , \22527 );
not \U$22283 ( \22529 , \22528 );
or \U$22284 ( \22530 , \22526 , \22529 );
not \U$22285 ( \22531 , \22524 );
not \U$22286 ( \22532 , \22527 );
or \U$22287 ( \22533 , \22531 , \22532 );
not \U$22288 ( \22534 , \22424 );
not \U$22289 ( \22535 , \22439 );
or \U$22290 ( \22536 , \22534 , \22535 );
not \U$22291 ( \22537 , \22433 );
not \U$22292 ( \22538 , \22427 );
or \U$22293 ( \22539 , \22537 , \22538 );
nand \U$22294 ( \22540 , \22539 , \22425 );
nand \U$22295 ( \22541 , \22536 , \22540 );
not \U$22296 ( \22542 , \22541 );
nand \U$22297 ( \22543 , \22533 , \22542 );
nand \U$22298 ( \22544 , \22530 , \22543 );
not \U$22299 ( \22545 , \22544 );
or \U$22300 ( \22546 , \22520 , \22545 );
xor \U$22301 ( \22547 , \18137 , \18140 );
xor \U$22302 ( \22548 , \22547 , \18135 );
not \U$22303 ( \22549 , \22548 );
xor \U$22304 ( \22550 , \22405 , \22409 );
and \U$22305 ( \22551 , \22550 , \22416 );
and \U$22306 ( \22552 , \22405 , \22409 );
or \U$22307 ( \22553 , \22551 , \22552 );
not \U$22308 ( \22554 , \22553 );
not \U$22309 ( \22555 , \22455 );
nand \U$22310 ( \22556 , \22555 , \22469 );
not \U$22311 ( \22557 , \22556 );
not \U$22312 ( \22558 , \22457 );
or \U$22313 ( \22559 , \22557 , \22558 );
not \U$22314 ( \22560 , \22469 );
nand \U$22315 ( \22561 , \22560 , \22455 );
nand \U$22316 ( \22562 , \22559 , \22561 );
not \U$22317 ( \22563 , \22562 );
and \U$22318 ( \22564 , \22554 , \22563 );
not \U$22319 ( \22565 , \22554 );
and \U$22320 ( \22566 , \22565 , \22562 );
nor \U$22321 ( \22567 , \22564 , \22566 );
not \U$22322 ( \22568 , \22567 );
or \U$22323 ( \22569 , \22549 , \22568 );
not \U$22324 ( \22570 , \22554 );
nand \U$22325 ( \22571 , \22570 , \22562 );
nand \U$22326 ( \22572 , \22569 , \22571 );
nand \U$22327 ( \22573 , \22546 , \22572 );
not \U$22328 ( \22574 , \22519 );
not \U$22329 ( \22575 , \22544 );
nand \U$22330 ( \22576 , \22574 , \22575 );
and \U$22331 ( \22577 , \22573 , \22576 );
xor \U$22332 ( \22578 , \22516 , \22577 );
nand \U$22333 ( \22579 , \18170 , \18172 );
and \U$22334 ( \22580 , \22579 , \18151 );
not \U$22335 ( \22581 , \22579 );
not \U$22336 ( \22582 , \18151 );
and \U$22337 ( \22583 , \22581 , \22582 );
nor \U$22338 ( \22584 , \22580 , \22583 );
xor \U$22339 ( \22585 , \22578 , \22584 );
not \U$22340 ( \22586 , \18149 );
not \U$22341 ( \22587 , \22586 );
not \U$22342 ( \22588 , \18122 );
not \U$22343 ( \22589 , \22588 );
or \U$22344 ( \22590 , \22587 , \22589 );
nand \U$22345 ( \22591 , \18149 , \18122 );
nand \U$22346 ( \22592 , \22590 , \22591 );
not \U$22347 ( \22593 , \22592 );
xor \U$22348 ( \22594 , \22518 , \22572 );
and \U$22349 ( \22595 , \22594 , \22575 );
not \U$22350 ( \22596 , \22594 );
and \U$22351 ( \22597 , \22596 , \22544 );
nor \U$22352 ( \22598 , \22595 , \22597 );
not \U$22353 ( \22599 , \22598 );
or \U$22354 ( \22600 , \22593 , \22599 );
or \U$22355 ( \22601 , \22598 , \22592 );
not \U$22356 ( \22602 , \22440 );
not \U$22357 ( \22603 , \22418 );
or \U$22358 ( \22604 , \22602 , \22603 );
nand \U$22359 ( \22605 , \22400 , \22417 );
nand \U$22360 ( \22606 , \22604 , \22605 );
not \U$22361 ( \22607 , \22606 );
not \U$22362 ( \22608 , \22471 );
and \U$22363 ( \22609 , \22489 , \22608 );
and \U$22364 ( \22610 , \22482 , \22488 );
nor \U$22365 ( \22611 , \22609 , \22610 );
not \U$22366 ( \22612 , \22611 );
not \U$22367 ( \22613 , \22548 );
not \U$22368 ( \22614 , \22567 );
not \U$22369 ( \22615 , \22614 );
or \U$22370 ( \22616 , \22613 , \22615 );
not \U$22371 ( \22617 , \22548 );
nand \U$22372 ( \22618 , \22617 , \22567 );
nand \U$22373 ( \22619 , \22616 , \22618 );
not \U$22374 ( \22620 , \22619 );
or \U$22375 ( \22621 , \22612 , \22620 );
or \U$22376 ( \22622 , \22619 , \22611 );
nand \U$22377 ( \22623 , \22621 , \22622 );
not \U$22378 ( \22624 , \22623 );
or \U$22379 ( \22625 , \22607 , \22624 );
not \U$22380 ( \22626 , \22611 );
nand \U$22381 ( \22627 , \22626 , \22619 );
nand \U$22382 ( \22628 , \22625 , \22627 );
nand \U$22383 ( \22629 , \22601 , \22628 );
nand \U$22384 ( \22630 , \22600 , \22629 );
not \U$22385 ( \22631 , \22630 );
nand \U$22386 ( \22632 , \22585 , \22631 );
not \U$22387 ( \22633 , \17515 );
and \U$22388 ( \22634 , \18298 , \22633 );
not \U$22389 ( \22635 , \18298 );
and \U$22390 ( \22636 , \22635 , \17515 );
nor \U$22391 ( \22637 , \22634 , \22636 );
xor \U$22392 ( \22638 , \22516 , \22577 );
and \U$22393 ( \22639 , \22638 , \22584 );
and \U$22394 ( \22640 , \22516 , \22577 );
or \U$22395 ( \22641 , \22639 , \22640 );
nand \U$22396 ( \22642 , \22637 , \22641 );
nand \U$22397 ( \22643 , \22632 , \22642 );
not \U$22398 ( \22644 , \22643 );
and \U$22399 ( \22645 , \22541 , \22525 );
not \U$22400 ( \22646 , \22541 );
and \U$22401 ( \22647 , \22646 , \22524 );
nor \U$22402 ( \22648 , \22645 , \22647 );
buf \U$22403 ( \22649 , \22528 );
not \U$22404 ( \22650 , \22649 );
and \U$22405 ( \22651 , \22648 , \22650 );
not \U$22406 ( \22652 , \22648 );
and \U$22407 ( \22653 , \22652 , \22649 );
nor \U$22408 ( \22654 , \22651 , \22653 );
not \U$22409 ( \22655 , \22499 );
not \U$22410 ( \22656 , \22655 );
not \U$22411 ( \22657 , \22510 );
or \U$22412 ( \22658 , \22656 , \22657 );
nand \U$22413 ( \22659 , \22658 , \22501 );
not \U$22414 ( \22660 , \22659 );
xor \U$22415 ( \22661 , \22654 , \22660 );
xor \U$22416 ( \22662 , \22611 , \22619 );
xor \U$22417 ( \22663 , \22662 , \22606 );
xor \U$22418 ( \22664 , \22661 , \22663 );
xor \U$22419 ( \22665 , \22441 , \22445 );
and \U$22420 ( \22666 , \22665 , \22511 );
and \U$22421 ( \22667 , \22441 , \22445 );
or \U$22422 ( \22668 , \22666 , \22667 );
nand \U$22423 ( \22669 , \22664 , \22668 );
xor \U$22424 ( \22670 , \22592 , \22598 );
xnor \U$22425 ( \22671 , \22670 , \22628 );
xor \U$22426 ( \22672 , \22654 , \22660 );
and \U$22427 ( \22673 , \22672 , \22663 );
and \U$22428 ( \22674 , \22654 , \22660 );
or \U$22429 ( \22675 , \22673 , \22674 );
nand \U$22430 ( \22676 , \22671 , \22675 );
nand \U$22431 ( \22677 , \22669 , \22676 );
not \U$22432 ( \22678 , \22677 );
and \U$22433 ( \22679 , \22160 , \22514 , \22644 , \22678 );
not \U$22434 ( \22680 , \22679 );
xor \U$22435 ( \22681 , RIbe29470_55, RIbe2aaf0_103);
not \U$22436 ( \22682 , \22681 );
not \U$22437 ( \22683 , \18832 );
or \U$22438 ( \22684 , \22682 , \22683 );
xor \U$22439 ( \22685 , RIbe294e8_56, RIbe2aaf0_103);
nand \U$22440 ( \22686 , \22685 , RIbe2ab68_104);
nand \U$22441 ( \22687 , \22684 , \22686 );
xor \U$22442 ( \22688 , RIbe27c88_4, RIbe2a190_83);
not \U$22443 ( \22689 , \22688 );
not \U$22444 ( \22690 , \10831 );
or \U$22445 ( \22691 , \22689 , \22690 );
xor \U$22446 ( \22692 , RIbe27df0_7, RIbe2a190_83);
nand \U$22447 ( \22693 , \10834 , \22692 );
nand \U$22448 ( \22694 , \22691 , \22693 );
buf \U$22449 ( \22695 , \22694 );
xor \U$22450 ( \22696 , \22687 , \22695 );
xor \U$22451 ( \22697 , RIbe29c68_72, RIbe2a898_98);
not \U$22452 ( \22698 , \22697 );
not \U$22453 ( \22699 , \7513 );
or \U$22454 ( \22700 , \22698 , \22699 );
xor \U$22455 ( \22701 , RIbe29c68_72, RIbe2aa00_101);
nand \U$22456 ( \22702 , \4580 , \22701 );
nand \U$22457 ( \22703 , \22700 , \22702 );
xnor \U$22458 ( \22704 , \22696 , \22703 );
not \U$22459 ( \22705 , \22704 );
not \U$22460 ( \22706 , \22705 );
and \U$22461 ( \22707 , \1263 , RIbe2ae38_110);
xor \U$22462 ( \22708 , RIbe29d58_74, RIbe2a2f8_86);
not \U$22463 ( \22709 , \22708 );
not \U$22464 ( \22710 , \10792 );
or \U$22465 ( \22711 , \22709 , \22710 );
xor \U$22466 ( \22712 , RIbe2a2f8_86, RIbe29ce0_73);
nand \U$22467 ( \22713 , \11094 , \22712 );
nand \U$22468 ( \22714 , \22711 , \22713 );
xor \U$22469 ( \22715 , \22707 , \22714 );
xor \U$22470 ( \22716 , RIbe28930_31, RIbe2b450_123);
not \U$22471 ( \22717 , \22716 );
or \U$22472 ( \22718 , \3949 , \22717 );
xor \U$22473 ( \22719 , RIbe28930_31, RIbe2a730_95);
not \U$22474 ( \22720 , \22719 );
or \U$22475 ( \22721 , \1200 , \22720 );
nand \U$22476 ( \22722 , \22718 , \22721 );
xor \U$22477 ( \22723 , \22715 , \22722 );
not \U$22478 ( \22724 , \22723 );
not \U$22479 ( \22725 , \22724 );
or \U$22480 ( \22726 , \22706 , \22725 );
nand \U$22481 ( \22727 , \22723 , \22704 );
nand \U$22482 ( \22728 , \22726 , \22727 );
xor \U$22483 ( \22729 , RIbe2a6b8_94, RIbe28390_19);
not \U$22484 ( \22730 , \22729 );
not \U$22485 ( \22731 , \3408 );
or \U$22486 ( \22732 , \22730 , \22731 );
xor \U$22487 ( \22733 , RIbe28390_19, RIbe2b4c8_124);
nand \U$22488 ( \22734 , \2648 , \22733 );
nand \U$22489 ( \22735 , \22732 , \22734 );
xor \U$22490 ( \22736 , RIbe285e8_24, RIbe2adc0_109);
not \U$22491 ( \22737 , \22736 );
not \U$22492 ( \22738 , \2890 );
or \U$22493 ( \22739 , \22737 , \22738 );
xor \U$22494 ( \22740 , RIbe285e8_24, RIbe2a460_89);
nand \U$22495 ( \22741 , \8270 , \22740 );
nand \U$22496 ( \22742 , \22739 , \22741 );
xor \U$22497 ( \22743 , \22735 , \22742 );
xor \U$22498 ( \22744 , RIbe2b540_125, RIbe28480_21);
not \U$22499 ( \22745 , \22744 );
not \U$22500 ( \22746 , \2519 );
or \U$22501 ( \22747 , \22745 , \22746 );
xor \U$22502 ( \22748 , RIbe2ad48_108, RIbe28480_21);
nand \U$22503 ( \22749 , \11263 , \22748 );
nand \U$22504 ( \22750 , \22747 , \22749 );
not \U$22505 ( \22751 , \22750 );
and \U$22506 ( \22752 , \22743 , \22751 );
not \U$22507 ( \22753 , \22743 );
and \U$22508 ( \22754 , \22753 , \22750 );
nor \U$22509 ( \22755 , \22752 , \22754 );
and \U$22510 ( \22756 , \22728 , \22755 );
not \U$22511 ( \22757 , \22728 );
not \U$22512 ( \22758 , \22755 );
and \U$22513 ( \22759 , \22757 , \22758 );
nor \U$22514 ( \22760 , \22756 , \22759 );
xor \U$22515 ( \22761 , RIbe297b8_62, RIbe2b018_114);
not \U$22516 ( \22762 , \22761 );
buf \U$22517 ( \22763 , \17570 );
not \U$22518 ( \22764 , \22763 );
or \U$22519 ( \22765 , \22762 , \22764 );
xnor \U$22520 ( \22766 , RIbe28138_14, RIbe2b018_114);
not \U$22521 ( \22767 , \22766 );
nand \U$22522 ( \22768 , \22767 , \19371 );
nand \U$22523 ( \22769 , \22765 , \22768 );
not \U$22524 ( \22770 , \22769 );
xor \U$22525 ( \22771 , RIbe29128_48, RIbe2b180_117);
not \U$22526 ( \22772 , \22771 );
not \U$22527 ( \22773 , \15353 );
or \U$22528 ( \22774 , \22772 , \22773 );
xor \U$22529 ( \22775 , RIbe2b180_117, RIbe291a0_49);
nand \U$22530 ( \22776 , \21759 , \22775 );
nand \U$22531 ( \22777 , \22774 , \22776 );
not \U$22532 ( \22778 , \22777 );
or \U$22533 ( \22779 , \22770 , \22778 );
not \U$22534 ( \22780 , \22769 );
not \U$22535 ( \22781 , \22780 );
not \U$22536 ( \22782 , \22777 );
not \U$22537 ( \22783 , \22782 );
or \U$22538 ( \22784 , \22781 , \22783 );
or \U$22539 ( \22785 , RIbe28930_31, RIbe29560_57);
nand \U$22540 ( \22786 , \22785 , RIbe2ae38_110);
nand \U$22541 ( \22787 , RIbe28930_31, RIbe29560_57);
and \U$22542 ( \22788 , \22786 , \22787 , RIbe28228_16);
xor \U$22543 ( \22789 , RIbe28930_31, RIbe2b3d8_122);
not \U$22544 ( \22790 , \22789 );
not \U$22545 ( \22791 , \965 );
or \U$22546 ( \22792 , \22790 , \22791 );
nand \U$22547 ( \22793 , \1199 , \22716 );
nand \U$22548 ( \22794 , \22792 , \22793 );
xor \U$22549 ( \22795 , \22788 , \22794 );
nand \U$22550 ( \22796 , \22784 , \22795 );
nand \U$22551 ( \22797 , \22779 , \22796 );
not \U$22552 ( \22798 , \22797 );
not \U$22553 ( \22799 , RIbe28a20_33);
not \U$22554 ( \22800 , RIbe2a7a8_96);
and \U$22555 ( \22801 , \22799 , \22800 );
and \U$22556 ( \22802 , RIbe28a20_33, RIbe2a7a8_96);
nor \U$22557 ( \22803 , \22801 , \22802 );
and \U$22558 ( \22804 , \1780 , \22803 );
xor \U$22559 ( \22805 , RIbe28a20_33, RIbe2abe0_105);
and \U$22560 ( \22806 , \1768 , \22805 );
nor \U$22561 ( \22807 , \22804 , \22806 );
xor \U$22562 ( \22808 , RIbe29740_61, RIbe2af28_112);
not \U$22563 ( \22809 , \22808 );
not \U$22564 ( \22810 , \16913 );
or \U$22565 ( \22811 , \22809 , \22810 );
not \U$22566 ( \22812 , RIbe297b8_62);
not \U$22567 ( \22813 , RIbe2af28_112);
and \U$22568 ( \22814 , \22812 , \22813 );
and \U$22569 ( \22815 , RIbe297b8_62, RIbe2af28_112);
nor \U$22570 ( \22816 , \22814 , \22815 );
nand \U$22571 ( \22817 , \17810 , \22816 );
nand \U$22572 ( \22818 , \22811 , \22817 );
not \U$22573 ( \22819 , \22818 );
xor \U$22574 ( \22820 , \22807 , \22819 );
xor \U$22575 ( \22821 , RIbe28f48_44, RIbe2a820_97);
and \U$22576 ( \22822 , \3249 , \22821 );
xor \U$22577 ( \22823 , RIbe28f48_44, RIbe2a118_82);
not \U$22578 ( \22824 , \22823 );
nor \U$22579 ( \22825 , \22824 , \13594 );
nor \U$22580 ( \22826 , \22822 , \22825 );
xor \U$22581 ( \22827 , \22820 , \22826 );
not \U$22582 ( \22828 , \22827 );
or \U$22583 ( \22829 , \22798 , \22828 );
or \U$22584 ( \22830 , \22827 , \22797 );
nand \U$22585 ( \22831 , \22829 , \22830 );
xor \U$22586 ( \22832 , RIbe27e68_8, RIbe2a4d8_90);
not \U$22587 ( \22833 , \22832 );
not \U$22588 ( \22834 , \2458 );
or \U$22589 ( \22835 , \22833 , \22834 );
xor \U$22590 ( \22836 , RIbe2b2e8_120, RIbe27e68_8);
nand \U$22591 ( \22837 , \13306 , \22836 );
nand \U$22592 ( \22838 , \22835 , \22837 );
xor \U$22593 ( \22839 , RIbe29b78_70, RIbe2a3e8_88);
not \U$22594 ( \22840 , \22839 );
not \U$22595 ( \22841 , \9262 );
or \U$22596 ( \22842 , \22840 , \22841 );
xor \U$22597 ( \22843 , RIbe27b20_1, RIbe2a3e8_88);
nand \U$22598 ( \22844 , \10476 , \22843 );
nand \U$22599 ( \22845 , \22842 , \22844 );
xor \U$22600 ( \22846 , \22838 , \22845 );
xor \U$22601 ( \22847 , RIbe29f38_78, RIbe2a028_80);
not \U$22602 ( \22848 , \22847 );
buf \U$22603 ( \22849 , \8168 );
not \U$22604 ( \22850 , \22849 );
or \U$22605 ( \22851 , \22848 , \22850 );
xor \U$22606 ( \22852 , RIbe29ec0_77, RIbe2a028_80);
nand \U$22607 ( \22853 , \9065 , \22852 );
nand \U$22608 ( \22854 , \22851 , \22853 );
xor \U$22609 ( \22855 , \22846 , \22854 );
not \U$22610 ( \22856 , \22855 );
and \U$22611 ( \22857 , \22831 , \22856 );
not \U$22612 ( \22858 , \22831 );
and \U$22613 ( \22859 , \22858 , \22855 );
nor \U$22614 ( \22860 , \22857 , \22859 );
or \U$22615 ( \22861 , \22760 , \22860 );
nand \U$22616 ( \22862 , \22760 , \22860 );
nand \U$22617 ( \22863 , \22861 , \22862 );
not \U$22618 ( \22864 , \22795 );
not \U$22619 ( \22865 , \22864 );
not \U$22620 ( \22866 , \22777 );
not \U$22621 ( \22867 , \22780 );
or \U$22622 ( \22868 , \22866 , \22867 );
or \U$22623 ( \22869 , \22777 , \22780 );
nand \U$22624 ( \22870 , \22868 , \22869 );
not \U$22625 ( \22871 , \22870 );
or \U$22626 ( \22872 , \22865 , \22871 );
or \U$22627 ( \22873 , \22870 , \22864 );
nand \U$22628 ( \22874 , \22872 , \22873 );
not \U$22629 ( \22875 , \22874 );
or \U$22630 ( \22876 , RIbe289a8_32, RIbe28a20_33);
nand \U$22631 ( \22877 , \22876 , RIbe2ae38_110);
nand \U$22632 ( \22878 , RIbe289a8_32, RIbe28a20_33);
and \U$22633 ( \22879 , \22877 , \22878 , RIbe28930_31);
xor \U$22634 ( \22880 , RIbe28a20_33, RIbe2b3d8_122);
not \U$22635 ( \22881 , \22880 );
not \U$22636 ( \22882 , \1780 );
or \U$22637 ( \22883 , \22881 , \22882 );
xor \U$22638 ( \22884 , RIbe28a20_33, RIbe2b450_123);
nand \U$22639 ( \22885 , \5055 , \22884 );
nand \U$22640 ( \22886 , \22883 , \22885 );
and \U$22641 ( \22887 , \22879 , \22886 );
xor \U$22642 ( \22888 , RIbe2a2f8_86, RIbe2b6a8_128);
not \U$22643 ( \22889 , \22888 );
not \U$22644 ( \22890 , \14827 );
or \U$22645 ( \22891 , \22889 , \22890 );
xor \U$22646 ( \22892 , RIbe29f38_78, RIbe2a2f8_86);
nand \U$22647 ( \22893 , \11094 , \22892 );
nand \U$22648 ( \22894 , \22891 , \22893 );
xor \U$22649 ( \22895 , RIbe27fd0_11, RIbe2a460_89);
not \U$22650 ( \22896 , \22895 );
not \U$22651 ( \22897 , \10466 );
or \U$22652 ( \22898 , \22896 , \22897 );
xor \U$22653 ( \22899 , RIbe27fd0_11, RIbe2a4d8_90);
nand \U$22654 ( \22900 , \2707 , \22899 );
nand \U$22655 ( \22901 , \22898 , \22900 );
or \U$22656 ( \22902 , \22894 , \22901 );
xor \U$22657 ( \22903 , RIbe2a910_99, RIbe29ce0_73);
not \U$22658 ( \22904 , \22903 );
not \U$22659 ( \22905 , \10987 );
or \U$22660 ( \22906 , \22904 , \22905 );
not \U$22661 ( \22907 , RIbe29b78_70);
not \U$22662 ( \22908 , RIbe2a910_99);
and \U$22663 ( \22909 , \22907 , \22908 );
and \U$22664 ( \22910 , RIbe29b78_70, RIbe2a910_99);
nor \U$22665 ( \22911 , \22909 , \22910 );
nand \U$22666 ( \22912 , \11456 , \22911 );
nand \U$22667 ( \22913 , \22906 , \22912 );
nand \U$22668 ( \22914 , \22902 , \22913 );
nand \U$22669 ( \22915 , \22894 , \22901 );
nand \U$22670 ( \22916 , \22914 , \22915 );
xor \U$22671 ( \22917 , \22887 , \22916 );
buf \U$22672 ( \22918 , \11399 );
not \U$22673 ( \22919 , \22918 );
xor \U$22674 ( \22920 , RIbe29998_66, RIbe2a190_83);
not \U$22675 ( \22921 , \22920 );
or \U$22676 ( \22922 , \22919 , \22921 );
xor \U$22677 ( \22923 , RIbe298a8_64, RIbe2a190_83);
not \U$22678 ( \22924 , \22923 );
or \U$22679 ( \22925 , \22924 , \10689 );
nand \U$22680 ( \22926 , \22922 , \22925 );
xor \U$22681 ( \22927 , RIbe29ec0_77, RIbe2a3e8_88);
not \U$22682 ( \22928 , \22927 );
not \U$22683 ( \22929 , \9263 );
or \U$22684 ( \22930 , \22928 , \22929 );
xor \U$22685 ( \22931 , RIbe2a3e8_88, RIbe29d58_74);
nand \U$22686 ( \22932 , \10476 , \22931 );
nand \U$22687 ( \22933 , \22930 , \22932 );
xor \U$22688 ( \22934 , \22926 , \22933 );
xor \U$22689 ( \22935 , RIbe28930_31, RIbe2ae38_110);
not \U$22690 ( \22936 , \22935 );
not \U$22691 ( \22937 , \1793 );
or \U$22692 ( \22938 , \22936 , \22937 );
xor \U$22693 ( \22939 , RIbe2aeb0_111, RIbe28930_31);
nand \U$22694 ( \22940 , \1797 , \22939 );
nand \U$22695 ( \22941 , \22938 , \22940 );
and \U$22696 ( \22942 , \22934 , \22941 );
and \U$22697 ( \22943 , \22926 , \22933 );
or \U$22698 ( \22944 , \22942 , \22943 );
and \U$22699 ( \22945 , \22917 , \22944 );
and \U$22700 ( \22946 , \22887 , \22916 );
or \U$22701 ( \22947 , \22945 , \22946 );
not \U$22702 ( \22948 , \22947 );
not \U$22703 ( \22949 , \22948 );
or \U$22704 ( \22950 , \22875 , \22949 );
or \U$22705 ( \22951 , \22948 , \22874 );
nand \U$22706 ( \22952 , \22950 , \22951 );
not \U$22707 ( \22953 , \22952 );
xor \U$22708 ( \22954 , RIbe2b360_121, RIbe28f48_44);
and \U$22709 ( \22955 , \3249 , \22954 );
xor \U$22710 ( \22956 , RIbe28f48_44, RIbe2b2e8_120);
not \U$22711 ( \22957 , \22956 );
nor \U$22712 ( \22958 , \22957 , \3257 );
nor \U$22713 ( \22959 , \22955 , \22958 );
not \U$22714 ( \22960 , \22959 );
not \U$22715 ( \22961 , \22960 );
xor \U$22716 ( \22962 , RIbe29a10_67, RIbe2b180_117);
not \U$22717 ( \22963 , \22962 );
not \U$22718 ( \22964 , \15353 );
or \U$22719 ( \22965 , \22963 , \22964 );
xor \U$22720 ( \22966 , RIbe29b00_69, RIbe2b180_117);
nand \U$22721 ( \22967 , \21759 , \22966 );
nand \U$22722 ( \22968 , \22965 , \22967 );
not \U$22723 ( \22969 , \22968 );
not \U$22724 ( \22970 , \12003 );
xor \U$22725 ( \22971 , RIbe2a550_91, RIbe28cf0_39);
not \U$22726 ( \22972 , \22971 );
not \U$22727 ( \22973 , \22972 );
and \U$22728 ( \22974 , \22970 , \22973 );
not \U$22729 ( \22975 , \15991 );
xor \U$22730 ( \22976 , RIbe2a550_91, RIbe27b20_1);
and \U$22731 ( \22977 , \22975 , \22976 );
nor \U$22732 ( \22978 , \22974 , \22977 );
not \U$22733 ( \22979 , \22978 );
or \U$22734 ( \22980 , \22969 , \22979 );
or \U$22735 ( \22981 , \22978 , \22968 );
nand \U$22736 ( \22982 , \22980 , \22981 );
not \U$22737 ( \22983 , \22982 );
or \U$22738 ( \22984 , \22961 , \22983 );
not \U$22739 ( \22985 , \22978 );
nand \U$22740 ( \22986 , \22985 , \22968 );
nand \U$22741 ( \22987 , \22984 , \22986 );
not \U$22742 ( \22988 , \22987 );
xor \U$22743 ( \22989 , RIbe295d8_58, RIbe2b018_114);
not \U$22744 ( \22990 , \22989 );
not \U$22745 ( \22991 , \15967 );
or \U$22746 ( \22992 , \22990 , \22991 );
not \U$22747 ( \22993 , RIbe29740_61);
not \U$22748 ( \22994 , RIbe2b018_114);
and \U$22749 ( \22995 , \22993 , \22994 );
and \U$22750 ( \22996 , RIbe29740_61, RIbe2b018_114);
nor \U$22751 ( \22997 , \22995 , \22996 );
nand \U$22752 ( \22998 , \15953 , \22997 );
nand \U$22753 ( \22999 , \22992 , \22998 );
not \U$22754 ( \23000 , \22999 );
xor \U$22755 ( \23001 , RIbe2ad48_108, RIbe27e68_8);
not \U$22756 ( \23002 , \23001 );
not \U$22757 ( \23003 , \2459 );
or \U$22758 ( \23004 , \23002 , \23003 );
xor \U$22759 ( \23005 , RIbe27e68_8, RIbe2adc0_109);
nand \U$22760 ( \23006 , \2603 , \23005 );
nand \U$22761 ( \23007 , \23004 , \23006 );
not \U$22762 ( \23008 , \23007 );
or \U$22763 ( \23009 , \23000 , \23008 );
or \U$22764 ( \23010 , \23007 , \22999 );
xor \U$22765 ( \23011 , RIbe27df0_7, RIbe2b108_116);
not \U$22766 ( \23012 , \23011 );
not \U$22767 ( \23013 , \13542 );
or \U$22768 ( \23014 , \23012 , \23013 );
buf \U$22769 ( \23015 , \16875 );
xor \U$22770 ( \23016 , RIbe29218_50, RIbe2b108_116);
nand \U$22771 ( \23017 , \23015 , \23016 );
nand \U$22772 ( \23018 , \23014 , \23017 );
nand \U$22773 ( \23019 , \23010 , \23018 );
nand \U$22774 ( \23020 , \23009 , \23019 );
not \U$22775 ( \23021 , \23020 );
xor \U$22776 ( \23022 , RIbe2a820_97, RIbe29e48_76);
not \U$22777 ( \23023 , \23022 );
not \U$22778 ( \23024 , \11039 );
or \U$22779 ( \23025 , \23023 , \23024 );
xor \U$22780 ( \23026 , RIbe29e48_76, RIbe2a898_98);
nand \U$22781 ( \23027 , \4850 , \23026 );
nand \U$22782 ( \23028 , \23025 , \23027 );
not \U$22783 ( \23029 , \23028 );
not \U$22784 ( \23030 , \19580 );
not \U$22785 ( \23031 , RIbe2aaf0_103);
not \U$22786 ( \23032 , RIbe297b8_62);
or \U$22787 ( \23033 , \23031 , \23032 );
or \U$22788 ( \23034 , RIbe297b8_62, RIbe2aaf0_103);
nand \U$22789 ( \23035 , \23033 , \23034 );
not \U$22790 ( \23036 , \23035 );
and \U$22791 ( \23037 , \23030 , \23036 );
xor \U$22792 ( \23038 , RIbe28138_14, RIbe2aaf0_103);
and \U$22793 ( \23039 , RIbe2ab68_104, \23038 );
nor \U$22794 ( \23040 , \23037 , \23039 );
not \U$22795 ( \23041 , \23040 );
and \U$22796 ( \23042 , \23029 , \23041 );
and \U$22797 ( \23043 , \23028 , \23040 );
nor \U$22798 ( \23044 , \23042 , \23043 );
xor \U$22799 ( \23045 , RIbe27c88_4, RIbe2a280_85);
and \U$22800 ( \23046 , \11348 , \23045 );
buf \U$22801 ( \23047 , \14942 );
not \U$22802 ( \23048 , RIbe28d68_40);
not \U$22803 ( \23049 , RIbe2a280_85);
and \U$22804 ( \23050 , \23048 , \23049 );
and \U$22805 ( \23051 , RIbe28d68_40, RIbe2a280_85);
nor \U$22806 ( \23052 , \23050 , \23051 );
and \U$22807 ( \23053 , \23047 , \23052 );
nor \U$22808 ( \23054 , \23046 , \23053 );
or \U$22809 ( \23055 , \23044 , \23054 );
not \U$22810 ( \23056 , \23028 );
or \U$22811 ( \23057 , \23056 , \23040 );
nand \U$22812 ( \23058 , \23055 , \23057 );
not \U$22813 ( \23059 , \23058 );
not \U$22814 ( \23060 , \23059 );
or \U$22815 ( \23061 , \23021 , \23060 );
or \U$22816 ( \23062 , \23059 , \23020 );
nand \U$22817 ( \23063 , \23061 , \23062 );
not \U$22818 ( \23064 , \23063 );
or \U$22819 ( \23065 , \22988 , \23064 );
nand \U$22820 ( \23066 , \23058 , \23020 );
nand \U$22821 ( \23067 , \23065 , \23066 );
not \U$22822 ( \23068 , \23067 );
or \U$22823 ( \23069 , \22953 , \23068 );
not \U$22824 ( \23070 , \22948 );
nand \U$22825 ( \23071 , \23070 , \22874 );
nand \U$22826 ( \23072 , \23069 , \23071 );
not \U$22827 ( \23073 , \23072 );
and \U$22828 ( \23074 , \22863 , \23073 );
not \U$22829 ( \23075 , \22863 );
and \U$22830 ( \23076 , \23075 , \23072 );
nor \U$22831 ( \23077 , \23074 , \23076 );
xor \U$22832 ( \23078 , RIbe28a20_33, RIbe2a730_95);
not \U$22833 ( \23079 , \23078 );
not \U$22834 ( \23080 , \1779 );
or \U$22835 ( \23081 , \23079 , \23080 );
nand \U$22836 ( \23082 , \5055 , \22803 );
nand \U$22837 ( \23083 , \23081 , \23082 );
not \U$22838 ( \23084 , \23083 );
xor \U$22839 ( \23085 , RIbe28b88_36, RIbe2abe0_105);
not \U$22840 ( \23086 , \23085 );
not \U$22841 ( \23087 , \2552 );
or \U$22842 ( \23088 , \23086 , \23087 );
xor \U$22843 ( \23089 , RIbe28b88_36, RIbe2ac58_106);
nand \U$22844 ( \23090 , \7549 , \23089 );
nand \U$22845 ( \23091 , \23088 , \23090 );
not \U$22846 ( \23092 , \23091 );
or \U$22847 ( \23093 , \23084 , \23092 );
or \U$22848 ( \23094 , \23091 , \23083 );
xor \U$22849 ( \23095 , RIbe2a0a0_81, RIbe28f48_44);
not \U$22850 ( \23096 , \23095 );
and \U$22851 ( \23097 , \3252 , \3253 );
not \U$22852 ( \23098 , \23097 );
or \U$22853 ( \23099 , \23096 , \23098 );
nand \U$22854 ( \23100 , \11201 , \22823 );
nand \U$22855 ( \23101 , \23099 , \23100 );
nand \U$22856 ( \23102 , \23094 , \23101 );
nand \U$22857 ( \23103 , \23093 , \23102 );
not \U$22858 ( \23104 , \23103 );
not \U$22859 ( \23105 , \23104 );
xor \U$22860 ( \23106 , RIbe27fd0_11, RIbe2b2e8_120);
not \U$22861 ( \23107 , \23106 );
not \U$22862 ( \23108 , \11366 );
or \U$22863 ( \23109 , \23107 , \23108 );
xor \U$22864 ( \23110 , RIbe27fd0_11, RIbe2b360_121);
nand \U$22865 ( \23111 , \2707 , \23110 );
nand \U$22866 ( \23112 , \23109 , \23111 );
not \U$22867 ( \23113 , \23112 );
xor \U$22868 ( \23114 , RIbe2b108_116, RIbe29a10_67);
not \U$22869 ( \23115 , \23114 );
not \U$22870 ( \23116 , \13527 );
or \U$22871 ( \23117 , \23115 , \23116 );
xor \U$22872 ( \23118 , RIbe2b108_116, RIbe29b00_69);
nand \U$22873 ( \23119 , \13533 , \23118 );
nand \U$22874 ( \23120 , \23117 , \23119 );
xor \U$22875 ( \23121 , RIbe27b20_1, RIbe2a910_99);
not \U$22876 ( \23122 , \23121 );
not \U$22877 ( \23123 , \9736 );
or \U$22878 ( \23124 , \23122 , \23123 );
xor \U$22879 ( \23125 , RIbe28cf0_39, RIbe2a910_99);
nand \U$22880 ( \23126 , \9725 , \23125 );
nand \U$22881 ( \23127 , \23124 , \23126 );
xor \U$22882 ( \23128 , \23120 , \23127 );
not \U$22883 ( \23129 , \23128 );
or \U$22884 ( \23130 , \23113 , \23129 );
nand \U$22885 ( \23131 , \23127 , \23120 );
nand \U$22886 ( \23132 , \23130 , \23131 );
not \U$22887 ( \23133 , \23132 );
or \U$22888 ( \23134 , \23105 , \23133 );
or \U$22889 ( \23135 , \23132 , \23104 );
nand \U$22890 ( \23136 , \23134 , \23135 );
xor \U$22891 ( \23137 , RIbe285e8_24, RIbe2ad48_108);
not \U$22892 ( \23138 , \23137 );
not \U$22893 ( \23139 , \2761 );
or \U$22894 ( \23140 , \23138 , \23139 );
nand \U$22895 ( \23141 , \2625 , \22736 );
nand \U$22896 ( \23142 , \23140 , \23141 );
xor \U$22897 ( \23143 , RIbe27df0_7, RIbe2a280_85);
not \U$22898 ( \23144 , \23143 );
not \U$22899 ( \23145 , \11345 );
or \U$22900 ( \23146 , \23144 , \23145 );
xor \U$22901 ( \23147 , RIbe29218_50, RIbe2a280_85);
nand \U$22902 ( \23148 , \14649 , \23147 );
nand \U$22903 ( \23149 , \23146 , \23148 );
xor \U$22904 ( \23150 , \23142 , \23149 );
xor \U$22905 ( \23151 , RIbe29e48_76, RIbe2aa00_101);
not \U$22906 ( \23152 , \23151 );
not \U$22907 ( \23153 , \7716 );
or \U$22908 ( \23154 , \23152 , \23153 );
xor \U$22909 ( \23155 , RIbe2aa78_102, RIbe29e48_76);
nand \U$22910 ( \23156 , \4851 , \23155 );
nand \U$22911 ( \23157 , \23154 , \23156 );
and \U$22912 ( \23158 , \23150 , \23157 );
and \U$22913 ( \23159 , \23142 , \23149 );
or \U$22914 ( \23160 , \23158 , \23159 );
not \U$22915 ( \23161 , \23160 );
and \U$22916 ( \23162 , \23136 , \23161 );
not \U$22917 ( \23163 , \23136 );
and \U$22918 ( \23164 , \23163 , \23160 );
nor \U$22919 ( \23165 , \23162 , \23164 );
not \U$22920 ( \23166 , \23165 );
xor \U$22921 ( \23167 , RIbe2aaf0_103, RIbe282a0_17);
not \U$22922 ( \23168 , \23167 );
not \U$22923 ( \23169 , \19580 );
not \U$22924 ( \23170 , \23169 );
or \U$22925 ( \23171 , \23168 , \23170 );
nand \U$22926 ( \23172 , \22681 , RIbe2ab68_104);
nand \U$22927 ( \23173 , \23171 , \23172 );
not \U$22928 ( \23174 , \23173 );
xor \U$22929 ( \23175 , RIbe28480_21, RIbe2b4c8_124);
not \U$22930 ( \23176 , \23175 );
not \U$22931 ( \23177 , \2518 );
or \U$22932 ( \23178 , \23176 , \23177 );
nand \U$22933 ( \23179 , \7483 , \22744 );
nand \U$22934 ( \23180 , \23178 , \23179 );
not \U$22935 ( \23181 , \23180 );
or \U$22936 ( \23182 , \23174 , \23181 );
or \U$22937 ( \23183 , \23180 , \23173 );
xor \U$22938 ( \23184 , RIbe28390_19, RIbe2a640_93);
not \U$22939 ( \23185 , \23184 );
not \U$22940 ( \23186 , \8651 );
or \U$22941 ( \23187 , \23185 , \23186 );
nand \U$22942 ( \23188 , \8654 , \22729 );
nand \U$22943 ( \23189 , \23187 , \23188 );
nand \U$22944 ( \23190 , \23183 , \23189 );
nand \U$22945 ( \23191 , \23182 , \23190 );
xor \U$22946 ( \23192 , RIbe27e68_8, RIbe2a460_89);
not \U$22947 ( \23193 , \23192 );
not \U$22948 ( \23194 , \4443 );
or \U$22949 ( \23195 , \23193 , \23194 );
nand \U$22950 ( \23196 , \2603 , \22832 );
nand \U$22951 ( \23197 , \23195 , \23196 );
not \U$22952 ( \23198 , \23197 );
xor \U$22953 ( \23199 , RIbe2af28_112, RIbe295d8_58);
not \U$22954 ( \23200 , \23199 );
not \U$22955 ( \23201 , \14423 );
or \U$22956 ( \23202 , \23200 , \23201 );
nand \U$22957 ( \23203 , \17809 , \22808 );
nand \U$22958 ( \23204 , \23202 , \23203 );
xor \U$22959 ( \23205 , RIbe29ce0_73, RIbe2a3e8_88);
not \U$22960 ( \23206 , \23205 );
not \U$22961 ( \23207 , \9262 );
or \U$22962 ( \23208 , \23206 , \23207 );
nand \U$22963 ( \23209 , \9089 , \22839 );
nand \U$22964 ( \23210 , \23208 , \23209 );
xor \U$22965 ( \23211 , \23204 , \23210 );
not \U$22966 ( \23212 , \23211 );
or \U$22967 ( \23213 , \23198 , \23212 );
nand \U$22968 ( \23214 , \23204 , \23210 );
nand \U$22969 ( \23215 , \23213 , \23214 );
xor \U$22970 ( \23216 , \23191 , \23215 );
xor \U$22971 ( \23217 , RIbe29ec0_77, RIbe2a2f8_86);
and \U$22972 ( \23218 , \10792 , \23217 );
and \U$22973 ( \23219 , \9379 , \22708 );
nor \U$22974 ( \23220 , \23218 , \23219 );
not \U$22975 ( \23221 , \23220 );
not \U$22976 ( \23222 , \23221 );
xor \U$22977 ( \23223 , RIbe2a550_91, RIbe298a8_64);
not \U$22978 ( \23224 , \23223 );
not \U$22979 ( \23225 , \11999 );
or \U$22980 ( \23226 , \23224 , \23225 );
xor \U$22981 ( \23227 , RIbe29998_66, RIbe2a550_91);
not \U$22982 ( \23228 , \23227 );
not \U$22983 ( \23229 , \23228 );
nand \U$22984 ( \23230 , \23229 , \11485 );
nand \U$22985 ( \23231 , \23226 , \23230 );
xor \U$22986 ( \23232 , RIbe28228_16, RIbe2ae38_110);
not \U$22987 ( \23233 , \23232 );
not \U$22988 ( \23234 , \15059 );
or \U$22989 ( \23235 , \23233 , \23234 );
xor \U$22990 ( \23236 , RIbe28228_16, RIbe2aeb0_111);
nand \U$22991 ( \23237 , \885 , \23236 );
nand \U$22992 ( \23238 , \23235 , \23237 );
and \U$22993 ( \23239 , \23231 , \23238 );
not \U$22994 ( \23240 , \23231 );
not \U$22995 ( \23241 , \23238 );
and \U$22996 ( \23242 , \23240 , \23241 );
nor \U$22997 ( \23243 , \23239 , \23242 );
not \U$22998 ( \23244 , \23243 );
or \U$22999 ( \23245 , \23222 , \23244 );
nand \U$23000 ( \23246 , \23231 , \23238 );
nand \U$23001 ( \23247 , \23245 , \23246 );
xor \U$23002 ( \23248 , \23216 , \23247 );
not \U$23003 ( \23249 , \23248 );
or \U$23004 ( \23250 , \23166 , \23249 );
or \U$23005 ( \23251 , \23248 , \23165 );
nand \U$23006 ( \23252 , \23250 , \23251 );
not \U$23007 ( \23253 , \23125 );
not \U$23008 ( \23254 , \9737 );
or \U$23009 ( \23255 , \23253 , \23254 );
xor \U$23010 ( \23256 , RIbe2a910_99, RIbe298a8_64);
nand \U$23011 ( \23257 , \9726 , \23256 );
nand \U$23012 ( \23258 , \23255 , \23257 );
not \U$23013 ( \23259 , \3377 );
not \U$23014 ( \23260 , \23110 );
or \U$23015 ( \23261 , \23259 , \23260 );
xor \U$23016 ( \23262 , RIbe2a0a0_81, RIbe27fd0_11);
nand \U$23017 ( \23263 , \2707 , \23262 );
nand \U$23018 ( \23264 , \23261 , \23263 );
nor \U$23019 ( \23265 , \23258 , \23264 );
not \U$23020 ( \23266 , \23265 );
nand \U$23021 ( \23267 , \23258 , \23264 );
nand \U$23022 ( \23268 , \23266 , \23267 );
not \U$23023 ( \23269 , \15968 );
not \U$23024 ( \23270 , \22766 );
and \U$23025 ( \23271 , \23269 , \23270 );
xor \U$23026 ( \23272 , RIbe282a0_17, RIbe2b018_114);
and \U$23027 ( \23273 , \15953 , \23272 );
nor \U$23028 ( \23274 , \23271 , \23273 );
not \U$23029 ( \23275 , \23274 );
and \U$23030 ( \23276 , \23268 , \23275 );
not \U$23031 ( \23277 , \23268 );
and \U$23032 ( \23278 , \23277 , \23274 );
nor \U$23033 ( \23279 , \23276 , \23278 );
not \U$23034 ( \23280 , \23279 );
not \U$23035 ( \23281 , \23118 );
not \U$23036 ( \23282 , \14297 );
or \U$23037 ( \23283 , \23281 , \23282 );
xor \U$23038 ( \23284 , RIbe2b108_116, RIbe29128_48);
nand \U$23039 ( \23285 , \13534 , \23284 );
nand \U$23040 ( \23286 , \23283 , \23285 );
not \U$23041 ( \23287 , \23147 );
not \U$23042 ( \23288 , \11345 );
or \U$23043 ( \23289 , \23287 , \23288 );
xor \U$23044 ( \23290 , RIbe2a280_85, RIbe29a10_67);
nand \U$23045 ( \23291 , \11348 , \23290 );
nand \U$23046 ( \23292 , \23289 , \23291 );
xor \U$23047 ( \23293 , \23286 , \23292 );
not \U$23048 ( \23294 , \23155 );
not \U$23049 ( \23295 , \4843 );
or \U$23050 ( \23296 , \23294 , \23295 );
xor \U$23051 ( \23297 , RIbe29e48_76, RIbe2b6a8_128);
nand \U$23052 ( \23298 , \7368 , \23297 );
nand \U$23053 ( \23299 , \23296 , \23298 );
xor \U$23054 ( \23300 , \23293 , \23299 );
not \U$23055 ( \23301 , \23300 );
or \U$23056 ( \23302 , \23280 , \23301 );
or \U$23057 ( \23303 , \23279 , \23300 );
nand \U$23058 ( \23304 , \23302 , \23303 );
or \U$23059 ( \23305 , \15991 , \23228 );
not \U$23060 ( \23306 , \10439 );
not \U$23061 ( \23307 , \23306 );
xor \U$23062 ( \23308 , RIbe28d68_40, RIbe2a550_91);
not \U$23063 ( \23309 , \23308 );
or \U$23064 ( \23310 , \23307 , \23309 );
nand \U$23065 ( \23311 , \23305 , \23310 );
not \U$23066 ( \23312 , \23311 );
not \U$23067 ( \23313 , \23089 );
not \U$23068 ( \23314 , \9052 );
or \U$23069 ( \23315 , \23313 , \23314 );
xor \U$23070 ( \23316 , RIbe2a640_93, RIbe28b88_36);
nand \U$23071 ( \23317 , \13250 , \23316 );
nand \U$23072 ( \23318 , \23315 , \23317 );
not \U$23073 ( \23319 , \23318 );
not \U$23074 ( \23320 , \23319 );
or \U$23075 ( \23321 , \23312 , \23320 );
not \U$23076 ( \23322 , \23311 );
nand \U$23077 ( \23323 , \23322 , \23318 );
nand \U$23078 ( \23324 , \23321 , \23323 );
not \U$23079 ( \23325 , \23236 );
not \U$23080 ( \23326 , \879 );
or \U$23081 ( \23327 , \23325 , \23326 );
xor \U$23082 ( \23328 , RIbe2b3d8_122, RIbe28228_16);
nand \U$23083 ( \23329 , \8680 , \23328 );
nand \U$23084 ( \23330 , \23327 , \23329 );
xnor \U$23085 ( \23331 , \23324 , \23330 );
not \U$23086 ( \23332 , \23331 );
and \U$23087 ( \23333 , \23304 , \23332 );
not \U$23088 ( \23334 , \23304 );
and \U$23089 ( \23335 , \23334 , \23331 );
nor \U$23090 ( \23336 , \23333 , \23335 );
xnor \U$23091 ( \23337 , \23252 , \23336 );
not \U$23092 ( \23338 , \23337 );
not \U$23093 ( \23339 , \23112 );
and \U$23094 ( \23340 , \23128 , \23339 );
not \U$23095 ( \23341 , \23128 );
and \U$23096 ( \23342 , \23341 , \23112 );
nor \U$23097 ( \23343 , \23340 , \23342 );
not \U$23098 ( \23344 , \23343 );
xor \U$23099 ( \23345 , RIbe28480_21, RIbe2a6b8_94);
not \U$23100 ( \23346 , \23345 );
not \U$23101 ( \23347 , \2518 );
or \U$23102 ( \23348 , \23346 , \23347 );
nand \U$23103 ( \23349 , \3074 , \23175 );
nand \U$23104 ( \23350 , \23348 , \23349 );
not \U$23105 ( \23351 , \23350 );
not \U$23106 ( \23352 , \23045 );
not \U$23107 ( \23353 , \11344 );
not \U$23108 ( \23354 , \23353 );
or \U$23109 ( \23355 , \23352 , \23354 );
nand \U$23110 ( \23356 , \14649 , \23143 );
nand \U$23111 ( \23357 , \23355 , \23356 );
not \U$23112 ( \23358 , \23357 );
nand \U$23113 ( \23359 , \23351 , \23358 );
not \U$23114 ( \23360 , \23359 );
not \U$23115 ( \23361 , \23026 );
not \U$23116 ( \23362 , \16652 );
or \U$23117 ( \23363 , \23361 , \23362 );
nand \U$23118 ( \23364 , \16655 , \23151 );
nand \U$23119 ( \23365 , \23363 , \23364 );
not \U$23120 ( \23366 , \23365 );
or \U$23121 ( \23367 , \23360 , \23366 );
nand \U$23122 ( \23368 , \23357 , \23350 );
nand \U$23123 ( \23369 , \23367 , \23368 );
not \U$23124 ( \23370 , \23369 );
not \U$23125 ( \23371 , \23370 );
or \U$23126 ( \23372 , \23344 , \23371 );
not \U$23127 ( \23373 , \22939 );
not \U$23128 ( \23374 , \3064 );
or \U$23129 ( \23375 , \23373 , \23374 );
nand \U$23130 ( \23376 , \1797 , \22789 );
nand \U$23131 ( \23377 , \23375 , \23376 );
not \U$23132 ( \23378 , \23377 );
xor \U$23133 ( \23379 , RIbe2ac58_106, RIbe28390_19);
not \U$23134 ( \23380 , \23379 );
not \U$23135 ( \23381 , \3712 );
or \U$23136 ( \23382 , \23380 , \23381 );
nand \U$23137 ( \23383 , \3714 , \23184 );
nand \U$23138 ( \23384 , \23382 , \23383 );
not \U$23139 ( \23385 , \23384 );
not \U$23140 ( \23386 , \22920 );
not \U$23141 ( \23387 , \10689 );
not \U$23142 ( \23388 , \23387 );
or \U$23143 ( \23389 , \23386 , \23388 );
xor \U$23144 ( \23390 , RIbe28d68_40, RIbe2a190_83);
nand \U$23145 ( \23391 , \13278 , \23390 );
nand \U$23146 ( \23392 , \23389 , \23391 );
not \U$23147 ( \23393 , \23392 );
not \U$23148 ( \23394 , \23393 );
or \U$23149 ( \23395 , \23385 , \23394 );
or \U$23150 ( \23396 , \23384 , \23393 );
nand \U$23151 ( \23397 , \23395 , \23396 );
not \U$23152 ( \23398 , \23397 );
or \U$23153 ( \23399 , \23378 , \23398 );
nand \U$23154 ( \23400 , \23392 , \23384 );
nand \U$23155 ( \23401 , \23399 , \23400 );
nand \U$23156 ( \23402 , \23372 , \23401 );
not \U$23157 ( \23403 , \23343 );
nand \U$23158 ( \23404 , \23369 , \23403 );
nand \U$23159 ( \23405 , \23402 , \23404 );
not \U$23160 ( \23406 , \23197 );
and \U$23161 ( \23407 , \23211 , \23406 );
not \U$23162 ( \23408 , \23211 );
and \U$23163 ( \23409 , \23408 , \23197 );
nor \U$23164 ( \23410 , \23407 , \23409 );
not \U$23165 ( \23411 , \23410 );
not \U$23166 ( \23412 , \23390 );
not \U$23167 ( \23413 , \10690 );
or \U$23168 ( \23414 , \23412 , \23413 );
nand \U$23169 ( \23415 , \10696 , \22688 );
nand \U$23170 ( \23416 , \23414 , \23415 );
xor \U$23171 ( \23417 , RIbe2a028_80, RIbe2b6a8_128);
not \U$23172 ( \23418 , \23417 );
not \U$23173 ( \23419 , \10674 );
or \U$23174 ( \23420 , \23418 , \23419 );
nand \U$23175 ( \23421 , \9065 , \22847 );
nand \U$23176 ( \23422 , \23420 , \23421 );
xor \U$23177 ( \23423 , \23416 , \23422 );
xor \U$23178 ( \23424 , RIbe29c68_72, RIbe2a820_97);
not \U$23179 ( \23425 , \23424 );
not \U$23180 ( \23426 , \4578 );
or \U$23181 ( \23427 , \23425 , \23426 );
nand \U$23182 ( \23428 , \7642 , \22697 );
nand \U$23183 ( \23429 , \23427 , \23428 );
xnor \U$23184 ( \23430 , \23423 , \23429 );
not \U$23185 ( \23431 , \23430 );
or \U$23186 ( \23432 , \23411 , \23431 );
xor \U$23187 ( \23433 , \23083 , \23091 );
and \U$23188 ( \23434 , \23433 , \23101 );
not \U$23189 ( \23435 , \23433 );
not \U$23190 ( \23436 , \23101 );
and \U$23191 ( \23437 , \23435 , \23436 );
nor \U$23192 ( \23438 , \23434 , \23437 );
nand \U$23193 ( \23439 , \23432 , \23438 );
not \U$23194 ( \23440 , \23410 );
not \U$23195 ( \23441 , \23430 );
nand \U$23196 ( \23442 , \23440 , \23441 );
nand \U$23197 ( \23443 , \23439 , \23442 );
xor \U$23198 ( \23444 , \23405 , \23443 );
not \U$23199 ( \23445 , \23220 );
not \U$23200 ( \23446 , \23243 );
or \U$23201 ( \23447 , \23445 , \23446 );
or \U$23202 ( \23448 , \23243 , \23220 );
nand \U$23203 ( \23449 , \23447 , \23448 );
not \U$23204 ( \23450 , \23449 );
xor \U$23205 ( \23451 , \23142 , \23149 );
xor \U$23206 ( \23452 , \23451 , \23157 );
not \U$23207 ( \23453 , \23452 );
nand \U$23208 ( \23454 , \23450 , \23453 );
nand \U$23209 ( \23455 , \23449 , \23452 );
xor \U$23210 ( \23456 , \23189 , \23173 );
not \U$23211 ( \23457 , \23180 );
and \U$23212 ( \23458 , \23456 , \23457 );
not \U$23213 ( \23459 , \23456 );
and \U$23214 ( \23460 , \23459 , \23180 );
nor \U$23215 ( \23461 , \23458 , \23460 );
nand \U$23216 ( \23462 , \23455 , \23461 );
and \U$23217 ( \23463 , \23454 , \23462 );
xor \U$23218 ( \23464 , \23444 , \23463 );
not \U$23219 ( \23465 , \23464 );
or \U$23220 ( \23466 , \23338 , \23465 );
or \U$23221 ( \23467 , \23464 , \23337 );
nand \U$23222 ( \23468 , \23466 , \23467 );
xor \U$23223 ( \23469 , \23077 , \23468 );
not \U$23224 ( \23470 , \23469 );
not \U$23225 ( \23471 , \13250 );
not \U$23226 ( \23472 , \23085 );
or \U$23227 ( \23473 , \23471 , \23472 );
xnor \U$23228 ( \23474 , RIbe28b88_36, RIbe2a7a8_96);
or \U$23229 ( \23475 , \8712 , \23474 );
nand \U$23230 ( \23476 , \23473 , \23475 );
not \U$23231 ( \23477 , \9374 );
not \U$23232 ( \23478 , \22892 );
or \U$23233 ( \23479 , \23477 , \23478 );
nand \U$23234 ( \23480 , \11094 , \23217 );
nand \U$23235 ( \23481 , \23479 , \23480 );
nor \U$23236 ( \23482 , \23476 , \23481 );
xor \U$23237 ( \23483 , RIbe2a118_82, RIbe29c68_72);
not \U$23238 ( \23484 , \23483 );
not \U$23239 ( \23485 , \8259 );
or \U$23240 ( \23486 , \23484 , \23485 );
nand \U$23241 ( \23487 , \7237 , \23424 );
nand \U$23242 ( \23488 , \23486 , \23487 );
not \U$23243 ( \23489 , \23488 );
or \U$23244 ( \23490 , \23482 , \23489 );
nand \U$23245 ( \23491 , \23476 , \23481 );
nand \U$23246 ( \23492 , \23490 , \23491 );
not \U$23247 ( \23493 , \22911 );
not \U$23248 ( \23494 , \15395 );
or \U$23249 ( \23495 , \23493 , \23494 );
nand \U$23250 ( \23496 , \9726 , \23121 );
nand \U$23251 ( \23497 , \23495 , \23496 );
not \U$23252 ( \23498 , \23497 );
not \U$23253 ( \23499 , \23038 );
not \U$23254 ( \23500 , \19581 );
or \U$23255 ( \23501 , \23499 , \23500 );
nand \U$23256 ( \23502 , \23167 , RIbe2ab68_104);
nand \U$23257 ( \23503 , \23501 , \23502 );
not \U$23258 ( \23504 , \22899 );
not \U$23259 ( \23505 , \4893 );
or \U$23260 ( \23506 , \23504 , \23505 );
nand \U$23261 ( \23507 , \2707 , \23106 );
nand \U$23262 ( \23508 , \23506 , \23507 );
xor \U$23263 ( \23509 , \23503 , \23508 );
not \U$23264 ( \23510 , \23509 );
or \U$23265 ( \23511 , \23498 , \23510 );
nand \U$23266 ( \23512 , \23508 , \23503 );
nand \U$23267 ( \23513 , \23511 , \23512 );
xor \U$23268 ( \23514 , \23492 , \23513 );
and \U$23269 ( \23515 , \9268 , \23205 );
not \U$23270 ( \23516 , \22931 );
nor \U$23271 ( \23517 , \23516 , \11544 );
nor \U$23272 ( \23518 , \23515 , \23517 );
not \U$23273 ( \23519 , \23518 );
not \U$23274 ( \23520 , \23519 );
nand \U$23275 ( \23521 , \885 , RIbe2ae38_110);
not \U$23276 ( \23522 , \23521 );
not \U$23277 ( \23523 , \22884 );
or \U$23278 ( \23524 , \12027 , \23523 );
nand \U$23279 ( \23525 , \5055 , \23078 );
nand \U$23280 ( \23526 , \23524 , \23525 );
not \U$23281 ( \23527 , \23526 );
or \U$23282 ( \23528 , \23522 , \23527 );
or \U$23283 ( \23529 , \23526 , \23521 );
nand \U$23284 ( \23530 , \23528 , \23529 );
not \U$23285 ( \23531 , \23530 );
or \U$23286 ( \23532 , \23520 , \23531 );
not \U$23287 ( \23533 , \23521 );
nand \U$23288 ( \23534 , \23533 , \23526 );
nand \U$23289 ( \23535 , \23532 , \23534 );
xor \U$23290 ( \23536 , \23514 , \23535 );
not \U$23291 ( \23537 , \23536 );
not \U$23292 ( \23538 , \23005 );
not \U$23293 ( \23539 , \2599 );
or \U$23294 ( \23540 , \23538 , \23539 );
nand \U$23295 ( \23541 , \13306 , \23192 );
nand \U$23296 ( \23542 , \23540 , \23541 );
xor \U$23297 ( \23543 , RIbe285e8_24, RIbe2b540_125);
not \U$23298 ( \23544 , \23543 );
not \U$23299 ( \23545 , \2618 );
or \U$23300 ( \23546 , \23544 , \23545 );
nand \U$23301 ( \23547 , \8270 , \23137 );
nand \U$23302 ( \23548 , \23546 , \23547 );
xor \U$23303 ( \23549 , \23542 , \23548 );
xor \U$23304 ( \23550 , RIbe2a028_80, RIbe2aa78_102);
not \U$23305 ( \23551 , \23550 );
not \U$23306 ( \23552 , \14513 );
or \U$23307 ( \23553 , \23551 , \23552 );
nand \U$23308 ( \23554 , \8172 , \23417 );
nand \U$23309 ( \23555 , \23553 , \23554 );
and \U$23310 ( \23556 , \23549 , \23555 );
and \U$23311 ( \23557 , \23542 , \23548 );
or \U$23312 ( \23558 , \23556 , \23557 );
xor \U$23313 ( \23559 , RIbe2af28_112, RIbe291a0_49);
not \U$23314 ( \23560 , \23559 );
not \U$23315 ( \23561 , \15345 );
or \U$23316 ( \23562 , \23560 , \23561 );
nand \U$23317 ( \23563 , \17811 , \23199 );
nand \U$23318 ( \23564 , \23562 , \23563 );
not \U$23319 ( \23565 , \23564 );
not \U$23320 ( \23566 , \22971 );
not \U$23321 ( \23567 , \10433 );
or \U$23322 ( \23568 , \23566 , \23567 );
nand \U$23323 ( \23569 , \20336 , \23223 );
nand \U$23324 ( \23570 , \23568 , \23569 );
not \U$23325 ( \23571 , \22966 );
not \U$23326 ( \23572 , \14852 );
or \U$23327 ( \23573 , \23571 , \23572 );
nand \U$23328 ( \23574 , \16646 , \22771 );
nand \U$23329 ( \23575 , \23573 , \23574 );
xor \U$23330 ( \23576 , \23570 , \23575 );
not \U$23331 ( \23577 , \23576 );
or \U$23332 ( \23578 , \23565 , \23577 );
nand \U$23333 ( \23579 , \23570 , \23575 );
nand \U$23334 ( \23580 , \23578 , \23579 );
xor \U$23335 ( \23581 , \23558 , \23580 );
buf \U$23336 ( \23582 , \13529 );
and \U$23337 ( \23583 , \23582 , \23016 );
not \U$23338 ( \23584 , \23114 );
nor \U$23339 ( \23585 , \23584 , \13538 );
nor \U$23340 ( \23586 , \23583 , \23585 );
not \U$23341 ( \23587 , \23586 );
not \U$23342 ( \23588 , \23587 );
not \U$23343 ( \23589 , \22954 );
not \U$23344 ( \23590 , \11461 );
or \U$23345 ( \23591 , \23589 , \23590 );
nand \U$23346 ( \23592 , \4180 , \23095 );
nand \U$23347 ( \23593 , \23591 , \23592 );
not \U$23348 ( \23594 , \22997 );
not \U$23349 ( \23595 , \20395 );
or \U$23350 ( \23596 , \23594 , \23595 );
nand \U$23351 ( \23597 , \15953 , \22761 );
nand \U$23352 ( \23598 , \23596 , \23597 );
and \U$23353 ( \23599 , \23593 , \23598 );
not \U$23354 ( \23600 , \23593 );
not \U$23355 ( \23601 , \23598 );
and \U$23356 ( \23602 , \23600 , \23601 );
nor \U$23357 ( \23603 , \23599 , \23602 );
not \U$23358 ( \23604 , \23603 );
or \U$23359 ( \23605 , \23588 , \23604 );
not \U$23360 ( \23606 , \23601 );
nand \U$23361 ( \23607 , \23606 , \23593 );
nand \U$23362 ( \23608 , \23605 , \23607 );
not \U$23363 ( \23609 , \23608 );
xor \U$23364 ( \23610 , \23581 , \23609 );
nand \U$23365 ( \23611 , \23537 , \23610 );
not \U$23366 ( \23612 , \23610 );
nand \U$23367 ( \23613 , \23612 , \23536 );
nand \U$23368 ( \23614 , \23611 , \23613 );
xor \U$23369 ( \23615 , \23365 , \23358 );
xnor \U$23370 ( \23616 , \23615 , \23350 );
not \U$23371 ( \23617 , \23616 );
not \U$23372 ( \23618 , \23530 );
not \U$23373 ( \23619 , \23518 );
and \U$23374 ( \23620 , \23618 , \23619 );
and \U$23375 ( \23621 , \23530 , \23518 );
nor \U$23376 ( \23622 , \23620 , \23621 );
not \U$23377 ( \23623 , \23622 );
or \U$23378 ( \23624 , \23617 , \23623 );
or \U$23379 ( \23625 , \23622 , \23616 );
nand \U$23380 ( \23626 , \23624 , \23625 );
not \U$23381 ( \23627 , \23626 );
xnor \U$23382 ( \23628 , \23509 , \23497 );
not \U$23383 ( \23629 , \23628 );
not \U$23384 ( \23630 , \23629 );
or \U$23385 ( \23631 , \23627 , \23630 );
not \U$23386 ( \23632 , \23622 );
nand \U$23387 ( \23633 , \23632 , \23616 );
nand \U$23388 ( \23634 , \23631 , \23633 );
xnor \U$23389 ( \23635 , \23614 , \23634 );
not \U$23390 ( \23636 , \23635 );
not \U$23391 ( \23637 , \23603 );
not \U$23392 ( \23638 , \23586 );
and \U$23393 ( \23639 , \23637 , \23638 );
and \U$23394 ( \23640 , \23603 , \23586 );
nor \U$23395 ( \23641 , \23639 , \23640 );
xor \U$23396 ( \23642 , \23542 , \23548 );
xor \U$23397 ( \23643 , \23642 , \23555 );
and \U$23398 ( \23644 , \23641 , \23643 );
not \U$23399 ( \23645 , \23641 );
not \U$23400 ( \23646 , \23643 );
and \U$23401 ( \23647 , \23645 , \23646 );
or \U$23402 ( \23648 , \23644 , \23647 );
not \U$23403 ( \23649 , \23397 );
not \U$23404 ( \23650 , \23377 );
not \U$23405 ( \23651 , \23650 );
and \U$23406 ( \23652 , \23649 , \23651 );
and \U$23407 ( \23653 , \23397 , \23650 );
nor \U$23408 ( \23654 , \23652 , \23653 );
buf \U$23409 ( \23655 , \23654 );
and \U$23410 ( \23656 , \23648 , \23655 );
not \U$23411 ( \23657 , \23648 );
not \U$23412 ( \23658 , \23655 );
and \U$23413 ( \23659 , \23657 , \23658 );
nor \U$23414 ( \23660 , \23656 , \23659 );
not \U$23415 ( \23661 , \23660 );
not \U$23416 ( \23662 , \23661 );
not \U$23417 ( \23663 , \23626 );
not \U$23418 ( \23664 , \23628 );
and \U$23419 ( \23665 , \23663 , \23664 );
and \U$23420 ( \23666 , \23626 , \23628 );
nor \U$23421 ( \23667 , \23665 , \23666 );
not \U$23422 ( \23668 , \23667 );
not \U$23423 ( \23669 , \23668 );
or \U$23424 ( \23670 , \23662 , \23669 );
not \U$23425 ( \23671 , \23660 );
not \U$23426 ( \23672 , \23667 );
or \U$23427 ( \23673 , \23671 , \23672 );
xor \U$23428 ( \23674 , \22879 , \22886 );
xor \U$23429 ( \23675 , RIbe2af28_112, RIbe29128_48);
not \U$23430 ( \23676 , \23675 );
not \U$23431 ( \23677 , \15345 );
or \U$23432 ( \23678 , \23676 , \23677 );
nand \U$23433 ( \23679 , \14413 , \23559 );
nand \U$23434 ( \23680 , \23678 , \23679 );
xor \U$23435 ( \23681 , \23674 , \23680 );
xor \U$23436 ( \23682 , RIbe27e68_8, RIbe2b540_125);
not \U$23437 ( \23683 , \23682 );
not \U$23438 ( \23684 , \2459 );
or \U$23439 ( \23685 , \23683 , \23684 );
nand \U$23440 ( \23686 , \4447 , \23001 );
nand \U$23441 ( \23687 , \23685 , \23686 );
not \U$23442 ( \23688 , \23687 );
xor \U$23443 ( \23689 , RIbe27fd0_11, RIbe2adc0_109);
not \U$23444 ( \23690 , \23689 );
not \U$23445 ( \23691 , \9825 );
or \U$23446 ( \23692 , \23690 , \23691 );
nand \U$23447 ( \23693 , \2707 , \22895 );
nand \U$23448 ( \23694 , \23692 , \23693 );
xor \U$23449 ( \23695 , RIbe29f38_78, RIbe2a3e8_88);
not \U$23450 ( \23696 , \23695 );
not \U$23451 ( \23697 , \9262 );
or \U$23452 ( \23698 , \23696 , \23697 );
nand \U$23453 ( \23699 , \8794 , \22927 );
nand \U$23454 ( \23700 , \23698 , \23699 );
nor \U$23455 ( \23701 , \23694 , \23700 );
not \U$23456 ( \23702 , \23701 );
not \U$23457 ( \23703 , \23702 );
or \U$23458 ( \23704 , \23688 , \23703 );
nand \U$23459 ( \23705 , \23694 , \23700 );
nand \U$23460 ( \23706 , \23704 , \23705 );
xor \U$23461 ( \23707 , \23681 , \23706 );
not \U$23462 ( \23708 , \23707 );
xor \U$23463 ( \23709 , RIbe2af28_112, RIbe29b00_69);
not \U$23464 ( \23710 , \23709 );
not \U$23465 ( \23711 , \15345 );
or \U$23466 ( \23712 , \23710 , \23711 );
nand \U$23467 ( \23713 , \17811 , \23675 );
nand \U$23468 ( \23714 , \23712 , \23713 );
not \U$23469 ( \23715 , \9379 );
not \U$23470 ( \23716 , \22888 );
or \U$23471 ( \23717 , \23715 , \23716 );
xnor \U$23472 ( \23718 , RIbe2a2f8_86, RIbe2aa78_102);
or \U$23473 ( \23719 , \8696 , \23718 );
nand \U$23474 ( \23720 , \23717 , \23719 );
nor \U$23475 ( \23721 , \23714 , \23720 );
not \U$23476 ( \23722 , \23721 );
not \U$23477 ( \23723 , \23722 );
not \U$23478 ( \23724 , \2559 );
xor \U$23479 ( \23725 , RIbe2b450_123, RIbe28b88_36);
not \U$23480 ( \23726 , \23725 );
or \U$23481 ( \23727 , \23724 , \23726 );
not \U$23482 ( \23728 , \2553 );
xor \U$23483 ( \23729 , RIbe28b88_36, RIbe2b3d8_122);
not \U$23484 ( \23730 , \23729 );
or \U$23485 ( \23731 , \23728 , \23730 );
nand \U$23486 ( \23732 , \23727 , \23731 );
or \U$23487 ( \23733 , RIbe28b88_36, RIbe29290_51);
nand \U$23488 ( \23734 , \23733 , RIbe2ae38_110);
nand \U$23489 ( \23735 , RIbe28b88_36, RIbe29290_51);
and \U$23490 ( \23736 , \23734 , \23735 , RIbe28a20_33);
nand \U$23491 ( \23737 , \23732 , \23736 );
not \U$23492 ( \23738 , \23737 );
not \U$23493 ( \23739 , \23738 );
or \U$23494 ( \23740 , \23723 , \23739 );
nand \U$23495 ( \23741 , \23714 , \23720 );
nand \U$23496 ( \23742 , \23740 , \23741 );
not \U$23497 ( \23743 , \23742 );
xor \U$23498 ( \23744 , RIbe2a0a0_81, RIbe29c68_72);
not \U$23499 ( \23745 , \23744 );
not \U$23500 ( \23746 , \8595 );
or \U$23501 ( \23747 , \23745 , \23746 );
nand \U$23502 ( \23748 , \4580 , \23483 );
nand \U$23503 ( \23749 , \23747 , \23748 );
xor \U$23504 ( \23750 , RIbe28b88_36, RIbe2a730_95);
not \U$23505 ( \23751 , \23750 );
not \U$23506 ( \23752 , \3401 );
or \U$23507 ( \23753 , \23751 , \23752 );
not \U$23508 ( \23754 , \23474 );
nand \U$23509 ( \23755 , \23754 , \2691 );
nand \U$23510 ( \23756 , \23753 , \23755 );
xor \U$23511 ( \23757 , \23749 , \23756 );
xor \U$23512 ( \23758 , RIbe2abe0_105, RIbe28390_19);
not \U$23513 ( \23759 , \23758 );
not \U$23514 ( \23760 , \2640 );
or \U$23515 ( \23761 , \23759 , \23760 );
nand \U$23516 ( \23762 , \2648 , \23379 );
nand \U$23517 ( \23763 , \23761 , \23762 );
xnor \U$23518 ( \23764 , \23757 , \23763 );
not \U$23519 ( \23765 , \23764 );
or \U$23520 ( \23766 , \23743 , \23765 );
or \U$23521 ( \23767 , \23764 , \23742 );
nand \U$23522 ( \23768 , \23766 , \23767 );
not \U$23523 ( \23769 , \23768 );
or \U$23524 ( \23770 , \23708 , \23769 );
not \U$23525 ( \23771 , \23764 );
nand \U$23526 ( \23772 , \23771 , \23742 );
nand \U$23527 ( \23773 , \23770 , \23772 );
nand \U$23528 ( \23774 , \23673 , \23773 );
nand \U$23529 ( \23775 , \23670 , \23774 );
not \U$23530 ( \23776 , \23775 );
and \U$23531 ( \23777 , \23370 , \23343 );
not \U$23532 ( \23778 , \23370 );
and \U$23533 ( \23779 , \23778 , \23403 );
nor \U$23534 ( \23780 , \23777 , \23779 );
not \U$23535 ( \23781 , \23401 );
and \U$23536 ( \23782 , \23780 , \23781 );
not \U$23537 ( \23783 , \23780 );
and \U$23538 ( \23784 , \23783 , \23401 );
nor \U$23539 ( \23785 , \23782 , \23784 );
not \U$23540 ( \23786 , \23785 );
not \U$23541 ( \23787 , \23786 );
not \U$23542 ( \23788 , \23646 );
not \U$23543 ( \23789 , \23654 );
or \U$23544 ( \23790 , \23788 , \23789 );
not \U$23545 ( \23791 , \23641 );
nand \U$23546 ( \23792 , \23790 , \23791 );
not \U$23547 ( \23793 , \23654 );
nand \U$23548 ( \23794 , \23793 , \23643 );
nand \U$23549 ( \23795 , \23792 , \23794 );
not \U$23550 ( \23796 , \23795 );
not \U$23551 ( \23797 , \23796 );
or \U$23552 ( \23798 , \23787 , \23797 );
nand \U$23553 ( \23799 , \23785 , \23795 );
nand \U$23554 ( \23800 , \23798 , \23799 );
not \U$23555 ( \23801 , \23749 );
not \U$23556 ( \23802 , \23756 );
or \U$23557 ( \23803 , \23801 , \23802 );
or \U$23558 ( \23804 , \23756 , \23749 );
nand \U$23559 ( \23805 , \23804 , \23763 );
nand \U$23560 ( \23806 , \23803 , \23805 );
not \U$23561 ( \23807 , \23806 );
not \U$23562 ( \23808 , \23576 );
not \U$23563 ( \23809 , \23564 );
not \U$23564 ( \23810 , \23809 );
and \U$23565 ( \23811 , \23808 , \23810 );
and \U$23566 ( \23812 , \23576 , \23809 );
nor \U$23567 ( \23813 , \23811 , \23812 );
not \U$23568 ( \23814 , \23813 );
not \U$23569 ( \23815 , \23814 );
xor \U$23570 ( \23816 , RIbe285e8_24, RIbe2b4c8_124);
not \U$23571 ( \23817 , \23816 );
not \U$23572 ( \23818 , \2890 );
or \U$23573 ( \23819 , \23817 , \23818 );
nand \U$23574 ( \23820 , \2626 , \23543 );
nand \U$23575 ( \23821 , \23819 , \23820 );
not \U$23576 ( \23822 , \23821 );
xor \U$23577 ( \23823 , RIbe28480_21, RIbe2a640_93);
not \U$23578 ( \23824 , \23823 );
not \U$23579 ( \23825 , \2518 );
or \U$23580 ( \23826 , \23824 , \23825 );
nand \U$23581 ( \23827 , \7483 , \23345 );
nand \U$23582 ( \23828 , \23826 , \23827 );
not \U$23583 ( \23829 , \23828 );
not \U$23584 ( \23830 , \23829 );
xor \U$23585 ( \23831 , RIbe2a028_80, RIbe2aa00_101);
not \U$23586 ( \23832 , \23831 );
not \U$23587 ( \23833 , \10674 );
or \U$23588 ( \23834 , \23832 , \23833 );
nand \U$23589 ( \23835 , \9065 , \23550 );
nand \U$23590 ( \23836 , \23834 , \23835 );
not \U$23591 ( \23837 , \23836 );
or \U$23592 ( \23838 , \23830 , \23837 );
or \U$23593 ( \23839 , \23836 , \23829 );
nand \U$23594 ( \23840 , \23838 , \23839 );
not \U$23595 ( \23841 , \23840 );
or \U$23596 ( \23842 , \23822 , \23841 );
not \U$23597 ( \23843 , \23829 );
nand \U$23598 ( \23844 , \23843 , \23836 );
nand \U$23599 ( \23845 , \23842 , \23844 );
not \U$23600 ( \23846 , \23845 );
not \U$23601 ( \23847 , \23846 );
or \U$23602 ( \23848 , \23815 , \23847 );
nand \U$23603 ( \23849 , \23813 , \23845 );
nand \U$23604 ( \23850 , \23848 , \23849 );
not \U$23605 ( \23851 , \23850 );
or \U$23606 ( \23852 , \23807 , \23851 );
nand \U$23607 ( \23853 , \23814 , \23845 );
nand \U$23608 ( \23854 , \23852 , \23853 );
not \U$23609 ( \23855 , \23854 );
and \U$23610 ( \23856 , \23800 , \23855 );
not \U$23611 ( \23857 , \23800 );
and \U$23612 ( \23858 , \23857 , \23854 );
nor \U$23613 ( \23859 , \23856 , \23858 );
not \U$23614 ( \23860 , \23859 );
or \U$23615 ( \23861 , \23776 , \23860 );
or \U$23616 ( \23862 , \23775 , \23859 );
nand \U$23617 ( \23863 , \23861 , \23862 );
not \U$23618 ( \23864 , \23863 );
or \U$23619 ( \23865 , \23636 , \23864 );
not \U$23620 ( \23866 , \23859 );
nand \U$23621 ( \23867 , \23866 , \23775 );
nand \U$23622 ( \23868 , \23865 , \23867 );
not \U$23623 ( \23869 , \23868 );
not \U$23624 ( \23870 , \23869 );
xor \U$23625 ( \23871 , \22887 , \22916 );
xor \U$23626 ( \23872 , \23871 , \22944 );
xor \U$23627 ( \23873 , \22926 , \22933 );
xor \U$23628 ( \23874 , \23873 , \22941 );
xor \U$23629 ( \23875 , \23821 , \23840 );
xor \U$23630 ( \23876 , \23874 , \23875 );
not \U$23631 ( \23877 , \22959 );
not \U$23632 ( \23878 , \22982 );
or \U$23633 ( \23879 , \23877 , \23878 );
or \U$23634 ( \23880 , \22982 , \22959 );
nand \U$23635 ( \23881 , \23879 , \23880 );
and \U$23636 ( \23882 , \23876 , \23881 );
and \U$23637 ( \23883 , \23874 , \23875 );
or \U$23638 ( \23884 , \23882 , \23883 );
xor \U$23639 ( \23885 , \23872 , \23884 );
and \U$23640 ( \23886 , \23063 , \22987 );
not \U$23641 ( \23887 , \23063 );
not \U$23642 ( \23888 , \22987 );
and \U$23643 ( \23889 , \23887 , \23888 );
nor \U$23644 ( \23890 , \23886 , \23889 );
xnor \U$23645 ( \23891 , \23885 , \23890 );
not \U$23646 ( \23892 , \23891 );
not \U$23647 ( \23893 , \23892 );
xor \U$23648 ( \23894 , \22894 , \22901 );
xor \U$23649 ( \23895 , \23894 , \22913 );
xor \U$23650 ( \23896 , \22999 , \23018 );
xnor \U$23651 ( \23897 , \23896 , \23007 );
xor \U$23652 ( \23898 , \23895 , \23897 );
xor \U$23653 ( \23899 , \23044 , \23054 );
xnor \U$23654 ( \23900 , \23898 , \23899 );
not \U$23655 ( \23901 , \23900 );
xor \U$23656 ( \23902 , \23874 , \23875 );
xor \U$23657 ( \23903 , \23902 , \23881 );
not \U$23658 ( \23904 , \23903 );
or \U$23659 ( \23905 , \23901 , \23904 );
or \U$23660 ( \23906 , \23903 , \23900 );
not \U$23661 ( \23907 , \23738 );
not \U$23662 ( \23908 , \23721 );
nand \U$23663 ( \23909 , \23908 , \23741 );
not \U$23664 ( \23910 , \23909 );
or \U$23665 ( \23911 , \23907 , \23910 );
or \U$23666 ( \23912 , \23909 , \23738 );
nand \U$23667 ( \23913 , \23911 , \23912 );
not \U$23668 ( \23914 , \23913 );
not \U$23669 ( \23915 , RIbe29e48_76);
not \U$23670 ( \23916 , RIbe2a118_82);
and \U$23671 ( \23917 , \23915 , \23916 );
and \U$23672 ( \23918 , RIbe29e48_76, RIbe2a118_82);
nor \U$23673 ( \23919 , \23917 , \23918 );
and \U$23674 ( \23920 , \11040 , \23919 );
and \U$23675 ( \23921 , \8245 , \23022 );
nor \U$23676 ( \23922 , \23920 , \23921 );
not \U$23677 ( \23923 , \23922 );
xor \U$23678 ( \23924 , RIbe29740_61, RIbe2aaf0_103);
and \U$23679 ( \23925 , \20574 , \23924 );
not \U$23680 ( \23926 , RIbe2ab68_104);
nor \U$23681 ( \23927 , \23926 , \23035 );
nor \U$23682 ( \23928 , \23925 , \23927 );
not \U$23683 ( \23929 , \23928 );
xor \U$23684 ( \23930 , RIbe2a7a8_96, RIbe28390_19);
not \U$23685 ( \23931 , \23930 );
not \U$23686 ( \23932 , \14806 );
or \U$23687 ( \23933 , \23931 , \23932 );
nand \U$23688 ( \23934 , \3714 , \23758 );
nand \U$23689 ( \23935 , \23933 , \23934 );
not \U$23690 ( \23936 , \23935 );
or \U$23691 ( \23937 , \23929 , \23936 );
or \U$23692 ( \23938 , \23935 , \23928 );
nand \U$23693 ( \23939 , \23937 , \23938 );
not \U$23694 ( \23940 , \23939 );
or \U$23695 ( \23941 , \23923 , \23940 );
or \U$23696 ( \23942 , \23939 , \23922 );
nand \U$23697 ( \23943 , \23941 , \23942 );
not \U$23698 ( \23944 , \23943 );
xor \U$23699 ( \23945 , RIbe29218_50, RIbe2b180_117);
not \U$23700 ( \23946 , \23945 );
not \U$23701 ( \23947 , \14852 );
or \U$23702 ( \23948 , \23946 , \23947 );
nand \U$23703 ( \23949 , \14966 , \22962 );
nand \U$23704 ( \23950 , \23948 , \23949 );
not \U$23705 ( \23951 , \23950 );
xor \U$23706 ( \23952 , RIbe28cf0_39, RIbe2a190_83);
not \U$23707 ( \23953 , \23952 );
not \U$23708 ( \23954 , \11396 );
or \U$23709 ( \23955 , \23953 , \23954 );
nand \U$23710 ( \23956 , \10696 , \22923 );
nand \U$23711 ( \23957 , \23955 , \23956 );
not \U$23712 ( \23958 , \23957 );
not \U$23713 ( \23959 , \23958 );
or \U$23714 ( \23960 , \23951 , \23959 );
not \U$23715 ( \23961 , \23950 );
nand \U$23716 ( \23962 , \23961 , \23957 );
nand \U$23717 ( \23963 , \23960 , \23962 );
xor \U$23718 ( \23964 , RIbe29c68_72, RIbe2b360_121);
not \U$23719 ( \23965 , \23964 );
not \U$23720 ( \23966 , \8595 );
or \U$23721 ( \23967 , \23965 , \23966 );
nand \U$23722 ( \23968 , \4580 , \23744 );
nand \U$23723 ( \23969 , \23967 , \23968 );
xnor \U$23724 ( \23970 , \23963 , \23969 );
not \U$23725 ( \23971 , \23970 );
and \U$23726 ( \23972 , \23944 , \23971 );
and \U$23727 ( \23973 , \23943 , \23970 );
nor \U$23728 ( \23974 , \23972 , \23973 );
not \U$23729 ( \23975 , \23974 );
not \U$23730 ( \23976 , \23975 );
or \U$23731 ( \23977 , \23914 , \23976 );
not \U$23732 ( \23978 , \23970 );
nand \U$23733 ( \23979 , \23978 , \23943 );
nand \U$23734 ( \23980 , \23977 , \23979 );
nand \U$23735 ( \23981 , \23906 , \23980 );
nand \U$23736 ( \23982 , \23905 , \23981 );
not \U$23737 ( \23983 , \23982 );
or \U$23738 ( \23984 , \23893 , \23983 );
not \U$23739 ( \23985 , \23982 );
not \U$23740 ( \23986 , \23985 );
not \U$23741 ( \23987 , \23891 );
or \U$23742 ( \23988 , \23986 , \23987 );
not \U$23743 ( \23989 , \23961 );
not \U$23744 ( \23990 , \23958 );
or \U$23745 ( \23991 , \23989 , \23990 );
nand \U$23746 ( \23992 , \23991 , \23969 );
not \U$23747 ( \23993 , \23958 );
nand \U$23748 ( \23994 , \23993 , \23950 );
nand \U$23749 ( \23995 , \23992 , \23994 );
and \U$23750 ( \23996 , RIbe29b78_70, RIbe2a550_91);
nor \U$23751 ( \23997 , RIbe29b78_70, RIbe2a550_91);
nor \U$23752 ( \23998 , \23996 , \23997 );
not \U$23753 ( \23999 , \23998 );
not \U$23754 ( \24000 , \10434 );
or \U$23755 ( \24001 , \23999 , \24000 );
nand \U$23756 ( \24002 , \11228 , \22976 );
nand \U$23757 ( \24003 , \24001 , \24002 );
not \U$23758 ( \24004 , \24003 );
xor \U$23759 ( \24005 , RIbe2a898_98, RIbe2a028_80);
not \U$23760 ( \24006 , \24005 );
not \U$23761 ( \24007 , \10674 );
or \U$23762 ( \24008 , \24006 , \24007 );
nand \U$23763 ( \24009 , \8930 , \23831 );
nand \U$23764 ( \24010 , \24008 , \24009 );
xor \U$23765 ( \24011 , RIbe28f48_44, RIbe2a4d8_90);
not \U$23766 ( \24012 , \24011 );
not \U$23767 ( \24013 , \8221 );
or \U$23768 ( \24014 , \24012 , \24013 );
nand \U$23769 ( \24015 , \11201 , \22956 );
nand \U$23770 ( \24016 , \24014 , \24015 );
and \U$23771 ( \24017 , \24010 , \24016 );
not \U$23772 ( \24018 , \24010 );
not \U$23773 ( \24019 , \24016 );
and \U$23774 ( \24020 , \24018 , \24019 );
nor \U$23775 ( \24021 , \24017 , \24020 );
not \U$23776 ( \24022 , \24021 );
or \U$23777 ( \24023 , \24004 , \24022 );
not \U$23778 ( \24024 , \24019 );
nand \U$23779 ( \24025 , \24024 , \24010 );
nand \U$23780 ( \24026 , \24023 , \24025 );
xor \U$23781 ( \24027 , \23995 , \24026 );
buf \U$23782 ( \24028 , \23353 );
buf \U$23783 ( \24029 , \24028 );
xor \U$23784 ( \24030 , RIbe2a280_85, RIbe29998_66);
and \U$23785 ( \24031 , \24029 , \24030 );
and \U$23786 ( \24032 , \11348 , \23052 );
nor \U$23787 ( \24033 , \24031 , \24032 );
not \U$23788 ( \24034 , \24033 );
not \U$23789 ( \24035 , \24034 );
xor \U$23790 ( \24036 , RIbe2ac58_106, RIbe28480_21);
not \U$23791 ( \24037 , \24036 );
not \U$23792 ( \24038 , \2518 );
or \U$23793 ( \24039 , \24037 , \24038 );
nand \U$23794 ( \24040 , \11263 , \23823 );
nand \U$23795 ( \24041 , \24039 , \24040 );
xor \U$23796 ( \24042 , RIbe2aeb0_111, RIbe28a20_33);
not \U$23797 ( \24043 , \24042 );
not \U$23798 ( \24044 , \1780 );
or \U$23799 ( \24045 , \24043 , \24044 );
nand \U$23800 ( \24046 , \2475 , \22880 );
nand \U$23801 ( \24047 , \24045 , \24046 );
xor \U$23802 ( \24048 , \24041 , \24047 );
not \U$23803 ( \24049 , \24048 );
or \U$23804 ( \24050 , \24035 , \24049 );
nand \U$23805 ( \24051 , \24047 , \24041 );
nand \U$23806 ( \24052 , \24050 , \24051 );
and \U$23807 ( \24053 , \24027 , \24052 );
and \U$23808 ( \24054 , \23995 , \24026 );
or \U$23809 ( \24055 , \24053 , \24054 );
not \U$23810 ( \24056 , \24055 );
not \U$23811 ( \24057 , \24056 );
not \U$23812 ( \24058 , \23895 );
not \U$23813 ( \24059 , \23897 );
not \U$23814 ( \24060 , \24059 );
or \U$23815 ( \24061 , \24058 , \24060 );
or \U$23816 ( \24062 , \24059 , \23895 );
nand \U$23817 ( \24063 , \24062 , \23899 );
nand \U$23818 ( \24064 , \24061 , \24063 );
not \U$23819 ( \24065 , \24064 );
or \U$23820 ( \24066 , \24057 , \24065 );
not \U$23821 ( \24067 , \24064 );
nand \U$23822 ( \24068 , \24055 , \24067 );
nand \U$23823 ( \24069 , \24066 , \24068 );
xor \U$23824 ( \24070 , \23850 , \23806 );
and \U$23825 ( \24071 , \24069 , \24070 );
not \U$23826 ( \24072 , \24069 );
not \U$23827 ( \24073 , \24070 );
and \U$23828 ( \24074 , \24072 , \24073 );
nor \U$23829 ( \24075 , \24071 , \24074 );
nand \U$23830 ( \24076 , \23988 , \24075 );
nand \U$23831 ( \24077 , \23984 , \24076 );
not \U$23832 ( \24078 , \24077 );
not \U$23833 ( \24079 , \23681 );
not \U$23834 ( \24080 , \23706 );
or \U$23835 ( \24081 , \24079 , \24080 );
nand \U$23836 ( \24082 , \23674 , \23680 );
nand \U$23837 ( \24083 , \24081 , \24082 );
not \U$23838 ( \24084 , \24083 );
not \U$23839 ( \24085 , \23482 );
nand \U$23840 ( \24086 , \24085 , \23491 );
xnor \U$23841 ( \24087 , \23489 , \24086 );
not \U$23842 ( \24088 , \24087 );
or \U$23843 ( \24089 , \24084 , \24088 );
or \U$23844 ( \24090 , \24083 , \24087 );
nand \U$23845 ( \24091 , \24089 , \24090 );
not \U$23846 ( \24092 , \24091 );
not \U$23847 ( \24093 , RIbe291a0_49);
not \U$23848 ( \24094 , RIbe2b018_114);
and \U$23849 ( \24095 , \24093 , \24094 );
and \U$23850 ( \24096 , RIbe291a0_49, RIbe2b018_114);
nor \U$23851 ( \24097 , \24095 , \24096 );
not \U$23852 ( \24098 , \24097 );
not \U$23853 ( \24099 , \22763 );
or \U$23854 ( \24100 , \24098 , \24099 );
nand \U$23855 ( \24101 , \20583 , \22989 );
nand \U$23856 ( \24102 , \24100 , \24101 );
not \U$23857 ( \24103 , \24102 );
xor \U$23858 ( \24104 , RIbe285e8_24, RIbe2a6b8_94);
not \U$23859 ( \24105 , \24104 );
not \U$23860 ( \24106 , \10863 );
or \U$23861 ( \24107 , \24105 , \24106 );
nand \U$23862 ( \24108 , \8270 , \23816 );
nand \U$23863 ( \24109 , \24107 , \24108 );
not \U$23864 ( \24110 , \24109 );
not \U$23865 ( \24111 , \24110 );
xor \U$23866 ( \24112 , RIbe27c88_4, RIbe2b108_116);
not \U$23867 ( \24113 , \24112 );
not \U$23868 ( \24114 , \14296 );
or \U$23869 ( \24115 , \24113 , \24114 );
nand \U$23870 ( \24116 , \13533 , \23011 );
nand \U$23871 ( \24117 , \24115 , \24116 );
not \U$23872 ( \24118 , \24117 );
or \U$23873 ( \24119 , \24111 , \24118 );
or \U$23874 ( \24120 , \24110 , \24117 );
nand \U$23875 ( \24121 , \24119 , \24120 );
not \U$23876 ( \24122 , \24121 );
or \U$23877 ( \24123 , \24103 , \24122 );
nand \U$23878 ( \24124 , \24117 , \24109 );
nand \U$23879 ( \24125 , \24123 , \24124 );
not \U$23880 ( \24126 , \23725 );
not \U$23881 ( \24127 , \9052 );
or \U$23882 ( \24128 , \24126 , \24127 );
nand \U$23883 ( \24129 , \23750 , \2559 );
nand \U$23884 ( \24130 , \24128 , \24129 );
and \U$23885 ( \24131 , \970 , RIbe2ae38_110);
or \U$23886 ( \24132 , \24130 , \24131 );
xor \U$23887 ( \24133 , RIbe2a910_99, RIbe29d58_74);
not \U$23888 ( \24134 , \24133 );
not \U$23889 ( \24135 , \9737 );
or \U$23890 ( \24136 , \24134 , \24135 );
nand \U$23891 ( \24137 , \11456 , \22903 );
nand \U$23892 ( \24138 , \24136 , \24137 );
nand \U$23893 ( \24139 , \24132 , \24138 );
nand \U$23894 ( \24140 , \24130 , \24131 );
nand \U$23895 ( \24141 , \24139 , \24140 );
or \U$23896 ( \24142 , \24125 , \24141 );
not \U$23897 ( \24143 , \23922 );
not \U$23898 ( \24144 , \24143 );
not \U$23899 ( \24145 , \23939 );
or \U$23900 ( \24146 , \24144 , \24145 );
not \U$23901 ( \24147 , \23928 );
nand \U$23902 ( \24148 , \24147 , \23935 );
nand \U$23903 ( \24149 , \24146 , \24148 );
nand \U$23904 ( \24150 , \24142 , \24149 );
nand \U$23905 ( \24151 , \24125 , \24141 );
nand \U$23906 ( \24152 , \24150 , \24151 );
not \U$23907 ( \24153 , \24152 );
or \U$23908 ( \24154 , \24092 , \24153 );
not \U$23909 ( \24155 , \24087 );
nand \U$23910 ( \24156 , \24155 , \24083 );
nand \U$23911 ( \24157 , \24154 , \24156 );
nand \U$23912 ( \24158 , \23454 , \23455 );
and \U$23913 ( \24159 , \24158 , \23461 );
not \U$23914 ( \24160 , \24158 );
not \U$23915 ( \24161 , \23461 );
and \U$23916 ( \24162 , \24160 , \24161 );
nor \U$23917 ( \24163 , \24159 , \24162 );
not \U$23918 ( \24164 , \24163 );
xor \U$23919 ( \24165 , \23438 , \23410 );
xor \U$23920 ( \24166 , \24165 , \23441 );
not \U$23921 ( \24167 , \24166 );
or \U$23922 ( \24168 , \24164 , \24167 );
or \U$23923 ( \24169 , \24163 , \24166 );
nand \U$23924 ( \24170 , \24168 , \24169 );
xor \U$23925 ( \24171 , \24157 , \24170 );
not \U$23926 ( \24172 , \24091 );
not \U$23927 ( \24173 , \24152 );
not \U$23928 ( \24174 , \24173 );
and \U$23929 ( \24175 , \24172 , \24174 );
and \U$23930 ( \24176 , \24173 , \24091 );
nor \U$23931 ( \24177 , \24175 , \24176 );
not \U$23932 ( \24178 , \24177 );
not \U$23933 ( \24179 , \24178 );
xor \U$23934 ( \24180 , \24125 , \24141 );
xnor \U$23935 ( \24181 , \24180 , \24149 );
xor \U$23936 ( \24182 , RIbe2af28_112, RIbe29a10_67);
not \U$23937 ( \24183 , \24182 );
not \U$23938 ( \24184 , \14423 );
or \U$23939 ( \24185 , \24183 , \24184 );
nand \U$23940 ( \24186 , \16728 , \23709 );
nand \U$23941 ( \24187 , \24185 , \24186 );
buf \U$23942 ( \24188 , \24187 );
xor \U$23943 ( \24189 , RIbe27b20_1, RIbe2a190_83);
and \U$23944 ( \24190 , \24189 , \10831 );
and \U$23945 ( \24191 , \10834 , \23952 );
nor \U$23946 ( \24192 , \24190 , \24191 );
not \U$23947 ( \24193 , \24192 );
or \U$23948 ( \24194 , \24188 , \24193 );
xor \U$23949 ( \24195 , RIbe2aa00_101, RIbe2a2f8_86);
not \U$23950 ( \24196 , \24195 );
not \U$23951 ( \24197 , \16714 );
or \U$23952 ( \24198 , \24196 , \24197 );
not \U$23953 ( \24199 , \23718 );
nand \U$23954 ( \24200 , \24199 , \9379 );
nand \U$23955 ( \24201 , \24198 , \24200 );
nand \U$23956 ( \24202 , \24194 , \24201 );
nand \U$23957 ( \24203 , \24188 , \24193 );
and \U$23958 ( \24204 , \24202 , \24203 );
not \U$23959 ( \24205 , \24204 );
xor \U$23960 ( \24206 , RIbe27fd0_11, RIbe2ad48_108);
not \U$23961 ( \24207 , \24206 );
not \U$23962 ( \24208 , \9082 );
or \U$23963 ( \24209 , \24207 , \24208 );
nand \U$23964 ( \24210 , \4897 , \23689 );
nand \U$23965 ( \24211 , \24209 , \24210 );
not \U$23966 ( \24212 , RIbe27df0_7);
not \U$23967 ( \24213 , RIbe2b180_117);
and \U$23968 ( \24214 , \24212 , \24213 );
and \U$23969 ( \24215 , RIbe27df0_7, RIbe2b180_117);
nor \U$23970 ( \24216 , \24214 , \24215 );
not \U$23971 ( \24217 , \24216 );
not \U$23972 ( \24218 , \17592 );
or \U$23973 ( \24219 , \24217 , \24218 );
nand \U$23974 ( \24220 , \14966 , \23945 );
nand \U$23975 ( \24221 , \24219 , \24220 );
xor \U$23976 ( \24222 , \24211 , \24221 );
xor \U$23977 ( \24223 , RIbe29c68_72, RIbe2b2e8_120);
not \U$23978 ( \24224 , \24223 );
not \U$23979 ( \24225 , \8594 );
or \U$23980 ( \24226 , \24224 , \24225 );
nand \U$23981 ( \24227 , \4580 , \23964 );
nand \U$23982 ( \24228 , \24226 , \24227 );
and \U$23983 ( \24229 , \24222 , \24228 );
and \U$23984 ( \24230 , \24211 , \24221 );
or \U$23985 ( \24231 , \24229 , \24230 );
not \U$23986 ( \24232 , \24231 );
not \U$23987 ( \24233 , \24232 );
or \U$23988 ( \24234 , \24205 , \24233 );
xor \U$23989 ( \24235 , RIbe2a3e8_88, RIbe2b6a8_128);
not \U$23990 ( \24236 , \24235 );
not \U$23991 ( \24237 , \8806 );
or \U$23992 ( \24238 , \24236 , \24237 );
nand \U$23993 ( \24239 , \9268 , \23695 );
nand \U$23994 ( \24240 , \24238 , \24239 );
xor \U$23995 ( \24241 , RIbe2b108_116, RIbe28d68_40);
not \U$23996 ( \24242 , \24241 );
not \U$23997 ( \24243 , \14297 );
or \U$23998 ( \24244 , \24242 , \24243 );
nand \U$23999 ( \24245 , \23015 , \24112 );
nand \U$24000 ( \24246 , \24244 , \24245 );
xor \U$24001 ( \24247 , \24240 , \24246 );
xor \U$24002 ( \24248 , RIbe2b4c8_124, RIbe27e68_8);
not \U$24003 ( \24249 , \24248 );
not \U$24004 ( \24250 , \2459 );
or \U$24005 ( \24251 , \24249 , \24250 );
nand \U$24006 ( \24252 , \2603 , \23682 );
nand \U$24007 ( \24253 , \24251 , \24252 );
and \U$24008 ( \24254 , \24247 , \24253 );
and \U$24009 ( \24255 , \24240 , \24246 );
or \U$24010 ( \24256 , \24254 , \24255 );
nand \U$24011 ( \24257 , \24234 , \24256 );
not \U$24012 ( \24258 , \24204 );
nand \U$24013 ( \24259 , \24258 , \24231 );
nand \U$24014 ( \24260 , \24257 , \24259 );
not \U$24015 ( \24261 , \24260 );
nand \U$24016 ( \24262 , \24181 , \24261 );
xor \U$24017 ( \24263 , RIbe28480_21, RIbe2abe0_105);
not \U$24018 ( \24264 , \24263 );
not \U$24019 ( \24265 , \3344 );
or \U$24020 ( \24266 , \24264 , \24265 );
nand \U$24021 ( \24267 , \7483 , \24036 );
nand \U$24022 ( \24268 , \24266 , \24267 );
not \U$24023 ( \24269 , \24268 );
xor \U$24024 ( \24270 , RIbe28390_19, RIbe2a730_95);
not \U$24025 ( \24271 , \24270 );
not \U$24026 ( \24272 , \8651 );
or \U$24027 ( \24273 , \24271 , \24272 );
nand \U$24028 ( \24274 , \8654 , \23930 );
nand \U$24029 ( \24275 , \24273 , \24274 );
not \U$24030 ( \24276 , \24275 );
or \U$24031 ( \24277 , \24269 , \24276 );
or \U$24032 ( \24278 , \24275 , \24268 );
xor \U$24033 ( \24279 , RIbe29e48_76, RIbe2a0a0_81);
not \U$24034 ( \24280 , \24279 );
not \U$24035 ( \24281 , \4843 );
or \U$24036 ( \24282 , \24280 , \24281 );
nand \U$24037 ( \24283 , \7368 , \23919 );
nand \U$24038 ( \24284 , \24282 , \24283 );
nand \U$24039 ( \24285 , \24278 , \24284 );
nand \U$24040 ( \24286 , \24277 , \24285 );
not \U$24041 ( \24287 , \24286 );
xor \U$24042 ( \24288 , RIbe295d8_58, RIbe2aaf0_103);
not \U$24043 ( \24289 , \24288 );
not \U$24044 ( \24290 , \20574 );
or \U$24045 ( \24291 , \24289 , \24290 );
nand \U$24046 ( \24292 , \23924 , RIbe2ab68_104);
nand \U$24047 ( \24293 , \24291 , \24292 );
xor \U$24048 ( \24294 , RIbe2a550_91, RIbe29ce0_73);
not \U$24049 ( \24295 , \24294 );
not \U$24050 ( \24296 , \12000 );
or \U$24051 ( \24297 , \24295 , \24296 );
nand \U$24052 ( \24298 , \15995 , \23998 );
nand \U$24053 ( \24299 , \24297 , \24298 );
xor \U$24054 ( \24300 , \24293 , \24299 );
xor \U$24055 ( \24301 , RIbe2a460_89, RIbe28f48_44);
not \U$24056 ( \24302 , \24301 );
not \U$24057 ( \24303 , \11461 );
or \U$24058 ( \24304 , \24302 , \24303 );
nand \U$24059 ( \24305 , \11201 , \24011 );
nand \U$24060 ( \24306 , \24304 , \24305 );
and \U$24061 ( \24307 , \24300 , \24306 );
and \U$24062 ( \24308 , \24293 , \24299 );
or \U$24063 ( \24309 , \24307 , \24308 );
not \U$24064 ( \24310 , \24309 );
not \U$24065 ( \24311 , \24310 );
xor \U$24066 ( \24312 , RIbe2ae38_110, RIbe28a20_33);
not \U$24067 ( \24313 , \24312 );
not \U$24068 ( \24314 , \9194 );
or \U$24069 ( \24315 , \24313 , \24314 );
nand \U$24070 ( \24316 , \2475 , \24042 );
nand \U$24071 ( \24317 , \24315 , \24316 );
not \U$24072 ( \24318 , \24317 );
not \U$24073 ( \24319 , \24318 );
xor \U$24074 ( \24320 , RIbe298a8_64, RIbe2a280_85);
not \U$24075 ( \24321 , \24320 );
not \U$24076 ( \24322 , \14942 );
or \U$24077 ( \24323 , \24321 , \24322 );
nand \U$24078 ( \24324 , \11348 , \24030 );
nand \U$24079 ( \24325 , \24323 , \24324 );
not \U$24080 ( \24326 , \24325 );
not \U$24081 ( \24327 , \24326 );
or \U$24082 ( \24328 , \24319 , \24327 );
xor \U$24083 ( \24329 , RIbe29ec0_77, RIbe2a910_99);
not \U$24084 ( \24330 , \24329 );
not \U$24085 ( \24331 , \13325 );
or \U$24086 ( \24332 , \24330 , \24331 );
nand \U$24087 ( \24333 , \11456 , \24133 );
nand \U$24088 ( \24334 , \24332 , \24333 );
nand \U$24089 ( \24335 , \24328 , \24334 );
nand \U$24090 ( \24336 , \24325 , \24317 );
nand \U$24091 ( \24337 , \24335 , \24336 );
not \U$24092 ( \24338 , \24337 );
or \U$24093 ( \24339 , \24311 , \24338 );
or \U$24094 ( \24340 , \24310 , \24337 );
nand \U$24095 ( \24341 , \24339 , \24340 );
not \U$24096 ( \24342 , \24341 );
or \U$24097 ( \24343 , \24287 , \24342 );
nand \U$24098 ( \24344 , \24337 , \24309 );
nand \U$24099 ( \24345 , \24343 , \24344 );
and \U$24100 ( \24346 , \24262 , \24345 );
nor \U$24101 ( \24347 , \24181 , \24261 );
nor \U$24102 ( \24348 , \24346 , \24347 );
not \U$24103 ( \24349 , \24348 );
not \U$24104 ( \24350 , \24349 );
or \U$24105 ( \24351 , \24179 , \24350 );
not \U$24106 ( \24352 , \24348 );
not \U$24107 ( \24353 , \24177 );
or \U$24108 ( \24354 , \24352 , \24353 );
xor \U$24109 ( \24355 , \23995 , \24026 );
xor \U$24110 ( \24356 , \24355 , \24052 );
not \U$24111 ( \24357 , \24356 );
xor \U$24112 ( \24358 , RIbe285e8_24, RIbe2a640_93);
not \U$24113 ( \24359 , \24358 );
not \U$24114 ( \24360 , \7618 );
or \U$24115 ( \24361 , \24359 , \24360 );
nand \U$24116 ( \24362 , \8270 , \24104 );
nand \U$24117 ( \24363 , \24361 , \24362 );
not \U$24118 ( \24364 , \24363 );
not \U$24119 ( \24365 , \24364 );
xor \U$24120 ( \24366 , RIbe29128_48, RIbe2b018_114);
not \U$24121 ( \24367 , \24366 );
not \U$24122 ( \24368 , \20395 );
or \U$24123 ( \24369 , \24367 , \24368 );
nand \U$24124 ( \24370 , \15953 , \24097 );
nand \U$24125 ( \24371 , \24369 , \24370 );
not \U$24126 ( \24372 , \24371 );
not \U$24127 ( \24373 , \24372 );
or \U$24128 ( \24374 , \24365 , \24373 );
xor \U$24129 ( \24375 , RIbe2a028_80, RIbe2a820_97);
not \U$24130 ( \24376 , \24375 );
not \U$24131 ( \24377 , \8169 );
or \U$24132 ( \24378 , \24376 , \24377 );
nand \U$24133 ( \24379 , \8172 , \24005 );
nand \U$24134 ( \24380 , \24378 , \24379 );
nand \U$24135 ( \24381 , \24374 , \24380 );
not \U$24136 ( \24382 , \24372 );
nand \U$24137 ( \24383 , \24382 , \24363 );
nand \U$24138 ( \24384 , \24381 , \24383 );
not \U$24139 ( \24385 , \24384 );
not \U$24140 ( \24386 , \24385 );
xor \U$24141 ( \24387 , \24131 , \24130 );
xnor \U$24142 ( \24388 , \24387 , \24138 );
not \U$24143 ( \24389 , \24388 );
or \U$24144 ( \24390 , \24386 , \24389 );
not \U$24145 ( \24391 , \24033 );
not \U$24146 ( \24392 , \24048 );
or \U$24147 ( \24393 , \24391 , \24392 );
or \U$24148 ( \24394 , \24048 , \24033 );
nand \U$24149 ( \24395 , \24393 , \24394 );
nand \U$24150 ( \24396 , \24390 , \24395 );
not \U$24151 ( \24397 , \24388 );
nand \U$24152 ( \24398 , \24397 , \24384 );
nand \U$24153 ( \24399 , \24396 , \24398 );
not \U$24154 ( \24400 , \24102 );
and \U$24155 ( \24401 , \24121 , \24400 );
not \U$24156 ( \24402 , \24121 );
and \U$24157 ( \24403 , \24402 , \24102 );
nor \U$24158 ( \24404 , \24401 , \24403 );
not \U$24159 ( \24405 , \24404 );
not \U$24160 ( \24406 , \23701 );
nand \U$24161 ( \24407 , \24406 , \23705 );
not \U$24162 ( \24408 , \24407 );
not \U$24163 ( \24409 , \23687 );
and \U$24164 ( \24410 , \24408 , \24409 );
and \U$24165 ( \24411 , \24407 , \23687 );
nor \U$24166 ( \24412 , \24410 , \24411 );
not \U$24167 ( \24413 , \24412 );
or \U$24168 ( \24414 , \24405 , \24413 );
xor \U$24169 ( \24415 , \24003 , \24021 );
nand \U$24170 ( \24416 , \24414 , \24415 );
not \U$24171 ( \24417 , \24412 );
not \U$24172 ( \24418 , \24404 );
nand \U$24173 ( \24419 , \24417 , \24418 );
nand \U$24174 ( \24420 , \24416 , \24419 );
and \U$24175 ( \24421 , \24399 , \24420 );
not \U$24176 ( \24422 , \24399 );
not \U$24177 ( \24423 , \24420 );
and \U$24178 ( \24424 , \24422 , \24423 );
nor \U$24179 ( \24425 , \24421 , \24424 );
not \U$24180 ( \24426 , \24425 );
or \U$24181 ( \24427 , \24357 , \24426 );
not \U$24182 ( \24428 , \24423 );
nand \U$24183 ( \24429 , \24428 , \24399 );
nand \U$24184 ( \24430 , \24427 , \24429 );
nand \U$24185 ( \24431 , \24354 , \24430 );
nand \U$24186 ( \24432 , \24351 , \24431 );
and \U$24187 ( \24433 , \24171 , \24432 );
not \U$24188 ( \24434 , \24171 );
not \U$24189 ( \24435 , \24432 );
and \U$24190 ( \24436 , \24434 , \24435 );
nor \U$24191 ( \24437 , \24433 , \24436 );
not \U$24192 ( \24438 , \24437 );
or \U$24193 ( \24439 , \24078 , \24438 );
nand \U$24194 ( \24440 , \24432 , \24171 );
nand \U$24195 ( \24441 , \24439 , \24440 );
not \U$24196 ( \24442 , \24441 );
or \U$24197 ( \24443 , \23870 , \24442 );
or \U$24198 ( \24444 , \23869 , \24441 );
nand \U$24199 ( \24445 , \24443 , \24444 );
not \U$24200 ( \24446 , \24445 );
or \U$24201 ( \24447 , \23470 , \24446 );
nand \U$24202 ( \24448 , \24441 , \23868 );
nand \U$24203 ( \24449 , \24447 , \24448 );
not \U$24204 ( \24450 , \15353 );
not \U$24205 ( \24451 , \24450 );
not \U$24206 ( \24452 , \22775 );
not \U$24207 ( \24453 , \24452 );
and \U$24208 ( \24454 , \24451 , \24453 );
xor \U$24209 ( \24455 , RIbe2b180_117, RIbe295d8_58);
not \U$24210 ( \24456 , \24455 );
nor \U$24211 ( \24457 , \24456 , \14846 );
nor \U$24212 ( \24458 , \24454 , \24457 );
nand \U$24213 ( \24459 , \22794 , \22788 );
or \U$24214 ( \24460 , \24458 , \24459 );
nand \U$24215 ( \24461 , \24459 , \24458 );
nand \U$24216 ( \24462 , \24460 , \24461 );
or \U$24217 ( \24463 , \23422 , \23416 );
nand \U$24218 ( \24464 , \24463 , \23429 );
nand \U$24219 ( \24465 , \23422 , \23416 );
nand \U$24220 ( \24466 , \24464 , \24465 );
not \U$24221 ( \24467 , \24466 );
and \U$24222 ( \24468 , \24462 , \24467 );
not \U$24223 ( \24469 , \24462 );
and \U$24224 ( \24470 , \24469 , \24466 );
nor \U$24225 ( \24471 , \24468 , \24470 );
not \U$24226 ( \24472 , \23558 );
not \U$24227 ( \24473 , \23608 );
or \U$24228 ( \24474 , \24472 , \24473 );
or \U$24229 ( \24475 , \23558 , \23608 );
nand \U$24230 ( \24476 , \24475 , \23580 );
nand \U$24231 ( \24477 , \24474 , \24476 );
xor \U$24232 ( \24478 , \24471 , \24477 );
xor \U$24233 ( \24479 , \23492 , \23513 );
and \U$24234 ( \24480 , \24479 , \23535 );
and \U$24235 ( \24481 , \23492 , \23513 );
or \U$24236 ( \24482 , \24480 , \24481 );
xor \U$24237 ( \24483 , \24478 , \24482 );
not \U$24238 ( \24484 , \24483 );
not \U$24239 ( \24485 , \23795 );
not \U$24240 ( \24486 , \23854 );
or \U$24241 ( \24487 , \24485 , \24486 );
not \U$24242 ( \24488 , \23796 );
not \U$24243 ( \24489 , \23855 );
or \U$24244 ( \24490 , \24488 , \24489 );
nand \U$24245 ( \24491 , \24490 , \23786 );
nand \U$24246 ( \24492 , \24487 , \24491 );
not \U$24247 ( \24493 , \24492 );
or \U$24248 ( \24494 , \24484 , \24493 );
or \U$24249 ( \24495 , \24492 , \24483 );
not \U$24250 ( \24496 , \23611 );
not \U$24251 ( \24497 , \23634 );
or \U$24252 ( \24498 , \24496 , \24497 );
nand \U$24253 ( \24499 , \24498 , \23613 );
nand \U$24254 ( \24500 , \24495 , \24499 );
nand \U$24255 ( \24501 , \24494 , \24500 );
not \U$24256 ( \24502 , \22719 );
not \U$24257 ( \24503 , \8887 );
or \U$24258 ( \24504 , \24502 , \24503 );
xor \U$24259 ( \24505 , RIbe28930_31, RIbe2a7a8_96);
nand \U$24260 ( \24506 , \1199 , \24505 );
nand \U$24261 ( \24507 , \24504 , \24506 );
not \U$24262 ( \24508 , \24507 );
not \U$24263 ( \24509 , \22805 );
not \U$24264 ( \24510 , \9192 );
or \U$24265 ( \24511 , \24509 , \24510 );
xor \U$24266 ( \24512 , RIbe28a20_33, RIbe2ac58_106);
nand \U$24267 ( \24513 , \1768 , \24512 );
nand \U$24268 ( \24514 , \24511 , \24513 );
not \U$24269 ( \24515 , \24514 );
not \U$24270 ( \24516 , \24515 );
or \U$24271 ( \24517 , \24508 , \24516 );
or \U$24272 ( \24518 , \24507 , \24515 );
nand \U$24273 ( \24519 , \24517 , \24518 );
not \U$24274 ( \24520 , \23262 );
not \U$24275 ( \24521 , \9825 );
or \U$24276 ( \24522 , \24520 , \24521 );
xor \U$24277 ( \24523 , RIbe2a118_82, RIbe27fd0_11);
nand \U$24278 ( \24524 , \4897 , \24523 );
nand \U$24279 ( \24525 , \24522 , \24524 );
xnor \U$24280 ( \24526 , \24519 , \24525 );
not \U$24281 ( \24527 , \22740 );
not \U$24282 ( \24528 , \8267 );
or \U$24283 ( \24529 , \24527 , \24528 );
xor \U$24284 ( \24530 , RIbe285e8_24, RIbe2a4d8_90);
nand \U$24285 ( \24531 , \8270 , \24530 );
nand \U$24286 ( \24532 , \24529 , \24531 );
not \U$24287 ( \24533 , \24532 );
not \U$24288 ( \24534 , \24533 );
not \U$24289 ( \24535 , \22712 );
not \U$24290 ( \24536 , \14826 );
or \U$24291 ( \24537 , \24535 , \24536 );
xor \U$24292 ( \24538 , RIbe2a2f8_86, RIbe29b78_70);
nand \U$24293 ( \24539 , \18963 , \24538 );
nand \U$24294 ( \24540 , \24537 , \24539 );
not \U$24295 ( \24541 , \24455 );
not \U$24296 ( \24542 , \17592 );
or \U$24297 ( \24543 , \24541 , \24542 );
xor \U$24298 ( \24544 , RIbe2b180_117, RIbe29740_61);
nand \U$24299 ( \24545 , \21759 , \24544 );
nand \U$24300 ( \24546 , \24543 , \24545 );
nor \U$24301 ( \24547 , \24540 , \24546 );
not \U$24302 ( \24548 , \24547 );
nand \U$24303 ( \24549 , \24546 , \24540 );
nand \U$24304 ( \24550 , \24548 , \24549 );
not \U$24305 ( \24551 , \24550 );
or \U$24306 ( \24552 , \24534 , \24551 );
or \U$24307 ( \24553 , \24550 , \24533 );
nand \U$24308 ( \24554 , \24552 , \24553 );
not \U$24309 ( \24555 , \22685 );
not \U$24310 ( \24556 , \18832 );
or \U$24311 ( \24557 , \24555 , \24556 );
xor \U$24312 ( \24558 , RIbe288b8_30, RIbe2aaf0_103);
nand \U$24313 ( \24559 , \24558 , RIbe2ab68_104);
nand \U$24314 ( \24560 , \24557 , \24559 );
not \U$24315 ( \24561 , \22852 );
not \U$24316 ( \24562 , \8168 );
or \U$24317 ( \24563 , \24561 , \24562 );
xor \U$24318 ( \24564 , RIbe29d58_74, RIbe2a028_80);
nand \U$24319 ( \24565 , \8930 , \24564 );
nand \U$24320 ( \24566 , \24563 , \24565 );
xor \U$24321 ( \24567 , \24560 , \24566 );
not \U$24322 ( \24568 , \22733 );
not \U$24323 ( \24569 , \3408 );
or \U$24324 ( \24570 , \24568 , \24569 );
xor \U$24325 ( \24571 , RIbe28390_19, RIbe2b540_125);
nand \U$24326 ( \24572 , \2777 , \24571 );
nand \U$24327 ( \24573 , \24570 , \24572 );
xnor \U$24328 ( \24574 , \24567 , \24573 );
nand \U$24329 ( \24575 , \24554 , \24574 );
not \U$24330 ( \24576 , \24554 );
not \U$24331 ( \24577 , \24574 );
nand \U$24332 ( \24578 , \24576 , \24577 );
nand \U$24333 ( \24579 , \24575 , \24578 );
xnor \U$24334 ( \24580 , \24526 , \24579 );
not \U$24335 ( \24581 , \24580 );
not \U$24336 ( \24582 , \23308 );
not \U$24337 ( \24583 , \15992 );
or \U$24338 ( \24584 , \24582 , \24583 );
xor \U$24339 ( \24585 , RIbe2a550_91, RIbe27c88_4);
nand \U$24340 ( \24586 , \15995 , \24585 );
nand \U$24341 ( \24587 , \24584 , \24586 );
not \U$24342 ( \24588 , \22821 );
not \U$24343 ( \24589 , \23097 );
or \U$24344 ( \24590 , \24588 , \24589 );
xor \U$24345 ( \24591 , RIbe28f48_44, RIbe2a898_98);
nand \U$24346 ( \24592 , \9523 , \24591 );
nand \U$24347 ( \24593 , \24590 , \24592 );
not \U$24348 ( \24594 , \24593 );
not \U$24349 ( \24595 , \24594 );
not \U$24350 ( \24596 , \22816 );
not \U$24351 ( \24597 , \14423 );
or \U$24352 ( \24598 , \24596 , \24597 );
xor \U$24353 ( \24599 , RIbe28138_14, RIbe2af28_112);
nand \U$24354 ( \24600 , \14413 , \24599 );
nand \U$24355 ( \24601 , \24598 , \24600 );
not \U$24356 ( \24602 , \24601 );
or \U$24357 ( \24603 , \24595 , \24602 );
or \U$24358 ( \24604 , \24601 , \24594 );
nand \U$24359 ( \24605 , \24603 , \24604 );
xnor \U$24360 ( \24606 , \24587 , \24605 );
not \U$24361 ( \24607 , \24606 );
not \U$24362 ( \24608 , \23297 );
not \U$24363 ( \24609 , \4842 );
or \U$24364 ( \24610 , \24608 , \24609 );
xor \U$24365 ( \24611 , RIbe29e48_76, RIbe29f38_78);
nand \U$24366 ( \24612 , \16655 , \24611 );
nand \U$24367 ( \24613 , \24610 , \24612 );
not \U$24368 ( \24614 , \22836 );
not \U$24369 ( \24615 , \2458 );
or \U$24370 ( \24616 , \24614 , \24615 );
xor \U$24371 ( \24617 , RIbe2b360_121, RIbe27e68_8);
nand \U$24372 ( \24618 , \2464 , \24617 );
nand \U$24373 ( \24619 , \24616 , \24618 );
xor \U$24374 ( \24620 , \24613 , \24619 );
not \U$24375 ( \24621 , \22701 );
not \U$24376 ( \24622 , \5024 );
or \U$24377 ( \24623 , \24621 , \24622 );
xor \U$24378 ( \24624 , RIbe2aa78_102, RIbe29c68_72);
nand \U$24379 ( \24625 , \4580 , \24624 );
nand \U$24380 ( \24626 , \24623 , \24625 );
xor \U$24381 ( \24627 , \24620 , \24626 );
not \U$24382 ( \24628 , \24627 );
or \U$24383 ( \24629 , \24607 , \24628 );
or \U$24384 ( \24630 , \24627 , \24606 );
nand \U$24385 ( \24631 , \24629 , \24630 );
xor \U$24386 ( \24632 , \23191 , \23215 );
and \U$24387 ( \24633 , \24632 , \23247 );
and \U$24388 ( \24634 , \23191 , \23215 );
or \U$24389 ( \24635 , \24633 , \24634 );
xor \U$24390 ( \24636 , \24631 , \24635 );
not \U$24391 ( \24637 , \24636 );
or \U$24392 ( \24638 , \24581 , \24637 );
or \U$24393 ( \24639 , \24636 , \24580 );
nand \U$24394 ( \24640 , \24638 , \24639 );
buf \U$24395 ( \24641 , \24640 );
xor \U$24396 ( \24642 , \24471 , \24477 );
and \U$24397 ( \24643 , \24642 , \24482 );
and \U$24398 ( \24644 , \24471 , \24477 );
or \U$24399 ( \24645 , \24643 , \24644 );
buf \U$24400 ( \24646 , \24645 );
and \U$24401 ( \24647 , \24641 , \24646 );
not \U$24402 ( \24648 , \24641 );
not \U$24403 ( \24649 , \24646 );
and \U$24404 ( \24650 , \24648 , \24649 );
nor \U$24405 ( \24651 , \24647 , \24650 );
and \U$24406 ( \24652 , \24501 , \24651 );
not \U$24407 ( \24653 , \24501 );
not \U$24408 ( \24654 , \24651 );
and \U$24409 ( \24655 , \24653 , \24654 );
nor \U$24410 ( \24656 , \24652 , \24655 );
buf \U$24411 ( \24657 , \24656 );
not \U$24412 ( \24658 , \24461 );
not \U$24413 ( \24659 , \24466 );
or \U$24414 ( \24660 , \24658 , \24659 );
nand \U$24415 ( \24661 , \24660 , \24460 );
not \U$24416 ( \24662 , \24661 );
and \U$24417 ( \24663 , \23136 , \23160 );
and \U$24418 ( \24664 , \23132 , \23103 );
nor \U$24419 ( \24665 , \24663 , \24664 );
not \U$24420 ( \24666 , \24665 );
or \U$24421 ( \24667 , \24662 , \24666 );
or \U$24422 ( \24668 , \24665 , \24661 );
nand \U$24423 ( \24669 , \24667 , \24668 );
not \U$24424 ( \24670 , \24669 );
not \U$24425 ( \24671 , \23286 );
not \U$24426 ( \24672 , \23292 );
or \U$24427 ( \24673 , \24671 , \24672 );
or \U$24428 ( \24674 , \23286 , \23292 );
nand \U$24429 ( \24675 , \24674 , \23299 );
nand \U$24430 ( \24676 , \24673 , \24675 );
or \U$24431 ( \24677 , \23274 , \23265 );
nand \U$24432 ( \24678 , \24677 , \23267 );
xor \U$24433 ( \24679 , \24676 , \24678 );
not \U$24434 ( \24680 , \22742 );
not \U$24435 ( \24681 , \22750 );
or \U$24436 ( \24682 , \24680 , \24681 );
or \U$24437 ( \24683 , \22750 , \22742 );
nand \U$24438 ( \24684 , \24683 , \22735 );
nand \U$24439 ( \24685 , \24682 , \24684 );
not \U$24440 ( \24686 , \24685 );
and \U$24441 ( \24687 , \24679 , \24686 );
not \U$24442 ( \24688 , \24679 );
and \U$24443 ( \24689 , \24688 , \24685 );
nor \U$24444 ( \24690 , \24687 , \24689 );
not \U$24445 ( \24691 , \24690 );
and \U$24446 ( \24692 , \24670 , \24691 );
and \U$24447 ( \24693 , \24669 , \24690 );
nor \U$24448 ( \24694 , \24692 , \24693 );
xor \U$24449 ( \24695 , \23405 , \23443 );
and \U$24450 ( \24696 , \24695 , \23463 );
and \U$24451 ( \24697 , \23405 , \23443 );
or \U$24452 ( \24698 , \24696 , \24697 );
not \U$24453 ( \24699 , \24698 );
and \U$24454 ( \24700 , \24694 , \24699 );
not \U$24455 ( \24701 , \24694 );
and \U$24456 ( \24702 , \24701 , \24698 );
nor \U$24457 ( \24703 , \24700 , \24702 );
buf \U$24458 ( \24704 , \24703 );
not \U$24459 ( \24705 , \23322 );
not \U$24460 ( \24706 , \23319 );
or \U$24461 ( \24707 , \24705 , \24706 );
nand \U$24462 ( \24708 , \24707 , \23330 );
nand \U$24463 ( \24709 , \23318 , \23311 );
nand \U$24464 ( \24710 , \24708 , \24709 );
not \U$24465 ( \24711 , \23328 );
not \U$24466 ( \24712 , \3056 );
or \U$24467 ( \24713 , \24711 , \24712 );
xor \U$24468 ( \24714 , RIbe28228_16, RIbe2b450_123);
nand \U$24469 ( \24715 , \885 , \24714 );
nand \U$24470 ( \24716 , \24713 , \24715 );
or \U$24471 ( \24717 , RIbe281b0_15, RIbe28228_16);
nand \U$24472 ( \24718 , \24717 , RIbe2ae38_110);
nand \U$24473 ( \24719 , RIbe281b0_15, RIbe28228_16);
and \U$24474 ( \24720 , \24718 , \24719 , RIbe280c0_13);
or \U$24475 ( \24721 , \24716 , \24720 );
nand \U$24476 ( \24722 , \24716 , \24720 );
nand \U$24477 ( \24723 , \24721 , \24722 );
not \U$24478 ( \24724 , \24723 );
nor \U$24479 ( \24725 , \24710 , \24724 );
not \U$24480 ( \24726 , \24725 );
nand \U$24481 ( \24727 , \24710 , \24724 );
nand \U$24482 ( \24728 , \24726 , \24727 );
not \U$24483 ( \24729 , \24728 );
xor \U$24484 ( \24730 , \22807 , \22819 );
and \U$24485 ( \24731 , \24730 , \22826 );
and \U$24486 ( \24732 , \22807 , \22819 );
or \U$24487 ( \24733 , \24731 , \24732 );
not \U$24488 ( \24734 , \24733 );
not \U$24489 ( \24735 , \24734 );
and \U$24490 ( \24736 , \24729 , \24735 );
and \U$24491 ( \24737 , \24728 , \24734 );
nor \U$24492 ( \24738 , \24736 , \24737 );
not \U$24493 ( \24739 , \24738 );
not \U$24494 ( \24740 , \24739 );
not \U$24495 ( \24741 , \23331 );
not \U$24496 ( \24742 , \23279 );
or \U$24497 ( \24743 , \24741 , \24742 );
nand \U$24498 ( \24744 , \24743 , \23300 );
not \U$24499 ( \24745 , \23279 );
nand \U$24500 ( \24746 , \24745 , \23332 );
nand \U$24501 ( \24747 , \24744 , \24746 );
not \U$24502 ( \24748 , \24747 );
not \U$24503 ( \24749 , \24748 );
or \U$24504 ( \24750 , \24740 , \24749 );
nand \U$24505 ( \24751 , \24738 , \24747 );
nand \U$24506 ( \24752 , \24750 , \24751 );
not \U$24507 ( \24753 , \22723 );
not \U$24508 ( \24754 , \22758 );
or \U$24509 ( \24755 , \24753 , \24754 );
not \U$24510 ( \24756 , \22755 );
not \U$24511 ( \24757 , \22724 );
or \U$24512 ( \24758 , \24756 , \24757 );
nand \U$24513 ( \24759 , \24758 , \22705 );
nand \U$24514 ( \24760 , \24755 , \24759 );
and \U$24515 ( \24761 , \24752 , \24760 );
not \U$24516 ( \24762 , \24752 );
not \U$24517 ( \24763 , \24760 );
and \U$24518 ( \24764 , \24762 , \24763 );
nor \U$24519 ( \24765 , \24761 , \24764 );
and \U$24520 ( \24766 , \24704 , \24765 );
not \U$24521 ( \24767 , \24704 );
not \U$24522 ( \24768 , \24765 );
and \U$24523 ( \24769 , \24767 , \24768 );
nor \U$24524 ( \24770 , \24766 , \24769 );
and \U$24525 ( \24771 , \24657 , \24770 );
not \U$24526 ( \24772 , \24657 );
not \U$24527 ( \24773 , \24770 );
and \U$24528 ( \24774 , \24772 , \24773 );
nor \U$24529 ( \24775 , \24771 , \24774 );
xor \U$24530 ( \24776 , \24449 , \24775 );
not \U$24531 ( \24777 , \24776 );
and \U$24532 ( \24778 , \24492 , \24483 );
not \U$24533 ( \24779 , \24492 );
not \U$24534 ( \24780 , \24483 );
and \U$24535 ( \24781 , \24779 , \24780 );
nor \U$24536 ( \24782 , \24778 , \24781 );
not \U$24537 ( \24783 , \24499 );
and \U$24538 ( \24784 , \24782 , \24783 );
not \U$24539 ( \24785 , \24782 );
and \U$24540 ( \24786 , \24785 , \24499 );
nor \U$24541 ( \24787 , \24784 , \24786 );
not \U$24542 ( \24788 , \24787 );
not \U$24543 ( \24789 , \24788 );
not \U$24544 ( \24790 , \23872 );
not \U$24545 ( \24791 , \23884 );
or \U$24546 ( \24792 , \24790 , \24791 );
or \U$24547 ( \24793 , \23884 , \23872 );
nand \U$24548 ( \24794 , \24793 , \23890 );
nand \U$24549 ( \24795 , \24792 , \24794 );
not \U$24550 ( \24796 , \24795 );
xnor \U$24551 ( \24797 , \23067 , \22952 );
not \U$24552 ( \24798 , \24797 );
not \U$24553 ( \24799 , \24067 );
not \U$24554 ( \24800 , \24056 );
or \U$24555 ( \24801 , \24799 , \24800 );
nand \U$24556 ( \24802 , \24801 , \24070 );
nand \U$24557 ( \24803 , \24055 , \24064 );
nand \U$24558 ( \24804 , \24802 , \24803 );
not \U$24559 ( \24805 , \24804 );
or \U$24560 ( \24806 , \24798 , \24805 );
or \U$24561 ( \24807 , \24797 , \24804 );
nand \U$24562 ( \24808 , \24806 , \24807 );
not \U$24563 ( \24809 , \24808 );
or \U$24564 ( \24810 , \24796 , \24809 );
not \U$24565 ( \24811 , \24797 );
nand \U$24566 ( \24812 , \24811 , \24804 );
nand \U$24567 ( \24813 , \24810 , \24812 );
not \U$24568 ( \24814 , \24813 );
not \U$24569 ( \24815 , \24157 );
not \U$24570 ( \24816 , \24170 );
or \U$24571 ( \24817 , \24815 , \24816 );
not \U$24572 ( \24818 , \24166 );
nand \U$24573 ( \24819 , \24818 , \24163 );
nand \U$24574 ( \24820 , \24817 , \24819 );
not \U$24575 ( \24821 , \24820 );
and \U$24576 ( \24822 , \24814 , \24821 );
not \U$24577 ( \24823 , \24814 );
and \U$24578 ( \24824 , \24823 , \24820 );
nor \U$24579 ( \24825 , \24822 , \24824 );
not \U$24580 ( \24826 , \24825 );
or \U$24581 ( \24827 , \24789 , \24826 );
not \U$24582 ( \24828 , \24814 );
nand \U$24583 ( \24829 , \24828 , \24820 );
nand \U$24584 ( \24830 , \24827 , \24829 );
not \U$24585 ( \24831 , \24830 );
not \U$24586 ( \24832 , \22862 );
not \U$24587 ( \24833 , \23072 );
or \U$24588 ( \24834 , \24832 , \24833 );
nand \U$24589 ( \24835 , \24834 , \22861 );
not \U$24590 ( \24836 , \24835 );
not \U$24591 ( \24837 , \23336 );
not \U$24592 ( \24838 , \23252 );
or \U$24593 ( \24839 , \24837 , \24838 );
not \U$24594 ( \24840 , \23165 );
nand \U$24595 ( \24841 , \24840 , \23248 );
nand \U$24596 ( \24842 , \24839 , \24841 );
not \U$24597 ( \24843 , \24842 );
not \U$24598 ( \24844 , \24843 );
or \U$24599 ( \24845 , \24836 , \24844 );
or \U$24600 ( \24846 , \24835 , \24843 );
nand \U$24601 ( \24847 , \24845 , \24846 );
buf \U$24602 ( \24848 , \24847 );
not \U$24603 ( \24849 , \22748 );
not \U$24604 ( \24850 , \2518 );
or \U$24605 ( \24851 , \24849 , \24850 );
xor \U$24606 ( \24852 , RIbe28480_21, RIbe2adc0_109);
nand \U$24607 ( \24853 , \7483 , \24852 );
nand \U$24608 ( \24854 , \24851 , \24853 );
not \U$24609 ( \24855 , \23316 );
not \U$24610 ( \24856 , \3401 );
or \U$24611 ( \24857 , \24855 , \24856 );
xor \U$24612 ( \24858 , RIbe28b88_36, RIbe2a6b8_94);
nand \U$24613 ( \24859 , \7550 , \24858 );
nand \U$24614 ( \24860 , \24857 , \24859 );
xor \U$24615 ( \24861 , \24854 , \24860 );
not \U$24616 ( \24862 , \22692 );
not \U$24617 ( \24863 , \15690 );
or \U$24618 ( \24864 , \24862 , \24863 );
xor \U$24619 ( \24865 , RIbe29218_50, RIbe2a190_83);
nand \U$24620 ( \24866 , \15693 , \24865 );
nand \U$24621 ( \24867 , \24864 , \24866 );
xnor \U$24622 ( \24868 , \24861 , \24867 );
and \U$24623 ( \24869 , RIbe280c0_13, RIbe2ae38_110);
not \U$24624 ( \24870 , RIbe280c0_13);
not \U$24625 ( \24871 , RIbe2ae38_110);
and \U$24626 ( \24872 , \24870 , \24871 );
nor \U$24627 ( \24873 , \24869 , \24872 );
not \U$24628 ( \24874 , \24873 );
not \U$24629 ( \24875 , \862 );
or \U$24630 ( \24876 , \24874 , \24875 );
xor \U$24631 ( \24877 , RIbe280c0_13, RIbe2aeb0_111);
nand \U$24632 ( \24878 , \2369 , \24877 );
nand \U$24633 ( \24879 , \24876 , \24878 );
not \U$24634 ( \24880 , \24879 );
not \U$24635 ( \24881 , \23256 );
not \U$24636 ( \24882 , \9737 );
or \U$24637 ( \24883 , \24881 , \24882 );
xor \U$24638 ( \24884 , RIbe2a910_99, RIbe29998_66);
nand \U$24639 ( \24885 , \10401 , \24884 );
nand \U$24640 ( \24886 , \24883 , \24885 );
not \U$24641 ( \24887 , \24886 );
not \U$24642 ( \24888 , \23284 );
not \U$24643 ( \24889 , \21852 );
or \U$24644 ( \24890 , \24888 , \24889 );
xor \U$24645 ( \24891 , RIbe291a0_49, RIbe2b108_116);
nand \U$24646 ( \24892 , \23015 , \24891 );
nand \U$24647 ( \24893 , \24890 , \24892 );
not \U$24648 ( \24894 , \24893 );
not \U$24649 ( \24895 , \24894 );
or \U$24650 ( \24896 , \24887 , \24895 );
or \U$24651 ( \24897 , \24886 , \24894 );
nand \U$24652 ( \24898 , \24896 , \24897 );
not \U$24653 ( \24899 , \24898 );
not \U$24654 ( \24900 , \24899 );
or \U$24655 ( \24901 , \24880 , \24900 );
not \U$24656 ( \24902 , \24879 );
nand \U$24657 ( \24903 , \24902 , \24898 );
nand \U$24658 ( \24904 , \24901 , \24903 );
not \U$24659 ( \24905 , \23272 );
not \U$24660 ( \24906 , \16811 );
or \U$24661 ( \24907 , \24905 , \24906 );
xor \U$24662 ( \24908 , RIbe29470_55, RIbe2b018_114);
nand \U$24663 ( \24909 , \18777 , \24908 );
nand \U$24664 ( \24910 , \24907 , \24909 );
not \U$24665 ( \24911 , \24910 );
not \U$24666 ( \24912 , \22843 );
not \U$24667 ( \24913 , \9262 );
or \U$24668 ( \24914 , \24912 , \24913 );
xor \U$24669 ( \24915 , RIbe28cf0_39, RIbe2a3e8_88);
nand \U$24670 ( \24916 , \8794 , \24915 );
nand \U$24671 ( \24917 , \24914 , \24916 );
not \U$24672 ( \24918 , \24917 );
and \U$24673 ( \24919 , \24911 , \24918 );
not \U$24674 ( \24920 , \24911 );
and \U$24675 ( \24921 , \24920 , \24917 );
nor \U$24676 ( \24922 , \24919 , \24921 );
not \U$24677 ( \24923 , \23290 );
not \U$24678 ( \24924 , \15793 );
or \U$24679 ( \24925 , \24923 , \24924 );
xor \U$24680 ( \24926 , RIbe29b00_69, RIbe2a280_85);
nand \U$24681 ( \24927 , \11348 , \24926 );
nand \U$24682 ( \24928 , \24925 , \24927 );
xor \U$24683 ( \24929 , \24922 , \24928 );
nor \U$24684 ( \24930 , \24904 , \24929 );
not \U$24685 ( \24931 , \24930 );
nand \U$24686 ( \24932 , \24904 , \24929 );
nand \U$24687 ( \24933 , \24931 , \24932 );
xor \U$24688 ( \24934 , \24868 , \24933 );
not \U$24689 ( \24935 , \22855 );
not \U$24690 ( \24936 , \22831 );
or \U$24691 ( \24937 , \24935 , \24936 );
not \U$24692 ( \24938 , \22827 );
nand \U$24693 ( \24939 , \24938 , \22797 );
nand \U$24694 ( \24940 , \24937 , \24939 );
or \U$24695 ( \24941 , \22694 , \22687 );
not \U$24696 ( \24942 , \24941 );
not \U$24697 ( \24943 , \22703 );
or \U$24698 ( \24944 , \24942 , \24943 );
nand \U$24699 ( \24945 , \22694 , \22687 );
nand \U$24700 ( \24946 , \24944 , \24945 );
not \U$24701 ( \24947 , \24946 );
xor \U$24702 ( \24948 , \22707 , \22714 );
and \U$24703 ( \24949 , \24948 , \22722 );
and \U$24704 ( \24950 , \22707 , \22714 );
or \U$24705 ( \24951 , \24949 , \24950 );
xor \U$24706 ( \24952 , \24947 , \24951 );
or \U$24707 ( \24953 , \22845 , \22838 );
nand \U$24708 ( \24954 , \24953 , \22854 );
nand \U$24709 ( \24955 , \22838 , \22845 );
and \U$24710 ( \24956 , \24954 , \24955 );
not \U$24711 ( \24957 , \24956 );
buf \U$24712 ( \24958 , \24957 );
xor \U$24713 ( \24959 , \24952 , \24958 );
and \U$24714 ( \24960 , \24940 , \24959 );
not \U$24715 ( \24961 , \24940 );
not \U$24716 ( \24962 , \24959 );
and \U$24717 ( \24963 , \24961 , \24962 );
or \U$24718 ( \24964 , \24960 , \24963 );
xor \U$24719 ( \24965 , \24934 , \24964 );
and \U$24720 ( \24966 , \24848 , \24965 );
not \U$24721 ( \24967 , \24848 );
not \U$24722 ( \24968 , \24965 );
and \U$24723 ( \24969 , \24967 , \24968 );
nor \U$24724 ( \24970 , \24966 , \24969 );
not \U$24725 ( \24971 , \24970 );
not \U$24726 ( \24972 , \23468 );
not \U$24727 ( \24973 , \23077 );
or \U$24728 ( \24974 , \24972 , \24973 );
not \U$24729 ( \24975 , \23337 );
nand \U$24730 ( \24976 , \24975 , \23464 );
nand \U$24731 ( \24977 , \24974 , \24976 );
not \U$24732 ( \24978 , \24977 );
not \U$24733 ( \24979 , \24978 );
and \U$24734 ( \24980 , \24971 , \24979 );
and \U$24735 ( \24981 , \24978 , \24970 );
nor \U$24736 ( \24982 , \24980 , \24981 );
not \U$24737 ( \24983 , \24982 );
and \U$24738 ( \24984 , \24831 , \24983 );
and \U$24739 ( \24985 , \24830 , \24982 );
nor \U$24740 ( \24986 , \24984 , \24985 );
not \U$24741 ( \24987 , \24986 );
or \U$24742 ( \24988 , \24777 , \24987 );
or \U$24743 ( \24989 , \24776 , \24986 );
nand \U$24744 ( \24990 , \24988 , \24989 );
buf \U$24745 ( \24991 , \24445 );
not \U$24746 ( \24992 , \23469 );
and \U$24747 ( \24993 , \24991 , \24992 );
not \U$24748 ( \24994 , \24991 );
and \U$24749 ( \24995 , \24994 , \23469 );
nor \U$24750 ( \24996 , \24993 , \24995 );
not \U$24751 ( \24997 , \24996 );
not \U$24752 ( \24998 , \24997 );
and \U$24753 ( \24999 , \24345 , \24261 );
not \U$24754 ( \25000 , \24345 );
and \U$24755 ( \25001 , \25000 , \24260 );
nor \U$24756 ( \25002 , \24999 , \25001 );
xor \U$24757 ( \25003 , \24181 , \25002 );
not \U$24758 ( \25004 , \25003 );
xnor \U$24759 ( \25005 , \24341 , \24286 );
not \U$24760 ( \25006 , \25005 );
not \U$24761 ( \25007 , \25006 );
xor \U$24762 ( \25008 , RIbe2a2f8_86, RIbe2a898_98);
not \U$24763 ( \25009 , \25008 );
not \U$24764 ( \25010 , \8697 );
or \U$24765 ( \25011 , \25009 , \25010 );
nand \U$24766 ( \25012 , \8706 , \24195 );
nand \U$24767 ( \25013 , \25011 , \25012 );
not \U$24768 ( \25014 , \25013 );
xor \U$24769 ( \25015 , RIbe28480_21, RIbe2a7a8_96);
not \U$24770 ( \25016 , \25015 );
not \U$24771 ( \25017 , \16953 );
or \U$24772 ( \25018 , \25016 , \25017 );
nand \U$24773 ( \25019 , \16676 , \24263 );
nand \U$24774 ( \25020 , \25018 , \25019 );
xor \U$24775 ( \25021 , RIbe2a028_80, RIbe2a118_82);
not \U$24776 ( \25022 , \25021 );
not \U$24777 ( \25023 , \8400 );
or \U$24778 ( \25024 , \25022 , \25023 );
nand \U$24779 ( \25025 , \8930 , \24375 );
nand \U$24780 ( \25026 , \25024 , \25025 );
xor \U$24781 ( \25027 , \25020 , \25026 );
not \U$24782 ( \25028 , \25027 );
or \U$24783 ( \25029 , \25014 , \25028 );
nand \U$24784 ( \25030 , \25026 , \25020 );
nand \U$24785 ( \25031 , \25029 , \25030 );
not \U$24786 ( \25032 , \10689 );
not \U$24787 ( \25033 , \25032 );
xor \U$24788 ( \25034 , RIbe29b78_70, RIbe2a190_83);
not \U$24789 ( \25035 , \25034 );
or \U$24790 ( \25036 , \25033 , \25035 );
nand \U$24791 ( \25037 , \15693 , \24189 );
nand \U$24792 ( \25038 , \25036 , \25037 );
not \U$24793 ( \25039 , \25038 );
xor \U$24794 ( \25040 , RIbe2a6b8_94, RIbe27e68_8);
not \U$24795 ( \25041 , \25040 );
not \U$24796 ( \25042 , \2600 );
or \U$24797 ( \25043 , \25041 , \25042 );
nand \U$24798 ( \25044 , \2464 , \24248 );
nand \U$24799 ( \25045 , \25043 , \25044 );
not \U$24800 ( \25046 , \25045 );
or \U$24801 ( \25047 , \25039 , \25046 );
or \U$24802 ( \25048 , \25038 , \25045 );
xor \U$24803 ( \25049 , RIbe2a4d8_90, RIbe29c68_72);
not \U$24804 ( \25050 , \25049 );
not \U$24805 ( \25051 , \4578 );
or \U$24806 ( \25052 , \25050 , \25051 );
nand \U$24807 ( \25053 , \4580 , \24223 );
nand \U$24808 ( \25054 , \25052 , \25053 );
nand \U$24809 ( \25055 , \25048 , \25054 );
nand \U$24810 ( \25056 , \25047 , \25055 );
nor \U$24811 ( \25057 , \25031 , \25056 );
xor \U$24812 ( \25058 , RIbe2b108_116, RIbe29998_66);
not \U$24813 ( \25059 , \25058 );
not \U$24814 ( \25060 , \21852 );
or \U$24815 ( \25061 , \25059 , \25060 );
nand \U$24816 ( \25062 , \23015 , \24241 );
nand \U$24817 ( \25063 , \25061 , \25062 );
not \U$24818 ( \25064 , \25063 );
xor \U$24819 ( \25065 , RIbe285e8_24, RIbe2ac58_106);
not \U$24820 ( \25066 , \25065 );
not \U$24821 ( \25067 , \8813 );
or \U$24822 ( \25068 , \25066 , \25067 );
nand \U$24823 ( \25069 , \8270 , \24358 );
nand \U$24824 ( \25070 , \25068 , \25069 );
xor \U$24825 ( \25071 , RIbe28b88_36, RIbe2aeb0_111);
not \U$24826 ( \25072 , \25071 );
not \U$24827 ( \25073 , \8711 );
or \U$24828 ( \25074 , \25072 , \25073 );
nand \U$24829 ( \25075 , \13250 , \23729 );
nand \U$24830 ( \25076 , \25074 , \25075 );
and \U$24831 ( \25077 , \25070 , \25076 );
not \U$24832 ( \25078 , \25070 );
not \U$24833 ( \25079 , \25076 );
and \U$24834 ( \25080 , \25078 , \25079 );
nor \U$24835 ( \25081 , \25077 , \25080 );
not \U$24836 ( \25082 , \25081 );
or \U$24837 ( \25083 , \25064 , \25082 );
not \U$24838 ( \25084 , \25079 );
nand \U$24839 ( \25085 , \25084 , \25070 );
nand \U$24840 ( \25086 , \25083 , \25085 );
not \U$24841 ( \25087 , \25086 );
or \U$24842 ( \25088 , \25057 , \25087 );
nand \U$24843 ( \25089 , \25031 , \25056 );
nand \U$24844 ( \25090 , \25088 , \25089 );
not \U$24845 ( \25091 , \25090 );
or \U$24846 ( \25092 , \23732 , \23736 );
nand \U$24847 ( \25093 , \25092 , \23737 );
not \U$24848 ( \25094 , \25093 );
xor \U$24849 ( \25095 , RIbe2af28_112, RIbe29218_50);
not \U$24850 ( \25096 , \25095 );
not \U$24851 ( \25097 , \15345 );
or \U$24852 ( \25098 , \25096 , \25097 );
nand \U$24853 ( \25099 , \19721 , \24182 );
nand \U$24854 ( \25100 , \25098 , \25099 );
not \U$24855 ( \25101 , \25100 );
xor \U$24856 ( \25102 , RIbe27fd0_11, RIbe2b540_125);
not \U$24857 ( \25103 , \25102 );
not \U$24858 ( \25104 , \9082 );
or \U$24859 ( \25105 , \25103 , \25104 );
nand \U$24860 ( \25106 , \4897 , \24206 );
nand \U$24861 ( \25107 , \25105 , \25106 );
not \U$24862 ( \25108 , \25107 );
not \U$24863 ( \25109 , \25108 );
xor \U$24864 ( \25110 , RIbe2adc0_109, RIbe28f48_44);
not \U$24865 ( \25111 , \25110 );
not \U$24866 ( \25112 , \12721 );
or \U$24867 ( \25113 , \25111 , \25112 );
nand \U$24868 ( \25114 , \4180 , \24301 );
nand \U$24869 ( \25115 , \25113 , \25114 );
not \U$24870 ( \25116 , \25115 );
or \U$24871 ( \25117 , \25109 , \25116 );
or \U$24872 ( \25118 , \25115 , \25108 );
nand \U$24873 ( \25119 , \25117 , \25118 );
not \U$24874 ( \25120 , \25119 );
or \U$24875 ( \25121 , \25101 , \25120 );
nand \U$24876 ( \25122 , \25115 , \25107 );
nand \U$24877 ( \25123 , \25121 , \25122 );
not \U$24878 ( \25124 , \25123 );
not \U$24879 ( \25125 , \25124 );
or \U$24880 ( \25126 , \25094 , \25125 );
not \U$24881 ( \25127 , RIbe29b00_69);
not \U$24882 ( \25128 , RIbe2b018_114);
and \U$24883 ( \25129 , \25127 , \25128 );
and \U$24884 ( \25130 , RIbe29b00_69, RIbe2b018_114);
nor \U$24885 ( \25131 , \25129 , \25130 );
not \U$24886 ( \25132 , \25131 );
not \U$24887 ( \25133 , \17571 );
or \U$24888 ( \25134 , \25132 , \25133 );
nand \U$24889 ( \25135 , \20583 , \24366 );
nand \U$24890 ( \25136 , \25134 , \25135 );
not \U$24891 ( \25137 , \25136 );
xor \U$24892 ( \25138 , RIbe28cf0_39, RIbe2a280_85);
not \U$24893 ( \25139 , \25138 );
not \U$24894 ( \25140 , \14382 );
or \U$24895 ( \25141 , \25139 , \25140 );
nand \U$24896 ( \25142 , \18667 , \24320 );
nand \U$24897 ( \25143 , \25141 , \25142 );
xor \U$24898 ( \25144 , RIbe29e48_76, RIbe2b360_121);
not \U$24899 ( \25145 , \25144 );
not \U$24900 ( \25146 , \4842 );
or \U$24901 ( \25147 , \25145 , \25146 );
nand \U$24902 ( \25148 , \4850 , \24279 );
nand \U$24903 ( \25149 , \25147 , \25148 );
and \U$24904 ( \25150 , \25143 , \25149 );
not \U$24905 ( \25151 , \25143 );
not \U$24906 ( \25152 , \25149 );
and \U$24907 ( \25153 , \25151 , \25152 );
nor \U$24908 ( \25154 , \25150 , \25153 );
not \U$24909 ( \25155 , \25154 );
or \U$24910 ( \25156 , \25137 , \25155 );
nand \U$24911 ( \25157 , \25149 , \25143 );
nand \U$24912 ( \25158 , \25156 , \25157 );
nand \U$24913 ( \25159 , \25126 , \25158 );
not \U$24914 ( \25160 , \25093 );
nand \U$24915 ( \25161 , \25160 , \25123 );
and \U$24916 ( \25162 , \25159 , \25161 );
not \U$24917 ( \25163 , \25162 );
or \U$24918 ( \25164 , \25091 , \25163 );
or \U$24919 ( \25165 , \25090 , \25162 );
nand \U$24920 ( \25166 , \25164 , \25165 );
not \U$24921 ( \25167 , \25166 );
or \U$24922 ( \25168 , \25007 , \25167 );
not \U$24923 ( \25169 , \25162 );
nand \U$24924 ( \25170 , \25169 , \25090 );
nand \U$24925 ( \25171 , \25168 , \25170 );
xor \U$24926 ( \25172 , \23768 , \23707 );
xor \U$24927 ( \25173 , \25171 , \25172 );
not \U$24928 ( \25174 , \25173 );
or \U$24929 ( \25175 , \25004 , \25174 );
nand \U$24930 ( \25176 , \25171 , \25172 );
nand \U$24931 ( \25177 , \25175 , \25176 );
not \U$24932 ( \25178 , \25177 );
and \U$24933 ( \25179 , \23773 , \23667 );
not \U$24934 ( \25180 , \23773 );
and \U$24935 ( \25181 , \25180 , \23668 );
or \U$24936 ( \25182 , \25179 , \25181 );
and \U$24937 ( \25183 , \25182 , \23661 );
not \U$24938 ( \25184 , \25182 );
and \U$24939 ( \25185 , \25184 , \23660 );
nor \U$24940 ( \25186 , \25183 , \25185 );
xor \U$24941 ( \25187 , \24232 , \24256 );
xor \U$24942 ( \25188 , \25187 , \24204 );
not \U$24943 ( \25189 , \25188 );
not \U$24944 ( \25190 , \23913 );
not \U$24945 ( \25191 , \23974 );
or \U$24946 ( \25192 , \25190 , \25191 );
or \U$24947 ( \25193 , \23974 , \23913 );
nand \U$24948 ( \25194 , \25192 , \25193 );
not \U$24949 ( \25195 , \25194 );
or \U$24950 ( \25196 , \25189 , \25195 );
or \U$24951 ( \25197 , \25194 , \25188 );
not \U$24952 ( \25198 , \24385 );
not \U$24953 ( \25199 , \24388 );
or \U$24954 ( \25200 , \25198 , \25199 );
nand \U$24955 ( \25201 , \25200 , \24398 );
xnor \U$24956 ( \25202 , \25201 , \24395 );
nand \U$24957 ( \25203 , \25197 , \25202 );
nand \U$24958 ( \25204 , \25196 , \25203 );
not \U$24959 ( \25205 , \25204 );
xor \U$24960 ( \25206 , \24425 , \24356 );
not \U$24961 ( \25207 , \25206 );
or \U$24962 ( \25208 , \25205 , \25207 );
or \U$24963 ( \25209 , \25206 , \25204 );
xor \U$24964 ( \25210 , \24192 , \24187 );
xnor \U$24965 ( \25211 , \25210 , \24201 );
xor \U$24966 ( \25212 , \24211 , \24221 );
xor \U$24967 ( \25213 , \25212 , \24228 );
nor \U$24968 ( \25214 , \25211 , \25213 );
xor \U$24969 ( \25215 , \24275 , \24268 );
xnor \U$24970 ( \25216 , \25215 , \24284 );
or \U$24971 ( \25217 , \25214 , \25216 );
nand \U$24972 ( \25218 , \25211 , \25213 );
nand \U$24973 ( \25219 , \25217 , \25218 );
not \U$24974 ( \25220 , \25219 );
xor \U$24975 ( \25221 , RIbe2a550_91, RIbe29d58_74);
not \U$24976 ( \25222 , \25221 );
not \U$24977 ( \25223 , \18635 );
or \U$24978 ( \25224 , \25222 , \25223 );
nand \U$24979 ( \25225 , \14612 , \24294 );
nand \U$24980 ( \25226 , \25224 , \25225 );
not \U$24981 ( \25227 , \25226 );
xor \U$24982 ( \25228 , RIbe28390_19, RIbe2b450_123);
not \U$24983 ( \25229 , \25228 );
not \U$24984 ( \25230 , \14806 );
or \U$24985 ( \25231 , \25229 , \25230 );
nand \U$24986 ( \25232 , \2647 , \24270 );
nand \U$24987 ( \25233 , \25231 , \25232 );
nand \U$24988 ( \25234 , \5055 , RIbe2ae38_110);
and \U$24989 ( \25235 , \25233 , \25234 );
not \U$24990 ( \25236 , \25233 );
not \U$24991 ( \25237 , \25234 );
and \U$24992 ( \25238 , \25236 , \25237 );
or \U$24993 ( \25239 , \25235 , \25238 );
not \U$24994 ( \25240 , \25239 );
or \U$24995 ( \25241 , \25227 , \25240 );
nand \U$24996 ( \25242 , \25233 , \25237 );
nand \U$24997 ( \25243 , \25241 , \25242 );
and \U$24998 ( \25244 , \24371 , \24364 );
not \U$24999 ( \25245 , \24371 );
and \U$25000 ( \25246 , \25245 , \24363 );
or \U$25001 ( \25247 , \25244 , \25246 );
xor \U$25002 ( \25248 , \25247 , \24380 );
xor \U$25003 ( \25249 , \25243 , \25248 );
xor \U$25004 ( \25250 , RIbe27c88_4, RIbe2b180_117);
not \U$25005 ( \25251 , \25250 );
nor \U$25006 ( \25252 , \25251 , \14853 );
not \U$25007 ( \25253 , \24216 );
not \U$25008 ( \25254 , \16646 );
nor \U$25009 ( \25255 , \25253 , \25254 );
nor \U$25010 ( \25256 , \25252 , \25255 );
not \U$25011 ( \25257 , \25256 );
not \U$25012 ( \25258 , \25257 );
not \U$25013 ( \25259 , \19580 );
not \U$25014 ( \25260 , RIbe291a0_49);
not \U$25015 ( \25261 , RIbe2aaf0_103);
and \U$25016 ( \25262 , \25260 , \25261 );
and \U$25017 ( \25263 , RIbe291a0_49, RIbe2aaf0_103);
nor \U$25018 ( \25264 , \25262 , \25263 );
not \U$25019 ( \25265 , \25264 );
not \U$25020 ( \25266 , \25265 );
and \U$25021 ( \25267 , \25259 , \25266 );
and \U$25022 ( \25268 , \24288 , RIbe2ab68_104);
nor \U$25023 ( \25269 , \25267 , \25268 );
not \U$25024 ( \25270 , \25269 );
xor \U$25025 ( \25271 , RIbe2a910_99, RIbe29f38_78);
not \U$25026 ( \25272 , \25271 );
not \U$25027 ( \25273 , \9737 );
or \U$25028 ( \25274 , \25272 , \25273 );
nand \U$25029 ( \25275 , \9726 , \24329 );
nand \U$25030 ( \25276 , \25274 , \25275 );
not \U$25031 ( \25277 , \25276 );
or \U$25032 ( \25278 , \25270 , \25277 );
or \U$25033 ( \25279 , \25276 , \25269 );
nand \U$25034 ( \25280 , \25278 , \25279 );
not \U$25035 ( \25281 , \25280 );
or \U$25036 ( \25282 , \25258 , \25281 );
not \U$25037 ( \25283 , \25269 );
nand \U$25038 ( \25284 , \25283 , \25276 );
nand \U$25039 ( \25285 , \25282 , \25284 );
and \U$25040 ( \25286 , \25249 , \25285 );
and \U$25041 ( \25287 , \25243 , \25248 );
or \U$25042 ( \25288 , \25286 , \25287 );
xor \U$25043 ( \25289 , \24293 , \24299 );
xor \U$25044 ( \25290 , \25289 , \24306 );
not \U$25045 ( \25291 , \25290 );
not \U$25046 ( \25292 , \24325 );
not \U$25047 ( \25293 , \24318 );
or \U$25048 ( \25294 , \25292 , \25293 );
nand \U$25049 ( \25295 , \24326 , \24317 );
nand \U$25050 ( \25296 , \25294 , \25295 );
xor \U$25051 ( \25297 , \25296 , \24334 );
not \U$25052 ( \25298 , \25297 );
or \U$25053 ( \25299 , \25291 , \25298 );
or \U$25054 ( \25300 , \25297 , \25290 );
xor \U$25055 ( \25301 , \24240 , \24246 );
xor \U$25056 ( \25302 , \25301 , \24253 );
nand \U$25057 ( \25303 , \25300 , \25302 );
nand \U$25058 ( \25304 , \25299 , \25303 );
xor \U$25059 ( \25305 , \25288 , \25304 );
not \U$25060 ( \25306 , \25305 );
or \U$25061 ( \25307 , \25220 , \25306 );
nand \U$25062 ( \25308 , \25288 , \25304 );
nand \U$25063 ( \25309 , \25307 , \25308 );
nand \U$25064 ( \25310 , \25209 , \25309 );
nand \U$25065 ( \25311 , \25208 , \25310 );
xor \U$25066 ( \25312 , \25186 , \25311 );
not \U$25067 ( \25313 , \25312 );
or \U$25068 ( \25314 , \25178 , \25313 );
nand \U$25069 ( \25315 , \25311 , \25186 );
nand \U$25070 ( \25316 , \25314 , \25315 );
not \U$25071 ( \25317 , \25316 );
not \U$25072 ( \25318 , \24808 );
not \U$25073 ( \25319 , \24795 );
not \U$25074 ( \25320 , \25319 );
and \U$25075 ( \25321 , \25318 , \25320 );
and \U$25076 ( \25322 , \25319 , \24808 );
nor \U$25077 ( \25323 , \25321 , \25322 );
not \U$25078 ( \25324 , \25323 );
xor \U$25079 ( \25325 , \23635 , \23863 );
not \U$25080 ( \25326 , \25325 );
or \U$25081 ( \25327 , \25324 , \25326 );
or \U$25082 ( \25328 , \25325 , \25323 );
nand \U$25083 ( \25329 , \25327 , \25328 );
not \U$25084 ( \25330 , \25329 );
or \U$25085 ( \25331 , \25317 , \25330 );
not \U$25086 ( \25332 , \25323 );
nand \U$25087 ( \25333 , \25332 , \25325 );
nand \U$25088 ( \25334 , \25331 , \25333 );
not \U$25089 ( \25335 , \24787 );
not \U$25090 ( \25336 , \24825 );
and \U$25091 ( \25337 , \25335 , \25336 );
and \U$25092 ( \25338 , \24787 , \24825 );
nor \U$25093 ( \25339 , \25337 , \25338 );
not \U$25094 ( \25340 , \25339 );
and \U$25095 ( \25341 , \25334 , \25340 );
not \U$25096 ( \25342 , \25334 );
and \U$25097 ( \25343 , \25342 , \25339 );
nor \U$25098 ( \25344 , \25341 , \25343 );
not \U$25099 ( \25345 , \25344 );
or \U$25100 ( \25346 , \24998 , \25345 );
nand \U$25101 ( \25347 , \25334 , \25340 );
nand \U$25102 ( \25348 , \25346 , \25347 );
nand \U$25103 ( \25349 , \24990 , \25348 );
not \U$25104 ( \25350 , \24996 );
not \U$25105 ( \25351 , \25344 );
or \U$25106 ( \25352 , \25350 , \25351 );
or \U$25107 ( \25353 , \25344 , \24996 );
nand \U$25108 ( \25354 , \25352 , \25353 );
xor \U$25109 ( \25355 , \24077 , \24437 );
xor \U$25110 ( \25356 , \24178 , \24349 );
xnor \U$25111 ( \25357 , \25356 , \24430 );
not \U$25112 ( \25358 , \25357 );
not \U$25113 ( \25359 , \23985 );
not \U$25114 ( \25360 , \23892 );
or \U$25115 ( \25361 , \25359 , \25360 );
nand \U$25116 ( \25362 , \23891 , \23982 );
nand \U$25117 ( \25363 , \25361 , \25362 );
xor \U$25118 ( \25364 , \25363 , \24075 );
not \U$25119 ( \25365 , \25364 );
or \U$25120 ( \25366 , \25358 , \25365 );
or \U$25121 ( \25367 , \25357 , \25364 );
nand \U$25122 ( \25368 , \25366 , \25367 );
not \U$25123 ( \25369 , \25368 );
not \U$25124 ( \25370 , \25312 );
not \U$25125 ( \25371 , \25177 );
not \U$25126 ( \25372 , \25371 );
or \U$25127 ( \25373 , \25370 , \25372 );
or \U$25128 ( \25374 , \25371 , \25312 );
nand \U$25129 ( \25375 , \25373 , \25374 );
not \U$25130 ( \25376 , \25375 );
or \U$25131 ( \25377 , \25369 , \25376 );
not \U$25132 ( \25378 , \25357 );
nand \U$25133 ( \25379 , \25378 , \25364 );
nand \U$25134 ( \25380 , \25377 , \25379 );
xor \U$25135 ( \25381 , \25355 , \25380 );
xor \U$25136 ( \25382 , \25316 , \25329 );
and \U$25137 ( \25383 , \25381 , \25382 );
and \U$25138 ( \25384 , \25355 , \25380 );
or \U$25139 ( \25385 , \25383 , \25384 );
nand \U$25140 ( \25386 , \25354 , \25385 );
nand \U$25141 ( \25387 , \25349 , \25386 );
not \U$25142 ( \25388 , \25387 );
nor \U$25143 ( \25389 , \24990 , \25348 );
not \U$25144 ( \25390 , \24631 );
not \U$25145 ( \25391 , \24635 );
or \U$25146 ( \25392 , \25390 , \25391 );
not \U$25147 ( \25393 , \24606 );
nand \U$25148 ( \25394 , \25393 , \24627 );
nand \U$25149 ( \25395 , \25392 , \25394 );
or \U$25150 ( \25396 , \24678 , \24676 );
nand \U$25151 ( \25397 , \25396 , \24685 );
nand \U$25152 ( \25398 , \24678 , \24676 );
nand \U$25153 ( \25399 , \25397 , \25398 );
not \U$25154 ( \25400 , \24611 );
not \U$25155 ( \25401 , \11039 );
or \U$25156 ( \25402 , \25400 , \25401 );
xor \U$25157 ( \25403 , RIbe29e48_76, RIbe29ec0_77);
nand \U$25158 ( \25404 , \7368 , \25403 );
nand \U$25159 ( \25405 , \25402 , \25404 );
not \U$25160 ( \25406 , \24915 );
not \U$25161 ( \25407 , \17060 );
or \U$25162 ( \25408 , \25406 , \25407 );
xor \U$25163 ( \25409 , RIbe298a8_64, RIbe2a3e8_88);
nand \U$25164 ( \25410 , \10476 , \25409 );
nand \U$25165 ( \25411 , \25408 , \25410 );
xor \U$25166 ( \25412 , \25405 , \25411 );
not \U$25167 ( \25413 , \24617 );
not \U$25168 ( \25414 , \2600 );
or \U$25169 ( \25415 , \25413 , \25414 );
xor \U$25170 ( \25416 , RIbe2a0a0_81, RIbe27e68_8);
nand \U$25171 ( \25417 , \2603 , \25416 );
nand \U$25172 ( \25418 , \25415 , \25417 );
xnor \U$25173 ( \25419 , \25412 , \25418 );
not \U$25174 ( \25420 , \25419 );
not \U$25175 ( \25421 , \25420 );
not \U$25176 ( \25422 , \24926 );
not \U$25177 ( \25423 , \11345 );
or \U$25178 ( \25424 , \25422 , \25423 );
xor \U$25179 ( \25425 , RIbe29128_48, RIbe2a280_85);
nand \U$25180 ( \25426 , \10849 , \25425 );
nand \U$25181 ( \25427 , \25424 , \25426 );
not \U$25182 ( \25428 , \25427 );
not \U$25183 ( \25429 , \24908 );
not \U$25184 ( \25430 , \16811 );
or \U$25185 ( \25431 , \25429 , \25430 );
xor \U$25186 ( \25432 , RIbe294e8_56, RIbe2b018_114);
nand \U$25187 ( \25433 , \15953 , \25432 );
nand \U$25188 ( \25434 , \25431 , \25433 );
not \U$25189 ( \25435 , \25434 );
not \U$25190 ( \25436 , \25435 );
or \U$25191 ( \25437 , \25428 , \25436 );
or \U$25192 ( \25438 , \25427 , \25435 );
nand \U$25193 ( \25439 , \25437 , \25438 );
not \U$25194 ( \25440 , \24722 );
and \U$25195 ( \25441 , \25439 , \25440 );
not \U$25196 ( \25442 , \25439 );
and \U$25197 ( \25443 , \25442 , \24722 );
nor \U$25198 ( \25444 , \25441 , \25443 );
not \U$25199 ( \25445 , \25444 );
not \U$25200 ( \25446 , \25445 );
or \U$25201 ( \25447 , \25421 , \25446 );
nand \U$25202 ( \25448 , \25444 , \25419 );
nand \U$25203 ( \25449 , \25447 , \25448 );
xor \U$25204 ( \25450 , \25399 , \25449 );
xor \U$25205 ( \25451 , \25395 , \25450 );
not \U$25206 ( \25452 , \24760 );
not \U$25207 ( \25453 , \24747 );
or \U$25208 ( \25454 , \25452 , \25453 );
or \U$25209 ( \25455 , \24747 , \24760 );
nand \U$25210 ( \25456 , \25455 , \24739 );
nand \U$25211 ( \25457 , \25454 , \25456 );
xnor \U$25212 ( \25458 , \25451 , \25457 );
not \U$25213 ( \25459 , \25458 );
not \U$25214 ( \25460 , \24703 );
not \U$25215 ( \25461 , \24765 );
or \U$25216 ( \25462 , \25460 , \25461 );
not \U$25217 ( \25463 , \24694 );
nand \U$25218 ( \25464 , \25463 , \24698 );
nand \U$25219 ( \25465 , \25462 , \25464 );
not \U$25220 ( \25466 , \25465 );
or \U$25221 ( \25467 , \25459 , \25466 );
or \U$25222 ( \25468 , \25465 , \25458 );
nand \U$25223 ( \25469 , \25467 , \25468 );
buf \U$25224 ( \25470 , \25469 );
not \U$25225 ( \25471 , \25470 );
or \U$25226 ( \25472 , \24725 , \24733 );
nand \U$25227 ( \25473 , \25472 , \24727 );
not \U$25228 ( \25474 , \24956 );
not \U$25229 ( \25475 , \24947 );
or \U$25230 ( \25476 , \25474 , \25475 );
nand \U$25231 ( \25477 , \25476 , \24951 );
nand \U$25232 ( \25478 , \24946 , \24957 );
nand \U$25233 ( \25479 , \25477 , \25478 );
and \U$25234 ( \25480 , \25473 , \25479 );
not \U$25235 ( \25481 , \25473 );
nand \U$25236 ( \25482 , \25477 , \25478 );
not \U$25237 ( \25483 , \25482 );
and \U$25238 ( \25484 , \25481 , \25483 );
nor \U$25239 ( \25485 , \25480 , \25484 );
not \U$25240 ( \25486 , \25485 );
or \U$25241 ( \25487 , \24566 , \24560 );
nand \U$25242 ( \25488 , \25487 , \24573 );
nand \U$25243 ( \25489 , \24566 , \24560 );
nand \U$25244 ( \25490 , \25488 , \25489 );
not \U$25245 ( \25491 , \24877 );
not \U$25246 ( \25492 , \1053 );
or \U$25247 ( \25493 , \25491 , \25492 );
xor \U$25248 ( \25494 , RIbe280c0_13, RIbe2b3d8_122);
nand \U$25249 ( \25495 , \1263 , \25494 );
nand \U$25250 ( \25496 , \25493 , \25495 );
not \U$25251 ( \25497 , \24512 );
not \U$25252 ( \25498 , \1780 );
or \U$25253 ( \25499 , \25497 , \25498 );
xor \U$25254 ( \25500 , RIbe28a20_33, RIbe2a640_93);
nand \U$25255 ( \25501 , \1769 , \25500 );
nand \U$25256 ( \25502 , \25499 , \25501 );
xor \U$25257 ( \25503 , \25496 , \25502 );
not \U$25258 ( \25504 , \24884 );
not \U$25259 ( \25505 , \10987 );
or \U$25260 ( \25506 , \25504 , \25505 );
xor \U$25261 ( \25507 , RIbe2a910_99, RIbe28d68_40);
nand \U$25262 ( \25508 , \11456 , \25507 );
nand \U$25263 ( \25509 , \25506 , \25508 );
xor \U$25264 ( \25510 , \25503 , \25509 );
xor \U$25265 ( \25511 , \25490 , \25510 );
not \U$25266 ( \25512 , \24867 );
not \U$25267 ( \25513 , \24861 );
or \U$25268 ( \25514 , \25512 , \25513 );
nand \U$25269 ( \25515 , \24860 , \24854 );
nand \U$25270 ( \25516 , \25514 , \25515 );
xor \U$25271 ( \25517 , \25511 , \25516 );
not \U$25272 ( \25518 , \25517 );
not \U$25273 ( \25519 , \25518 );
and \U$25274 ( \25520 , \25486 , \25519 );
and \U$25275 ( \25521 , \25485 , \25518 );
nor \U$25276 ( \25522 , \25520 , \25521 );
not \U$25277 ( \25523 , \25522 );
not \U$25278 ( \25524 , \24690 );
not \U$25279 ( \25525 , \25524 );
not \U$25280 ( \25526 , \24669 );
or \U$25281 ( \25527 , \25525 , \25526 );
not \U$25282 ( \25528 , \24665 );
nand \U$25283 ( \25529 , \25528 , \24661 );
nand \U$25284 ( \25530 , \25527 , \25529 );
not \U$25285 ( \25531 , \25530 );
or \U$25286 ( \25532 , \25523 , \25531 );
or \U$25287 ( \25533 , \25530 , \25522 );
nand \U$25288 ( \25534 , \25532 , \25533 );
not \U$25289 ( \25535 , \24934 );
not \U$25290 ( \25536 , \24964 );
or \U$25291 ( \25537 , \25535 , \25536 );
nand \U$25292 ( \25538 , \24940 , \24962 );
nand \U$25293 ( \25539 , \25537 , \25538 );
xor \U$25294 ( \25540 , \25534 , \25539 );
not \U$25295 ( \25541 , \25540 );
not \U$25296 ( \25542 , \25541 );
and \U$25297 ( \25543 , \25471 , \25542 );
and \U$25298 ( \25544 , \25470 , \25541 );
nor \U$25299 ( \25545 , \25543 , \25544 );
not \U$25300 ( \25546 , \24965 );
not \U$25301 ( \25547 , \24847 );
or \U$25302 ( \25548 , \25546 , \25547 );
nand \U$25303 ( \25549 , \24835 , \24842 );
nand \U$25304 ( \25550 , \25548 , \25549 );
not \U$25305 ( \25551 , \25550 );
not \U$25306 ( \25552 , \24526 );
nand \U$25307 ( \25553 , \25552 , \24575 );
nand \U$25308 ( \25554 , \25553 , \24578 );
not \U$25309 ( \25555 , \24918 );
not \U$25310 ( \25556 , \24911 );
or \U$25311 ( \25557 , \25555 , \25556 );
nand \U$25312 ( \25558 , \25557 , \24928 );
nand \U$25313 ( \25559 , \24910 , \24917 );
nand \U$25314 ( \25560 , \25558 , \25559 );
xor \U$25315 ( \25561 , \24613 , \24619 );
and \U$25316 ( \25562 , \25561 , \24626 );
and \U$25317 ( \25563 , \24613 , \24619 );
or \U$25318 ( \25564 , \25562 , \25563 );
xor \U$25319 ( \25565 , \25560 , \25564 );
not \U$25320 ( \25566 , \24525 );
not \U$25321 ( \25567 , \24519 );
or \U$25322 ( \25568 , \25566 , \25567 );
nand \U$25323 ( \25569 , \24514 , \24507 );
nand \U$25324 ( \25570 , \25568 , \25569 );
xor \U$25325 ( \25571 , \25565 , \25570 );
xor \U$25326 ( \25572 , \25554 , \25571 );
or \U$25327 ( \25573 , \24930 , \24868 );
nand \U$25328 ( \25574 , \25573 , \24932 );
xor \U$25329 ( \25575 , \25572 , \25574 );
or \U$25330 ( \25576 , \24547 , \24533 );
nand \U$25331 ( \25577 , \25576 , \24549 );
not \U$25332 ( \25578 , \25577 );
not \U$25333 ( \25579 , \24587 );
not \U$25334 ( \25580 , \24605 );
or \U$25335 ( \25581 , \25579 , \25580 );
nand \U$25336 ( \25582 , \24601 , \24593 );
nand \U$25337 ( \25583 , \25581 , \25582 );
not \U$25338 ( \25584 , \25583 );
not \U$25339 ( \25585 , \25584 );
or \U$25340 ( \25586 , \25578 , \25585 );
or \U$25341 ( \25587 , \25584 , \25577 );
nand \U$25342 ( \25588 , \25586 , \25587 );
not \U$25343 ( \25589 , \24879 );
not \U$25344 ( \25590 , \24898 );
or \U$25345 ( \25591 , \25589 , \25590 );
nand \U$25346 ( \25592 , \24893 , \24886 );
nand \U$25347 ( \25593 , \25591 , \25592 );
not \U$25348 ( \25594 , \25593 );
and \U$25349 ( \25595 , \25588 , \25594 );
not \U$25350 ( \25596 , \25588 );
and \U$25351 ( \25597 , \25596 , \25593 );
nor \U$25352 ( \25598 , \25595 , \25597 );
not \U$25353 ( \25599 , \25598 );
nand \U$25354 ( \25600 , \907 , RIbe2ae38_110);
not \U$25355 ( \25601 , \25600 );
not \U$25356 ( \25602 , \24714 );
not \U$25357 ( \25603 , \15059 );
or \U$25358 ( \25604 , \25602 , \25603 );
xor \U$25359 ( \25605 , RIbe28228_16, RIbe2a730_95);
nand \U$25360 ( \25606 , \885 , \25605 );
nand \U$25361 ( \25607 , \25604 , \25606 );
not \U$25362 ( \25608 , \25607 );
or \U$25363 ( \25609 , \25601 , \25608 );
or \U$25364 ( \25610 , \25607 , \25600 );
nand \U$25365 ( \25611 , \25609 , \25610 );
not \U$25366 ( \25612 , \25611 );
not \U$25367 ( \25613 , \16897 );
xnor \U$25368 ( \25614 , RIbe295d8_58, RIbe2b108_116);
not \U$25369 ( \25615 , \25614 );
and \U$25370 ( \25616 , \25613 , \25615 );
buf \U$25371 ( \25617 , \14296 );
buf \U$25372 ( \25618 , \25617 );
and \U$25373 ( \25619 , \25618 , \24891 );
nor \U$25374 ( \25620 , \25616 , \25619 );
not \U$25375 ( \25621 , \25620 );
or \U$25376 ( \25622 , \25612 , \25621 );
or \U$25377 ( \25623 , \25611 , \25620 );
nand \U$25378 ( \25624 , \25622 , \25623 );
not \U$25379 ( \25625 , \25624 );
not \U$25380 ( \25626 , \25625 );
not \U$25381 ( \25627 , \24865 );
not \U$25382 ( \25628 , \10831 );
or \U$25383 ( \25629 , \25627 , \25628 );
xor \U$25384 ( \25630 , RIbe29a10_67, RIbe2a190_83);
nand \U$25385 ( \25631 , \10695 , \25630 );
nand \U$25386 ( \25632 , \25629 , \25631 );
not \U$25387 ( \25633 , \24858 );
not \U$25388 ( \25634 , \2552 );
or \U$25389 ( \25635 , \25633 , \25634 );
xor \U$25390 ( \25636 , RIbe28b88_36, RIbe2b4c8_124);
nand \U$25391 ( \25637 , \7549 , \25636 );
nand \U$25392 ( \25638 , \25635 , \25637 );
xor \U$25393 ( \25639 , \25632 , \25638 );
not \U$25394 ( \25640 , \24624 );
not \U$25395 ( \25641 , \7513 );
or \U$25396 ( \25642 , \25640 , \25641 );
xor \U$25397 ( \25643 , RIbe29c68_72, RIbe2b6a8_128);
nand \U$25398 ( \25644 , \4580 , \25643 );
nand \U$25399 ( \25645 , \25642 , \25644 );
xnor \U$25400 ( \25646 , \25639 , \25645 );
not \U$25401 ( \25647 , \25646 );
not \U$25402 ( \25648 , \25647 );
or \U$25403 ( \25649 , \25626 , \25648 );
nand \U$25404 ( \25650 , \25646 , \25624 );
nand \U$25405 ( \25651 , \25649 , \25650 );
not \U$25406 ( \25652 , \24571 );
not \U$25407 ( \25653 , \14806 );
or \U$25408 ( \25654 , \25652 , \25653 );
xor \U$25409 ( \25655 , RIbe28390_19, RIbe2ad48_108);
nand \U$25410 ( \25656 , \8654 , \25655 );
nand \U$25411 ( \25657 , \25654 , \25656 );
not \U$25412 ( \25658 , \24558 );
not \U$25413 ( \25659 , \20574 );
or \U$25414 ( \25660 , \25658 , \25659 );
xor \U$25415 ( \25661 , RIbe28a98_34, RIbe2aaf0_103);
nand \U$25416 ( \25662 , \25661 , RIbe2ab68_104);
nand \U$25417 ( \25663 , \25660 , \25662 );
xor \U$25418 ( \25664 , \25657 , \25663 );
not \U$25419 ( \25665 , \24852 );
not \U$25420 ( \25666 , \3344 );
or \U$25421 ( \25667 , \25665 , \25666 );
xor \U$25422 ( \25668 , RIbe2a460_89, RIbe28480_21);
nand \U$25423 ( \25669 , \11263 , \25668 );
nand \U$25424 ( \25670 , \25667 , \25669 );
xnor \U$25425 ( \25671 , \25664 , \25670 );
not \U$25426 ( \25672 , \25671 );
and \U$25427 ( \25673 , \25651 , \25672 );
not \U$25428 ( \25674 , \25651 );
and \U$25429 ( \25675 , \25674 , \25671 );
nor \U$25430 ( \25676 , \25673 , \25675 );
not \U$25431 ( \25677 , \25676 );
or \U$25432 ( \25678 , \25599 , \25677 );
or \U$25433 ( \25679 , \25598 , \25676 );
nand \U$25434 ( \25680 , \25678 , \25679 );
not \U$25435 ( \25681 , \24538 );
not \U$25436 ( \25682 , \9374 );
or \U$25437 ( \25683 , \25681 , \25682 );
xor \U$25438 ( \25684 , RIbe27b20_1, RIbe2a2f8_86);
nand \U$25439 ( \25685 , \8705 , \25684 );
nand \U$25440 ( \25686 , \25683 , \25685 );
not \U$25441 ( \25687 , \24530 );
not \U$25442 ( \25688 , \7618 );
or \U$25443 ( \25689 , \25687 , \25688 );
xor \U$25444 ( \25690 , RIbe285e8_24, RIbe2b2e8_120);
nand \U$25445 ( \25691 , \8270 , \25690 );
nand \U$25446 ( \25692 , \25689 , \25691 );
xor \U$25447 ( \25693 , \25686 , \25692 );
not \U$25448 ( \25694 , \24599 );
not \U$25449 ( \25695 , \16913 );
or \U$25450 ( \25696 , \25694 , \25695 );
xor \U$25451 ( \25697 , RIbe282a0_17, RIbe2af28_112);
nand \U$25452 ( \25698 , \17810 , \25697 );
nand \U$25453 ( \25699 , \25696 , \25698 );
xor \U$25454 ( \25700 , \25693 , \25699 );
not \U$25455 ( \25701 , \25700 );
not \U$25456 ( \25702 , \25701 );
not \U$25457 ( \25703 , \24544 );
not \U$25458 ( \25704 , \14852 );
or \U$25459 ( \25705 , \25703 , \25704 );
xor \U$25460 ( \25706 , RIbe2b180_117, RIbe297b8_62);
nand \U$25461 ( \25707 , \14966 , \25706 );
nand \U$25462 ( \25708 , \25705 , \25707 );
not \U$25463 ( \25709 , \25708 );
not \U$25464 ( \25710 , \24523 );
not \U$25465 ( \25711 , \9825 );
or \U$25466 ( \25712 , \25710 , \25711 );
xor \U$25467 ( \25713 , RIbe2a820_97, RIbe27fd0_11);
nand \U$25468 ( \25714 , \4897 , \25713 );
nand \U$25469 ( \25715 , \25712 , \25714 );
not \U$25470 ( \25716 , \25715 );
and \U$25471 ( \25717 , \25709 , \25716 );
not \U$25472 ( \25718 , \25709 );
and \U$25473 ( \25719 , \25718 , \25715 );
nor \U$25474 ( \25720 , \25717 , \25719 );
not \U$25475 ( \25721 , \24505 );
not \U$25476 ( \25722 , \966 );
or \U$25477 ( \25723 , \25721 , \25722 );
xor \U$25478 ( \25724 , RIbe28930_31, RIbe2abe0_105);
nand \U$25479 ( \25725 , \1199 , \25724 );
nand \U$25480 ( \25726 , \25723 , \25725 );
not \U$25481 ( \25727 , \25726 );
and \U$25482 ( \25728 , \25720 , \25727 );
not \U$25483 ( \25729 , \25720 );
and \U$25484 ( \25730 , \25729 , \25726 );
nor \U$25485 ( \25731 , \25728 , \25730 );
not \U$25486 ( \25732 , \25731 );
not \U$25487 ( \25733 , \25732 );
or \U$25488 ( \25734 , \25702 , \25733 );
nand \U$25489 ( \25735 , \25731 , \25700 );
nand \U$25490 ( \25736 , \25734 , \25735 );
not \U$25491 ( \25737 , \24585 );
not \U$25492 ( \25738 , \10433 );
or \U$25493 ( \25739 , \25737 , \25738 );
xor \U$25494 ( \25740 , RIbe2a550_91, RIbe27df0_7);
nand \U$25495 ( \25741 , \14612 , \25740 );
nand \U$25496 ( \25742 , \25739 , \25741 );
not \U$25497 ( \25743 , \24564 );
not \U$25498 ( \25744 , \8400 );
or \U$25499 ( \25745 , \25743 , \25744 );
xor \U$25500 ( \25746 , RIbe2a028_80, RIbe29ce0_73);
nand \U$25501 ( \25747 , \8930 , \25746 );
nand \U$25502 ( \25748 , \25745 , \25747 );
xor \U$25503 ( \25749 , \25742 , \25748 );
not \U$25504 ( \25750 , \24591 );
not \U$25505 ( \25751 , \7609 );
or \U$25506 ( \25752 , \25750 , \25751 );
xor \U$25507 ( \25753 , RIbe28f48_44, RIbe2aa00_101);
nand \U$25508 ( \25754 , \4180 , \25753 );
nand \U$25509 ( \25755 , \25752 , \25754 );
not \U$25510 ( \25756 , \25755 );
xor \U$25511 ( \25757 , \25749 , \25756 );
not \U$25512 ( \25758 , \25757 );
and \U$25513 ( \25759 , \25736 , \25758 );
not \U$25514 ( \25760 , \25736 );
and \U$25515 ( \25761 , \25760 , \25757 );
nor \U$25516 ( \25762 , \25759 , \25761 );
and \U$25517 ( \25763 , \25680 , \25762 );
not \U$25518 ( \25764 , \25680 );
not \U$25519 ( \25765 , \25762 );
and \U$25520 ( \25766 , \25764 , \25765 );
nor \U$25521 ( \25767 , \25763 , \25766 );
xor \U$25522 ( \25768 , \25575 , \25767 );
not \U$25523 ( \25769 , \24645 );
not \U$25524 ( \25770 , \24640 );
or \U$25525 ( \25771 , \25769 , \25770 );
not \U$25526 ( \25772 , \24580 );
nand \U$25527 ( \25773 , \25772 , \24636 );
nand \U$25528 ( \25774 , \25771 , \25773 );
xor \U$25529 ( \25775 , \25768 , \25774 );
xor \U$25530 ( \25776 , \25551 , \25775 );
not \U$25531 ( \25777 , \24770 );
not \U$25532 ( \25778 , \24656 );
or \U$25533 ( \25779 , \25777 , \25778 );
nand \U$25534 ( \25780 , \24501 , \24651 );
nand \U$25535 ( \25781 , \25779 , \25780 );
xnor \U$25536 ( \25782 , \25776 , \25781 );
xor \U$25537 ( \25783 , \25545 , \25782 );
not \U$25538 ( \25784 , \24982 );
not \U$25539 ( \25785 , \25784 );
not \U$25540 ( \25786 , \24830 );
or \U$25541 ( \25787 , \25785 , \25786 );
nand \U$25542 ( \25788 , \24970 , \24977 );
nand \U$25543 ( \25789 , \25787 , \25788 );
xnor \U$25544 ( \25790 , \25783 , \25789 );
not \U$25545 ( \25791 , \24986 );
not \U$25546 ( \25792 , \25791 );
not \U$25547 ( \25793 , \24776 );
or \U$25548 ( \25794 , \25792 , \25793 );
nand \U$25549 ( \25795 , \24449 , \24775 );
nand \U$25550 ( \25796 , \25794 , \25795 );
nor \U$25551 ( \25797 , \25790 , \25796 );
nor \U$25552 ( \25798 , \25389 , \25797 );
not \U$25553 ( \25799 , \25798 );
or \U$25554 ( \25800 , \25388 , \25799 );
nand \U$25555 ( \25801 , \25796 , \25790 );
not \U$25556 ( \25802 , \25545 );
not \U$25557 ( \25803 , \25802 );
not \U$25558 ( \25804 , \25782 );
or \U$25559 ( \25805 , \25803 , \25804 );
not \U$25560 ( \25806 , \25789 );
nand \U$25561 ( \25807 , \25805 , \25806 );
not \U$25562 ( \25808 , \25782 );
nand \U$25563 ( \25809 , \25808 , \25545 );
nand \U$25564 ( \25810 , \25807 , \25809 );
not \U$25565 ( \25811 , \25810 );
not \U$25566 ( \25812 , \25539 );
not \U$25567 ( \25813 , \25534 );
or \U$25568 ( \25814 , \25812 , \25813 );
not \U$25569 ( \25815 , \25522 );
nand \U$25570 ( \25816 , \25815 , \25530 );
nand \U$25571 ( \25817 , \25814 , \25816 );
not \U$25572 ( \25818 , \25817 );
not \U$25573 ( \25819 , \25399 );
not \U$25574 ( \25820 , \25449 );
or \U$25575 ( \25821 , \25819 , \25820 );
nand \U$25576 ( \25822 , \25444 , \25420 );
nand \U$25577 ( \25823 , \25821 , \25822 );
xor \U$25578 ( \25824 , \25554 , \25571 );
and \U$25579 ( \25825 , \25824 , \25574 );
and \U$25580 ( \25826 , \25554 , \25571 );
or \U$25581 ( \25827 , \25825 , \25826 );
xor \U$25582 ( \25828 , \25823 , \25827 );
not \U$25583 ( \25829 , \25828 );
not \U$25584 ( \25830 , \25517 );
not \U$25585 ( \25831 , \25485 );
or \U$25586 ( \25832 , \25830 , \25831 );
nand \U$25587 ( \25833 , \25473 , \25482 );
nand \U$25588 ( \25834 , \25832 , \25833 );
not \U$25589 ( \25835 , \25834 );
not \U$25590 ( \25836 , \25835 );
and \U$25591 ( \25837 , \25829 , \25836 );
and \U$25592 ( \25838 , \25828 , \25835 );
nor \U$25593 ( \25839 , \25837 , \25838 );
not \U$25594 ( \25840 , \25839 );
or \U$25595 ( \25841 , \25818 , \25840 );
or \U$25596 ( \25842 , \25839 , \25817 );
nand \U$25597 ( \25843 , \25841 , \25842 );
not \U$25598 ( \25844 , \25767 );
not \U$25599 ( \25845 , \25575 );
not \U$25600 ( \25846 , \25845 );
not \U$25601 ( \25847 , \25774 );
or \U$25602 ( \25848 , \25846 , \25847 );
or \U$25603 ( \25849 , \25774 , \25845 );
nand \U$25604 ( \25850 , \25848 , \25849 );
not \U$25605 ( \25851 , \25850 );
or \U$25606 ( \25852 , \25844 , \25851 );
nand \U$25607 ( \25853 , \25774 , \25575 );
nand \U$25608 ( \25854 , \25852 , \25853 );
xor \U$25609 ( \25855 , \25843 , \25854 );
not \U$25610 ( \25856 , \25540 );
not \U$25611 ( \25857 , \25469 );
or \U$25612 ( \25858 , \25856 , \25857 );
not \U$25613 ( \25859 , \25458 );
nand \U$25614 ( \25860 , \25859 , \25465 );
nand \U$25615 ( \25861 , \25858 , \25860 );
not \U$25616 ( \25862 , \25440 );
not \U$25617 ( \25863 , \25439 );
or \U$25618 ( \25864 , \25862 , \25863 );
not \U$25619 ( \25865 , \25435 );
nand \U$25620 ( \25866 , \25865 , \25427 );
nand \U$25621 ( \25867 , \25864 , \25866 );
not \U$25622 ( \25868 , \25867 );
not \U$25623 ( \25869 , \25868 );
xor \U$25624 ( \25870 , \25560 , \25564 );
and \U$25625 ( \25871 , \25870 , \25570 );
and \U$25626 ( \25872 , \25560 , \25564 );
or \U$25627 ( \25873 , \25871 , \25872 );
not \U$25628 ( \25874 , \25873 );
or \U$25629 ( \25875 , \25869 , \25874 );
or \U$25630 ( \25876 , \25873 , \25868 );
nand \U$25631 ( \25877 , \25875 , \25876 );
not \U$25632 ( \25878 , \25494 );
not \U$25633 ( \25879 , \860 );
or \U$25634 ( \25880 , \25878 , \25879 );
xor \U$25635 ( \25881 , RIbe280c0_13, RIbe2b450_123);
nand \U$25636 ( \25882 , \869 , \25881 );
nand \U$25637 ( \25883 , \25880 , \25882 );
or \U$25638 ( \25884 , RIbe280c0_13, RIbe29830_63);
nand \U$25639 ( \25885 , \25884 , RIbe2ae38_110);
nand \U$25640 ( \25886 , RIbe280c0_13, RIbe29830_63);
and \U$25641 ( \25887 , \25885 , \25886 , RIbe296c8_60);
or \U$25642 ( \25888 , \25883 , \25887 );
nand \U$25643 ( \25889 , \25883 , \25887 );
nand \U$25644 ( \25890 , \25888 , \25889 );
not \U$25645 ( \25891 , \19371 );
not \U$25646 ( \25892 , \25891 );
xor \U$25647 ( \25893 , RIbe288b8_30, RIbe2b018_114);
not \U$25648 ( \25894 , \25893 );
not \U$25649 ( \25895 , \25894 );
and \U$25650 ( \25896 , \25892 , \25895 );
buf \U$25651 ( \25897 , \17571 );
and \U$25652 ( \25898 , \25897 , \25432 );
nor \U$25653 ( \25899 , \25896 , \25898 );
or \U$25654 ( \25900 , \25890 , \25899 );
nand \U$25655 ( \25901 , \25890 , \25899 );
and \U$25656 ( \25902 , \25900 , \25901 );
not \U$25657 ( \25903 , \25418 );
not \U$25658 ( \25904 , \25411 );
or \U$25659 ( \25905 , \25903 , \25904 );
or \U$25660 ( \25906 , \25411 , \25418 );
nand \U$25661 ( \25907 , \25906 , \25405 );
nand \U$25662 ( \25908 , \25905 , \25907 );
buf \U$25663 ( \25909 , \25908 );
xor \U$25664 ( \25910 , \25902 , \25909 );
and \U$25665 ( \25911 , \25877 , \25910 );
not \U$25666 ( \25912 , \25877 );
not \U$25667 ( \25913 , \25910 );
and \U$25668 ( \25914 , \25912 , \25913 );
nor \U$25669 ( \25915 , \25911 , \25914 );
not \U$25670 ( \25916 , \25632 );
not \U$25671 ( \25917 , \25638 );
or \U$25672 ( \25918 , \25916 , \25917 );
or \U$25673 ( \25919 , \25638 , \25632 );
nand \U$25674 ( \25920 , \25919 , \25645 );
nand \U$25675 ( \25921 , \25918 , \25920 );
not \U$25676 ( \25922 , \25708 );
not \U$25677 ( \25923 , \25715 );
or \U$25678 ( \25924 , \25922 , \25923 );
not \U$25679 ( \25925 , \25716 );
not \U$25680 ( \25926 , \25709 );
or \U$25681 ( \25927 , \25925 , \25926 );
nand \U$25682 ( \25928 , \25927 , \25726 );
nand \U$25683 ( \25929 , \25924 , \25928 );
not \U$25684 ( \25930 , \25929 );
not \U$25685 ( \25931 , \25620 );
not \U$25686 ( \25932 , \25931 );
not \U$25687 ( \25933 , \25611 );
or \U$25688 ( \25934 , \25932 , \25933 );
not \U$25689 ( \25935 , \25600 );
nand \U$25690 ( \25936 , \25935 , \25607 );
nand \U$25691 ( \25937 , \25934 , \25936 );
not \U$25692 ( \25938 , \25937 );
not \U$25693 ( \25939 , \25938 );
or \U$25694 ( \25940 , \25930 , \25939 );
or \U$25695 ( \25941 , \25938 , \25929 );
nand \U$25696 ( \25942 , \25940 , \25941 );
xor \U$25697 ( \25943 , \25921 , \25942 );
not \U$25698 ( \25944 , \25943 );
not \U$25699 ( \25945 , \25944 );
not \U$25700 ( \25946 , \25672 );
not \U$25701 ( \25947 , \25647 );
or \U$25702 ( \25948 , \25946 , \25947 );
not \U$25703 ( \25949 , \25646 );
not \U$25704 ( \25950 , \25671 );
or \U$25705 ( \25951 , \25949 , \25950 );
nand \U$25706 ( \25952 , \25951 , \25624 );
nand \U$25707 ( \25953 , \25948 , \25952 );
not \U$25708 ( \25954 , \25953 );
or \U$25709 ( \25955 , \25748 , \25742 );
nand \U$25710 ( \25956 , \25955 , \25755 );
nand \U$25711 ( \25957 , \25748 , \25742 );
nand \U$25712 ( \25958 , \25956 , \25957 );
xor \U$25713 ( \25959 , \25496 , \25502 );
and \U$25714 ( \25960 , \25959 , \25509 );
and \U$25715 ( \25961 , \25496 , \25502 );
or \U$25716 ( \25962 , \25960 , \25961 );
xor \U$25717 ( \25963 , \25958 , \25962 );
or \U$25718 ( \25964 , \25699 , \25692 );
nand \U$25719 ( \25965 , \25964 , \25686 );
nand \U$25720 ( \25966 , \25699 , \25692 );
nand \U$25721 ( \25967 , \25965 , \25966 );
xnor \U$25722 ( \25968 , \25963 , \25967 );
not \U$25723 ( \25969 , \25968 );
or \U$25724 ( \25970 , \25954 , \25969 );
or \U$25725 ( \25971 , \25953 , \25968 );
nand \U$25726 ( \25972 , \25970 , \25971 );
not \U$25727 ( \25973 , \25972 );
or \U$25728 ( \25974 , \25945 , \25973 );
or \U$25729 ( \25975 , \25972 , \25944 );
nand \U$25730 ( \25976 , \25974 , \25975 );
xor \U$25731 ( \25977 , \25915 , \25976 );
not \U$25732 ( \25978 , \25758 );
not \U$25733 ( \25979 , \25700 );
or \U$25734 ( \25980 , \25978 , \25979 );
not \U$25735 ( \25981 , \25757 );
not \U$25736 ( \25982 , \25701 );
or \U$25737 ( \25983 , \25981 , \25982 );
nand \U$25738 ( \25984 , \25983 , \25732 );
nand \U$25739 ( \25985 , \25980 , \25984 );
xor \U$25740 ( \25986 , \25490 , \25510 );
and \U$25741 ( \25987 , \25986 , \25516 );
and \U$25742 ( \25988 , \25490 , \25510 );
or \U$25743 ( \25989 , \25987 , \25988 );
xor \U$25744 ( \25990 , \25985 , \25989 );
not \U$25745 ( \25991 , \25593 );
not \U$25746 ( \25992 , \25588 );
or \U$25747 ( \25993 , \25991 , \25992 );
not \U$25748 ( \25994 , \25584 );
nand \U$25749 ( \25995 , \25994 , \25577 );
nand \U$25750 ( \25996 , \25993 , \25995 );
xor \U$25751 ( \25997 , \25990 , \25996 );
xor \U$25752 ( \25998 , \25977 , \25997 );
not \U$25753 ( \25999 , \25998 );
not \U$25754 ( \26000 , \25762 );
not \U$25755 ( \26001 , \25680 );
or \U$25756 ( \26002 , \26000 , \26001 );
not \U$25757 ( \26003 , \25598 );
nand \U$25758 ( \26004 , \26003 , \25676 );
nand \U$25759 ( \26005 , \26002 , \26004 );
not \U$25760 ( \26006 , \26005 );
not \U$25761 ( \26007 , \26006 );
not \U$25762 ( \26008 , \25670 );
not \U$25763 ( \26009 , \25664 );
or \U$25764 ( \26010 , \26008 , \26009 );
nand \U$25765 ( \26011 , \25657 , \25663 );
nand \U$25766 ( \26012 , \26010 , \26011 );
not \U$25767 ( \26013 , \25643 );
not \U$25768 ( \26014 , \14971 );
or \U$25769 ( \26015 , \26013 , \26014 );
xor \U$25770 ( \26016 , RIbe29c68_72, RIbe29f38_78);
nand \U$25771 ( \26017 , \4580 , \26016 );
nand \U$25772 ( \26018 , \26015 , \26017 );
not \U$25773 ( \26019 , \25630 );
not \U$25774 ( \26020 , \10831 );
or \U$25775 ( \26021 , \26019 , \26020 );
xor \U$25776 ( \26022 , RIbe2a190_83, RIbe29b00_69);
nand \U$25777 ( \26023 , \22918 , \26022 );
nand \U$25778 ( \26024 , \26021 , \26023 );
xor \U$25779 ( \26025 , \26018 , \26024 );
not \U$25780 ( \26026 , \25684 );
not \U$25781 ( \26027 , \9375 );
or \U$25782 ( \26028 , \26026 , \26027 );
xor \U$25783 ( \26029 , RIbe28cf0_39, RIbe2a2f8_86);
nand \U$25784 ( \26030 , \8706 , \26029 );
nand \U$25785 ( \26031 , \26028 , \26030 );
and \U$25786 ( \26032 , \26025 , \26031 );
not \U$25787 ( \26033 , \26025 );
not \U$25788 ( \26034 , \26031 );
and \U$25789 ( \26035 , \26033 , \26034 );
nor \U$25790 ( \26036 , \26032 , \26035 );
xor \U$25791 ( \26037 , \26012 , \26036 );
not \U$25792 ( \26038 , \25425 );
not \U$25793 ( \26039 , \20237 );
or \U$25794 ( \26040 , \26038 , \26039 );
xor \U$25795 ( \26041 , RIbe291a0_49, RIbe2a280_85);
nand \U$25796 ( \26042 , \18667 , \26041 );
nand \U$25797 ( \26043 , \26040 , \26042 );
not \U$25798 ( \26044 , \25409 );
not \U$25799 ( \26045 , \8806 );
or \U$25800 ( \26046 , \26044 , \26045 );
xor \U$25801 ( \26047 , RIbe29998_66, RIbe2a3e8_88);
nand \U$25802 ( \26048 , \8794 , \26047 );
nand \U$25803 ( \26049 , \26046 , \26048 );
xor \U$25804 ( \26050 , \26043 , \26049 );
xor \U$25805 ( \26051 , RIbe296c8_60, RIbe2ae38_110);
not \U$25806 ( \26052 , \26051 );
not \U$25807 ( \26053 , \2875 );
or \U$25808 ( \26054 , \26052 , \26053 );
xor \U$25809 ( \26055 , RIbe2aeb0_111, RIbe296c8_60);
nand \U$25810 ( \26056 , \1137 , \26055 );
nand \U$25811 ( \26057 , \26054 , \26056 );
xor \U$25812 ( \26058 , \26050 , \26057 );
xor \U$25813 ( \26059 , \26037 , \26058 );
not \U$25814 ( \26060 , \26059 );
not \U$25815 ( \26061 , \25746 );
not \U$25816 ( \26062 , \8400 );
or \U$25817 ( \26063 , \26061 , \26062 );
xor \U$25818 ( \26064 , RIbe2a028_80, RIbe29b78_70);
nand \U$25819 ( \26065 , \8172 , \26064 );
nand \U$25820 ( \26066 , \26063 , \26065 );
or \U$25821 ( \26067 , \13540 , \25614 );
and \U$25822 ( \26068 , RIbe2b108_116, RIbe29740_61);
not \U$25823 ( \26069 , RIbe2b108_116);
and \U$25824 ( \26070 , \26069 , \3185 );
nor \U$25825 ( \26071 , \26068 , \26070 );
not \U$25826 ( \26072 , \26071 );
or \U$25827 ( \26073 , \16897 , \26072 );
nand \U$25828 ( \26074 , \26067 , \26073 );
xor \U$25829 ( \26075 , \26066 , \26074 );
not \U$25830 ( \26076 , \25668 );
not \U$25831 ( \26077 , \2518 );
or \U$25832 ( \26078 , \26076 , \26077 );
xor \U$25833 ( \26079 , RIbe28480_21, RIbe2a4d8_90);
nand \U$25834 ( \26080 , \7483 , \26079 );
nand \U$25835 ( \26081 , \26078 , \26080 );
not \U$25836 ( \26082 , \26081 );
and \U$25837 ( \26083 , \26075 , \26082 );
not \U$25838 ( \26084 , \26075 );
and \U$25839 ( \26085 , \26084 , \26081 );
nor \U$25840 ( \26086 , \26083 , \26085 );
not \U$25841 ( \26087 , \26086 );
not \U$25842 ( \26088 , \26087 );
not \U$25843 ( \26089 , \25636 );
nor \U$25844 ( \26090 , \26089 , \23728 );
xor \U$25845 ( \26091 , RIbe28b88_36, RIbe2b540_125);
and \U$25846 ( \26092 , \7550 , \26091 );
nor \U$25847 ( \26093 , \26090 , \26092 );
not \U$25848 ( \26094 , \25403 );
not \U$25849 ( \26095 , \14307 );
or \U$25850 ( \26096 , \26094 , \26095 );
xor \U$25851 ( \26097 , RIbe29d58_74, RIbe29e48_76);
nand \U$25852 ( \26098 , \4849 , \26097 );
nand \U$25853 ( \26099 , \26096 , \26098 );
not \U$25854 ( \26100 , \26099 );
not \U$25855 ( \26101 , \26100 );
not \U$25856 ( \26102 , \25697 );
not \U$25857 ( \26103 , \14423 );
or \U$25858 ( \26104 , \26102 , \26103 );
xor \U$25859 ( \26105 , RIbe29470_55, RIbe2af28_112);
nand \U$25860 ( \26106 , \14413 , \26105 );
nand \U$25861 ( \26107 , \26104 , \26106 );
not \U$25862 ( \26108 , \26107 );
or \U$25863 ( \26109 , \26101 , \26108 );
or \U$25864 ( \26110 , \26107 , \26100 );
nand \U$25865 ( \26111 , \26109 , \26110 );
xnor \U$25866 ( \26112 , \26093 , \26111 );
not \U$25867 ( \26113 , \26112 );
not \U$25868 ( \26114 , \26113 );
or \U$25869 ( \26115 , \26088 , \26114 );
nand \U$25870 ( \26116 , \26112 , \26086 );
nand \U$25871 ( \26117 , \26115 , \26116 );
not \U$25872 ( \26118 , \25706 );
not \U$25873 ( \26119 , \15353 );
or \U$25874 ( \26120 , \26118 , \26119 );
xor \U$25875 ( \26121 , RIbe2b180_117, RIbe28138_14);
nand \U$25876 ( \26122 , \16646 , \26121 );
nand \U$25877 ( \26123 , \26120 , \26122 );
not \U$25878 ( \26124 , \25713 );
not \U$25879 ( \26125 , \10466 );
or \U$25880 ( \26126 , \26124 , \26125 );
xor \U$25881 ( \26127 , RIbe27fd0_11, RIbe2a898_98);
nand \U$25882 ( \26128 , \4897 , \26127 );
nand \U$25883 ( \26129 , \26126 , \26128 );
xor \U$25884 ( \26130 , \26123 , \26129 );
not \U$25885 ( \26131 , \25507 );
not \U$25886 ( \26132 , \12716 );
or \U$25887 ( \26133 , \26131 , \26132 );
xor \U$25888 ( \26134 , RIbe27c88_4, RIbe2a910_99);
nand \U$25889 ( \26135 , \9726 , \26134 );
nand \U$25890 ( \26136 , \26133 , \26135 );
xor \U$25891 ( \26137 , \26130 , \26136 );
not \U$25892 ( \26138 , \26137 );
and \U$25893 ( \26139 , \26117 , \26138 );
not \U$25894 ( \26140 , \26117 );
and \U$25895 ( \26141 , \26140 , \26137 );
nor \U$25896 ( \26142 , \26139 , \26141 );
not \U$25897 ( \26143 , \26142 );
or \U$25898 ( \26144 , \26060 , \26143 );
or \U$25899 ( \26145 , \26142 , \26059 );
nand \U$25900 ( \26146 , \26144 , \26145 );
xor \U$25901 ( \26147 , RIbe293f8_54, RIbe2aaf0_103);
not \U$25902 ( \26148 , \26147 );
not \U$25903 ( \26149 , RIbe2ab68_104);
or \U$25904 ( \26150 , \26148 , \26149 );
not \U$25905 ( \26151 , \25661 );
or \U$25906 ( \26152 , \19580 , \26151 );
nand \U$25907 ( \26153 , \26150 , \26152 );
not \U$25908 ( \26154 , \26153 );
not \U$25909 ( \26155 , \25753 );
not \U$25910 ( \26156 , \11461 );
or \U$25911 ( \26157 , \26155 , \26156 );
xor \U$25912 ( \26158 , RIbe28f48_44, RIbe2aa78_102);
nand \U$25913 ( \26159 , \11201 , \26158 );
nand \U$25914 ( \26160 , \26157 , \26159 );
not \U$25915 ( \26161 , \26160 );
not \U$25916 ( \26162 , \26161 );
or \U$25917 ( \26163 , \26154 , \26162 );
not \U$25918 ( \26164 , \26153 );
nand \U$25919 ( \26165 , \26164 , \26160 );
nand \U$25920 ( \26166 , \26163 , \26165 );
not \U$25921 ( \26167 , \25690 );
not \U$25922 ( \26168 , \2618 );
or \U$25923 ( \26169 , \26167 , \26168 );
xor \U$25924 ( \26170 , RIbe285e8_24, RIbe2b360_121);
nand \U$25925 ( \26171 , \2758 , \26170 );
nand \U$25926 ( \26172 , \26169 , \26171 );
not \U$25927 ( \26173 , \26172 );
and \U$25928 ( \26174 , \26166 , \26173 );
not \U$25929 ( \26175 , \26166 );
and \U$25930 ( \26176 , \26175 , \26172 );
nor \U$25931 ( \26177 , \26174 , \26176 );
not \U$25932 ( \26178 , \26177 );
not \U$25933 ( \26179 , \25724 );
not \U$25934 ( \26180 , \965 );
or \U$25935 ( \26181 , \26179 , \26180 );
xor \U$25936 ( \26182 , RIbe28930_31, RIbe2ac58_106);
nand \U$25937 ( \26183 , \1199 , \26182 );
nand \U$25938 ( \26184 , \26181 , \26183 );
not \U$25939 ( \26185 , \25416 );
not \U$25940 ( \26186 , \4443 );
or \U$25941 ( \26187 , \26185 , \26186 );
xor \U$25942 ( \26188 , RIbe2a118_82, RIbe27e68_8);
nand \U$25943 ( \26189 , \2603 , \26188 );
nand \U$25944 ( \26190 , \26187 , \26189 );
xor \U$25945 ( \26191 , \26184 , \26190 );
not \U$25946 ( \26192 , \25605 );
not \U$25947 ( \26193 , \879 );
or \U$25948 ( \26194 , \26192 , \26193 );
xor \U$25949 ( \26195 , RIbe28228_16, RIbe2a7a8_96);
nand \U$25950 ( \26196 , \8680 , \26195 );
nand \U$25951 ( \26197 , \26194 , \26196 );
xor \U$25952 ( \26198 , \26191 , \26197 );
not \U$25953 ( \26199 , \26198 );
or \U$25954 ( \26200 , \26178 , \26199 );
or \U$25955 ( \26201 , \26198 , \26177 );
nand \U$25956 ( \26202 , \26200 , \26201 );
not \U$25957 ( \26203 , \25740 );
not \U$25958 ( \26204 , \11999 );
or \U$25959 ( \26205 , \26203 , \26204 );
xor \U$25960 ( \26206 , RIbe2a550_91, RIbe29218_50);
nand \U$25961 ( \26207 , \20336 , \26206 );
nand \U$25962 ( \26208 , \26205 , \26207 );
not \U$25963 ( \26209 , \25500 );
not \U$25964 ( \26210 , \1780 );
or \U$25965 ( \26211 , \26209 , \26210 );
xor \U$25966 ( \26212 , RIbe28a20_33, RIbe2a6b8_94);
nand \U$25967 ( \26213 , \5055 , \26212 );
nand \U$25968 ( \26214 , \26211 , \26213 );
xor \U$25969 ( \26215 , \26208 , \26214 );
not \U$25970 ( \26216 , \25655 );
not \U$25971 ( \26217 , \8651 );
or \U$25972 ( \26218 , \26216 , \26217 );
xor \U$25973 ( \26219 , RIbe2adc0_109, RIbe28390_19);
nand \U$25974 ( \26220 , \8868 , \26219 );
nand \U$25975 ( \26221 , \26218 , \26220 );
xnor \U$25976 ( \26222 , \26215 , \26221 );
and \U$25977 ( \26223 , \26202 , \26222 );
not \U$25978 ( \26224 , \26202 );
not \U$25979 ( \26225 , \26222 );
and \U$25980 ( \26226 , \26224 , \26225 );
nor \U$25981 ( \26227 , \26223 , \26226 );
and \U$25982 ( \26228 , \26146 , \26227 );
not \U$25983 ( \26229 , \26146 );
not \U$25984 ( \26230 , \26227 );
and \U$25985 ( \26231 , \26229 , \26230 );
nor \U$25986 ( \26232 , \26228 , \26231 );
not \U$25987 ( \26233 , \26232 );
not \U$25988 ( \26234 , \26233 );
or \U$25989 ( \26235 , \26007 , \26234 );
nand \U$25990 ( \26236 , \26232 , \26005 );
nand \U$25991 ( \26237 , \26235 , \26236 );
not \U$25992 ( \26238 , \26237 );
not \U$25993 ( \26239 , \25457 );
not \U$25994 ( \26240 , \25451 );
or \U$25995 ( \26241 , \26239 , \26240 );
nand \U$25996 ( \26242 , \25450 , \25395 );
nand \U$25997 ( \26243 , \26241 , \26242 );
not \U$25998 ( \26244 , \26243 );
not \U$25999 ( \26245 , \26244 );
or \U$26000 ( \26246 , \26238 , \26245 );
or \U$26001 ( \26247 , \26244 , \26237 );
nand \U$26002 ( \26248 , \26246 , \26247 );
not \U$26003 ( \26249 , \26248 );
not \U$26004 ( \26250 , \26249 );
or \U$26005 ( \26251 , \25999 , \26250 );
not \U$26006 ( \26252 , \25998 );
nand \U$26007 ( \26253 , \26252 , \26248 );
nand \U$26008 ( \26254 , \26251 , \26253 );
and \U$26009 ( \26255 , \25861 , \26254 );
not \U$26010 ( \26256 , \25861 );
not \U$26011 ( \26257 , \26254 );
and \U$26012 ( \26258 , \26256 , \26257 );
nor \U$26013 ( \26259 , \26255 , \26258 );
xor \U$26014 ( \26260 , \25855 , \26259 );
not \U$26015 ( \26261 , \25781 );
not \U$26016 ( \26262 , \25775 );
not \U$26017 ( \26263 , \25551 );
or \U$26018 ( \26264 , \26262 , \26263 );
or \U$26019 ( \26265 , \25775 , \25551 );
nand \U$26020 ( \26266 , \26264 , \26265 );
not \U$26021 ( \26267 , \26266 );
or \U$26022 ( \26268 , \26261 , \26267 );
not \U$26023 ( \26269 , \25551 );
nand \U$26024 ( \26270 , \26269 , \25775 );
nand \U$26025 ( \26271 , \26268 , \26270 );
xor \U$26026 ( \26272 , \26260 , \26271 );
nand \U$26027 ( \26273 , \25811 , \26272 );
and \U$26028 ( \26274 , \25801 , \26273 );
nand \U$26029 ( \26275 , \25800 , \26274 );
not \U$26030 ( \26276 , \26275 );
and \U$26031 ( \26277 , \19163 , \26219 );
xor \U$26032 ( \26278 , RIbe2a460_89, RIbe28390_19);
and \U$26033 ( \26279 , \2776 , \26278 );
nor \U$26034 ( \26280 , \26277 , \26279 );
not \U$26035 ( \26281 , \26280 );
not \U$26036 ( \26282 , \26091 );
not \U$26037 ( \26283 , \2552 );
or \U$26038 ( \26284 , \26282 , \26283 );
xor \U$26039 ( \26285 , RIbe28b88_36, RIbe2ad48_108);
nand \U$26040 ( \26286 , \2558 , \26285 );
nand \U$26041 ( \26287 , \26284 , \26286 );
not \U$26042 ( \26288 , \26287 );
or \U$26043 ( \26289 , \26281 , \26288 );
or \U$26044 ( \26290 , \26287 , \26280 );
nand \U$26045 ( \26291 , \26289 , \26290 );
not \U$26046 ( \26292 , \19978 );
not \U$26047 ( \26293 , \26097 );
or \U$26048 ( \26294 , \26292 , \26293 );
xor \U$26049 ( \26295 , RIbe29e48_76, RIbe29ce0_73);
nand \U$26050 ( \26296 , \4850 , \26295 );
nand \U$26051 ( \26297 , \26294 , \26296 );
xor \U$26052 ( \26298 , \26291 , \26297 );
not \U$26053 ( \26299 , \26016 );
not \U$26054 ( \26300 , \8595 );
or \U$26055 ( \26301 , \26299 , \26300 );
xor \U$26056 ( \26302 , RIbe29c68_72, RIbe29ec0_77);
nand \U$26057 ( \26303 , \4580 , \26302 );
nand \U$26058 ( \26304 , \26301 , \26303 );
not \U$26059 ( \26305 , \26147 );
not \U$26060 ( \26306 , \23169 );
or \U$26061 ( \26307 , \26305 , \26306 );
xor \U$26062 ( \26308 , RIbe29308_52, RIbe2aaf0_103);
nand \U$26063 ( \26309 , \26308 , RIbe2ab68_104);
nand \U$26064 ( \26310 , \26307 , \26309 );
not \U$26065 ( \26311 , \26170 );
not \U$26066 ( \26312 , \10863 );
or \U$26067 ( \26313 , \26311 , \26312 );
xor \U$26068 ( \26314 , RIbe285e8_24, RIbe2a0a0_81);
nand \U$26069 ( \26315 , \2625 , \26314 );
nand \U$26070 ( \26316 , \26313 , \26315 );
xor \U$26071 ( \26317 , \26310 , \26316 );
xor \U$26072 ( \26318 , \26304 , \26317 );
xor \U$26073 ( \26319 , \26298 , \26318 );
not \U$26074 ( \26320 , \26121 );
not \U$26075 ( \26321 , \15353 );
or \U$26076 ( \26322 , \26320 , \26321 );
xor \U$26077 ( \26323 , RIbe282a0_17, RIbe2b180_117);
nand \U$26078 ( \26324 , \14966 , \26323 );
nand \U$26079 ( \26325 , \26322 , \26324 );
not \U$26080 ( \26326 , \26079 );
not \U$26081 ( \26327 , \2518 );
or \U$26082 ( \26328 , \26326 , \26327 );
xor \U$26083 ( \26329 , RIbe28480_21, RIbe2b2e8_120);
nand \U$26084 ( \26330 , \3074 , \26329 );
nand \U$26085 ( \26331 , \26328 , \26330 );
not \U$26086 ( \26332 , \26331 );
not \U$26087 ( \26333 , \26332 );
not \U$26088 ( \26334 , \26064 );
not \U$26089 ( \26335 , \8400 );
or \U$26090 ( \26336 , \26334 , \26335 );
xor \U$26091 ( \26337 , RIbe27b20_1, RIbe2a028_80);
nand \U$26092 ( \26338 , \8930 , \26337 );
nand \U$26093 ( \26339 , \26336 , \26338 );
not \U$26094 ( \26340 , \26339 );
or \U$26095 ( \26341 , \26333 , \26340 );
or \U$26096 ( \26342 , \26339 , \26332 );
nand \U$26097 ( \26343 , \26341 , \26342 );
xor \U$26098 ( \26344 , \26325 , \26343 );
and \U$26099 ( \26345 , \26319 , \26344 );
and \U$26100 ( \26346 , \26298 , \26318 );
or \U$26101 ( \26347 , \26345 , \26346 );
not \U$26102 ( \26348 , \26188 );
not \U$26103 ( \26349 , \2457 );
or \U$26104 ( \26350 , \26348 , \26349 );
xor \U$26105 ( \26351 , RIbe2a820_97, RIbe27e68_8);
nand \U$26106 ( \26352 , \2463 , \26351 );
nand \U$26107 ( \26353 , \26350 , \26352 );
not \U$26108 ( \26354 , \26353 );
not \U$26109 ( \26355 , \26354 );
not \U$26110 ( \26356 , \26071 );
not \U$26111 ( \26357 , \14296 );
or \U$26112 ( \26358 , \26356 , \26357 );
xor \U$26113 ( \26359 , RIbe297b8_62, RIbe2b108_116);
nand \U$26114 ( \26360 , \13533 , \26359 );
nand \U$26115 ( \26361 , \26358 , \26360 );
not \U$26116 ( \26362 , \26361 );
or \U$26117 ( \26363 , \26355 , \26362 );
or \U$26118 ( \26364 , \26361 , \26354 );
nand \U$26119 ( \26365 , \26363 , \26364 );
not \U$26120 ( \26366 , \26195 );
not \U$26121 ( \26367 , \879 );
or \U$26122 ( \26368 , \26366 , \26367 );
xor \U$26123 ( \26369 , RIbe28228_16, RIbe2abe0_105);
nand \U$26124 ( \26370 , \885 , \26369 );
nand \U$26125 ( \26371 , \26368 , \26370 );
and \U$26126 ( \26372 , \26365 , \26371 );
not \U$26127 ( \26373 , \26365 );
not \U$26128 ( \26374 , \26371 );
and \U$26129 ( \26375 , \26373 , \26374 );
nor \U$26130 ( \26376 , \26372 , \26375 );
not \U$26131 ( \26377 , \26376 );
not \U$26132 ( \26378 , \26127 );
not \U$26133 ( \26379 , \9082 );
or \U$26134 ( \26380 , \26378 , \26379 );
xor \U$26135 ( \26381 , RIbe27fd0_11, RIbe2aa00_101);
nand \U$26136 ( \26382 , \2707 , \26381 );
nand \U$26137 ( \26383 , \26380 , \26382 );
not \U$26138 ( \26384 , \26134 );
not \U$26139 ( \26385 , \9736 );
or \U$26140 ( \26386 , \26384 , \26385 );
xor \U$26141 ( \26387 , RIbe27df0_7, RIbe2a910_99);
nand \U$26142 ( \26388 , \9725 , \26387 );
nand \U$26143 ( \26389 , \26386 , \26388 );
xor \U$26144 ( \26390 , \26383 , \26389 );
not \U$26145 ( \26391 , \26105 );
not \U$26146 ( \26392 , \16913 );
or \U$26147 ( \26393 , \26391 , \26392 );
xor \U$26148 ( \26394 , RIbe2af28_112, RIbe294e8_56);
nand \U$26149 ( \26395 , \16728 , \26394 );
nand \U$26150 ( \26396 , \26393 , \26395 );
not \U$26151 ( \26397 , \26396 );
and \U$26152 ( \26398 , \26390 , \26397 );
not \U$26153 ( \26399 , \26390 );
and \U$26154 ( \26400 , \26399 , \26396 );
nor \U$26155 ( \26401 , \26398 , \26400 );
not \U$26156 ( \26402 , \26401 );
not \U$26157 ( \26403 , \26402 );
or \U$26158 ( \26404 , \26377 , \26403 );
or \U$26159 ( \26405 , \26402 , \26376 );
not \U$26160 ( \26406 , \26158 );
not \U$26161 ( \26407 , \23097 );
or \U$26162 ( \26408 , \26406 , \26407 );
xor \U$26163 ( \26409 , RIbe28f48_44, RIbe2b6a8_128);
nand \U$26164 ( \26410 , \4180 , \26409 );
nand \U$26165 ( \26411 , \26408 , \26410 );
not \U$26166 ( \26412 , \26411 );
not \U$26167 ( \26413 , \26412 );
not \U$26168 ( \26414 , \26206 );
not \U$26169 ( \26415 , \15991 );
not \U$26170 ( \26416 , \26415 );
or \U$26171 ( \26417 , \26414 , \26416 );
xor \U$26172 ( \26418 , RIbe29a10_67, RIbe2a550_91);
nand \U$26173 ( \26419 , \23306 , \26418 );
nand \U$26174 ( \26420 , \26417 , \26419 );
not \U$26175 ( \26421 , \26420 );
or \U$26176 ( \26422 , \26413 , \26421 );
or \U$26177 ( \26423 , \26420 , \26412 );
nand \U$26178 ( \26424 , \26422 , \26423 );
not \U$26179 ( \26425 , \26212 );
not \U$26180 ( \26426 , \1781 );
or \U$26181 ( \26427 , \26425 , \26426 );
xor \U$26182 ( \26428 , RIbe28a20_33, RIbe2b4c8_124);
nand \U$26183 ( \26429 , \5055 , \26428 );
nand \U$26184 ( \26430 , \26427 , \26429 );
and \U$26185 ( \26431 , \26424 , \26430 );
not \U$26186 ( \26432 , \26424 );
not \U$26187 ( \26433 , \26430 );
and \U$26188 ( \26434 , \26432 , \26433 );
nor \U$26189 ( \26435 , \26431 , \26434 );
nand \U$26190 ( \26436 , \26405 , \26435 );
nand \U$26191 ( \26437 , \26404 , \26436 );
buf \U$26192 ( \26438 , \26437 );
nor \U$26193 ( \26439 , \26347 , \26438 );
not \U$26194 ( \26440 , \25893 );
not \U$26195 ( \26441 , \19855 );
or \U$26196 ( \26442 , \26440 , \26441 );
xor \U$26197 ( \26443 , RIbe28a98_34, RIbe2b018_114);
nand \U$26198 ( \26444 , \15952 , \26443 );
nand \U$26199 ( \26445 , \26442 , \26444 );
not \U$26200 ( \26446 , \26022 );
not \U$26201 ( \26447 , \10831 );
or \U$26202 ( \26448 , \26446 , \26447 );
xor \U$26203 ( \26449 , RIbe29128_48, RIbe2a190_83);
nand \U$26204 ( \26450 , \10695 , \26449 );
nand \U$26205 ( \26451 , \26448 , \26450 );
xor \U$26206 ( \26452 , \26445 , \26451 );
not \U$26207 ( \26453 , \26029 );
not \U$26208 ( \26454 , \14827 );
or \U$26209 ( \26455 , \26453 , \26454 );
xor \U$26210 ( \26456 , RIbe298a8_64, RIbe2a2f8_86);
nand \U$26211 ( \26457 , \11094 , \26456 );
nand \U$26212 ( \26458 , \26455 , \26457 );
and \U$26213 ( \26459 , \26452 , \26458 );
and \U$26214 ( \26460 , \26445 , \26451 );
or \U$26215 ( \26461 , \26459 , \26460 );
not \U$26216 ( \26462 , \26297 );
not \U$26217 ( \26463 , \26291 );
or \U$26218 ( \26464 , \26462 , \26463 );
not \U$26219 ( \26465 , \26280 );
nand \U$26220 ( \26466 , \26465 , \26287 );
nand \U$26221 ( \26467 , \26464 , \26466 );
xor \U$26222 ( \26468 , \26461 , \26467 );
not \U$26223 ( \26469 , \26430 );
not \U$26224 ( \26470 , \26424 );
or \U$26225 ( \26471 , \26469 , \26470 );
nand \U$26226 ( \26472 , \26420 , \26411 );
nand \U$26227 ( \26473 , \26471 , \26472 );
and \U$26228 ( \26474 , \26468 , \26473 );
not \U$26229 ( \26475 , \26468 );
not \U$26230 ( \26476 , \26473 );
and \U$26231 ( \26477 , \26475 , \26476 );
nor \U$26232 ( \26478 , \26474 , \26477 );
not \U$26233 ( \26479 , \26478 );
or \U$26234 ( \26480 , \26439 , \26479 );
nand \U$26235 ( \26481 , \26347 , \26438 );
nand \U$26236 ( \26482 , \26480 , \26481 );
not \U$26237 ( \26483 , \26409 );
not \U$26238 ( \26484 , \12721 );
or \U$26239 ( \26485 , \26483 , \26484 );
xor \U$26240 ( \26486 , RIbe28f48_44, RIbe29f38_78);
nand \U$26241 ( \26487 , \9524 , \26486 );
nand \U$26242 ( \26488 , \26485 , \26487 );
not \U$26243 ( \26489 , \26488 );
not \U$26244 ( \26490 , \26449 );
not \U$26245 ( \26491 , \11396 );
or \U$26246 ( \26492 , \26490 , \26491 );
xor \U$26247 ( \26493 , RIbe291a0_49, RIbe2a190_83);
nand \U$26248 ( \26494 , \22918 , \26493 );
nand \U$26249 ( \26495 , \26492 , \26494 );
not \U$26250 ( \26496 , \26495 );
nand \U$26251 ( \26497 , \26489 , \26496 );
not \U$26252 ( \26498 , \26497 );
xor \U$26253 ( \26499 , RIbe2b3d8_122, RIbe296c8_60);
not \U$26254 ( \26500 , \26499 );
not \U$26255 ( \26501 , \8531 );
or \U$26256 ( \26502 , \26500 , \26501 );
xor \U$26257 ( \26503 , RIbe296c8_60, RIbe2b450_123);
nand \U$26258 ( \26504 , \907 , \26503 );
nand \U$26259 ( \26505 , \26502 , \26504 );
or \U$26260 ( \26506 , RIbe29650_59, RIbe296c8_60);
nand \U$26261 ( \26507 , \26506 , RIbe2ae38_110);
nand \U$26262 ( \26508 , RIbe29650_59, RIbe296c8_60);
and \U$26263 ( \26509 , \26507 , \26508 , RIbe29038_46);
nor \U$26264 ( \26510 , \26505 , \26509 );
not \U$26265 ( \26511 , \26510 );
nand \U$26266 ( \26512 , \26505 , \26509 );
nand \U$26267 ( \26513 , \26511 , \26512 );
not \U$26268 ( \26514 , \26513 );
not \U$26269 ( \26515 , \26514 );
or \U$26270 ( \26516 , \26498 , \26515 );
nand \U$26271 ( \26517 , \26488 , \26495 );
nand \U$26272 ( \26518 , \26516 , \26517 );
not \U$26273 ( \26519 , RIbe28cf0_39);
not \U$26274 ( \26520 , RIbe2a028_80);
and \U$26275 ( \26521 , \26519 , \26520 );
and \U$26276 ( \26522 , RIbe28cf0_39, RIbe2a028_80);
nor \U$26277 ( \26523 , \26521 , \26522 );
not \U$26278 ( \26524 , \26523 );
not \U$26279 ( \26525 , \9530 );
or \U$26280 ( \26526 , \26524 , \26525 );
xor \U$26281 ( \26527 , RIbe298a8_64, RIbe2a028_80);
nand \U$26282 ( \26528 , \8930 , \26527 );
nand \U$26283 ( \26529 , \26526 , \26528 );
xor \U$26284 ( \26530 , RIbe29b00_69, RIbe2a550_91);
not \U$26285 ( \26531 , \26530 );
not \U$26286 ( \26532 , \12000 );
or \U$26287 ( \26533 , \26531 , \26532 );
xor \U$26288 ( \26534 , RIbe29128_48, RIbe2a550_91);
nand \U$26289 ( \26535 , \12004 , \26534 );
nand \U$26290 ( \26536 , \26533 , \26535 );
nor \U$26291 ( \26537 , \26529 , \26536 );
not \U$26292 ( \26538 , \26537 );
nand \U$26293 ( \26539 , \26529 , \26536 );
nand \U$26294 ( \26540 , \26538 , \26539 );
not \U$26295 ( \26541 , \26486 );
nor \U$26296 ( \26542 , \26541 , \3257 );
xor \U$26297 ( \26543 , RIbe29ec0_77, RIbe28f48_44);
and \U$26298 ( \26544 , \9524 , \26543 );
nor \U$26299 ( \26545 , \26542 , \26544 );
not \U$26300 ( \26546 , \26545 );
and \U$26301 ( \26547 , \26540 , \26546 );
not \U$26302 ( \26548 , \26540 );
and \U$26303 ( \26549 , \26548 , \26545 );
nor \U$26304 ( \26550 , \26547 , \26549 );
and \U$26305 ( \26551 , \26518 , \26550 );
not \U$26306 ( \26552 , \26518 );
not \U$26307 ( \26553 , \26550 );
and \U$26308 ( \26554 , \26552 , \26553 );
or \U$26309 ( \26555 , \26551 , \26554 );
not \U$26310 ( \26556 , \26493 );
not \U$26311 ( \26557 , \15690 );
or \U$26312 ( \26558 , \26556 , \26557 );
xor \U$26313 ( \26559 , RIbe295d8_58, RIbe2a190_83);
nand \U$26314 ( \26560 , \11400 , \26559 );
nand \U$26315 ( \26561 , \26558 , \26560 );
not \U$26316 ( \26562 , \26561 );
not \U$26317 ( \26563 , \26512 );
or \U$26318 ( \26564 , \26562 , \26563 );
or \U$26319 ( \26565 , \26512 , \26561 );
nand \U$26320 ( \26566 , \26564 , \26565 );
not \U$26321 ( \26567 , \26566 );
xor \U$26322 ( \26568 , RIbe28d68_40, RIbe2a3e8_88);
not \U$26323 ( \26569 , \26568 );
not \U$26324 ( \26570 , \9262 );
or \U$26325 ( \26571 , \26569 , \26570 );
not \U$26326 ( \26572 , \8793 );
not \U$26327 ( \26573 , \26572 );
xor \U$26328 ( \26574 , RIbe27c88_4, RIbe2a3e8_88);
nand \U$26329 ( \26575 , \26573 , \26574 );
nand \U$26330 ( \26576 , \26571 , \26575 );
not \U$26331 ( \26577 , \26351 );
not \U$26332 ( \26578 , \2599 );
or \U$26333 ( \26579 , \26577 , \26578 );
xor \U$26334 ( \26580 , RIbe27e68_8, RIbe2a898_98);
nand \U$26335 ( \26581 , \2464 , \26580 );
nand \U$26336 ( \26582 , \26579 , \26581 );
xor \U$26337 ( \26583 , \26576 , \26582 );
not \U$26338 ( \26584 , \14296 );
not \U$26339 ( \26585 , \26359 );
or \U$26340 ( \26586 , \26584 , \26585 );
xnor \U$26341 ( \26587 , RIbe28138_14, RIbe2b108_116);
or \U$26342 ( \26588 , \16897 , \26587 );
nand \U$26343 ( \26589 , \26586 , \26588 );
and \U$26344 ( \26590 , \26583 , \26589 );
and \U$26345 ( \26591 , \26576 , \26582 );
or \U$26346 ( \26592 , \26590 , \26591 );
not \U$26347 ( \26593 , \26592 );
or \U$26348 ( \26594 , \26567 , \26593 );
or \U$26349 ( \26595 , \26592 , \26566 );
nand \U$26350 ( \26596 , \26594 , \26595 );
not \U$26351 ( \26597 , \26596 );
xor \U$26352 ( \26598 , \26555 , \26597 );
nor \U$26353 ( \26599 , \26482 , \26598 );
not \U$26354 ( \26600 , \26599 );
nand \U$26355 ( \26601 , \26482 , \26598 );
nand \U$26356 ( \26602 , \26600 , \26601 );
xor \U$26357 ( \26603 , \26445 , \26451 );
xor \U$26358 ( \26604 , \26603 , \26458 );
not \U$26359 ( \26605 , \26604 );
not \U$26360 ( \26606 , \26605 );
xor \U$26361 ( \26607 , RIbe28930_31, RIbe2a640_93);
and \U$26362 ( \26608 , \970 , \26607 );
not \U$26363 ( \26609 , \970 );
and \U$26364 ( \26610 , \961 , \26182 );
and \U$26365 ( \26611 , \26609 , \26610 );
nor \U$26366 ( \26612 , \26608 , \26611 );
not \U$26367 ( \26613 , \26612 );
not \U$26368 ( \26614 , \26055 );
not \U$26369 ( \26615 , \9793 );
or \U$26370 ( \26616 , \26614 , \26615 );
nand \U$26371 ( \26617 , \1937 , \26499 );
nand \U$26372 ( \26618 , \26616 , \26617 );
not \U$26373 ( \26619 , \26618 );
or \U$26374 ( \26620 , \26613 , \26619 );
or \U$26375 ( \26621 , \26618 , \26612 );
nand \U$26376 ( \26622 , \26620 , \26621 );
not \U$26377 ( \26623 , \26622 );
and \U$26378 ( \26624 , \8794 , \26568 );
not \U$26379 ( \26625 , \26047 );
nor \U$26380 ( \26626 , \26625 , \17059 );
nor \U$26381 ( \26627 , \26624 , \26626 );
not \U$26382 ( \26628 , \26627 );
and \U$26383 ( \26629 , \26623 , \26628 );
and \U$26384 ( \26630 , \26622 , \26627 );
nor \U$26385 ( \26631 , \26629 , \26630 );
not \U$26386 ( \26632 , \26631 );
or \U$26387 ( \26633 , \26606 , \26632 );
and \U$26388 ( \26634 , \1583 , RIbe2ae38_110);
not \U$26389 ( \26635 , \25881 );
not \U$26390 ( \26636 , \860 );
or \U$26391 ( \26637 , \26635 , \26636 );
xor \U$26392 ( \26638 , RIbe280c0_13, RIbe2a730_95);
nand \U$26393 ( \26639 , \1263 , \26638 );
nand \U$26394 ( \26640 , \26637 , \26639 );
xor \U$26395 ( \26641 , \26634 , \26640 );
not \U$26396 ( \26642 , \26041 );
not \U$26397 ( \26643 , \15793 );
or \U$26398 ( \26644 , \26642 , \26643 );
xor \U$26399 ( \26645 , RIbe295d8_58, RIbe2a280_85);
nand \U$26400 ( \26646 , \11348 , \26645 );
nand \U$26401 ( \26647 , \26644 , \26646 );
xor \U$26402 ( \26648 , \26641 , \26647 );
nand \U$26403 ( \26649 , \26633 , \26648 );
not \U$26404 ( \26650 , \26631 );
nand \U$26405 ( \26651 , \26650 , \26604 );
nand \U$26406 ( \26652 , \26649 , \26651 );
not \U$26407 ( \26653 , \26396 );
not \U$26408 ( \26654 , \26390 );
or \U$26409 ( \26655 , \26653 , \26654 );
nand \U$26410 ( \26656 , \26389 , \26383 );
nand \U$26411 ( \26657 , \26655 , \26656 );
not \U$26412 ( \26658 , \26657 );
not \U$26413 ( \26659 , \26371 );
not \U$26414 ( \26660 , \26365 );
or \U$26415 ( \26661 , \26659 , \26660 );
nand \U$26416 ( \26662 , \26361 , \26353 );
nand \U$26417 ( \26663 , \26661 , \26662 );
not \U$26418 ( \26664 , \26663 );
not \U$26419 ( \26665 , \26664 );
or \U$26420 ( \26666 , \26658 , \26665 );
not \U$26421 ( \26667 , \26657 );
nand \U$26422 ( \26668 , \26667 , \26663 );
nand \U$26423 ( \26669 , \26666 , \26668 );
not \U$26424 ( \26670 , \26325 );
not \U$26425 ( \26671 , \26343 );
or \U$26426 ( \26672 , \26670 , \26671 );
nand \U$26427 ( \26673 , \26339 , \26331 );
nand \U$26428 ( \26674 , \26672 , \26673 );
and \U$26429 ( \26675 , \26669 , \26674 );
not \U$26430 ( \26676 , \26669 );
not \U$26431 ( \26677 , \26674 );
and \U$26432 ( \26678 , \26676 , \26677 );
nor \U$26433 ( \26679 , \26675 , \26678 );
xor \U$26434 ( \26680 , \26652 , \26679 );
not \U$26435 ( \26681 , \26304 );
not \U$26436 ( \26682 , \26317 );
or \U$26437 ( \26683 , \26681 , \26682 );
nand \U$26438 ( \26684 , \26316 , \26310 );
nand \U$26439 ( \26685 , \26683 , \26684 );
xor \U$26440 ( \26686 , \26634 , \26640 );
and \U$26441 ( \26687 , \26686 , \26647 );
and \U$26442 ( \26688 , \26634 , \26640 );
or \U$26443 ( \26689 , \26687 , \26688 );
xor \U$26444 ( \26690 , \26685 , \26689 );
not \U$26445 ( \26691 , \26627 );
not \U$26446 ( \26692 , \26691 );
not \U$26447 ( \26693 , \26622 );
or \U$26448 ( \26694 , \26692 , \26693 );
not \U$26449 ( \26695 , \26612 );
nand \U$26450 ( \26696 , \26695 , \26618 );
nand \U$26451 ( \26697 , \26694 , \26696 );
and \U$26452 ( \26698 , \26690 , \26697 );
not \U$26453 ( \26699 , \26690 );
not \U$26454 ( \26700 , \26697 );
and \U$26455 ( \26701 , \26699 , \26700 );
nor \U$26456 ( \26702 , \26698 , \26701 );
and \U$26457 ( \26703 , \26680 , \26702 );
and \U$26458 ( \26704 , \26652 , \26679 );
or \U$26459 ( \26705 , \26703 , \26704 );
and \U$26460 ( \26706 , \26602 , \26705 );
not \U$26461 ( \26707 , \26602 );
not \U$26462 ( \26708 , \26705 );
and \U$26463 ( \26709 , \26707 , \26708 );
nor \U$26464 ( \26710 , \26706 , \26709 );
not \U$26465 ( \26711 , \26710 );
not \U$26466 ( \26712 , \26711 );
xor \U$26467 ( \26713 , \26652 , \26679 );
xor \U$26468 ( \26714 , \26713 , \26702 );
not \U$26469 ( \26715 , \26714 );
not \U$26470 ( \26716 , \26715 );
not \U$26471 ( \26717 , \26716 );
xor \U$26472 ( \26718 , \26437 , \26478 );
xnor \U$26473 ( \26719 , \26718 , \26347 );
not \U$26474 ( \26720 , \26719 );
not \U$26475 ( \26721 , \26720 );
or \U$26476 ( \26722 , \26717 , \26721 );
or \U$26477 ( \26723 , \26043 , \26049 );
nand \U$26478 ( \26724 , \26723 , \26057 );
nand \U$26479 ( \26725 , \26043 , \26049 );
nand \U$26480 ( \26726 , \26724 , \26725 );
xor \U$26481 ( \26727 , \26184 , \26190 );
and \U$26482 ( \26728 , \26727 , \26197 );
and \U$26483 ( \26729 , \26184 , \26190 );
or \U$26484 ( \26730 , \26728 , \26729 );
xor \U$26485 ( \26731 , \26726 , \26730 );
not \U$26486 ( \26732 , \26031 );
not \U$26487 ( \26733 , \26025 );
or \U$26488 ( \26734 , \26732 , \26733 );
nand \U$26489 ( \26735 , \26018 , \26024 );
nand \U$26490 ( \26736 , \26734 , \26735 );
xor \U$26491 ( \26737 , \26731 , \26736 );
not \U$26492 ( \26738 , \26137 );
not \U$26493 ( \26739 , \26117 );
or \U$26494 ( \26740 , \26738 , \26739 );
not \U$26495 ( \26741 , \26113 );
nand \U$26496 ( \26742 , \26741 , \26087 );
nand \U$26497 ( \26743 , \26740 , \26742 );
xor \U$26498 ( \26744 , \26737 , \26743 );
not \U$26499 ( \26745 , \26129 );
not \U$26500 ( \26746 , \26123 );
or \U$26501 ( \26747 , \26745 , \26746 );
or \U$26502 ( \26748 , \26123 , \26129 );
nand \U$26503 ( \26749 , \26748 , \26136 );
nand \U$26504 ( \26750 , \26747 , \26749 );
buf \U$26505 ( \26751 , \26750 );
not \U$26506 ( \26752 , \26093 );
not \U$26507 ( \26753 , \26752 );
not \U$26508 ( \26754 , \26111 );
or \U$26509 ( \26755 , \26753 , \26754 );
nand \U$26510 ( \26756 , \26107 , \26099 );
nand \U$26511 ( \26757 , \26755 , \26756 );
not \U$26512 ( \26758 , \26074 );
not \U$26513 ( \26759 , \26066 );
or \U$26514 ( \26760 , \26758 , \26759 );
or \U$26515 ( \26761 , \26066 , \26074 );
nand \U$26516 ( \26762 , \26761 , \26081 );
nand \U$26517 ( \26763 , \26760 , \26762 );
xnor \U$26518 ( \26764 , \26757 , \26763 );
not \U$26519 ( \26765 , \26764 );
xor \U$26520 ( \26766 , \26751 , \26765 );
and \U$26521 ( \26767 , \26744 , \26766 );
and \U$26522 ( \26768 , \26743 , \26737 );
nor \U$26523 ( \26769 , \26767 , \26768 );
not \U$26524 ( \26770 , \26769 );
nand \U$26525 ( \26771 , \26719 , \26715 );
nand \U$26526 ( \26772 , \26770 , \26771 );
nand \U$26527 ( \26773 , \26722 , \26772 );
not \U$26528 ( \26774 , \26773 );
not \U$26529 ( \26775 , \26774 );
or \U$26530 ( \26776 , \26712 , \26775 );
nand \U$26531 ( \26777 , \26773 , \26710 );
nand \U$26532 ( \26778 , \26776 , \26777 );
not \U$26533 ( \26779 , \26369 );
not \U$26534 ( \26780 , \3056 );
or \U$26535 ( \26781 , \26779 , \26780 );
xor \U$26536 ( \26782 , RIbe28228_16, RIbe2ac58_106);
nand \U$26537 ( \26783 , \26782 , \885 );
nand \U$26538 ( \26784 , \26781 , \26783 );
not \U$26539 ( \26785 , \26784 );
and \U$26540 ( \26786 , \26314 , \7618 );
xor \U$26541 ( \26787 , RIbe285e8_24, RIbe2a118_82);
and \U$26542 ( \26788 , \8270 , \26787 );
nor \U$26543 ( \26789 , \26786 , \26788 );
nand \U$26544 ( \26790 , \26785 , \26789 );
not \U$26545 ( \26791 , \26790 );
not \U$26546 ( \26792 , \26638 );
not \U$26547 ( \26793 , \2380 );
or \U$26548 ( \26794 , \26792 , \26793 );
xor \U$26549 ( \26795 , RIbe2a7a8_96, RIbe280c0_13);
nand \U$26550 ( \26796 , \869 , \26795 );
nand \U$26551 ( \26797 , \26794 , \26796 );
not \U$26552 ( \26798 , \26797 );
or \U$26553 ( \26799 , \26791 , \26798 );
not \U$26554 ( \26800 , \26789 );
nand \U$26555 ( \26801 , \26800 , \26784 );
nand \U$26556 ( \26802 , \26799 , \26801 );
not \U$26557 ( \26803 , \26456 );
not \U$26558 ( \26804 , \10446 );
or \U$26559 ( \26805 , \26803 , \26804 );
xor \U$26560 ( \26806 , RIbe29998_66, RIbe2a2f8_86);
nand \U$26561 ( \26807 , \9379 , \26806 );
nand \U$26562 ( \26808 , \26805 , \26807 );
not \U$26563 ( \26809 , \26808 );
not \U$26564 ( \26810 , \26302 );
not \U$26565 ( \26811 , \14971 );
or \U$26566 ( \26812 , \26810 , \26811 );
xor \U$26567 ( \26813 , RIbe29c68_72, RIbe29d58_74);
nand \U$26568 ( \26814 , \4580 , \26813 );
nand \U$26569 ( \26815 , \26812 , \26814 );
not \U$26570 ( \26816 , \26815 );
xor \U$26571 ( \26817 , RIbe29038_46, RIbe2ae38_110);
not \U$26572 ( \26818 , \26817 );
not \U$26573 ( \26819 , \16854 );
or \U$26574 ( \26820 , \26818 , \26819 );
xor \U$26575 ( \26821 , RIbe29038_46, RIbe2aeb0_111);
nand \U$26576 ( \26822 , \1583 , \26821 );
nand \U$26577 ( \26823 , \26820 , \26822 );
not \U$26578 ( \26824 , \26823 );
not \U$26579 ( \26825 , \26824 );
or \U$26580 ( \26826 , \26816 , \26825 );
or \U$26581 ( \26827 , \26824 , \26815 );
nand \U$26582 ( \26828 , \26826 , \26827 );
not \U$26583 ( \26829 , \26828 );
or \U$26584 ( \26830 , \26809 , \26829 );
nand \U$26585 ( \26831 , \26823 , \26815 );
nand \U$26586 ( \26832 , \26830 , \26831 );
xor \U$26587 ( \26833 , \26802 , \26832 );
not \U$26588 ( \26834 , \26337 );
not \U$26589 ( \26835 , \8170 );
or \U$26590 ( \26836 , \26834 , \26835 );
nand \U$26591 ( \26837 , \8172 , \26523 );
nand \U$26592 ( \26838 , \26836 , \26837 );
not \U$26593 ( \26839 , \26838 );
and \U$26594 ( \26840 , \19581 , \26308 );
xor \U$26595 ( \26841 , RIbe28c00_37, RIbe2aaf0_103);
and \U$26596 ( \26842 , \26841 , RIbe2ab68_104);
nor \U$26597 ( \26843 , \26840 , \26842 );
not \U$26598 ( \26844 , \26843 );
not \U$26599 ( \26845 , \26418 );
not \U$26600 ( \26846 , \10433 );
or \U$26601 ( \26847 , \26845 , \26846 );
nand \U$26602 ( \26848 , \23306 , \26530 );
nand \U$26603 ( \26849 , \26847 , \26848 );
not \U$26604 ( \26850 , \26849 );
or \U$26605 ( \26851 , \26844 , \26850 );
or \U$26606 ( \26852 , \26849 , \26843 );
nand \U$26607 ( \26853 , \26851 , \26852 );
not \U$26608 ( \26854 , \26853 );
or \U$26609 ( \26855 , \26839 , \26854 );
not \U$26610 ( \26856 , \26843 );
nand \U$26611 ( \26857 , \26856 , \26849 );
nand \U$26612 ( \26858 , \26855 , \26857 );
xor \U$26613 ( \26859 , \26833 , \26858 );
not \U$26614 ( \26860 , \26394 );
not \U$26615 ( \26861 , \15345 );
or \U$26616 ( \26862 , \26860 , \26861 );
not \U$26617 ( \26863 , RIbe288b8_30);
not \U$26618 ( \26864 , RIbe2af28_112);
and \U$26619 ( \26865 , \26863 , \26864 );
and \U$26620 ( \26866 , RIbe288b8_30, RIbe2af28_112);
nor \U$26621 ( \26867 , \26865 , \26866 );
nand \U$26622 ( \26868 , \17811 , \26867 );
nand \U$26623 ( \26869 , \26862 , \26868 );
not \U$26624 ( \26870 , \26869 );
not \U$26625 ( \26871 , \26323 );
not \U$26626 ( \26872 , \14852 );
or \U$26627 ( \26873 , \26871 , \26872 );
xor \U$26628 ( \26874 , RIbe29470_55, RIbe2b180_117);
nand \U$26629 ( \26875 , \16646 , \26874 );
nand \U$26630 ( \26876 , \26873 , \26875 );
not \U$26631 ( \26877 , \26876 );
not \U$26632 ( \26878 , \26428 );
not \U$26633 ( \26879 , \1780 );
or \U$26634 ( \26880 , \26878 , \26879 );
xnor \U$26635 ( \26881 , RIbe28a20_33, RIbe2b540_125);
not \U$26636 ( \26882 , \26881 );
nand \U$26637 ( \26883 , \26882 , \2475 );
nand \U$26638 ( \26884 , \26880 , \26883 );
not \U$26639 ( \26885 , \26884 );
not \U$26640 ( \26886 , \26885 );
or \U$26641 ( \26887 , \26877 , \26886 );
or \U$26642 ( \26888 , \26885 , \26876 );
nand \U$26643 ( \26889 , \26887 , \26888 );
not \U$26644 ( \26890 , \26889 );
or \U$26645 ( \26891 , \26870 , \26890 );
nand \U$26646 ( \26892 , \26884 , \26876 );
nand \U$26647 ( \26893 , \26891 , \26892 );
not \U$26648 ( \26894 , \26295 );
not \U$26649 ( \26895 , \9252 );
or \U$26650 ( \26896 , \26894 , \26895 );
and \U$26651 ( \26897 , RIbe29b78_70, RIbe29e48_76);
nor \U$26652 ( \26898 , RIbe29b78_70, RIbe29e48_76);
nor \U$26653 ( \26899 , \26897 , \26898 );
nand \U$26654 ( \26900 , \8245 , \26899 );
nand \U$26655 ( \26901 , \26896 , \26900 );
not \U$26656 ( \26902 , \26901 );
not \U$26657 ( \26903 , \26329 );
not \U$26658 ( \26904 , \2518 );
or \U$26659 ( \26905 , \26903 , \26904 );
and \U$26660 ( \26906 , RIbe28480_21, RIbe2b360_121);
not \U$26661 ( \26907 , RIbe28480_21);
not \U$26662 ( \26908 , RIbe2b360_121);
and \U$26663 ( \26909 , \26907 , \26908 );
nor \U$26664 ( \26910 , \26906 , \26909 );
nand \U$26665 ( \26911 , \16676 , \26910 );
nand \U$26666 ( \26912 , \26905 , \26911 );
not \U$26667 ( \26913 , \26381 );
not \U$26668 ( \26914 , \3377 );
or \U$26669 ( \26915 , \26913 , \26914 );
xor \U$26670 ( \26916 , RIbe27fd0_11, RIbe2aa78_102);
nand \U$26671 ( \26917 , \7709 , \26916 );
nand \U$26672 ( \26918 , \26915 , \26917 );
xor \U$26673 ( \26919 , \26912 , \26918 );
not \U$26674 ( \26920 , \26919 );
or \U$26675 ( \26921 , \26902 , \26920 );
nand \U$26676 ( \26922 , \26912 , \26918 );
nand \U$26677 ( \26923 , \26921 , \26922 );
not \U$26678 ( \26924 , \26923 );
and \U$26679 ( \26925 , \26893 , \26924 );
not \U$26680 ( \26926 , \26893 );
and \U$26681 ( \26927 , \26926 , \26923 );
nor \U$26682 ( \26928 , \26925 , \26927 );
not \U$26683 ( \26929 , \26285 );
not \U$26684 ( \26930 , \2552 );
or \U$26685 ( \26931 , \26929 , \26930 );
xor \U$26686 ( \26932 , RIbe28b88_36, RIbe2adc0_109);
nand \U$26687 ( \26933 , \7549 , \26932 );
nand \U$26688 ( \26934 , \26931 , \26933 );
not \U$26689 ( \26935 , \26934 );
not \U$26690 ( \26936 , \26935 );
not \U$26691 ( \26937 , \26387 );
not \U$26692 ( \26938 , \9737 );
or \U$26693 ( \26939 , \26937 , \26938 );
xor \U$26694 ( \26940 , RIbe29218_50, RIbe2a910_99);
nand \U$26695 ( \26941 , \9726 , \26940 );
nand \U$26696 ( \26942 , \26939 , \26941 );
buf \U$26697 ( \26943 , \26942 );
not \U$26698 ( \26944 , \26943 );
not \U$26699 ( \26945 , \26944 );
or \U$26700 ( \26946 , \26936 , \26945 );
not \U$26701 ( \26947 , \26607 );
not \U$26702 ( \26948 , \11374 );
or \U$26703 ( \26949 , \26947 , \26948 );
xor \U$26704 ( \26950 , RIbe28930_31, RIbe2a6b8_94);
nand \U$26705 ( \26951 , \1797 , \26950 );
nand \U$26706 ( \26952 , \26949 , \26951 );
nand \U$26707 ( \26953 , \26946 , \26952 );
nand \U$26708 ( \26954 , \26943 , \26934 );
nand \U$26709 ( \26955 , \26953 , \26954 );
buf \U$26710 ( \26956 , \26955 );
not \U$26711 ( \26957 , \26956 );
and \U$26712 ( \26958 , \26928 , \26957 );
not \U$26713 ( \26959 , \26928 );
and \U$26714 ( \26960 , \26959 , \26956 );
nor \U$26715 ( \26961 , \26958 , \26960 );
xor \U$26716 ( \26962 , \26859 , \26961 );
and \U$26717 ( \26963 , \26919 , \26901 );
not \U$26718 ( \26964 , \26919 );
not \U$26719 ( \26965 , \26901 );
and \U$26720 ( \26966 , \26964 , \26965 );
nor \U$26721 ( \26967 , \26963 , \26966 );
not \U$26722 ( \26968 , \26967 );
not \U$26723 ( \26969 , \26784 );
not \U$26724 ( \26970 , \26789 );
or \U$26725 ( \26971 , \26969 , \26970 );
or \U$26726 ( \26972 , \26784 , \26789 );
nand \U$26727 ( \26973 , \26971 , \26972 );
not \U$26728 ( \26974 , \26797 );
and \U$26729 ( \26975 , \26973 , \26974 );
not \U$26730 ( \26976 , \26973 );
and \U$26731 ( \26977 , \26976 , \26797 );
nor \U$26732 ( \26978 , \26975 , \26977 );
not \U$26733 ( \26979 , \26978 );
xor \U$26734 ( \26980 , \26838 , \26853 );
not \U$26735 ( \26981 , \26980 );
or \U$26736 ( \26982 , \26979 , \26981 );
or \U$26737 ( \26983 , \26980 , \26978 );
nand \U$26738 ( \26984 , \26982 , \26983 );
not \U$26739 ( \26985 , \26984 );
or \U$26740 ( \26986 , \26968 , \26985 );
not \U$26741 ( \26987 , \26978 );
nand \U$26742 ( \26988 , \26980 , \26987 );
nand \U$26743 ( \26989 , \26986 , \26988 );
not \U$26744 ( \26990 , \26989 );
and \U$26745 ( \26991 , \26962 , \26990 );
not \U$26746 ( \26992 , \26962 );
and \U$26747 ( \26993 , \26992 , \26989 );
nor \U$26748 ( \26994 , \26991 , \26993 );
not \U$26749 ( \26995 , \26994 );
not \U$26750 ( \26996 , \26669 );
not \U$26751 ( \26997 , \26674 );
or \U$26752 ( \26998 , \26996 , \26997 );
nand \U$26753 ( \26999 , \26663 , \26657 );
nand \U$26754 ( \27000 , \26998 , \26999 );
not \U$26755 ( \27001 , \27000 );
not \U$26756 ( \27002 , \26473 );
not \U$26757 ( \27003 , \26468 );
or \U$26758 ( \27004 , \27002 , \27003 );
nand \U$26759 ( \27005 , \26467 , \26461 );
nand \U$26760 ( \27006 , \27004 , \27005 );
not \U$26761 ( \27007 , \27006 );
not \U$26762 ( \27008 , \27007 );
or \U$26763 ( \27009 , \27001 , \27008 );
or \U$26764 ( \27010 , \27007 , \27000 );
nand \U$26765 ( \27011 , \27009 , \27010 );
not \U$26766 ( \27012 , \26697 );
not \U$26767 ( \27013 , \26690 );
or \U$26768 ( \27014 , \27012 , \27013 );
nand \U$26769 ( \27015 , \26685 , \26689 );
nand \U$26770 ( \27016 , \27014 , \27015 );
not \U$26771 ( \27017 , \27016 );
and \U$26772 ( \27018 , \27011 , \27017 );
not \U$26773 ( \27019 , \27011 );
and \U$26774 ( \27020 , \27019 , \27016 );
nor \U$26775 ( \27021 , \27018 , \27020 );
xor \U$26776 ( \27022 , \26576 , \26582 );
xor \U$26777 ( \27023 , \27022 , \26589 );
xor \U$26778 ( \27024 , \26808 , \26828 );
xor \U$26779 ( \27025 , \27023 , \27024 );
and \U$26780 ( \27026 , \26488 , \26495 );
not \U$26781 ( \27027 , \26488 );
and \U$26782 ( \27028 , \27027 , \26496 );
or \U$26783 ( \27029 , \27026 , \27028 );
xor \U$26784 ( \27030 , \27029 , \26513 );
xor \U$26785 ( \27031 , \27025 , \27030 );
not \U$26786 ( \27032 , \26443 );
not \U$26787 ( \27033 , \17570 );
or \U$26788 ( \27034 , \27032 , \27033 );
xor \U$26789 ( \27035 , RIbe293f8_54, RIbe2b018_114);
nand \U$26790 ( \27036 , \18777 , \27035 );
nand \U$26791 ( \27037 , \27034 , \27036 );
not \U$26792 ( \27038 , \26645 );
not \U$26793 ( \27039 , \20237 );
or \U$26794 ( \27040 , \27038 , \27039 );
xor \U$26795 ( \27041 , RIbe29740_61, RIbe2a280_85);
nand \U$26796 ( \27042 , \11348 , \27041 );
nand \U$26797 ( \27043 , \27040 , \27042 );
xor \U$26798 ( \27044 , \27037 , \27043 );
not \U$26799 ( \27045 , \26278 );
not \U$26800 ( \27046 , \2639 );
or \U$26801 ( \27047 , \27045 , \27046 );
xor \U$26802 ( \27048 , RIbe28390_19, RIbe2a4d8_90);
nand \U$26803 ( \27049 , \8654 , \27048 );
nand \U$26804 ( \27050 , \27047 , \27049 );
xor \U$26805 ( \27051 , \27044 , \27050 );
not \U$26806 ( \27052 , \27051 );
not \U$26807 ( \27053 , \27052 );
not \U$26808 ( \27054 , \26935 );
not \U$26809 ( \27055 , \26942 );
or \U$26810 ( \27056 , \27054 , \27055 );
or \U$26811 ( \27057 , \26942 , \26935 );
nand \U$26812 ( \27058 , \27056 , \27057 );
not \U$26813 ( \27059 , \27058 );
not \U$26814 ( \27060 , \26952 );
not \U$26815 ( \27061 , \27060 );
and \U$26816 ( \27062 , \27059 , \27061 );
and \U$26817 ( \27063 , \27058 , \27060 );
nor \U$26818 ( \27064 , \27062 , \27063 );
not \U$26819 ( \27065 , \27064 );
not \U$26820 ( \27066 , \27065 );
or \U$26821 ( \27067 , \27053 , \27066 );
nand \U$26822 ( \27068 , \27064 , \27051 );
nand \U$26823 ( \27069 , \27067 , \27068 );
and \U$26824 ( \27070 , \26889 , \26869 );
not \U$26825 ( \27071 , \26889 );
not \U$26826 ( \27072 , \26869 );
and \U$26827 ( \27073 , \27071 , \27072 );
nor \U$26828 ( \27074 , \27070 , \27073 );
and \U$26829 ( \27075 , \27069 , \27074 );
not \U$26830 ( \27076 , \27069 );
not \U$26831 ( \27077 , \27074 );
and \U$26832 ( \27078 , \27076 , \27077 );
nor \U$26833 ( \27079 , \27075 , \27078 );
xor \U$26834 ( \27080 , \27031 , \27079 );
xor \U$26835 ( \27081 , \26967 , \26987 );
xor \U$26836 ( \27082 , \27081 , \26980 );
and \U$26837 ( \27083 , \27080 , \27082 );
and \U$26838 ( \27084 , \27031 , \27079 );
or \U$26839 ( \27085 , \27083 , \27084 );
xnor \U$26840 ( \27086 , \27021 , \27085 );
not \U$26841 ( \27087 , \27086 );
or \U$26842 ( \27088 , \26995 , \27087 );
or \U$26843 ( \27089 , \27086 , \26994 );
nand \U$26844 ( \27090 , \27088 , \27089 );
not \U$26845 ( \27091 , \27090 );
and \U$26846 ( \27092 , \26778 , \27091 );
not \U$26847 ( \27093 , \26778 );
and \U$26848 ( \27094 , \27093 , \27090 );
nor \U$26849 ( \27095 , \27092 , \27094 );
not \U$26850 ( \27096 , \27095 );
not \U$26851 ( \27097 , \27064 );
or \U$26852 ( \27098 , \27051 , \27097 );
nand \U$26853 ( \27099 , \27098 , \27074 );
nand \U$26854 ( \27100 , \27097 , \27051 );
nand \U$26855 ( \27101 , \27099 , \27100 );
not \U$26856 ( \27102 , \26841 );
not \U$26857 ( \27103 , \18832 );
or \U$26858 ( \27104 , \27102 , \27103 );
xor \U$26859 ( \27105 , RIbe2aaf0_103, RIbe28c78_38);
nand \U$26860 ( \27106 , \27105 , RIbe2ab68_104);
nand \U$26861 ( \27107 , \27104 , \27106 );
not \U$26862 ( \27108 , \27107 );
not \U$26863 ( \27109 , \27108 );
not \U$26864 ( \27110 , \26910 );
not \U$26865 ( \27111 , \16953 );
or \U$26866 ( \27112 , \27110 , \27111 );
xor \U$26867 ( \27113 , RIbe28480_21, RIbe2a0a0_81);
nand \U$26868 ( \27114 , \27113 , \16676 );
nand \U$26869 ( \27115 , \27112 , \27114 );
not \U$26870 ( \27116 , \27115 );
or \U$26871 ( \27117 , \27109 , \27116 );
or \U$26872 ( \27118 , \27115 , \27108 );
nand \U$26873 ( \27119 , \27117 , \27118 );
not \U$26874 ( \27120 , \26899 );
not \U$26875 ( \27121 , \16652 );
or \U$26876 ( \27122 , \27120 , \27121 );
xor \U$26877 ( \27123 , RIbe29e48_76, RIbe27b20_1);
nand \U$26878 ( \27124 , \4851 , \27123 );
nand \U$26879 ( \27125 , \27122 , \27124 );
xor \U$26880 ( \27126 , \27119 , \27125 );
xor \U$26881 ( \27127 , \27037 , \27043 );
and \U$26882 ( \27128 , \27127 , \27050 );
and \U$26883 ( \27129 , \27037 , \27043 );
or \U$26884 ( \27130 , \27128 , \27129 );
xor \U$26885 ( \27131 , \27126 , \27130 );
not \U$26886 ( \27132 , \26821 );
not \U$26887 ( \27133 , \281 );
or \U$26888 ( \27134 , \27132 , \27133 );
xor \U$26889 ( \27135 , RIbe29038_46, RIbe2b3d8_122);
nand \U$26890 ( \27136 , \1583 , \27135 );
nand \U$26891 ( \27137 , \27134 , \27136 );
not \U$26892 ( \27138 , \26806 );
not \U$26893 ( \27139 , \16714 );
or \U$26894 ( \27140 , \27138 , \27139 );
xor \U$26895 ( \27141 , RIbe28d68_40, RIbe2a2f8_86);
nand \U$26896 ( \27142 , \8705 , \27141 );
nand \U$26897 ( \27143 , \27140 , \27142 );
and \U$26898 ( \27144 , \27137 , \27143 );
not \U$26899 ( \27145 , \27137 );
not \U$26900 ( \27146 , \27143 );
and \U$26901 ( \27147 , \27145 , \27146 );
nor \U$26902 ( \27148 , \27144 , \27147 );
not \U$26903 ( \27149 , \26782 );
not \U$26904 ( \27150 , \879 );
or \U$26905 ( \27151 , \27149 , \27150 );
xor \U$26906 ( \27152 , RIbe2a640_93, RIbe28228_16);
nand \U$26907 ( \27153 , \885 , \27152 );
nand \U$26908 ( \27154 , \27151 , \27153 );
xor \U$26909 ( \27155 , \27148 , \27154 );
xor \U$26910 ( \27156 , \27131 , \27155 );
xor \U$26911 ( \27157 , \27101 , \27156 );
not \U$26912 ( \27158 , \7794 );
not \U$26913 ( \27159 , \26881 );
and \U$26914 ( \27160 , \27158 , \27159 );
xor \U$26915 ( \27161 , RIbe28a20_33, RIbe2ad48_108);
and \U$26916 ( \27162 , \27161 , \5055 );
nor \U$26917 ( \27163 , \27160 , \27162 );
not \U$26918 ( \27164 , \27163 );
not \U$26919 ( \27165 , \26932 );
not \U$26920 ( \27166 , \3401 );
or \U$26921 ( \27167 , \27165 , \27166 );
xor \U$26922 ( \27168 , RIbe28b88_36, RIbe2a460_89);
nand \U$26923 ( \27169 , \2559 , \27168 );
nand \U$26924 ( \27170 , \27167 , \27169 );
not \U$26925 ( \27171 , \27170 );
or \U$26926 ( \27172 , \27164 , \27171 );
or \U$26927 ( \27173 , \27163 , \27170 );
nand \U$26928 ( \27174 , \27172 , \27173 );
not \U$26929 ( \27175 , \26867 );
not \U$26930 ( \27176 , \15345 );
or \U$26931 ( \27177 , \27175 , \27176 );
xor \U$26932 ( \27178 , RIbe2af28_112, RIbe28a98_34);
nand \U$26933 ( \27179 , \19721 , \27178 );
nand \U$26934 ( \27180 , \27177 , \27179 );
xor \U$26935 ( \27181 , \27174 , \27180 );
not \U$26936 ( \27182 , \27035 );
not \U$26937 ( \27183 , \16811 );
or \U$26938 ( \27184 , \27182 , \27183 );
xor \U$26939 ( \27185 , RIbe29308_52, RIbe2b018_114);
nand \U$26940 ( \27186 , \15953 , \27185 );
nand \U$26941 ( \27187 , \27184 , \27186 );
not \U$26942 ( \27188 , \26787 );
not \U$26943 ( \27189 , \8813 );
or \U$26944 ( \27190 , \27188 , \27189 );
xor \U$26945 ( \27191 , RIbe285e8_24, RIbe2a820_97);
nand \U$26946 ( \27192 , \2758 , \27191 );
nand \U$26947 ( \27193 , \27190 , \27192 );
and \U$26948 ( \27194 , \27187 , \27193 );
not \U$26949 ( \27195 , \27187 );
not \U$26950 ( \27196 , \27193 );
and \U$26951 ( \27197 , \27195 , \27196 );
nor \U$26952 ( \27198 , \27194 , \27197 );
not \U$26953 ( \27199 , \26795 );
not \U$26954 ( \27200 , \861 );
or \U$26955 ( \27201 , \27199 , \27200 );
xor \U$26956 ( \27202 , RIbe280c0_13, RIbe2abe0_105);
nand \U$26957 ( \27203 , \869 , \27202 );
nand \U$26958 ( \27204 , \27201 , \27203 );
xnor \U$26959 ( \27205 , \27198 , \27204 );
not \U$26960 ( \27206 , \27205 );
xor \U$26961 ( \27207 , \27181 , \27206 );
not \U$26962 ( \27208 , \11768 );
not \U$26963 ( \27209 , \26916 );
not \U$26964 ( \27210 , \27209 );
and \U$26965 ( \27211 , \27208 , \27210 );
xor \U$26966 ( \27212 , RIbe2b6a8_128, RIbe27fd0_11);
and \U$26967 ( \27213 , \2707 , \27212 );
nor \U$26968 ( \27214 , \27211 , \27213 );
not \U$26969 ( \27215 , \26940 );
not \U$26970 ( \27216 , \10987 );
or \U$26971 ( \27217 , \27215 , \27216 );
xor \U$26972 ( \27218 , RIbe29a10_67, RIbe2a910_99);
nand \U$26973 ( \27219 , \11456 , \27218 );
nand \U$26974 ( \27220 , \27217 , \27219 );
not \U$26975 ( \27221 , \27220 );
not \U$26976 ( \27222 , \26950 );
not \U$26977 ( \27223 , \965 );
or \U$26978 ( \27224 , \27222 , \27223 );
xor \U$26979 ( \27225 , RIbe28930_31, RIbe2b4c8_124);
nand \U$26980 ( \27226 , \1797 , \27225 );
nand \U$26981 ( \27227 , \27224 , \27226 );
not \U$26982 ( \27228 , \27227 );
not \U$26983 ( \27229 , \27228 );
or \U$26984 ( \27230 , \27221 , \27229 );
or \U$26985 ( \27231 , \27220 , \27228 );
nand \U$26986 ( \27232 , \27230 , \27231 );
not \U$26987 ( \27233 , \27232 );
xor \U$26988 ( \27234 , \27214 , \27233 );
buf \U$26989 ( \27235 , \27234 );
xor \U$26990 ( \27236 , \27207 , \27235 );
xnor \U$26991 ( \27237 , \27157 , \27236 );
not \U$26992 ( \27238 , \27237 );
not \U$26993 ( \27239 , \27238 );
not \U$26994 ( \27240 , \25889 );
not \U$26995 ( \27241 , \26208 );
not \U$26996 ( \27242 , \26214 );
or \U$26997 ( \27243 , \27241 , \27242 );
or \U$26998 ( \27244 , \26214 , \26208 );
nand \U$26999 ( \27245 , \27244 , \26221 );
nand \U$27000 ( \27246 , \27243 , \27245 );
xor \U$27001 ( \27247 , \27240 , \27246 );
not \U$27002 ( \27248 , \26172 );
not \U$27003 ( \27249 , \26166 );
or \U$27004 ( \27250 , \27248 , \27249 );
nand \U$27005 ( \27251 , \26160 , \26153 );
nand \U$27006 ( \27252 , \27250 , \27251 );
and \U$27007 ( \27253 , \27247 , \27252 );
and \U$27008 ( \27254 , \27240 , \27246 );
or \U$27009 ( \27255 , \27253 , \27254 );
or \U$27010 ( \27256 , \26750 , \26763 );
nand \U$27011 ( \27257 , \27256 , \26757 );
nand \U$27012 ( \27258 , \26751 , \26763 );
nand \U$27013 ( \27259 , \27257 , \27258 );
nor \U$27014 ( \27260 , \27255 , \27259 );
xor \U$27015 ( \27261 , \26726 , \26730 );
and \U$27016 ( \27262 , \27261 , \26736 );
and \U$27017 ( \27263 , \26726 , \26730 );
or \U$27018 ( \27264 , \27262 , \27263 );
not \U$27019 ( \27265 , \27264 );
or \U$27020 ( \27266 , \27260 , \27265 );
nand \U$27021 ( \27267 , \27255 , \27259 );
nand \U$27022 ( \27268 , \27266 , \27267 );
not \U$27023 ( \27269 , \27268 );
not \U$27024 ( \27270 , \27041 );
not \U$27025 ( \27271 , \10845 );
or \U$27026 ( \27272 , \27270 , \27271 );
xor \U$27027 ( \27273 , RIbe297b8_62, RIbe2a280_85);
nand \U$27028 ( \27274 , \18667 , \27273 );
nand \U$27029 ( \27275 , \27272 , \27274 );
or \U$27030 ( \27276 , \13528 , \26587 );
xor \U$27031 ( \27277 , RIbe282a0_17, RIbe2b108_116);
not \U$27032 ( \27278 , \27277 );
or \U$27033 ( \27279 , \19967 , \27278 );
nand \U$27034 ( \27280 , \27276 , \27279 );
xor \U$27035 ( \27281 , \27275 , \27280 );
not \U$27036 ( \27282 , \27048 );
not \U$27037 ( \27283 , \8651 );
or \U$27038 ( \27284 , \27282 , \27283 );
xor \U$27039 ( \27285 , RIbe28390_19, RIbe2b2e8_120);
nand \U$27040 ( \27286 , \8868 , \27285 );
nand \U$27041 ( \27287 , \27284 , \27286 );
not \U$27042 ( \27288 , \27287 );
and \U$27043 ( \27289 , \27281 , \27288 );
not \U$27044 ( \27290 , \27281 );
and \U$27045 ( \27291 , \27290 , \27287 );
nor \U$27046 ( \27292 , \27289 , \27291 );
not \U$27047 ( \27293 , \27292 );
and \U$27048 ( \27294 , \26874 , \17592 );
xor \U$27049 ( \27295 , RIbe294e8_56, RIbe2b180_117);
and \U$27050 ( \27296 , \16646 , \27295 );
nor \U$27051 ( \27297 , \27294 , \27296 );
not \U$27052 ( \27298 , \26574 );
not \U$27053 ( \27299 , \9262 );
or \U$27054 ( \27300 , \27298 , \27299 );
xor \U$27055 ( \27301 , RIbe27df0_7, RIbe2a3e8_88);
nand \U$27056 ( \27302 , \8793 , \27301 );
nand \U$27057 ( \27303 , \27300 , \27302 );
not \U$27058 ( \27304 , \27303 );
and \U$27059 ( \27305 , \27297 , \27304 );
not \U$27060 ( \27306 , \27297 );
and \U$27061 ( \27307 , \27306 , \27303 );
nor \U$27062 ( \27308 , \27305 , \27307 );
not \U$27063 ( \27309 , \26580 );
not \U$27064 ( \27310 , \2458 );
or \U$27065 ( \27311 , \27309 , \27310 );
xor \U$27066 ( \27312 , RIbe2aa00_101, RIbe27e68_8);
nand \U$27067 ( \27313 , \2464 , \27312 );
nand \U$27068 ( \27314 , \27311 , \27313 );
not \U$27069 ( \27315 , \27314 );
and \U$27070 ( \27316 , \27308 , \27315 );
not \U$27071 ( \27317 , \27308 );
and \U$27072 ( \27318 , \27317 , \27314 );
nor \U$27073 ( \27319 , \27316 , \27318 );
not \U$27074 ( \27320 , \27319 );
nand \U$27075 ( \27321 , \27293 , \27320 );
nand \U$27076 ( \27322 , \27292 , \27319 );
nand \U$27077 ( \27323 , \27321 , \27322 );
nor \U$27078 ( \27324 , \468 , \24871 );
not \U$27079 ( \27325 , \26503 );
not \U$27080 ( \27326 , \1129 );
or \U$27081 ( \27327 , \27325 , \27326 );
xor \U$27082 ( \27328 , RIbe2a730_95, RIbe296c8_60);
nand \U$27083 ( \27329 , \907 , \27328 );
nand \U$27084 ( \27330 , \27327 , \27329 );
xor \U$27085 ( \27331 , \27324 , \27330 );
not \U$27086 ( \27332 , \10720 );
not \U$27087 ( \27333 , \26813 );
or \U$27088 ( \27334 , \27332 , \27333 );
xor \U$27089 ( \27335 , RIbe29c68_72, RIbe29ce0_73);
not \U$27090 ( \27336 , \27335 );
or \U$27091 ( \27337 , \4581 , \27336 );
nand \U$27092 ( \27338 , \27334 , \27337 );
xor \U$27093 ( \27339 , \27331 , \27338 );
xor \U$27094 ( \27340 , \27323 , \27339 );
not \U$27095 ( \27341 , \27340 );
xor \U$27096 ( \27342 , \27023 , \27024 );
and \U$27097 ( \27343 , \27342 , \27030 );
and \U$27098 ( \27344 , \27023 , \27024 );
or \U$27099 ( \27345 , \27343 , \27344 );
not \U$27100 ( \27346 , \27345 );
and \U$27101 ( \27347 , \27341 , \27346 );
and \U$27102 ( \27348 , \27345 , \27340 );
nor \U$27103 ( \27349 , \27347 , \27348 );
not \U$27104 ( \27350 , \27349 );
or \U$27105 ( \27351 , \27269 , \27350 );
or \U$27106 ( \27352 , \27349 , \27268 );
nand \U$27107 ( \27353 , \27351 , \27352 );
not \U$27108 ( \27354 , \27353 );
not \U$27109 ( \27355 , \27354 );
or \U$27110 ( \27356 , \27239 , \27355 );
nand \U$27111 ( \27357 , \27353 , \27237 );
nand \U$27112 ( \27358 , \27356 , \27357 );
not \U$27113 ( \27359 , \27265 );
not \U$27114 ( \27360 , \27260 );
nand \U$27115 ( \27361 , \27360 , \27267 );
not \U$27116 ( \27362 , \27361 );
or \U$27117 ( \27363 , \27359 , \27362 );
or \U$27118 ( \27364 , \27361 , \27265 );
nand \U$27119 ( \27365 , \27363 , \27364 );
not \U$27120 ( \27366 , \25921 );
not \U$27121 ( \27367 , \25942 );
or \U$27122 ( \27368 , \27366 , \27367 );
nand \U$27123 ( \27369 , \25937 , \25929 );
nand \U$27124 ( \27370 , \27368 , \27369 );
not \U$27125 ( \27371 , \27370 );
not \U$27126 ( \27372 , \25901 );
not \U$27127 ( \27373 , \25908 );
or \U$27128 ( \27374 , \27372 , \27373 );
nand \U$27129 ( \27375 , \27374 , \25900 );
not \U$27130 ( \27376 , \27375 );
not \U$27131 ( \27377 , \27376 );
or \U$27132 ( \27378 , \25967 , \25958 );
not \U$27133 ( \27379 , \27378 );
not \U$27134 ( \27380 , \25962 );
or \U$27135 ( \27381 , \27379 , \27380 );
nand \U$27136 ( \27382 , \25967 , \25958 );
nand \U$27137 ( \27383 , \27381 , \27382 );
not \U$27138 ( \27384 , \27383 );
or \U$27139 ( \27385 , \27377 , \27384 );
or \U$27140 ( \27386 , \27383 , \27376 );
nand \U$27141 ( \27387 , \27385 , \27386 );
not \U$27142 ( \27388 , \27387 );
or \U$27143 ( \27389 , \27371 , \27388 );
nand \U$27144 ( \27390 , \27383 , \27375 );
nand \U$27145 ( \27391 , \27389 , \27390 );
not \U$27146 ( \27392 , \26225 );
not \U$27147 ( \27393 , \26177 );
not \U$27148 ( \27394 , \27393 );
or \U$27149 ( \27395 , \27392 , \27394 );
not \U$27150 ( \27396 , \26222 );
not \U$27151 ( \27397 , \26177 );
or \U$27152 ( \27398 , \27396 , \27397 );
nand \U$27153 ( \27399 , \27398 , \26198 );
nand \U$27154 ( \27400 , \27395 , \27399 );
xor \U$27155 ( \27401 , \27240 , \27246 );
xor \U$27156 ( \27402 , \27401 , \27252 );
nor \U$27157 ( \27403 , \27400 , \27402 );
xor \U$27158 ( \27404 , \26012 , \26036 );
and \U$27159 ( \27405 , \27404 , \26058 );
and \U$27160 ( \27406 , \26012 , \26036 );
or \U$27161 ( \27407 , \27405 , \27406 );
not \U$27162 ( \27408 , \27407 );
or \U$27163 ( \27409 , \27403 , \27408 );
nand \U$27164 ( \27410 , \27400 , \27402 );
nand \U$27165 ( \27411 , \27409 , \27410 );
nor \U$27166 ( \27412 , \27391 , \27411 );
or \U$27167 ( \27413 , \27365 , \27412 );
nand \U$27168 ( \27414 , \27391 , \27411 );
nand \U$27169 ( \27415 , \27413 , \27414 );
not \U$27170 ( \27416 , \27415 );
and \U$27171 ( \27417 , \27358 , \27416 );
not \U$27172 ( \27418 , \27358 );
and \U$27173 ( \27419 , \27418 , \27415 );
nor \U$27174 ( \27420 , \27417 , \27419 );
not \U$27175 ( \27421 , \27420 );
not \U$27176 ( \27422 , \27421 );
xor \U$27177 ( \27423 , \27031 , \27079 );
xor \U$27178 ( \27424 , \27423 , \27082 );
xor \U$27179 ( \27425 , \26298 , \26318 );
xor \U$27180 ( \27426 , \27425 , \26344 );
not \U$27181 ( \27427 , \27426 );
not \U$27182 ( \27428 , \26376 );
not \U$27183 ( \27429 , \27428 );
not \U$27184 ( \27430 , \26402 );
or \U$27185 ( \27431 , \27429 , \27430 );
nand \U$27186 ( \27432 , \26401 , \26376 );
nand \U$27187 ( \27433 , \27431 , \27432 );
and \U$27188 ( \27434 , \27433 , \26435 );
not \U$27189 ( \27435 , \27433 );
not \U$27190 ( \27436 , \26435 );
and \U$27191 ( \27437 , \27435 , \27436 );
nor \U$27192 ( \27438 , \27434 , \27437 );
not \U$27193 ( \27439 , \27438 );
not \U$27194 ( \27440 , \27439 );
xor \U$27195 ( \27441 , \26604 , \26650 );
xnor \U$27196 ( \27442 , \27441 , \26648 );
not \U$27197 ( \27443 , \27442 );
not \U$27198 ( \27444 , \27443 );
or \U$27199 ( \27445 , \27440 , \27444 );
nand \U$27200 ( \27446 , \27442 , \27438 );
nand \U$27201 ( \27447 , \27445 , \27446 );
not \U$27202 ( \27448 , \27447 );
or \U$27203 ( \27449 , \27427 , \27448 );
nand \U$27204 ( \27450 , \27443 , \27438 );
nand \U$27205 ( \27451 , \27449 , \27450 );
and \U$27206 ( \27452 , \27424 , \27451 );
not \U$27207 ( \27453 , \27424 );
not \U$27208 ( \27454 , \27451 );
and \U$27209 ( \27455 , \27453 , \27454 );
nor \U$27210 ( \27456 , \27452 , \27455 );
not \U$27211 ( \27457 , \25910 );
not \U$27212 ( \27458 , \25877 );
or \U$27213 ( \27459 , \27457 , \27458 );
not \U$27214 ( \27460 , \25868 );
nand \U$27215 ( \27461 , \27460 , \25873 );
nand \U$27216 ( \27462 , \27459 , \27461 );
xor \U$27217 ( \27463 , \27387 , \27370 );
nand \U$27218 ( \27464 , \27462 , \27463 );
not \U$27219 ( \27465 , \25943 );
not \U$27220 ( \27466 , \25953 );
nand \U$27221 ( \27467 , \27466 , \25968 );
not \U$27222 ( \27468 , \27467 );
or \U$27223 ( \27469 , \27465 , \27468 );
not \U$27224 ( \27470 , \25968 );
nand \U$27225 ( \27471 , \27470 , \25953 );
nand \U$27226 ( \27472 , \27469 , \27471 );
nand \U$27227 ( \27473 , \27463 , \27472 );
nand \U$27228 ( \27474 , \27462 , \27472 );
nand \U$27229 ( \27475 , \27464 , \27473 , \27474 );
nand \U$27230 ( \27476 , \27456 , \27475 );
nand \U$27231 ( \27477 , \27424 , \27451 );
and \U$27232 ( \27478 , \27476 , \27477 );
not \U$27233 ( \27479 , \27478 );
or \U$27234 ( \27480 , \27422 , \27479 );
not \U$27235 ( \27481 , \27477 );
not \U$27236 ( \27482 , \27476 );
or \U$27237 ( \27483 , \27481 , \27482 );
nand \U$27238 ( \27484 , \27483 , \27420 );
nand \U$27239 ( \27485 , \27480 , \27484 );
not \U$27240 ( \27486 , \27412 );
nand \U$27241 ( \27487 , \27486 , \27414 );
not \U$27242 ( \27488 , \27365 );
and \U$27243 ( \27489 , \27487 , \27488 );
not \U$27244 ( \27490 , \27487 );
and \U$27245 ( \27491 , \27490 , \27365 );
nor \U$27246 ( \27492 , \27489 , \27491 );
not \U$27247 ( \27493 , \27492 );
not \U$27248 ( \27494 , \27493 );
not \U$27249 ( \27495 , \26714 );
not \U$27250 ( \27496 , \26719 );
or \U$27251 ( \27497 , \27495 , \27496 );
or \U$27252 ( \27498 , \26719 , \26714 );
nand \U$27253 ( \27499 , \27497 , \27498 );
xor \U$27254 ( \27500 , \27499 , \26769 );
not \U$27255 ( \27501 , \27500 );
not \U$27256 ( \27502 , \27501 );
or \U$27257 ( \27503 , \27494 , \27502 );
not \U$27258 ( \27504 , \27492 );
not \U$27259 ( \27505 , \27500 );
or \U$27260 ( \27506 , \27504 , \27505 );
not \U$27261 ( \27507 , \26059 );
not \U$27262 ( \27508 , \26230 );
or \U$27263 ( \27509 , \27507 , \27508 );
not \U$27264 ( \27510 , \26142 );
not \U$27265 ( \27511 , \26059 );
nand \U$27266 ( \27512 , \26227 , \27511 );
nand \U$27267 ( \27513 , \27510 , \27512 );
nand \U$27268 ( \27514 , \27509 , \27513 );
not \U$27269 ( \27515 , \25985 );
xor \U$27270 ( \27516 , \25989 , \25996 );
not \U$27271 ( \27517 , \27516 );
or \U$27272 ( \27518 , \27515 , \27517 );
nand \U$27273 ( \27519 , \25996 , \25989 );
nand \U$27274 ( \27520 , \27518 , \27519 );
and \U$27275 ( \27521 , \27514 , \27520 );
not \U$27276 ( \27522 , \27514 );
not \U$27277 ( \27523 , \27520 );
and \U$27278 ( \27524 , \27522 , \27523 );
nor \U$27279 ( \27525 , \27521 , \27524 );
not \U$27280 ( \27526 , \27525 );
xor \U$27281 ( \27527 , \26744 , \26766 );
not \U$27282 ( \27528 , \27527 );
or \U$27283 ( \27529 , \27526 , \27528 );
nand \U$27284 ( \27530 , \27520 , \27514 );
nand \U$27285 ( \27531 , \27529 , \27530 );
nand \U$27286 ( \27532 , \27506 , \27531 );
nand \U$27287 ( \27533 , \27503 , \27532 );
and \U$27288 ( \27534 , \27485 , \27533 );
not \U$27289 ( \27535 , \27485 );
not \U$27290 ( \27536 , \27533 );
and \U$27291 ( \27537 , \27535 , \27536 );
nor \U$27292 ( \27538 , \27534 , \27537 );
not \U$27293 ( \27539 , \27538 );
or \U$27294 ( \27540 , \27096 , \27539 );
or \U$27295 ( \27541 , \27095 , \27538 );
nand \U$27296 ( \27542 , \27540 , \27541 );
not \U$27297 ( \27543 , \27542 );
xor \U$27298 ( \27544 , \27525 , \27527 );
not \U$27299 ( \27545 , \27544 );
xor \U$27300 ( \27546 , \27472 , \27462 );
buf \U$27301 ( \27547 , \27463 );
not \U$27302 ( \27548 , \27547 );
and \U$27303 ( \27549 , \27546 , \27548 );
not \U$27304 ( \27550 , \27546 );
and \U$27305 ( \27551 , \27550 , \27547 );
nor \U$27306 ( \27552 , \27549 , \27551 );
not \U$27307 ( \27553 , \27552 );
xor \U$27308 ( \27554 , \25915 , \25976 );
and \U$27309 ( \27555 , \27554 , \25997 );
and \U$27310 ( \27556 , \25915 , \25976 );
or \U$27311 ( \27557 , \27555 , \27556 );
not \U$27312 ( \27558 , \27557 );
or \U$27313 ( \27559 , \27553 , \27558 );
or \U$27314 ( \27560 , \27557 , \27552 );
nand \U$27315 ( \27561 , \27559 , \27560 );
not \U$27316 ( \27562 , \27561 );
or \U$27317 ( \27563 , \27545 , \27562 );
not \U$27318 ( \27564 , \27552 );
nand \U$27319 ( \27565 , \27564 , \27557 );
nand \U$27320 ( \27566 , \27563 , \27565 );
not \U$27321 ( \27567 , \27566 );
buf \U$27322 ( \27568 , \27456 );
buf \U$27323 ( \27569 , \27475 );
not \U$27324 ( \27570 , \27569 );
and \U$27325 ( \27571 , \27568 , \27570 );
not \U$27326 ( \27572 , \27568 );
and \U$27327 ( \27573 , \27572 , \27569 );
nor \U$27328 ( \27574 , \27571 , \27573 );
not \U$27329 ( \27575 , \27574 );
not \U$27330 ( \27576 , \25828 );
not \U$27331 ( \27577 , \25834 );
or \U$27332 ( \27578 , \27576 , \27577 );
nand \U$27333 ( \27579 , \25827 , \25823 );
nand \U$27334 ( \27580 , \27578 , \27579 );
not \U$27335 ( \27581 , \27580 );
xor \U$27336 ( \27582 , \27402 , \27407 );
xor \U$27337 ( \27583 , \27582 , \27400 );
and \U$27338 ( \27584 , \27447 , \27426 );
not \U$27339 ( \27585 , \27447 );
not \U$27340 ( \27586 , \27426 );
and \U$27341 ( \27587 , \27585 , \27586 );
nor \U$27342 ( \27588 , \27584 , \27587 );
xnor \U$27343 ( \27589 , \27583 , \27588 );
not \U$27344 ( \27590 , \27589 );
not \U$27345 ( \27591 , \27590 );
or \U$27346 ( \27592 , \27581 , \27591 );
nand \U$27347 ( \27593 , \27588 , \27583 );
nand \U$27348 ( \27594 , \27592 , \27593 );
not \U$27349 ( \27595 , \27594 );
and \U$27350 ( \27596 , \27575 , \27595 );
and \U$27351 ( \27597 , \27594 , \27574 );
nor \U$27352 ( \27598 , \27596 , \27597 );
not \U$27353 ( \27599 , \27598 );
not \U$27354 ( \27600 , \27599 );
or \U$27355 ( \27601 , \27567 , \27600 );
not \U$27356 ( \27602 , \27574 );
nand \U$27357 ( \27603 , \27602 , \27594 );
nand \U$27358 ( \27604 , \27601 , \27603 );
not \U$27359 ( \27605 , \27604 );
not \U$27360 ( \27606 , \27605 );
and \U$27361 ( \27607 , \27543 , \27606 );
and \U$27362 ( \27608 , \27542 , \27605 );
nor \U$27363 ( \27609 , \27607 , \27608 );
xor \U$27364 ( \27610 , \27531 , \27493 );
and \U$27365 ( \27611 , \27610 , \27501 );
not \U$27366 ( \27612 , \27610 );
and \U$27367 ( \27613 , \27612 , \27500 );
nor \U$27368 ( \27614 , \27611 , \27613 );
not \U$27369 ( \27615 , \27614 );
not \U$27370 ( \27616 , \26243 );
not \U$27371 ( \27617 , \26237 );
or \U$27372 ( \27618 , \27616 , \27617 );
nand \U$27373 ( \27619 , \26233 , \26005 );
nand \U$27374 ( \27620 , \27618 , \27619 );
not \U$27375 ( \27621 , \27620 );
not \U$27376 ( \27622 , \27621 );
or \U$27377 ( \27623 , \27580 , \27589 );
nand \U$27378 ( \27624 , \27580 , \27589 );
nand \U$27379 ( \27625 , \27623 , \27624 );
not \U$27380 ( \27626 , \27625 );
or \U$27381 ( \27627 , \27622 , \27626 );
or \U$27382 ( \27628 , \27621 , \27625 );
nand \U$27383 ( \27629 , \27627 , \27628 );
not \U$27384 ( \27630 , \25854 );
not \U$27385 ( \27631 , \25843 );
or \U$27386 ( \27632 , \27630 , \27631 );
not \U$27387 ( \27633 , \25839 );
nand \U$27388 ( \27634 , \27633 , \25817 );
nand \U$27389 ( \27635 , \27632 , \27634 );
nand \U$27390 ( \27636 , \27629 , \27635 );
not \U$27391 ( \27637 , \27621 );
nand \U$27392 ( \27638 , \27637 , \27625 );
nand \U$27393 ( \27639 , \27636 , \27638 );
not \U$27394 ( \27640 , \27639 );
not \U$27395 ( \27641 , \27640 );
or \U$27396 ( \27642 , \27615 , \27641 );
not \U$27397 ( \27643 , \27638 );
not \U$27398 ( \27644 , \27636 );
or \U$27399 ( \27645 , \27643 , \27644 );
not \U$27400 ( \27646 , \27614 );
nand \U$27401 ( \27647 , \27645 , \27646 );
nand \U$27402 ( \27648 , \27642 , \27647 );
not \U$27403 ( \27649 , \27599 );
not \U$27404 ( \27650 , \27566 );
not \U$27405 ( \27651 , \27650 );
or \U$27406 ( \27652 , \27649 , \27651 );
nand \U$27407 ( \27653 , \27598 , \27566 );
nand \U$27408 ( \27654 , \27652 , \27653 );
nand \U$27409 ( \27655 , \27648 , \27654 );
not \U$27410 ( \27656 , \27638 );
not \U$27411 ( \27657 , \27636 );
or \U$27412 ( \27658 , \27656 , \27657 );
nand \U$27413 ( \27659 , \27658 , \27614 );
nand \U$27414 ( \27660 , \27609 , \27655 , \27659 );
not \U$27415 ( \27661 , \27604 );
not \U$27416 ( \27662 , \27542 );
or \U$27417 ( \27663 , \27661 , \27662 );
not \U$27418 ( \27664 , \27095 );
nand \U$27419 ( \27665 , \27538 , \27664 );
nand \U$27420 ( \27666 , \27663 , \27665 );
not \U$27421 ( \27667 , \27666 );
not \U$27422 ( \27668 , \26561 );
nand \U$27423 ( \27669 , \27668 , \26512 );
not \U$27424 ( \27670 , \27669 );
not \U$27425 ( \27671 , \26592 );
or \U$27426 ( \27672 , \27670 , \27671 );
not \U$27427 ( \27673 , \26512 );
nand \U$27428 ( \27674 , \27673 , \26561 );
nand \U$27429 ( \27675 , \27672 , \27674 );
not \U$27430 ( \27676 , \26527 );
not \U$27431 ( \27677 , \8169 );
or \U$27432 ( \27678 , \27676 , \27677 );
xor \U$27433 ( \27679 , RIbe2a028_80, RIbe29998_66);
nand \U$27434 ( \27680 , \8172 , \27679 );
nand \U$27435 ( \27681 , \27678 , \27680 );
not \U$27436 ( \27682 , \26543 );
not \U$27437 ( \27683 , \7609 );
or \U$27438 ( \27684 , \27682 , \27683 );
xor \U$27439 ( \27685 , RIbe29d58_74, RIbe28f48_44);
nand \U$27440 ( \27686 , \11201 , \27685 );
nand \U$27441 ( \27687 , \27684 , \27686 );
xor \U$27442 ( \27688 , \27681 , \27687 );
xor \U$27443 ( \27689 , RIbe290b0_47, RIbe2ae38_110);
not \U$27444 ( \27690 , \27689 );
not \U$27445 ( \27691 , \2730 );
or \U$27446 ( \27692 , \27690 , \27691 );
xor \U$27447 ( \27693 , RIbe290b0_47, RIbe2aeb0_111);
nand \U$27448 ( \27694 , \399 , \27693 );
nand \U$27449 ( \27695 , \27692 , \27694 );
not \U$27450 ( \27696 , \27695 );
and \U$27451 ( \27697 , \27688 , \27696 );
not \U$27452 ( \27698 , \27688 );
and \U$27453 ( \27699 , \27698 , \27695 );
nor \U$27454 ( \27700 , \27697 , \27699 );
not \U$27455 ( \27701 , \27700 );
and \U$27456 ( \27702 , \27675 , \27701 );
not \U$27457 ( \27703 , \27675 );
and \U$27458 ( \27704 , \27703 , \27700 );
nor \U$27459 ( \27705 , \27702 , \27704 );
not \U$27460 ( \27706 , \26923 );
not \U$27461 ( \27707 , \26955 );
or \U$27462 ( \27708 , \27706 , \27707 );
or \U$27463 ( \27709 , \26955 , \26923 );
nand \U$27464 ( \27710 , \27709 , \26893 );
nand \U$27465 ( \27711 , \27708 , \27710 );
and \U$27466 ( \27712 , \27705 , \27711 );
not \U$27467 ( \27713 , \27705 );
not \U$27468 ( \27714 , \27711 );
and \U$27469 ( \27715 , \27713 , \27714 );
nor \U$27470 ( \27716 , \27712 , \27715 );
or \U$27471 ( \27717 , \26989 , \26859 );
nand \U$27472 ( \27718 , \27717 , \26961 );
nand \U$27473 ( \27719 , \26989 , \26859 );
nand \U$27474 ( \27720 , \27718 , \27719 );
xor \U$27475 ( \27721 , \27716 , \27720 );
not \U$27476 ( \27722 , \27322 );
not \U$27477 ( \27723 , \27339 );
or \U$27478 ( \27724 , \27722 , \27723 );
nand \U$27479 ( \27725 , \27724 , \27321 );
xor \U$27480 ( \27726 , \27126 , \27130 );
and \U$27481 ( \27727 , \27726 , \27155 );
and \U$27482 ( \27728 , \27126 , \27130 );
or \U$27483 ( \27729 , \27727 , \27728 );
xnor \U$27484 ( \27730 , \27725 , \27729 );
not \U$27485 ( \27731 , \27181 );
xnor \U$27486 ( \27732 , \27205 , \27234 );
not \U$27487 ( \27733 , \27732 );
or \U$27488 ( \27734 , \27731 , \27733 );
nand \U$27489 ( \27735 , \27235 , \27206 );
nand \U$27490 ( \27736 , \27734 , \27735 );
xor \U$27491 ( \27737 , \27730 , \27736 );
xnor \U$27492 ( \27738 , \27721 , \27737 );
not \U$27493 ( \27739 , \26994 );
not \U$27494 ( \27740 , \27739 );
not \U$27495 ( \27741 , \27086 );
or \U$27496 ( \27742 , \27740 , \27741 );
not \U$27497 ( \27743 , \27021 );
nand \U$27498 ( \27744 , \27743 , \27085 );
nand \U$27499 ( \27745 , \27742 , \27744 );
xor \U$27500 ( \27746 , \27738 , \27745 );
or \U$27501 ( \27747 , \27156 , \27236 );
nand \U$27502 ( \27748 , \27747 , \27101 );
nand \U$27503 ( \27749 , \27236 , \27156 );
nand \U$27504 ( \27750 , \27748 , \27749 );
xor \U$27505 ( \27751 , \26802 , \26832 );
and \U$27506 ( \27752 , \27751 , \26858 );
and \U$27507 ( \27753 , \26802 , \26832 );
or \U$27508 ( \27754 , \27752 , \27753 );
not \U$27509 ( \27755 , \27135 );
not \U$27510 ( \27756 , \282 );
or \U$27511 ( \27757 , \27755 , \27756 );
xor \U$27512 ( \27758 , RIbe29038_46, RIbe2b450_123);
nand \U$27513 ( \27759 , \1583 , \27758 );
nand \U$27514 ( \27760 , \27757 , \27759 );
or \U$27515 ( \27761 , RIbe28fc0_45, RIbe29038_46);
nand \U$27516 ( \27762 , \27761 , RIbe2ae38_110);
nand \U$27517 ( \27763 , RIbe28fc0_45, RIbe29038_46);
and \U$27518 ( \27764 , \27762 , \27763 , RIbe290b0_47);
or \U$27519 ( \27765 , \27760 , \27764 );
nand \U$27520 ( \27766 , \27760 , \27764 );
nand \U$27521 ( \27767 , \27765 , \27766 );
not \U$27522 ( \27768 , \27767 );
buf \U$27523 ( \27769 , \27280 );
not \U$27524 ( \27770 , \27769 );
not \U$27525 ( \27771 , \27275 );
or \U$27526 ( \27772 , \27770 , \27771 );
or \U$27527 ( \27773 , \27769 , \27275 );
nand \U$27528 ( \27774 , \27773 , \27287 );
nand \U$27529 ( \27775 , \27772 , \27774 );
not \U$27530 ( \27776 , \27775 );
or \U$27531 ( \27777 , \27768 , \27776 );
or \U$27532 ( \27778 , \27775 , \27767 );
nand \U$27533 ( \27779 , \27777 , \27778 );
buf \U$27534 ( \27780 , \27303 );
not \U$27535 ( \27781 , \27780 );
not \U$27536 ( \27782 , \27314 );
or \U$27537 ( \27783 , \27781 , \27782 );
or \U$27538 ( \27784 , \27780 , \27314 );
not \U$27539 ( \27785 , \27297 );
nand \U$27540 ( \27786 , \27784 , \27785 );
nand \U$27541 ( \27787 , \27783 , \27786 );
and \U$27542 ( \27788 , \27779 , \27787 );
not \U$27543 ( \27789 , \27779 );
not \U$27544 ( \27790 , \27787 );
and \U$27545 ( \27791 , \27789 , \27790 );
nor \U$27546 ( \27792 , \27788 , \27791 );
nor \U$27547 ( \27793 , \27754 , \27792 );
not \U$27548 ( \27794 , \27793 );
nand \U$27549 ( \27795 , \27754 , \27792 );
nand \U$27550 ( \27796 , \27794 , \27795 );
not \U$27551 ( \27797 , \27180 );
not \U$27552 ( \27798 , \27174 );
or \U$27553 ( \27799 , \27797 , \27798 );
not \U$27554 ( \27800 , \27163 );
nand \U$27555 ( \27801 , \27800 , \27170 );
nand \U$27556 ( \27802 , \27799 , \27801 );
not \U$27557 ( \27803 , \27125 );
not \U$27558 ( \27804 , \27119 );
or \U$27559 ( \27805 , \27803 , \27804 );
nand \U$27560 ( \27806 , \27115 , \27107 );
nand \U$27561 ( \27807 , \27805 , \27806 );
xor \U$27562 ( \27808 , \27802 , \27807 );
not \U$27563 ( \27809 , \27214 );
not \U$27564 ( \27810 , \27809 );
not \U$27565 ( \27811 , \27232 );
or \U$27566 ( \27812 , \27810 , \27811 );
nand \U$27567 ( \27813 , \27220 , \27227 );
nand \U$27568 ( \27814 , \27812 , \27813 );
not \U$27569 ( \27815 , \27814 );
and \U$27570 ( \27816 , \27808 , \27815 );
not \U$27571 ( \27817 , \27808 );
and \U$27572 ( \27818 , \27817 , \27814 );
nor \U$27573 ( \27819 , \27816 , \27818 );
xor \U$27574 ( \27820 , \27796 , \27819 );
xor \U$27575 ( \27821 , \27750 , \27820 );
not \U$27576 ( \27822 , \27268 );
not \U$27577 ( \27823 , \27349 );
not \U$27578 ( \27824 , \27823 );
or \U$27579 ( \27825 , \27822 , \27824 );
not \U$27580 ( \27826 , \27340 );
nand \U$27581 ( \27827 , \27826 , \27345 );
nand \U$27582 ( \27828 , \27825 , \27827 );
xor \U$27583 ( \27829 , \27821 , \27828 );
xor \U$27584 ( \27830 , \27746 , \27829 );
nand \U$27585 ( \27831 , \27485 , \27533 );
or \U$27586 ( \27832 , \27478 , \27420 );
nand \U$27587 ( \27833 , \27831 , \27832 );
and \U$27588 ( \27834 , \27830 , \27833 );
not \U$27589 ( \27835 , \27830 );
and \U$27590 ( \27836 , \27832 , \27831 );
and \U$27591 ( \27837 , \27835 , \27836 );
nor \U$27592 ( \27838 , \27834 , \27837 );
buf \U$27593 ( \27839 , \27353 );
not \U$27594 ( \27840 , \27839 );
not \U$27595 ( \27841 , \27237 );
not \U$27596 ( \27842 , \27841 );
and \U$27597 ( \27843 , \27840 , \27842 );
nand \U$27598 ( \27844 , \27839 , \27841 );
and \U$27599 ( \27845 , \27844 , \27416 );
nor \U$27600 ( \27846 , \27843 , \27845 );
not \U$27601 ( \27847 , \27137 );
not \U$27602 ( \27848 , \27143 );
or \U$27603 ( \27849 , \27847 , \27848 );
not \U$27604 ( \27850 , \27146 );
not \U$27605 ( \27851 , \27137 );
not \U$27606 ( \27852 , \27851 );
or \U$27607 ( \27853 , \27850 , \27852 );
nand \U$27608 ( \27854 , \27853 , \27154 );
nand \U$27609 ( \27855 , \27849 , \27854 );
xor \U$27610 ( \27856 , \27324 , \27330 );
and \U$27611 ( \27857 , \27856 , \27338 );
and \U$27612 ( \27858 , \27324 , \27330 );
or \U$27613 ( \27859 , \27857 , \27858 );
xor \U$27614 ( \27860 , \27855 , \27859 );
or \U$27615 ( \27861 , \26537 , \26545 );
nand \U$27616 ( \27862 , \27861 , \26539 );
xor \U$27617 ( \27863 , \27860 , \27862 );
not \U$27618 ( \27864 , \27202 );
not \U$27619 ( \27865 , \8624 );
or \U$27620 ( \27866 , \27864 , \27865 );
xor \U$27621 ( \27867 , RIbe280c0_13, RIbe2ac58_106);
nand \U$27622 ( \27868 , \1263 , \27867 );
nand \U$27623 ( \27869 , \27866 , \27868 );
not \U$27624 ( \27870 , \27869 );
not \U$27625 ( \27871 , \27328 );
not \U$27626 ( \27872 , \10812 );
or \U$27627 ( \27873 , \27871 , \27872 );
xor \U$27628 ( \27874 , RIbe296c8_60, RIbe2a7a8_96);
nand \U$27629 ( \27875 , \907 , \27874 );
nand \U$27630 ( \27876 , \27873 , \27875 );
not \U$27631 ( \27877 , \27876 );
not \U$27632 ( \27878 , \27877 );
or \U$27633 ( \27879 , \27870 , \27878 );
not \U$27634 ( \27880 , \27869 );
nand \U$27635 ( \27881 , \27880 , \27876 );
nand \U$27636 ( \27882 , \27879 , \27881 );
not \U$27637 ( \27883 , \27113 );
not \U$27638 ( \27884 , \2519 );
or \U$27639 ( \27885 , \27883 , \27884 );
xor \U$27640 ( \27886 , RIbe2a118_82, RIbe28480_21);
nand \U$27641 ( \27887 , \11263 , \27886 );
nand \U$27642 ( \27888 , \27885 , \27887 );
xor \U$27643 ( \27889 , \27882 , \27888 );
buf \U$27644 ( \27890 , \27889 );
not \U$27645 ( \27891 , \27890 );
not \U$27646 ( \27892 , \27187 );
not \U$27647 ( \27893 , \27193 );
or \U$27648 ( \27894 , \27892 , \27893 );
not \U$27649 ( \27895 , \27187 );
not \U$27650 ( \27896 , \27895 );
not \U$27651 ( \27897 , \27196 );
or \U$27652 ( \27898 , \27896 , \27897 );
nand \U$27653 ( \27899 , \27898 , \27204 );
nand \U$27654 ( \27900 , \27894 , \27899 );
not \U$27655 ( \27901 , \18831 );
not \U$27656 ( \27902 , \27105 );
not \U$27657 ( \27903 , \27902 );
and \U$27658 ( \27904 , \27901 , \27903 );
xor \U$27659 ( \27905 , RIbe2aaf0_103, RIbe28318_18);
and \U$27660 ( \27906 , \27905 , RIbe2ab68_104);
nor \U$27661 ( \27907 , \27904 , \27906 );
not \U$27662 ( \27908 , \27907 );
not \U$27663 ( \27909 , \26534 );
not \U$27664 ( \27910 , \10433 );
or \U$27665 ( \27911 , \27909 , \27910 );
xor \U$27666 ( \27912 , RIbe291a0_49, RIbe2a550_91);
nand \U$27667 ( \27913 , \20336 , \27912 );
nand \U$27668 ( \27914 , \27911 , \27913 );
not \U$27669 ( \27915 , \27914 );
or \U$27670 ( \27916 , \27908 , \27915 );
or \U$27671 ( \27917 , \27914 , \27907 );
nand \U$27672 ( \27918 , \27916 , \27917 );
not \U$27673 ( \27919 , \27212 );
not \U$27674 ( \27920 , \4893 );
or \U$27675 ( \27921 , \27919 , \27920 );
nand \U$27676 ( \27922 , \2707 , \21975 );
nand \U$27677 ( \27923 , \27921 , \27922 );
and \U$27678 ( \27924 , \27918 , \27923 );
not \U$27679 ( \27925 , \27918 );
not \U$27680 ( \27926 , \27923 );
and \U$27681 ( \27927 , \27925 , \27926 );
nor \U$27682 ( \27928 , \27924 , \27927 );
xnor \U$27683 ( \27929 , \27900 , \27928 );
not \U$27684 ( \27930 , \27929 );
or \U$27685 ( \27931 , \27891 , \27930 );
or \U$27686 ( \27932 , \27929 , \27890 );
nand \U$27687 ( \27933 , \27931 , \27932 );
xor \U$27688 ( \27934 , \27863 , \27933 );
not \U$27689 ( \27935 , \27301 );
not \U$27690 ( \27936 , \8806 );
or \U$27691 ( \27937 , \27935 , \27936 );
nand \U$27692 ( \27938 , \8794 , \22004 );
nand \U$27693 ( \27939 , \27937 , \27938 );
not \U$27694 ( \27940 , \27161 );
not \U$27695 ( \27941 , \1780 );
or \U$27696 ( \27942 , \27940 , \27941 );
nand \U$27697 ( \27943 , \2475 , \22028 );
nand \U$27698 ( \27944 , \27942 , \27943 );
xor \U$27699 ( \27945 , \27939 , \27944 );
not \U$27700 ( \27946 , \27152 );
not \U$27701 ( \27947 , \879 );
or \U$27702 ( \27948 , \27946 , \27947 );
nand \U$27703 ( \27949 , \8680 , \22018 );
nand \U$27704 ( \27950 , \27948 , \27949 );
xor \U$27705 ( \27951 , \27945 , \27950 );
not \U$27706 ( \27952 , \27312 );
not \U$27707 ( \27953 , \2457 );
or \U$27708 ( \27954 , \27952 , \27953 );
nand \U$27709 ( \27955 , \2463 , \22010 );
nand \U$27710 ( \27956 , \27954 , \27955 );
not \U$27711 ( \27957 , \27178 );
not \U$27712 ( \27958 , \14423 );
or \U$27713 ( \27959 , \27957 , \27958 );
xor \U$27714 ( \27960 , RIbe293f8_54, RIbe2af28_112);
nand \U$27715 ( \27961 , \16917 , \27960 );
nand \U$27716 ( \27962 , \27959 , \27961 );
xor \U$27717 ( \27963 , \27956 , \27962 );
not \U$27718 ( \27964 , \27285 );
not \U$27719 ( \27965 , \3408 );
or \U$27720 ( \27966 , \27964 , \27965 );
xor \U$27721 ( \27967 , RIbe2b360_121, RIbe28390_19);
nand \U$27722 ( \27968 , \2777 , \27967 );
nand \U$27723 ( \27969 , \27966 , \27968 );
xor \U$27724 ( \27970 , \27963 , \27969 );
xor \U$27725 ( \27971 , \27951 , \27970 );
not \U$27726 ( \27972 , \26559 );
not \U$27727 ( \27973 , \17563 );
or \U$27728 ( \27974 , \27972 , \27973 );
xor \U$27729 ( \27975 , RIbe29740_61, RIbe2a190_83);
nand \U$27730 ( \27976 , \11400 , \27975 );
nand \U$27731 ( \27977 , \27974 , \27976 );
not \U$27732 ( \27978 , \27977 );
not \U$27733 ( \27979 , \27168 );
not \U$27734 ( \27980 , \3401 );
or \U$27735 ( \27981 , \27979 , \27980 );
xor \U$27736 ( \27982 , RIbe2a4d8_90, RIbe28b88_36);
nand \U$27737 ( \27983 , \13250 , \27982 );
nand \U$27738 ( \27984 , \27981 , \27983 );
not \U$27739 ( \27985 , \27984 );
not \U$27740 ( \27986 , \27985 );
or \U$27741 ( \27987 , \27978 , \27986 );
not \U$27742 ( \27988 , \27977 );
nand \U$27743 ( \27989 , \27984 , \27988 );
nand \U$27744 ( \27990 , \27987 , \27989 );
not \U$27745 ( \27991 , \27273 );
not \U$27746 ( \27992 , \11344 );
buf \U$27747 ( \27993 , \27992 );
not \U$27748 ( \27994 , \27993 );
or \U$27749 ( \27995 , \27991 , \27994 );
xor \U$27750 ( \27996 , RIbe28138_14, RIbe2a280_85);
nand \U$27751 ( \27997 , \11348 , \27996 );
nand \U$27752 ( \27998 , \27995 , \27997 );
and \U$27753 ( \27999 , \27990 , \27998 );
not \U$27754 ( \28000 , \27990 );
not \U$27755 ( \28001 , \27998 );
and \U$27756 ( \28002 , \28000 , \28001 );
nor \U$27757 ( \28003 , \27999 , \28002 );
xor \U$27758 ( \28004 , \27971 , \28003 );
xor \U$27759 ( \28005 , \27934 , \28004 );
or \U$27760 ( \28006 , \26708 , \26599 );
nand \U$27761 ( \28007 , \28006 , \26601 );
xor \U$27762 ( \28008 , \28005 , \28007 );
not \U$27763 ( \28009 , \27016 );
not \U$27764 ( \28010 , \27011 );
or \U$27765 ( \28011 , \28009 , \28010 );
nand \U$27766 ( \28012 , \27006 , \27000 );
nand \U$27767 ( \28013 , \28011 , \28012 );
not \U$27768 ( \28014 , \27225 );
not \U$27769 ( \28015 , \1793 );
or \U$27770 ( \28016 , \28014 , \28015 );
nand \U$27771 ( \28017 , \970 , \22041 );
nand \U$27772 ( \28018 , \28016 , \28017 );
not \U$27773 ( \28019 , \27277 );
not \U$27774 ( \28020 , \13529 );
or \U$27775 ( \28021 , \28019 , \28020 );
xor \U$27776 ( \28022 , RIbe29470_55, RIbe2b108_116);
nand \U$27777 ( \28023 , \16875 , \28022 );
nand \U$27778 ( \28024 , \28021 , \28023 );
not \U$27779 ( \28025 , \27295 );
not \U$27780 ( \28026 , \17592 );
or \U$27781 ( \28027 , \28025 , \28026 );
nand \U$27782 ( \28028 , \16646 , \22034 );
nand \U$27783 ( \28029 , \28027 , \28028 );
and \U$27784 ( \28030 , \28024 , \28029 );
not \U$27785 ( \28031 , \28024 );
not \U$27786 ( \28032 , \28029 );
and \U$27787 ( \28033 , \28031 , \28032 );
nor \U$27788 ( \28034 , \28030 , \28033 );
xor \U$27789 ( \28035 , \28018 , \28034 );
not \U$27790 ( \28036 , \27185 );
not \U$27791 ( \28037 , \25897 );
or \U$27792 ( \28038 , \28036 , \28037 );
xor \U$27793 ( \28039 , RIbe28c00_37, RIbe2b018_114);
nand \U$27794 ( \28040 , \20583 , \28039 );
nand \U$27795 ( \28041 , \28038 , \28040 );
not \U$27796 ( \28042 , \27191 );
or \U$27797 ( \28043 , \2891 , \28042 );
xor \U$27798 ( \28044 , RIbe285e8_24, RIbe2a898_98);
nand \U$27799 ( \28045 , \8270 , \28044 );
nand \U$27800 ( \28046 , \28043 , \28045 );
not \U$27801 ( \28047 , \27141 );
not \U$27802 ( \28048 , \8697 );
or \U$27803 ( \28049 , \28047 , \28048 );
xor \U$27804 ( \28050 , RIbe27c88_4, RIbe2a2f8_86);
nand \U$27805 ( \28051 , \11094 , \28050 );
nand \U$27806 ( \28052 , \28049 , \28051 );
xor \U$27807 ( \28053 , \28046 , \28052 );
xor \U$27808 ( \28054 , \28041 , \28053 );
xor \U$27809 ( \28055 , \28035 , \28054 );
not \U$27810 ( \28056 , \27123 );
not \U$27811 ( \28057 , \10938 );
or \U$27812 ( \28058 , \28056 , \28057 );
nand \U$27813 ( \28059 , \8245 , \21982 );
nand \U$27814 ( \28060 , \28058 , \28059 );
not \U$27815 ( \28061 , \27335 );
not \U$27816 ( \28062 , \7513 );
or \U$27817 ( \28063 , \28061 , \28062 );
xor \U$27818 ( \28064 , RIbe29b78_70, RIbe29c68_72);
nand \U$27819 ( \28065 , \4580 , \28064 );
nand \U$27820 ( \28066 , \28063 , \28065 );
not \U$27821 ( \28067 , \28066 );
not \U$27822 ( \28068 , \28067 );
not \U$27823 ( \28069 , \27218 );
not \U$27824 ( \28070 , \11453 );
or \U$27825 ( \28071 , \28069 , \28070 );
nand \U$27826 ( \28072 , \10401 , \21987 );
nand \U$27827 ( \28073 , \28071 , \28072 );
not \U$27828 ( \28074 , \28073 );
or \U$27829 ( \28075 , \28068 , \28074 );
or \U$27830 ( \28076 , \28073 , \28067 );
nand \U$27831 ( \28077 , \28075 , \28076 );
xor \U$27832 ( \28078 , \28060 , \28077 );
xor \U$27833 ( \28079 , \28055 , \28078 );
not \U$27834 ( \28080 , \26596 );
not \U$27835 ( \28081 , \26550 );
or \U$27836 ( \28082 , \28080 , \28081 );
nand \U$27837 ( \28083 , \28082 , \26518 );
nand \U$27838 ( \28084 , \26597 , \26553 );
nand \U$27839 ( \28085 , \28083 , \28084 );
xor \U$27840 ( \28086 , \28079 , \28085 );
xor \U$27841 ( \28087 , \28013 , \28086 );
xor \U$27842 ( \28088 , \28008 , \28087 );
xor \U$27843 ( \28089 , \27846 , \28088 );
not \U$27844 ( \28090 , \27090 );
not \U$27845 ( \28091 , \26778 );
or \U$27846 ( \28092 , \28090 , \28091 );
nand \U$27847 ( \28093 , \26773 , \26711 );
nand \U$27848 ( \28094 , \28092 , \28093 );
xor \U$27849 ( \28095 , \28089 , \28094 );
not \U$27850 ( \28096 , \28095 );
and \U$27851 ( \28097 , \27838 , \28096 );
not \U$27852 ( \28098 , \27838 );
and \U$27853 ( \28099 , \28098 , \28095 );
nor \U$27854 ( \28100 , \28097 , \28099 );
nand \U$27855 ( \28101 , \27667 , \28100 );
not \U$27856 ( \28102 , \26272 );
nand \U$27857 ( \28103 , \28102 , \25810 );
nand \U$27858 ( \28104 , \27660 , \28101 , \28103 );
not \U$27859 ( \28105 , \27629 );
not \U$27860 ( \28106 , \28105 );
not \U$27861 ( \28107 , \27635 );
and \U$27862 ( \28108 , \28106 , \28107 );
and \U$27863 ( \28109 , \27635 , \28105 );
nor \U$27864 ( \28110 , \28108 , \28109 );
not \U$27865 ( \28111 , \28110 );
not \U$27866 ( \28112 , \27544 );
not \U$27867 ( \28113 , \28112 );
not \U$27868 ( \28114 , \27561 );
or \U$27869 ( \28115 , \28113 , \28114 );
or \U$27870 ( \28116 , \28112 , \27561 );
nand \U$27871 ( \28117 , \28115 , \28116 );
not \U$27872 ( \28118 , \28117 );
and \U$27873 ( \28119 , \25861 , \26254 );
nand \U$27874 ( \28120 , \26248 , \25998 );
not \U$27875 ( \28121 , \28120 );
nor \U$27876 ( \28122 , \28119 , \28121 );
not \U$27877 ( \28123 , \28122 );
or \U$27878 ( \28124 , \28118 , \28123 );
not \U$27879 ( \28125 , \28120 );
nand \U$27880 ( \28126 , \25861 , \26254 );
not \U$27881 ( \28127 , \28126 );
or \U$27882 ( \28128 , \28125 , \28127 );
not \U$27883 ( \28129 , \28117 );
nand \U$27884 ( \28130 , \28128 , \28129 );
nand \U$27885 ( \28131 , \28124 , \28130 );
not \U$27886 ( \28132 , \28131 );
or \U$27887 ( \28133 , \28111 , \28132 );
or \U$27888 ( \28134 , \28131 , \28110 );
nand \U$27889 ( \28135 , \28133 , \28134 );
xor \U$27890 ( \28136 , \25855 , \26259 );
and \U$27891 ( \28137 , \28136 , \26271 );
and \U$27892 ( \28138 , \25855 , \26259 );
or \U$27893 ( \28139 , \28137 , \28138 );
or \U$27894 ( \28140 , \28135 , \28139 );
and \U$27895 ( \28141 , \27648 , \27654 );
not \U$27896 ( \28142 , \27648 );
not \U$27897 ( \28143 , \27654 );
and \U$27898 ( \28144 , \28142 , \28143 );
nor \U$27899 ( \28145 , \28141 , \28144 );
not \U$27900 ( \28146 , \28145 );
not \U$27901 ( \28147 , \28110 );
not \U$27902 ( \28148 , \28147 );
not \U$27903 ( \28149 , \28131 );
or \U$27904 ( \28150 , \28148 , \28149 );
or \U$27905 ( \28151 , \28122 , \28129 );
nand \U$27906 ( \28152 , \28150 , \28151 );
not \U$27907 ( \28153 , \28152 );
nand \U$27908 ( \28154 , \28146 , \28153 );
nand \U$27909 ( \28155 , \28140 , \28154 );
nor \U$27910 ( \28156 , \28104 , \28155 );
not \U$27911 ( \28157 , \28156 );
or \U$27912 ( \28158 , \26276 , \28157 );
nand \U$27913 ( \28159 , \28145 , \28152 );
nand \U$27914 ( \28160 , \28135 , \28139 );
nand \U$27915 ( \28161 , \28159 , \28160 );
and \U$27916 ( \28162 , \28161 , \28154 );
not \U$27917 ( \28163 , \27660 );
not \U$27918 ( \28164 , \28101 );
nor \U$27919 ( \28165 , \28163 , \28164 );
and \U$27920 ( \28166 , \28162 , \28165 );
not \U$27921 ( \28167 , \28100 );
nand \U$27922 ( \28168 , \28167 , \27666 );
not \U$27923 ( \28169 , \28168 );
not \U$27924 ( \28170 , \27659 );
not \U$27925 ( \28171 , \27655 );
or \U$27926 ( \28172 , \28170 , \28171 );
not \U$27927 ( \28173 , \27609 );
nand \U$27928 ( \28174 , \28172 , \28173 );
not \U$27929 ( \28175 , \28174 );
or \U$27930 ( \28176 , \28169 , \28175 );
nand \U$27931 ( \28177 , \28176 , \28101 );
not \U$27932 ( \28178 , \28177 );
nor \U$27933 ( \28179 , \28166 , \28178 );
nand \U$27934 ( \28180 , \28158 , \28179 );
not \U$27935 ( \28181 , \28180 );
xor \U$27936 ( \28182 , \21696 , \21697 );
xor \U$27937 ( \28183 , \28182 , \21920 );
xor \U$27938 ( \28184 , \21915 , \21733 );
not \U$27939 ( \28185 , \28184 );
and \U$27940 ( \28186 , \21904 , \21848 );
not \U$27941 ( \28187 , \21904 );
not \U$27942 ( \28188 , \21848 );
and \U$27943 ( \28189 , \28187 , \28188 );
nor \U$27944 ( \28190 , \28186 , \28189 );
not \U$27945 ( \28191 , \28190 );
not \U$27946 ( \28192 , \27874 );
not \U$27947 ( \28193 , \900 );
or \U$27948 ( \28194 , \28192 , \28193 );
nand \U$27949 ( \28195 , \908 , \21561 );
nand \U$27950 ( \28196 , \28194 , \28195 );
not \U$27951 ( \28197 , \27975 );
not \U$27952 ( \28198 , \10690 );
or \U$27953 ( \28199 , \28197 , \28198 );
nand \U$27954 ( \28200 , \13278 , \21887 );
nand \U$27955 ( \28201 , \28199 , \28200 );
or \U$27956 ( \28202 , \28196 , \28201 );
not \U$27957 ( \28203 , \27886 );
not \U$27958 ( \28204 , \3483 );
or \U$27959 ( \28205 , \28203 , \28204 );
nand \U$27960 ( \28206 , \2527 , \21896 );
nand \U$27961 ( \28207 , \28205 , \28206 );
nand \U$27962 ( \28208 , \28202 , \28207 );
nand \U$27963 ( \28209 , \28196 , \28201 );
nand \U$27964 ( \28210 , \28208 , \28209 );
not \U$27965 ( \28211 , \28210 );
not \U$27966 ( \28212 , \28044 );
not \U$27967 ( \28213 , \7618 );
or \U$27968 ( \28214 , \28212 , \28213 );
nand \U$27969 ( \28215 , \2625 , \21738 );
nand \U$27970 ( \28216 , \28214 , \28215 );
not \U$27971 ( \28217 , \28216 );
not \U$27972 ( \28218 , \28217 );
not \U$27973 ( \28219 , \28050 );
not \U$27974 ( \28220 , \9374 );
or \U$27975 ( \28221 , \28219 , \28220 );
nand \U$27976 ( \28222 , \8705 , \21787 );
nand \U$27977 ( \28223 , \28221 , \28222 );
not \U$27978 ( \28224 , \28223 );
not \U$27979 ( \28225 , \28224 );
or \U$27980 ( \28226 , \28218 , \28225 );
not \U$27981 ( \28227 , \28022 );
not \U$27982 ( \28228 , \21852 );
or \U$27983 ( \28229 , \28227 , \28228 );
nand \U$27984 ( \28230 , \13534 , \21850 );
nand \U$27985 ( \28231 , \28229 , \28230 );
nand \U$27986 ( \28232 , \28226 , \28231 );
nand \U$27987 ( \28233 , \28216 , \28223 );
nand \U$27988 ( \28234 , \28232 , \28233 );
not \U$27989 ( \28235 , \28039 );
not \U$27990 ( \28236 , \17570 );
or \U$27991 ( \28237 , \28235 , \28236 );
nand \U$27992 ( \28238 , \21442 , \21864 );
nand \U$27993 ( \28239 , \28237 , \28238 );
not \U$27994 ( \28240 , \28239 );
not \U$27995 ( \28241 , \27982 );
not \U$27996 ( \28242 , \2553 );
or \U$27997 ( \28243 , \28241 , \28242 );
nand \U$27998 ( \28244 , \2559 , \21746 );
nand \U$27999 ( \28245 , \28243 , \28244 );
not \U$28000 ( \28246 , \28245 );
or \U$28001 ( \28247 , \28240 , \28246 );
or \U$28002 ( \28248 , \28239 , \28245 );
not \U$28003 ( \28249 , \27996 );
not \U$28004 ( \28250 , \13268 );
or \U$28005 ( \28251 , \28249 , \28250 );
nand \U$28006 ( \28252 , \18667 , \21777 );
nand \U$28007 ( \28253 , \28251 , \28252 );
nand \U$28008 ( \28254 , \28248 , \28253 );
nand \U$28009 ( \28255 , \28247 , \28254 );
xor \U$28010 ( \28256 , \28234 , \28255 );
not \U$28011 ( \28257 , \28256 );
or \U$28012 ( \28258 , \28211 , \28257 );
nand \U$28013 ( \28259 , \28234 , \28255 );
nand \U$28014 ( \28260 , \28258 , \28259 );
not \U$28015 ( \28261 , \27679 );
not \U$28016 ( \28262 , \22849 );
or \U$28017 ( \28263 , \28261 , \28262 );
nand \U$28018 ( \28264 , \8930 , \21880 );
nand \U$28019 ( \28265 , \28263 , \28264 );
not \U$28020 ( \28266 , \27693 );
not \U$28021 ( \28267 , \10567 );
or \U$28022 ( \28268 , \28266 , \28267 );
nand \U$28023 ( \28269 , \398 , \21547 );
nand \U$28024 ( \28270 , \28268 , \28269 );
or \U$28025 ( \28271 , \28265 , \28270 );
not \U$28026 ( \28272 , \27867 );
not \U$28027 ( \28273 , \10542 );
or \U$28028 ( \28274 , \28272 , \28273 );
nand \U$28029 ( \28275 , \1265 , \21801 );
nand \U$28030 ( \28276 , \28274 , \28275 );
nand \U$28031 ( \28277 , \28271 , \28276 );
nand \U$28032 ( \28278 , \28265 , \28270 );
nand \U$28033 ( \28279 , \28277 , \28278 );
not \U$28034 ( \28280 , \28279 );
xor \U$28035 ( \28281 , RIbe284f8_22, RIbe2aaf0_103);
not \U$28036 ( \28282 , \19580 );
and \U$28037 ( \28283 , \28281 , \28282 );
and \U$28038 ( \28284 , \21346 , RIbe2ab68_104);
nor \U$28039 ( \28285 , \28283 , \28284 );
xor \U$28040 ( \28286 , \28285 , \21558 );
xnor \U$28041 ( \28287 , \28286 , \21552 );
not \U$28042 ( \28288 , \28287 );
or \U$28043 ( \28289 , \28280 , \28288 );
not \U$28044 ( \28290 , \28285 );
xor \U$28045 ( \28291 , \21558 , \21552 );
nand \U$28046 ( \28292 , \28290 , \28291 );
nand \U$28047 ( \28293 , \28289 , \28292 );
xor \U$28048 ( \28294 , \28260 , \28293 );
not \U$28049 ( \28295 , \28294 );
or \U$28050 ( \28296 , \28191 , \28295 );
nand \U$28051 ( \28297 , \28260 , \28293 );
nand \U$28052 ( \28298 , \28296 , \28297 );
xor \U$28053 ( \28299 , \21704 , \21709 );
xor \U$28054 ( \28300 , \28299 , \21711 );
xor \U$28055 ( \28301 , \21793 , \21807 );
not \U$28056 ( \28302 , \28301 );
not \U$28057 ( \28303 , \27912 );
not \U$28058 ( \28304 , \12000 );
or \U$28059 ( \28305 , \28303 , \28304 );
nand \U$28060 ( \28306 , \11485 , \21825 );
nand \U$28061 ( \28307 , \28305 , \28306 );
not \U$28062 ( \28308 , \27905 );
not \U$28063 ( \28309 , \28282 );
or \U$28064 ( \28310 , \28308 , \28309 );
nand \U$28065 ( \28311 , \28281 , RIbe2ab68_104);
nand \U$28066 ( \28312 , \28310 , \28311 );
nor \U$28067 ( \28313 , \28307 , \28312 );
or \U$28068 ( \28314 , \28313 , \27766 );
nand \U$28069 ( \28315 , \28307 , \28312 );
nand \U$28070 ( \28316 , \28314 , \28315 );
not \U$28071 ( \28317 , \28316 );
not \U$28072 ( \28318 , \28317 );
and \U$28073 ( \28319 , \21874 , \21856 );
not \U$28074 ( \28320 , \21874 );
not \U$28075 ( \28321 , \21856 );
and \U$28076 ( \28322 , \28320 , \28321 );
nor \U$28077 ( \28323 , \28319 , \28322 );
not \U$28078 ( \28324 , \28323 );
or \U$28079 ( \28325 , \28318 , \28324 );
or \U$28080 ( \28326 , \28323 , \28317 );
nand \U$28081 ( \28327 , \28325 , \28326 );
not \U$28082 ( \28328 , \28327 );
or \U$28083 ( \28329 , \28302 , \28328 );
nand \U$28084 ( \28330 , \28323 , \28316 );
nand \U$28085 ( \28331 , \28329 , \28330 );
nor \U$28086 ( \28332 , \28300 , \28331 );
xor \U$28087 ( \28333 , \22078 , \22086 );
xor \U$28088 ( \28334 , \28333 , \22080 );
or \U$28089 ( \28335 , \28332 , \28334 );
nand \U$28090 ( \28336 , \28300 , \28331 );
nand \U$28091 ( \28337 , \28335 , \28336 );
xor \U$28092 ( \28338 , \28298 , \28337 );
xor \U$28093 ( \28339 , \22069 , \22089 );
xor \U$28094 ( \28340 , \28339 , \22132 );
and \U$28095 ( \28341 , \28338 , \28340 );
and \U$28096 ( \28342 , \28298 , \28337 );
or \U$28097 ( \28343 , \28341 , \28342 );
xor \U$28098 ( \28344 , \21522 , \21593 );
xor \U$28099 ( \28345 , \21588 , \21545 );
xor \U$28100 ( \28346 , \21529 , \21535 );
xor \U$28101 ( \28347 , \28346 , \21542 );
not \U$28102 ( \28348 , \28347 );
not \U$28103 ( \28349 , \22098 );
not \U$28104 ( \28350 , \22116 );
not \U$28105 ( \28351 , \28350 );
or \U$28106 ( \28352 , \28349 , \28351 );
not \U$28107 ( \28353 , \22098 );
nand \U$28108 ( \28354 , \28353 , \22116 );
nand \U$28109 ( \28355 , \28352 , \28354 );
not \U$28110 ( \28356 , \28355 );
or \U$28111 ( \28357 , \28348 , \28356 );
or \U$28112 ( \28358 , \28355 , \28347 );
xor \U$28113 ( \28359 , \21573 , \21566 );
xor \U$28114 ( \28360 , \28359 , \21582 );
nand \U$28115 ( \28361 , \28358 , \28360 );
nand \U$28116 ( \28362 , \28357 , \28361 );
or \U$28117 ( \28363 , \28345 , \28362 );
xor \U$28118 ( \28364 , \21763 , \21785 );
xor \U$28119 ( \28365 , \28364 , \21811 );
nand \U$28120 ( \28366 , \28363 , \28365 );
nand \U$28121 ( \28367 , \28345 , \28362 );
nand \U$28122 ( \28368 , \28366 , \28367 );
xor \U$28123 ( \28369 , \28344 , \28368 );
xor \U$28124 ( \28370 , \21814 , \21816 );
xor \U$28125 ( \28371 , \28370 , \21908 );
and \U$28126 ( \28372 , \28369 , \28371 );
and \U$28127 ( \28373 , \28344 , \28368 );
or \U$28128 ( \28374 , \28372 , \28373 );
xor \U$28129 ( \28375 , \28343 , \28374 );
not \U$28130 ( \28376 , \28375 );
or \U$28131 ( \28377 , \28185 , \28376 );
nand \U$28132 ( \28378 , \28343 , \28374 );
nand \U$28133 ( \28379 , \28377 , \28378 );
xor \U$28134 ( \28380 , \28183 , \28379 );
not \U$28135 ( \28381 , \22064 );
not \U$28136 ( \28382 , \28381 );
not \U$28137 ( \28383 , \22139 );
or \U$28138 ( \28384 , \28382 , \28383 );
not \U$28139 ( \28385 , \22139 );
nand \U$28140 ( \28386 , \28385 , \22064 );
nand \U$28141 ( \28387 , \28384 , \28386 );
not \U$28142 ( \28388 , \28387 );
xor \U$28143 ( \28389 , \21714 , \21728 );
xor \U$28144 ( \28390 , \21761 , \21751 );
buf \U$28145 ( \28391 , \21744 );
xnor \U$28146 ( \28392 , \28390 , \28391 );
not \U$28147 ( \28393 , \28392 );
not \U$28148 ( \28394 , \28393 );
not \U$28149 ( \28395 , \21830 );
not \U$28150 ( \28396 , \21823 );
not \U$28151 ( \28397 , \28396 );
or \U$28152 ( \28398 , \28395 , \28397 );
or \U$28153 ( \28399 , \21835 , \21830 );
nand \U$28154 ( \28400 , \28398 , \28399 );
xor \U$28155 ( \28401 , \28400 , \21845 );
not \U$28156 ( \28402 , \28401 );
xor \U$28157 ( \28403 , \21769 , \21775 );
xor \U$28158 ( \28404 , \28403 , \21782 );
not \U$28159 ( \28405 , \28404 );
or \U$28160 ( \28406 , \28402 , \28405 );
or \U$28161 ( \28407 , \28404 , \28401 );
nand \U$28162 ( \28408 , \28406 , \28407 );
not \U$28163 ( \28409 , \28408 );
or \U$28164 ( \28410 , \28394 , \28409 );
not \U$28165 ( \28411 , \28401 );
nand \U$28166 ( \28412 , \28411 , \28404 );
nand \U$28167 ( \28413 , \28410 , \28412 );
not \U$28168 ( \28414 , \28413 );
xor \U$28169 ( \28415 , \22092 , \22127 );
xor \U$28170 ( \28416 , \28415 , \22120 );
xor \U$28171 ( \28417 , \21901 , \21892 );
not \U$28172 ( \28418 , \21885 );
and \U$28173 ( \28419 , \28417 , \28418 );
not \U$28174 ( \28420 , \28417 );
and \U$28175 ( \28421 , \28420 , \21885 );
nor \U$28176 ( \28422 , \28419 , \28421 );
not \U$28177 ( \28423 , \28422 );
not \U$28178 ( \28424 , \28423 );
not \U$28179 ( \28425 , \27960 );
not \U$28180 ( \28426 , \14423 );
or \U$28181 ( \28427 , \28425 , \28426 );
nand \U$28182 ( \28428 , \16728 , \21770 );
nand \U$28183 ( \28429 , \28427 , \28428 );
not \U$28184 ( \28430 , \28064 );
not \U$28185 ( \28431 , \10720 );
or \U$28186 ( \28432 , \28430 , \28431 );
nand \U$28187 ( \28433 , \4580 , \22100 );
nand \U$28188 ( \28434 , \28432 , \28433 );
nor \U$28189 ( \28435 , \28429 , \28434 );
not \U$28190 ( \28436 , \27967 );
not \U$28191 ( \28437 , \3408 );
or \U$28192 ( \28438 , \28436 , \28437 );
nand \U$28193 ( \28439 , \8654 , \21577 );
nand \U$28194 ( \28440 , \28438 , \28439 );
not \U$28195 ( \28441 , \28440 );
or \U$28196 ( \28442 , \28435 , \28441 );
nand \U$28197 ( \28443 , \28429 , \28434 );
nand \U$28198 ( \28444 , \28442 , \28443 );
not \U$28199 ( \28445 , \27685 );
not \U$28200 ( \28446 , \11461 );
or \U$28201 ( \28447 , \28445 , \28446 );
not \U$28202 ( \28448 , \21843 );
nand \U$28203 ( \28449 , \28448 , \9524 );
nand \U$28204 ( \28450 , \28447 , \28449 );
not \U$28205 ( \28451 , \28450 );
and \U$28206 ( \28452 , \10752 , RIbe2ae38_110);
not \U$28207 ( \28453 , \27758 );
not \U$28208 ( \28454 , \16854 );
or \U$28209 ( \28455 , \28453 , \28454 );
nand \U$28210 ( \28456 , \1583 , \21568 );
nand \U$28211 ( \28457 , \28455 , \28456 );
xor \U$28212 ( \28458 , \28452 , \28457 );
not \U$28213 ( \28459 , \28458 );
or \U$28214 ( \28460 , \28451 , \28459 );
nand \U$28215 ( \28461 , \28457 , \28452 );
nand \U$28216 ( \28462 , \28460 , \28461 );
xor \U$28217 ( \28463 , \28444 , \28462 );
not \U$28218 ( \28464 , \28463 );
or \U$28219 ( \28465 , \28424 , \28464 );
nand \U$28220 ( \28466 , \28462 , \28444 );
nand \U$28221 ( \28467 , \28465 , \28466 );
not \U$28222 ( \28468 , \28467 );
not \U$28223 ( \28469 , \28468 );
xor \U$28224 ( \28470 , \28416 , \28469 );
not \U$28225 ( \28471 , \28470 );
or \U$28226 ( \28472 , \28414 , \28471 );
not \U$28227 ( \28473 , \28468 );
and \U$28228 ( \28474 , \28416 , \28473 );
not \U$28229 ( \28475 , \28474 );
nand \U$28230 ( \28476 , \28472 , \28475 );
xor \U$28231 ( \28477 , \28389 , \28476 );
not \U$28232 ( \28478 , \22059 );
not \U$28233 ( \28479 , \21961 );
or \U$28234 ( \28480 , \28478 , \28479 );
or \U$28235 ( \28481 , \22059 , \21961 );
nand \U$28236 ( \28482 , \28480 , \28481 );
and \U$28237 ( \28483 , \28477 , \28482 );
and \U$28238 ( \28484 , \28389 , \28476 );
or \U$28239 ( \28485 , \28483 , \28484 );
not \U$28240 ( \28486 , \28485 );
or \U$28241 ( \28487 , \28388 , \28486 );
or \U$28242 ( \28488 , \28485 , \28387 );
xor \U$28243 ( \28489 , \21689 , \21691 );
xor \U$28244 ( \28490 , \28489 , \21693 );
nand \U$28245 ( \28491 , \28488 , \28490 );
nand \U$28246 ( \28492 , \28487 , \28491 );
and \U$28247 ( \28493 , \28380 , \28492 );
and \U$28248 ( \28494 , \28183 , \28379 );
or \U$28249 ( \28495 , \28493 , \28494 );
not \U$28250 ( \28496 , \28495 );
not \U$28251 ( \28497 , \28496 );
not \U$28252 ( \28498 , \21647 );
not \U$28253 ( \28499 , \21504 );
and \U$28254 ( \28500 , \28498 , \28499 );
and \U$28255 ( \28501 , \21647 , \21504 );
nor \U$28256 ( \28502 , \28500 , \28501 );
xor \U$28257 ( \28503 , \22147 , \28502 );
and \U$28258 ( \28504 , \21930 , \21935 );
not \U$28259 ( \28505 , \21930 );
and \U$28260 ( \28506 , \28505 , \21923 );
nor \U$28261 ( \28507 , \28504 , \28506 );
xnor \U$28262 ( \28508 , \28503 , \28507 );
not \U$28263 ( \28509 , \28508 );
or \U$28264 ( \28510 , \28497 , \28509 );
or \U$28265 ( \28511 , \28508 , \28496 );
nand \U$28266 ( \28512 , \28510 , \28511 );
xor \U$28267 ( \28513 , \21947 , \21948 );
xor \U$28268 ( \28514 , \28513 , \22144 );
xor \U$28269 ( \28515 , \28253 , \28239 );
xnor \U$28270 ( \28516 , \28515 , \28245 );
not \U$28271 ( \28517 , \28516 );
not \U$28272 ( \28518 , \28517 );
not \U$28273 ( \28519 , \22009 );
not \U$28274 ( \28520 , \22024 );
or \U$28275 ( \28521 , \28519 , \28520 );
not \U$28276 ( \28522 , \22009 );
nand \U$28277 ( \28523 , \28522 , \22023 );
nand \U$28278 ( \28524 , \28521 , \28523 );
not \U$28279 ( \28525 , \22016 );
and \U$28280 ( \28526 , \28524 , \28525 );
not \U$28281 ( \28527 , \28524 );
and \U$28282 ( \28528 , \28527 , \22016 );
nor \U$28283 ( \28529 , \28526 , \28528 );
not \U$28284 ( \28530 , \28529 );
not \U$28285 ( \28531 , \28530 );
or \U$28286 ( \28532 , \28518 , \28531 );
not \U$28287 ( \28533 , \28529 );
not \U$28288 ( \28534 , \28516 );
or \U$28289 ( \28535 , \28533 , \28534 );
not \U$28290 ( \28536 , \28434 );
not \U$28291 ( \28537 , \28429 );
or \U$28292 ( \28538 , \28536 , \28537 );
or \U$28293 ( \28539 , \28429 , \28434 );
nand \U$28294 ( \28540 , \28538 , \28539 );
and \U$28295 ( \28541 , \28540 , \28441 );
not \U$28296 ( \28542 , \28540 );
and \U$28297 ( \28543 , \28542 , \28440 );
nor \U$28298 ( \28544 , \28541 , \28543 );
nand \U$28299 ( \28545 , \28535 , \28544 );
nand \U$28300 ( \28546 , \28532 , \28545 );
not \U$28301 ( \28547 , \28450 );
and \U$28302 ( \28548 , \28458 , \28547 );
not \U$28303 ( \28549 , \28458 );
and \U$28304 ( \28550 , \28549 , \28450 );
nor \U$28305 ( \28551 , \28548 , \28550 );
not \U$28306 ( \28552 , \28551 );
xor \U$28307 ( \28553 , \28270 , \28265 );
xnor \U$28308 ( \28554 , \28553 , \28276 );
not \U$28309 ( \28555 , \28554 );
or \U$28310 ( \28556 , \28552 , \28555 );
xor \U$28311 ( \28557 , \28207 , \28201 );
xor \U$28312 ( \28558 , \28557 , \28196 );
nand \U$28313 ( \28559 , \28556 , \28558 );
not \U$28314 ( \28560 , \28554 );
not \U$28315 ( \28561 , \28551 );
nand \U$28316 ( \28562 , \28560 , \28561 );
nand \U$28317 ( \28563 , \28559 , \28562 );
xor \U$28318 ( \28564 , \28546 , \28563 );
not \U$28319 ( \28565 , \28422 );
not \U$28320 ( \28566 , \28463 );
or \U$28321 ( \28567 , \28565 , \28566 );
or \U$28322 ( \28568 , \28463 , \28422 );
nand \U$28323 ( \28569 , \28567 , \28568 );
and \U$28324 ( \28570 , \28564 , \28569 );
and \U$28325 ( \28571 , \28546 , \28563 );
or \U$28326 ( \28572 , \28570 , \28571 );
not \U$28327 ( \28573 , \28572 );
xor \U$28328 ( \28574 , \28210 , \28256 );
not \U$28329 ( \28575 , \28574 );
not \U$28330 ( \28576 , \22002 );
not \U$28331 ( \28577 , \28576 );
not \U$28332 ( \28578 , \22050 );
and \U$28333 ( \28579 , \28577 , \28578 );
and \U$28334 ( \28580 , \22050 , \28576 );
nor \U$28335 ( \28581 , \28579 , \28580 );
nand \U$28336 ( \28582 , \28575 , \28581 );
not \U$28337 ( \28583 , \28582 );
not \U$28338 ( \28584 , \28041 );
not \U$28339 ( \28585 , \28053 );
or \U$28340 ( \28586 , \28584 , \28585 );
nand \U$28341 ( \28587 , \28052 , \28046 );
nand \U$28342 ( \28588 , \28586 , \28587 );
not \U$28343 ( \28589 , \28588 );
not \U$28344 ( \28590 , \27876 );
not \U$28345 ( \28591 , \27869 );
or \U$28346 ( \28592 , \28590 , \28591 );
not \U$28347 ( \28593 , \27880 );
not \U$28348 ( \28594 , \27877 );
or \U$28349 ( \28595 , \28593 , \28594 );
nand \U$28350 ( \28596 , \28595 , \27888 );
nand \U$28351 ( \28597 , \28592 , \28596 );
not \U$28352 ( \28598 , \27984 );
not \U$28353 ( \28599 , \27977 );
or \U$28354 ( \28600 , \28598 , \28599 );
not \U$28355 ( \28601 , \27988 );
not \U$28356 ( \28602 , \27985 );
or \U$28357 ( \28603 , \28601 , \28602 );
nand \U$28358 ( \28604 , \28603 , \27998 );
nand \U$28359 ( \28605 , \28600 , \28604 );
xor \U$28360 ( \28606 , \28597 , \28605 );
not \U$28361 ( \28607 , \28606 );
or \U$28362 ( \28608 , \28589 , \28607 );
nand \U$28363 ( \28609 , \28605 , \28597 );
nand \U$28364 ( \28610 , \28608 , \28609 );
not \U$28365 ( \28611 , \28610 );
or \U$28366 ( \28612 , \28583 , \28611 );
not \U$28367 ( \28613 , \28581 );
nand \U$28368 ( \28614 , \28613 , \28574 );
nand \U$28369 ( \28615 , \28612 , \28614 );
not \U$28370 ( \28616 , \28615 );
or \U$28371 ( \28617 , \28573 , \28616 );
or \U$28372 ( \28618 , \28615 , \28572 );
not \U$28373 ( \28619 , \28392 );
not \U$28374 ( \28620 , \28408 );
or \U$28375 ( \28621 , \28619 , \28620 );
or \U$28376 ( \28622 , \28408 , \28392 );
nand \U$28377 ( \28623 , \28621 , \28622 );
xor \U$28378 ( \28624 , \22039 , \22033 );
xor \U$28379 ( \28625 , \28624 , \22046 );
xor \U$28380 ( \28626 , \28216 , \28223 );
xor \U$28381 ( \28627 , \28626 , \28231 );
or \U$28382 ( \28628 , \28625 , \28627 );
and \U$28383 ( \28629 , \21997 , \21980 );
not \U$28384 ( \28630 , \21997 );
not \U$28385 ( \28631 , \21980 );
and \U$28386 ( \28632 , \28630 , \28631 );
nor \U$28387 ( \28633 , \28629 , \28632 );
nand \U$28388 ( \28634 , \28628 , \28633 );
nand \U$28389 ( \28635 , \28625 , \28627 );
nand \U$28390 ( \28636 , \28634 , \28635 );
or \U$28391 ( \28637 , \28623 , \28636 );
not \U$28392 ( \28638 , \28327 );
and \U$28393 ( \28639 , \28301 , \28638 );
not \U$28394 ( \28640 , \28301 );
and \U$28395 ( \28641 , \28640 , \28327 );
or \U$28396 ( \28642 , \28639 , \28641 );
nand \U$28397 ( \28643 , \28637 , \28642 );
nand \U$28398 ( \28644 , \28623 , \28636 );
nand \U$28399 ( \28645 , \28643 , \28644 );
nand \U$28400 ( \28646 , \28618 , \28645 );
nand \U$28401 ( \28647 , \28617 , \28646 );
xor \U$28402 ( \28648 , \28344 , \28368 );
xor \U$28403 ( \28649 , \28648 , \28371 );
xor \U$28404 ( \28650 , \28647 , \28649 );
not \U$28405 ( \28651 , \28294 );
not \U$28406 ( \28652 , \28190 );
not \U$28407 ( \28653 , \28652 );
and \U$28408 ( \28654 , \28651 , \28653 );
and \U$28409 ( \28655 , \28294 , \28652 );
nor \U$28410 ( \28656 , \28654 , \28655 );
not \U$28411 ( \28657 , \28656 );
not \U$28412 ( \28658 , \28657 );
not \U$28413 ( \28659 , \21973 );
not \U$28414 ( \28660 , \28659 );
not \U$28415 ( \28661 , \22054 );
or \U$28416 ( \28662 , \28660 , \28661 );
or \U$28417 ( \28663 , \22054 , \28659 );
nand \U$28418 ( \28664 , \28662 , \28663 );
not \U$28419 ( \28665 , \28664 );
xor \U$28420 ( \28666 , \27939 , \27944 );
and \U$28421 ( \28667 , \28666 , \27950 );
and \U$28422 ( \28668 , \27939 , \27944 );
or \U$28423 ( \28669 , \28667 , \28668 );
not \U$28424 ( \28670 , \28669 );
not \U$28425 ( \28671 , \27962 );
not \U$28426 ( \28672 , \27956 );
or \U$28427 ( \28673 , \28671 , \28672 );
or \U$28428 ( \28674 , \27956 , \27962 );
nand \U$28429 ( \28675 , \28674 , \27969 );
nand \U$28430 ( \28676 , \28673 , \28675 );
not \U$28431 ( \28677 , \28676 );
or \U$28432 ( \28678 , \28024 , \28029 );
nand \U$28433 ( \28679 , \28678 , \28018 );
nand \U$28434 ( \28680 , \28024 , \28029 );
nand \U$28435 ( \28681 , \28679 , \28680 );
not \U$28436 ( \28682 , \28681 );
not \U$28437 ( \28683 , \28682 );
or \U$28438 ( \28684 , \28677 , \28683 );
or \U$28439 ( \28685 , \28682 , \28676 );
nand \U$28440 ( \28686 , \28684 , \28685 );
not \U$28441 ( \28687 , \28686 );
or \U$28442 ( \28688 , \28670 , \28687 );
nand \U$28443 ( \28689 , \28676 , \28681 );
nand \U$28444 ( \28690 , \28688 , \28689 );
not \U$28445 ( \28691 , \28690 );
not \U$28446 ( \28692 , \27923 );
not \U$28447 ( \28693 , \27918 );
or \U$28448 ( \28694 , \28692 , \28693 );
not \U$28449 ( \28695 , \27907 );
nand \U$28450 ( \28696 , \28695 , \27914 );
nand \U$28451 ( \28697 , \28694 , \28696 );
not \U$28452 ( \28698 , \27687 );
not \U$28453 ( \28699 , \27681 );
or \U$28454 ( \28700 , \28698 , \28699 );
or \U$28455 ( \28701 , \27681 , \27687 );
nand \U$28456 ( \28702 , \28701 , \27695 );
nand \U$28457 ( \28703 , \28700 , \28702 );
or \U$28458 ( \28704 , \28697 , \28703 );
not \U$28459 ( \28705 , \28060 );
not \U$28460 ( \28706 , \28077 );
or \U$28461 ( \28707 , \28705 , \28706 );
nand \U$28462 ( \28708 , \28073 , \28066 );
nand \U$28463 ( \28709 , \28707 , \28708 );
nand \U$28464 ( \28710 , \28704 , \28709 );
nand \U$28465 ( \28711 , \28697 , \28703 );
and \U$28466 ( \28712 , \28710 , \28711 );
nand \U$28467 ( \28713 , \28691 , \28712 );
xor \U$28468 ( \28714 , \28279 , \28287 );
buf \U$28469 ( \28715 , \28714 );
and \U$28470 ( \28716 , \28713 , \28715 );
nor \U$28471 ( \28717 , \28691 , \28712 );
nor \U$28472 ( \28718 , \28716 , \28717 );
not \U$28473 ( \28719 , \28718 );
or \U$28474 ( \28720 , \28665 , \28719 );
or \U$28475 ( \28721 , \28718 , \28664 );
nand \U$28476 ( \28722 , \28720 , \28721 );
not \U$28477 ( \28723 , \28722 );
or \U$28478 ( \28724 , \28658 , \28723 );
not \U$28479 ( \28725 , \28718 );
nand \U$28480 ( \28726 , \28725 , \28664 );
nand \U$28481 ( \28727 , \28724 , \28726 );
and \U$28482 ( \28728 , \28650 , \28727 );
and \U$28483 ( \28729 , \28647 , \28649 );
or \U$28484 ( \28730 , \28728 , \28729 );
xor \U$28485 ( \28731 , \28298 , \28337 );
xor \U$28486 ( \28732 , \28731 , \28340 );
not \U$28487 ( \28733 , \28345 );
xnor \U$28488 ( \28734 , \28365 , \28362 );
not \U$28489 ( \28735 , \28734 );
or \U$28490 ( \28736 , \28733 , \28735 );
or \U$28491 ( \28737 , \28734 , \28345 );
nand \U$28492 ( \28738 , \28736 , \28737 );
not \U$28493 ( \28739 , \28331 );
not \U$28494 ( \28740 , \28300 );
or \U$28495 ( \28741 , \28739 , \28740 );
or \U$28496 ( \28742 , \28300 , \28331 );
nand \U$28497 ( \28743 , \28741 , \28742 );
xor \U$28498 ( \28744 , \28743 , \28334 );
xor \U$28499 ( \28745 , \28738 , \28744 );
xor \U$28500 ( \28746 , \28467 , \28413 );
xor \U$28501 ( \28747 , \28746 , \28416 );
and \U$28502 ( \28748 , \28745 , \28747 );
and \U$28503 ( \28749 , \28738 , \28744 );
or \U$28504 ( \28750 , \28748 , \28749 );
xor \U$28505 ( \28751 , \28732 , \28750 );
xor \U$28506 ( \28752 , \28482 , \28389 );
xor \U$28507 ( \28753 , \28752 , \28476 );
and \U$28508 ( \28754 , \28751 , \28753 );
and \U$28509 ( \28755 , \28732 , \28750 );
or \U$28510 ( \28756 , \28754 , \28755 );
xor \U$28511 ( \28757 , \28730 , \28756 );
xor \U$28512 ( \28758 , \28184 , \28375 );
and \U$28513 ( \28759 , \28757 , \28758 );
and \U$28514 ( \28760 , \28730 , \28756 );
or \U$28515 ( \28761 , \28759 , \28760 );
xor \U$28516 ( \28762 , \28514 , \28761 );
xor \U$28517 ( \28763 , \28183 , \28379 );
xor \U$28518 ( \28764 , \28763 , \28492 );
and \U$28519 ( \28765 , \28762 , \28764 );
and \U$28520 ( \28766 , \28514 , \28761 );
or \U$28521 ( \28767 , \28765 , \28766 );
not \U$28522 ( \28768 , \28767 );
nand \U$28523 ( \28769 , \28512 , \28768 );
xor \U$28524 ( \28770 , \28514 , \28761 );
xor \U$28525 ( \28771 , \28770 , \28764 );
not \U$28526 ( \28772 , \28771 );
xor \U$28527 ( \28773 , \28490 , \28387 );
xnor \U$28528 ( \28774 , \28773 , \28485 );
not \U$28529 ( \28775 , \28774 );
not \U$28530 ( \28776 , \28775 );
xor \U$28531 ( \28777 , \28636 , \28642 );
xor \U$28532 ( \28778 , \28777 , \28623 );
not \U$28533 ( \28779 , \28778 );
xor \U$28534 ( \28780 , \28574 , \28581 );
xnor \U$28535 ( \28781 , \28780 , \28610 );
and \U$28536 ( \28782 , \28544 , \28517 );
not \U$28537 ( \28783 , \28544 );
and \U$28538 ( \28784 , \28783 , \28516 );
or \U$28539 ( \28785 , \28782 , \28784 );
and \U$28540 ( \28786 , \28785 , \28529 );
not \U$28541 ( \28787 , \28785 );
and \U$28542 ( \28788 , \28787 , \28530 );
nor \U$28543 ( \28789 , \28786 , \28788 );
xor \U$28544 ( \28790 , \28703 , \28697 );
xor \U$28545 ( \28791 , \28790 , \28709 );
or \U$28546 ( \28792 , \28789 , \28791 );
or \U$28547 ( \28793 , \28625 , \28627 );
nand \U$28548 ( \28794 , \28793 , \28635 );
not \U$28549 ( \28795 , \28633 );
and \U$28550 ( \28796 , \28794 , \28795 );
not \U$28551 ( \28797 , \28794 );
and \U$28552 ( \28798 , \28797 , \28633 );
nor \U$28553 ( \28799 , \28796 , \28798 );
nand \U$28554 ( \28800 , \28792 , \28799 );
nand \U$28555 ( \28801 , \28789 , \28791 );
nand \U$28556 ( \28802 , \28800 , \28801 );
and \U$28557 ( \28803 , \28781 , \28802 );
not \U$28558 ( \28804 , \28781 );
not \U$28559 ( \28805 , \28802 );
and \U$28560 ( \28806 , \28804 , \28805 );
nor \U$28561 ( \28807 , \28803 , \28806 );
not \U$28562 ( \28808 , \28807 );
or \U$28563 ( \28809 , \28779 , \28808 );
not \U$28564 ( \28810 , \28805 );
nand \U$28565 ( \28811 , \28810 , \28781 );
nand \U$28566 ( \28812 , \28809 , \28811 );
xor \U$28567 ( \28813 , \28572 , \28615 );
buf \U$28568 ( \28814 , \28645 );
and \U$28569 ( \28815 , \28813 , \28814 );
not \U$28570 ( \28816 , \28813 );
not \U$28571 ( \28817 , \28814 );
and \U$28572 ( \28818 , \28816 , \28817 );
nor \U$28573 ( \28819 , \28815 , \28818 );
xor \U$28574 ( \28820 , \28812 , \28819 );
xor \U$28575 ( \28821 , \28738 , \28744 );
xor \U$28576 ( \28822 , \28821 , \28747 );
and \U$28577 ( \28823 , \28820 , \28822 );
and \U$28578 ( \28824 , \28812 , \28819 );
nor \U$28579 ( \28825 , \28823 , \28824 );
not \U$28580 ( \28826 , \28825 );
not \U$28581 ( \28827 , \27970 );
not \U$28582 ( \28828 , \27951 );
or \U$28583 ( \28829 , \28827 , \28828 );
or \U$28584 ( \28830 , \27951 , \27970 );
nand \U$28585 ( \28831 , \28830 , \28003 );
nand \U$28586 ( \28832 , \28829 , \28831 );
not \U$28587 ( \28833 , \28832 );
not \U$28588 ( \28834 , \27900 );
not \U$28589 ( \28835 , \27889 );
or \U$28590 ( \28836 , \28834 , \28835 );
or \U$28591 ( \28837 , \27889 , \27900 );
nand \U$28592 ( \28838 , \28837 , \27928 );
nand \U$28593 ( \28839 , \28836 , \28838 );
not \U$28594 ( \28840 , \28839 );
or \U$28595 ( \28841 , \28833 , \28840 );
not \U$28596 ( \28842 , \28839 );
not \U$28597 ( \28843 , \28842 );
not \U$28598 ( \28844 , \28832 );
not \U$28599 ( \28845 , \28844 );
or \U$28600 ( \28846 , \28843 , \28845 );
xor \U$28601 ( \28847 , \28035 , \28054 );
and \U$28602 ( \28848 , \28847 , \28078 );
and \U$28603 ( \28849 , \28035 , \28054 );
or \U$28604 ( \28850 , \28848 , \28849 );
nand \U$28605 ( \28851 , \28846 , \28850 );
nand \U$28606 ( \28852 , \28841 , \28851 );
not \U$28607 ( \28853 , \28852 );
not \U$28608 ( \28854 , \28588 );
not \U$28609 ( \28855 , \28854 );
not \U$28610 ( \28856 , \28606 );
or \U$28611 ( \28857 , \28855 , \28856 );
or \U$28612 ( \28858 , \28606 , \28854 );
nand \U$28613 ( \28859 , \28857 , \28858 );
not \U$28614 ( \28860 , \28859 );
nor \U$28615 ( \28861 , \27787 , \27775 );
or \U$28616 ( \28862 , \28861 , \27767 );
nand \U$28617 ( \28863 , \27787 , \27775 );
nand \U$28618 ( \28864 , \28862 , \28863 );
not \U$28619 ( \28865 , \28864 );
not \U$28620 ( \28866 , \28669 );
and \U$28621 ( \28867 , \28686 , \28866 );
not \U$28622 ( \28868 , \28686 );
and \U$28623 ( \28869 , \28868 , \28669 );
nor \U$28624 ( \28870 , \28867 , \28869 );
nand \U$28625 ( \28871 , \28865 , \28870 );
not \U$28626 ( \28872 , \28871 );
or \U$28627 ( \28873 , \28860 , \28872 );
not \U$28628 ( \28874 , \28870 );
nand \U$28629 ( \28875 , \28874 , \28864 );
nand \U$28630 ( \28876 , \28873 , \28875 );
not \U$28631 ( \28877 , \28876 );
or \U$28632 ( \28878 , \28853 , \28877 );
or \U$28633 ( \28879 , \28876 , \28852 );
xor \U$28634 ( \28880 , \28546 , \28563 );
xor \U$28635 ( \28881 , \28880 , \28569 );
nand \U$28636 ( \28882 , \28879 , \28881 );
nand \U$28637 ( \28883 , \28878 , \28882 );
not \U$28638 ( \28884 , \28883 );
not \U$28639 ( \28885 , \28722 );
not \U$28640 ( \28886 , \28656 );
and \U$28641 ( \28887 , \28885 , \28886 );
and \U$28642 ( \28888 , \28722 , \28656 );
nor \U$28643 ( \28889 , \28887 , \28888 );
xor \U$28644 ( \28890 , \28884 , \28889 );
xor \U$28645 ( \28891 , \28355 , \28360 );
xor \U$28646 ( \28892 , \28891 , \28347 );
xor \U$28647 ( \28893 , \27855 , \27859 );
and \U$28648 ( \28894 , \28893 , \27862 );
and \U$28649 ( \28895 , \27855 , \27859 );
or \U$28650 ( \28896 , \28894 , \28895 );
not \U$28651 ( \28897 , \28896 );
xor \U$28652 ( \28898 , \28312 , \28307 );
xnor \U$28653 ( \28899 , \28898 , \27766 );
not \U$28654 ( \28900 , \28899 );
not \U$28655 ( \28901 , \28900 );
not \U$28656 ( \28902 , \27808 );
not \U$28657 ( \28903 , \27814 );
or \U$28658 ( \28904 , \28902 , \28903 );
nand \U$28659 ( \28905 , \27802 , \27807 );
nand \U$28660 ( \28906 , \28904 , \28905 );
not \U$28661 ( \28907 , \28906 );
or \U$28662 ( \28908 , \28901 , \28907 );
or \U$28663 ( \28909 , \28906 , \28900 );
nand \U$28664 ( \28910 , \28908 , \28909 );
not \U$28665 ( \28911 , \28910 );
or \U$28666 ( \28912 , \28897 , \28911 );
nand \U$28667 ( \28913 , \28906 , \28899 );
nand \U$28668 ( \28914 , \28912 , \28913 );
xor \U$28669 ( \28915 , \28892 , \28914 );
xor \U$28670 ( \28916 , \28714 , \28691 );
xor \U$28671 ( \28917 , \28916 , \28712 );
and \U$28672 ( \28918 , \28915 , \28917 );
and \U$28673 ( \28919 , \28892 , \28914 );
nor \U$28674 ( \28920 , \28918 , \28919 );
and \U$28675 ( \28921 , \28890 , \28920 );
and \U$28676 ( \28922 , \28884 , \28889 );
or \U$28677 ( \28923 , \28921 , \28922 );
not \U$28678 ( \28924 , \28923 );
not \U$28679 ( \28925 , \28924 );
xor \U$28680 ( \28926 , \28647 , \28649 );
xor \U$28681 ( \28927 , \28926 , \28727 );
not \U$28682 ( \28928 , \28927 );
not \U$28683 ( \28929 , \28928 );
or \U$28684 ( \28930 , \28925 , \28929 );
nand \U$28685 ( \28931 , \28923 , \28927 );
nand \U$28686 ( \28932 , \28930 , \28931 );
not \U$28687 ( \28933 , \28932 );
or \U$28688 ( \28934 , \28826 , \28933 );
not \U$28689 ( \28935 , \28927 );
nand \U$28690 ( \28936 , \28935 , \28923 );
nand \U$28691 ( \28937 , \28934 , \28936 );
not \U$28692 ( \28938 , \28937 );
not \U$28693 ( \28939 , \28938 );
or \U$28694 ( \28940 , \28776 , \28939 );
not \U$28695 ( \28941 , \28774 );
not \U$28696 ( \28942 , \28937 );
or \U$28697 ( \28943 , \28941 , \28942 );
xor \U$28698 ( \28944 , \28730 , \28756 );
xor \U$28699 ( \28945 , \28944 , \28758 );
nand \U$28700 ( \28946 , \28943 , \28945 );
nand \U$28701 ( \28947 , \28940 , \28946 );
not \U$28702 ( \28948 , \28947 );
nand \U$28703 ( \28949 , \28772 , \28948 );
not \U$28704 ( \28950 , \22155 );
not \U$28705 ( \28951 , \22151 );
not \U$28706 ( \28952 , \22149 );
or \U$28707 ( \28953 , \28951 , \28952 );
or \U$28708 ( \28954 , \22149 , \22151 );
nand \U$28709 ( \28955 , \28953 , \28954 );
not \U$28710 ( \28956 , \28955 );
or \U$28711 ( \28957 , \28950 , \28956 );
or \U$28712 ( \28958 , \22155 , \28955 );
nand \U$28713 ( \28959 , \28957 , \28958 );
not \U$28714 ( \28960 , \28495 );
not \U$28715 ( \28961 , \22147 );
not \U$28716 ( \28962 , \28961 );
not \U$28717 ( \28963 , \28507 );
or \U$28718 ( \28964 , \28962 , \28963 );
or \U$28719 ( \28965 , \28961 , \28507 );
nand \U$28720 ( \28966 , \28964 , \28965 );
nand \U$28721 ( \28967 , \28966 , \28502 );
not \U$28722 ( \28968 , \28967 );
or \U$28723 ( \28969 , \28960 , \28968 );
not \U$28724 ( \28970 , \28966 );
not \U$28725 ( \28971 , \28502 );
nand \U$28726 ( \28972 , \28970 , \28971 );
nand \U$28727 ( \28973 , \28969 , \28972 );
not \U$28728 ( \28974 , \28973 );
nand \U$28729 ( \28975 , \28959 , \28974 );
not \U$28730 ( \28976 , \28932 );
not \U$28731 ( \28977 , \28825 );
not \U$28732 ( \28978 , \28977 );
and \U$28733 ( \28979 , \28976 , \28978 );
and \U$28734 ( \28980 , \28977 , \28932 );
nor \U$28735 ( \28981 , \28979 , \28980 );
not \U$28736 ( \28982 , \28881 );
not \U$28737 ( \28983 , \28982 );
xor \U$28738 ( \28984 , \28852 , \28876 );
not \U$28739 ( \28985 , \28984 );
or \U$28740 ( \28986 , \28983 , \28985 );
or \U$28741 ( \28987 , \28984 , \28982 );
nand \U$28742 ( \28988 , \28986 , \28987 );
not \U$28743 ( \28989 , \28791 );
not \U$28744 ( \28990 , \28989 );
not \U$28745 ( \28991 , \28789 );
not \U$28746 ( \28992 , \28991 );
or \U$28747 ( \28993 , \28990 , \28992 );
nand \U$28748 ( \28994 , \28993 , \28801 );
not \U$28749 ( \28995 , \28799 );
and \U$28750 ( \28996 , \28994 , \28995 );
not \U$28751 ( \28997 , \28994 );
and \U$28752 ( \28998 , \28997 , \28799 );
nor \U$28753 ( \28999 , \28996 , \28998 );
not \U$28754 ( \29000 , \28999 );
nand \U$28755 ( \29001 , \28875 , \28871 );
xor \U$28756 ( \29002 , \29001 , \28859 );
not \U$28757 ( \29003 , \29002 );
xor \U$28758 ( \29004 , \27863 , \27933 );
and \U$28759 ( \29005 , \29004 , \28004 );
and \U$28760 ( \29006 , \27863 , \27933 );
or \U$28761 ( \29007 , \29005 , \29006 );
not \U$28762 ( \29008 , \29007 );
or \U$28763 ( \29009 , \29003 , \29008 );
or \U$28764 ( \29010 , \29007 , \29002 );
nand \U$28765 ( \29011 , \29009 , \29010 );
not \U$28766 ( \29012 , \29011 );
or \U$28767 ( \29013 , \29000 , \29012 );
not \U$28768 ( \29014 , \29002 );
nand \U$28769 ( \29015 , \29014 , \29007 );
nand \U$28770 ( \29016 , \29013 , \29015 );
xor \U$28771 ( \29017 , \28988 , \29016 );
xor \U$28772 ( \29018 , \28778 , \28807 );
and \U$28773 ( \29019 , \29017 , \29018 );
and \U$28774 ( \29020 , \28988 , \29016 );
or \U$28775 ( \29021 , \29019 , \29020 );
not \U$28776 ( \29022 , \29021 );
xor \U$28777 ( \29023 , \28884 , \28889 );
xor \U$28778 ( \29024 , \29023 , \28920 );
not \U$28779 ( \29025 , \29024 );
not \U$28780 ( \29026 , \29025 );
or \U$28781 ( \29027 , \29022 , \29026 );
not \U$28782 ( \29028 , \27700 );
not \U$28783 ( \29029 , \27675 );
not \U$28784 ( \29030 , \29029 );
or \U$28785 ( \29031 , \29028 , \29030 );
nand \U$28786 ( \29032 , \29031 , \27711 );
nand \U$28787 ( \29033 , \27675 , \27701 );
and \U$28788 ( \29034 , \29032 , \29033 );
not \U$28789 ( \29035 , \28551 );
not \U$28790 ( \29036 , \28554 );
or \U$28791 ( \29037 , \29035 , \29036 );
nand \U$28792 ( \29038 , \29037 , \28562 );
not \U$28793 ( \29039 , \28558 );
and \U$28794 ( \29040 , \29038 , \29039 );
not \U$28795 ( \29041 , \29038 );
and \U$28796 ( \29042 , \29041 , \28558 );
nor \U$28797 ( \29043 , \29040 , \29042 );
xor \U$28798 ( \29044 , \29034 , \29043 );
not \U$28799 ( \29045 , \29044 );
not \U$28800 ( \29046 , \29045 );
not \U$28801 ( \29047 , \28896 );
xor \U$28802 ( \29048 , \28899 , \29047 );
xnor \U$28803 ( \29049 , \29048 , \28906 );
not \U$28804 ( \29050 , \29049 );
or \U$28805 ( \29051 , \29046 , \29050 );
not \U$28806 ( \29052 , \29034 );
nand \U$28807 ( \29053 , \29052 , \29043 );
nand \U$28808 ( \29054 , \29051 , \29053 );
and \U$28809 ( \29055 , \28844 , \28842 );
not \U$28810 ( \29056 , \28844 );
and \U$28811 ( \29057 , \29056 , \28839 );
nor \U$28812 ( \29058 , \29055 , \29057 );
xor \U$28813 ( \29059 , \28850 , \29058 );
not \U$28814 ( \29060 , \29059 );
or \U$28815 ( \29061 , \27725 , \27729 );
not \U$28816 ( \29062 , \29061 );
not \U$28817 ( \29063 , \27736 );
or \U$28818 ( \29064 , \29062 , \29063 );
nand \U$28819 ( \29065 , \27725 , \27729 );
nand \U$28820 ( \29066 , \29064 , \29065 );
or \U$28821 ( \29067 , \27793 , \27819 );
nand \U$28822 ( \29068 , \29067 , \27795 );
and \U$28823 ( \29069 , \29066 , \29068 );
not \U$28824 ( \29070 , \29066 );
not \U$28825 ( \29071 , \29068 );
and \U$28826 ( \29072 , \29070 , \29071 );
nor \U$28827 ( \29073 , \29069 , \29072 );
not \U$28828 ( \29074 , \29073 );
or \U$28829 ( \29075 , \29060 , \29074 );
not \U$28830 ( \29076 , \29071 );
nand \U$28831 ( \29077 , \29076 , \29066 );
nand \U$28832 ( \29078 , \29075 , \29077 );
and \U$28833 ( \29079 , \29054 , \29078 );
not \U$28834 ( \29080 , \29079 );
not \U$28835 ( \29081 , \29080 );
xor \U$28836 ( \29082 , \28892 , \28914 );
xor \U$28837 ( \29083 , \29082 , \28917 );
xor \U$28838 ( \29084 , \29054 , \29078 );
and \U$28839 ( \29085 , \29083 , \29084 );
not \U$28840 ( \29086 , \29085 );
not \U$28841 ( \29087 , \29086 );
or \U$28842 ( \29088 , \29081 , \29087 );
or \U$28843 ( \29089 , \29025 , \29021 );
nand \U$28844 ( \29090 , \29088 , \29089 );
nand \U$28845 ( \29091 , \29027 , \29090 );
or \U$28846 ( \29092 , \28981 , \29091 );
xor \U$28847 ( \29093 , \28732 , \28750 );
xor \U$28848 ( \29094 , \29093 , \28753 );
nand \U$28849 ( \29095 , \29092 , \29094 );
nand \U$28850 ( \29096 , \28981 , \29091 );
nand \U$28851 ( \29097 , \29095 , \29096 );
not \U$28852 ( \29098 , \29097 );
xor \U$28853 ( \29099 , \28774 , \28937 );
xnor \U$28854 ( \29100 , \29099 , \28945 );
nand \U$28855 ( \29101 , \29098 , \29100 );
and \U$28856 ( \29102 , \28769 , \28949 , \28975 , \29101 );
not \U$28857 ( \29103 , \29021 );
and \U$28858 ( \29104 , \28820 , \28822 );
not \U$28859 ( \29105 , \28820 );
not \U$28860 ( \29106 , \28822 );
and \U$28861 ( \29107 , \29105 , \29106 );
nor \U$28862 ( \29108 , \29104 , \29107 );
xor \U$28863 ( \29109 , \29103 , \29108 );
nor \U$28864 ( \29110 , \29085 , \29079 );
not \U$28865 ( \29111 , \29110 );
not \U$28866 ( \29112 , \29025 );
or \U$28867 ( \29113 , \29111 , \29112 );
not \U$28868 ( \29114 , \29080 );
not \U$28869 ( \29115 , \29086 );
or \U$28870 ( \29116 , \29114 , \29115 );
nand \U$28871 ( \29117 , \29116 , \29024 );
nand \U$28872 ( \29118 , \29113 , \29117 );
xnor \U$28873 ( \29119 , \29109 , \29118 );
xor \U$28874 ( \29120 , \27750 , \27820 );
and \U$28875 ( \29121 , \29120 , \27828 );
and \U$28876 ( \29122 , \27750 , \27820 );
or \U$28877 ( \29123 , \29121 , \29122 );
not \U$28878 ( \29124 , \29123 );
buf \U$28879 ( \29125 , \29073 );
not \U$28880 ( \29126 , \29059 );
and \U$28881 ( \29127 , \29125 , \29126 );
not \U$28882 ( \29128 , \29125 );
and \U$28883 ( \29129 , \29128 , \29059 );
nor \U$28884 ( \29130 , \29127 , \29129 );
not \U$28885 ( \29131 , \29130 );
not \U$28886 ( \29132 , \29131 );
xor \U$28887 ( \29133 , \28999 , \29011 );
not \U$28888 ( \29134 , \29133 );
not \U$28889 ( \29135 , \29134 );
or \U$28890 ( \29136 , \29132 , \29135 );
nand \U$28891 ( \29137 , \29133 , \29130 );
nand \U$28892 ( \29138 , \29136 , \29137 );
not \U$28893 ( \29139 , \29138 );
or \U$28894 ( \29140 , \29124 , \29139 );
nand \U$28895 ( \29141 , \29133 , \29131 );
nand \U$28896 ( \29142 , \29140 , \29141 );
not \U$28897 ( \29143 , \29142 );
nor \U$28898 ( \29144 , \27720 , \27716 );
or \U$28899 ( \29145 , \27737 , \29144 );
nand \U$28900 ( \29146 , \27720 , \27716 );
nand \U$28901 ( \29147 , \29145 , \29146 );
not \U$28902 ( \29148 , \29147 );
not \U$28903 ( \29149 , \29044 );
not \U$28904 ( \29150 , \29049 );
and \U$28905 ( \29151 , \29149 , \29150 );
and \U$28906 ( \29152 , \29049 , \29044 );
nor \U$28907 ( \29153 , \29151 , \29152 );
not \U$28908 ( \29154 , \29153 );
not \U$28909 ( \29155 , \29154 );
not \U$28910 ( \29156 , \28086 );
not \U$28911 ( \29157 , \28013 );
or \U$28912 ( \29158 , \29156 , \29157 );
nand \U$28913 ( \29159 , \28079 , \28085 );
nand \U$28914 ( \29160 , \29158 , \29159 );
not \U$28915 ( \29161 , \29160 );
not \U$28916 ( \29162 , \29161 );
or \U$28917 ( \29163 , \29155 , \29162 );
nand \U$28918 ( \29164 , \29153 , \29160 );
nand \U$28919 ( \29165 , \29163 , \29164 );
not \U$28920 ( \29166 , \29165 );
or \U$28921 ( \29167 , \29148 , \29166 );
nand \U$28922 ( \29168 , \29154 , \29160 );
nand \U$28923 ( \29169 , \29167 , \29168 );
not \U$28924 ( \29170 , \29169 );
xor \U$28925 ( \29171 , \29083 , \29084 );
xnor \U$28926 ( \29172 , \29170 , \29171 );
not \U$28927 ( \29173 , \29172 );
or \U$28928 ( \29174 , \29143 , \29173 );
not \U$28929 ( \29175 , \29170 );
nand \U$28930 ( \29176 , \29175 , \29171 );
nand \U$28931 ( \29177 , \29174 , \29176 );
not \U$28932 ( \29178 , \29177 );
and \U$28933 ( \29179 , \29119 , \29178 );
not \U$28934 ( \29180 , \29119 );
and \U$28935 ( \29181 , \29180 , \29177 );
nor \U$28936 ( \29182 , \29179 , \29181 );
xor \U$28937 ( \29183 , \27738 , \27745 );
and \U$28938 ( \29184 , \29183 , \27829 );
and \U$28939 ( \29185 , \27738 , \27745 );
or \U$28940 ( \29186 , \29184 , \29185 );
not \U$28941 ( \29187 , \29186 );
not \U$28942 ( \29188 , \29147 );
xor \U$28943 ( \29189 , \29188 , \29165 );
xor \U$28944 ( \29190 , \28005 , \28007 );
and \U$28945 ( \29191 , \29190 , \28087 );
and \U$28946 ( \29192 , \28005 , \28007 );
or \U$28947 ( \29193 , \29191 , \29192 );
xnor \U$28948 ( \29194 , \29189 , \29193 );
not \U$28949 ( \29195 , \29194 );
or \U$28950 ( \29196 , \29187 , \29195 );
nand \U$28951 ( \29197 , \29165 , \29188 );
not \U$28952 ( \29198 , \29197 );
not \U$28953 ( \29199 , \29165 );
nand \U$28954 ( \29200 , \29199 , \29147 );
not \U$28955 ( \29201 , \29200 );
or \U$28956 ( \29202 , \29198 , \29201 );
nand \U$28957 ( \29203 , \29202 , \29193 );
nand \U$28958 ( \29204 , \29196 , \29203 );
not \U$28959 ( \29205 , \29204 );
not \U$28960 ( \29206 , \29205 );
xor \U$28961 ( \29207 , \28988 , \29016 );
xor \U$28962 ( \29208 , \29207 , \29018 );
nand \U$28963 ( \29209 , \29206 , \29208 );
not \U$28964 ( \29210 , \29209 );
xor \U$28965 ( \29211 , \29170 , \29171 );
xnor \U$28966 ( \29212 , \29211 , \29142 );
not \U$28967 ( \29213 , \29212 );
not \U$28968 ( \29214 , \29213 );
or \U$28969 ( \29215 , \29210 , \29214 );
or \U$28970 ( \29216 , \29206 , \29208 );
nand \U$28971 ( \29217 , \29215 , \29216 );
nand \U$28972 ( \29218 , \29182 , \29217 );
not \U$28973 ( \29219 , \29103 );
not \U$28974 ( \29220 , \29219 );
not \U$28975 ( \29221 , \29118 );
or \U$28976 ( \29222 , \29220 , \29221 );
or \U$28977 ( \29223 , \29118 , \29219 );
nand \U$28978 ( \29224 , \29222 , \29223 );
not \U$28979 ( \29225 , \29224 );
not \U$28980 ( \29226 , \29225 );
not \U$28981 ( \29227 , \29108 );
not \U$28982 ( \29228 , \29227 );
not \U$28983 ( \29229 , \29228 );
or \U$28984 ( \29230 , \29226 , \29229 );
not \U$28985 ( \29231 , \29224 );
not \U$28986 ( \29232 , \29227 );
or \U$28987 ( \29233 , \29231 , \29232 );
nand \U$28988 ( \29234 , \29233 , \29177 );
nand \U$28989 ( \29235 , \29230 , \29234 );
not \U$28990 ( \29236 , \29235 );
xor \U$28991 ( \29237 , \29094 , \29091 );
xnor \U$28992 ( \29238 , \29237 , \28981 );
nand \U$28993 ( \29239 , \29236 , \29238 );
and \U$28994 ( \29240 , \29208 , \29204 );
not \U$28995 ( \29241 , \29208 );
and \U$28996 ( \29242 , \29241 , \29205 );
nor \U$28997 ( \29243 , \29240 , \29242 );
not \U$28998 ( \29244 , \29243 );
not \U$28999 ( \29245 , \29213 );
or \U$29000 ( \29246 , \29244 , \29245 );
not \U$29001 ( \29247 , \29243 );
nand \U$29002 ( \29248 , \29247 , \29212 );
nand \U$29003 ( \29249 , \29246 , \29248 );
not \U$29004 ( \29250 , \29249 );
xor \U$29005 ( \29251 , \27846 , \28088 );
and \U$29006 ( \29252 , \29251 , \28094 );
and \U$29007 ( \29253 , \27846 , \28088 );
or \U$29008 ( \29254 , \29252 , \29253 );
xor \U$29009 ( \29255 , \29123 , \29138 );
xor \U$29010 ( \29256 , \29254 , \29255 );
xor \U$29011 ( \29257 , \29194 , \29186 );
and \U$29012 ( \29258 , \29256 , \29257 );
and \U$29013 ( \29259 , \29254 , \29255 );
or \U$29014 ( \29260 , \29258 , \29259 );
not \U$29015 ( \29261 , \29260 );
nand \U$29016 ( \29262 , \29250 , \29261 );
xor \U$29017 ( \29263 , \29254 , \29255 );
xor \U$29018 ( \29264 , \29263 , \29257 );
not \U$29019 ( \29265 , \29264 );
nand \U$29020 ( \29266 , \27838 , \28095 );
nand \U$29021 ( \29267 , \27830 , \27833 );
and \U$29022 ( \29268 , \29266 , \29267 );
nand \U$29023 ( \29269 , \29265 , \29268 );
and \U$29024 ( \29270 , \29218 , \29239 , \29262 , \29269 );
nand \U$29025 ( \29271 , \29102 , \29270 );
nor \U$29026 ( \29272 , \28181 , \29271 );
not \U$29027 ( \29273 , \29102 );
not \U$29028 ( \29274 , \29260 );
not \U$29029 ( \29275 , \29249 );
or \U$29030 ( \29276 , \29274 , \29275 );
not \U$29031 ( \29277 , \29267 );
not \U$29032 ( \29278 , \29266 );
or \U$29033 ( \29279 , \29277 , \29278 );
nand \U$29034 ( \29280 , \29279 , \29264 );
nand \U$29035 ( \29281 , \29276 , \29280 );
nand \U$29036 ( \29282 , \29281 , \29218 , \29239 , \29262 );
nor \U$29037 ( \29283 , \29182 , \29217 );
and \U$29038 ( \29284 , \29239 , \29283 );
not \U$29039 ( \29285 , \29238 );
nand \U$29040 ( \29286 , \29285 , \29235 );
not \U$29041 ( \29287 , \29286 );
nor \U$29042 ( \29288 , \29284 , \29287 );
nand \U$29043 ( \29289 , \29282 , \29288 );
not \U$29044 ( \29290 , \29289 );
or \U$29045 ( \29291 , \29273 , \29290 );
not \U$29046 ( \29292 , \29100 );
nand \U$29047 ( \29293 , \29292 , \29097 );
nand \U$29048 ( \29294 , \28771 , \28947 );
and \U$29049 ( \29295 , \29293 , \29294 );
nand \U$29050 ( \29296 , \28949 , \28769 );
nor \U$29051 ( \29297 , \29295 , \29296 );
not \U$29052 ( \29298 , \28512 );
nand \U$29053 ( \29299 , \29298 , \28767 );
or \U$29054 ( \29300 , \28959 , \28974 );
nand \U$29055 ( \29301 , \29299 , \29300 );
or \U$29056 ( \29302 , \29297 , \29301 );
buf \U$29057 ( \29303 , \28975 );
nand \U$29058 ( \29304 , \29302 , \29303 );
nand \U$29059 ( \29305 , \29291 , \29304 );
nor \U$29060 ( \29306 , \29272 , \29305 );
xor \U$29061 ( \29307 , RIbe2a640_93, RIbe27e68_8);
not \U$29062 ( \29308 , \29307 );
not \U$29063 ( \29309 , \2459 );
or \U$29064 ( \29310 , \29308 , \29309 );
nand \U$29065 ( \29311 , \4447 , \25040 );
nand \U$29066 ( \29312 , \29310 , \29311 );
not \U$29067 ( \29313 , \29312 );
xor \U$29068 ( \29314 , RIbe28d68_40, RIbe2b180_117);
not \U$29069 ( \29315 , \29314 );
not \U$29070 ( \29316 , \15353 );
or \U$29071 ( \29317 , \29315 , \29316 );
nand \U$29072 ( \29318 , \16646 , \25250 );
nand \U$29073 ( \29319 , \29317 , \29318 );
xor \U$29074 ( \29320 , RIbe29128_48, RIbe2aaf0_103);
not \U$29075 ( \29321 , \29320 );
not \U$29076 ( \29322 , \28282 );
or \U$29077 ( \29323 , \29321 , \29322 );
nand \U$29078 ( \29324 , \25264 , RIbe2ab68_104);
nand \U$29079 ( \29325 , \29323 , \29324 );
xor \U$29080 ( \29326 , \29319 , \29325 );
not \U$29081 ( \29327 , \29326 );
or \U$29082 ( \29328 , \29313 , \29327 );
nand \U$29083 ( \29329 , \29319 , \29325 );
nand \U$29084 ( \29330 , \29328 , \29329 );
xor \U$29085 ( \29331 , RIbe2a550_91, RIbe29ec0_77);
not \U$29086 ( \29332 , \29331 );
not \U$29087 ( \29333 , \11999 );
or \U$29088 ( \29334 , \29332 , \29333 );
nand \U$29089 ( \29335 , \23306 , \25221 );
nand \U$29090 ( \29336 , \29334 , \29335 );
not \U$29091 ( \29337 , \29336 );
xor \U$29092 ( \29338 , RIbe2ae38_110, RIbe28b88_36);
not \U$29093 ( \29339 , \29338 );
not \U$29094 ( \29340 , \2553 );
or \U$29095 ( \29341 , \29339 , \29340 );
nand \U$29096 ( \29342 , \2559 , \25071 );
nand \U$29097 ( \29343 , \29341 , \29342 );
not \U$29098 ( \29344 , \29343 );
or \U$29099 ( \29345 , \29337 , \29344 );
or \U$29100 ( \29346 , \29343 , \29336 );
xor \U$29101 ( \29347 , RIbe2b108_116, RIbe298a8_64);
not \U$29102 ( \29348 , \29347 );
not \U$29103 ( \29349 , \25617 );
or \U$29104 ( \29350 , \29348 , \29349 );
nand \U$29105 ( \29351 , \23015 , \25058 );
nand \U$29106 ( \29352 , \29350 , \29351 );
nand \U$29107 ( \29353 , \29346 , \29352 );
nand \U$29108 ( \29354 , \29345 , \29353 );
nand \U$29109 ( \29355 , \29330 , \29354 );
not \U$29110 ( \29356 , \29355 );
not \U$29111 ( \29357 , \29330 );
not \U$29112 ( \29358 , \29354 );
and \U$29113 ( \29359 , \29357 , \29358 );
not \U$29114 ( \29360 , \25136 );
and \U$29115 ( \29361 , \25154 , \29360 );
not \U$29116 ( \29362 , \25154 );
and \U$29117 ( \29363 , \29362 , \25136 );
nor \U$29118 ( \29364 , \29361 , \29363 );
nor \U$29119 ( \29365 , \29359 , \29364 );
nor \U$29120 ( \29366 , \29356 , \29365 );
xor \U$29121 ( \29367 , \25243 , \25248 );
xor \U$29122 ( \29368 , \29367 , \25285 );
xor \U$29123 ( \29369 , \29366 , \29368 );
xor \U$29124 ( \29370 , \25038 , \25045 );
xor \U$29125 ( \29371 , \29370 , \25054 );
not \U$29126 ( \29372 , \29371 );
not \U$29127 ( \29373 , \25239 );
not \U$29128 ( \29374 , \25226 );
not \U$29129 ( \29375 , \29374 );
and \U$29130 ( \29376 , \29373 , \29375 );
and \U$29131 ( \29377 , \25239 , \29374 );
nor \U$29132 ( \29378 , \29376 , \29377 );
not \U$29133 ( \29379 , \29378 );
not \U$29134 ( \29380 , \29379 );
not \U$29135 ( \29381 , \25256 );
not \U$29136 ( \29382 , \25280 );
or \U$29137 ( \29383 , \29381 , \29382 );
or \U$29138 ( \29384 , \25280 , \25256 );
nand \U$29139 ( \29385 , \29383 , \29384 );
not \U$29140 ( \29386 , \29385 );
not \U$29141 ( \29387 , \29386 );
or \U$29142 ( \29388 , \29380 , \29387 );
nand \U$29143 ( \29389 , \29385 , \29378 );
nand \U$29144 ( \29390 , \29388 , \29389 );
not \U$29145 ( \29391 , \29390 );
or \U$29146 ( \29392 , \29372 , \29391 );
nand \U$29147 ( \29393 , \29385 , \29379 );
nand \U$29148 ( \29394 , \29392 , \29393 );
xor \U$29149 ( \29395 , \29369 , \29394 );
not \U$29150 ( \29396 , \29395 );
not \U$29151 ( \29397 , RIbe27c88_4);
not \U$29152 ( \29398 , RIbe2af28_112);
and \U$29153 ( \29399 , \29397 , \29398 );
and \U$29154 ( \29400 , RIbe27c88_4, RIbe2af28_112);
nor \U$29155 ( \29401 , \29399 , \29400 );
not \U$29156 ( \29402 , \29401 );
not \U$29157 ( \29403 , \15345 );
or \U$29158 ( \29404 , \29402 , \29403 );
and \U$29159 ( \29405 , RIbe27df0_7, RIbe2af28_112);
nor \U$29160 ( \29406 , RIbe27df0_7, RIbe2af28_112);
nor \U$29161 ( \29407 , \29405 , \29406 );
nand \U$29162 ( \29408 , \17811 , \29407 );
nand \U$29163 ( \29409 , \29404 , \29408 );
not \U$29164 ( \29410 , \29409 );
xor \U$29165 ( \29411 , RIbe2b540_125, RIbe28f48_44);
not \U$29166 ( \29412 , \29411 );
not \U$29167 ( \29413 , \8221 );
or \U$29168 ( \29414 , \29412 , \29413 );
xor \U$29169 ( \29415 , RIbe28f48_44, RIbe2ad48_108);
nand \U$29170 ( \29416 , \3249 , \29415 );
nand \U$29171 ( \29417 , \29414 , \29416 );
xor \U$29172 ( \29418 , RIbe2a550_91, RIbe29f38_78);
not \U$29173 ( \29419 , \29418 );
not \U$29174 ( \29420 , \10433 );
or \U$29175 ( \29421 , \29419 , \29420 );
nand \U$29176 ( \29422 , \11227 , \29331 );
nand \U$29177 ( \29423 , \29421 , \29422 );
xor \U$29178 ( \29424 , \29417 , \29423 );
not \U$29179 ( \29425 , \29424 );
or \U$29180 ( \29426 , \29410 , \29425 );
nand \U$29181 ( \29427 , \29423 , \29417 );
nand \U$29182 ( \29428 , \29426 , \29427 );
not \U$29183 ( \29429 , \29428 );
xor \U$29184 ( \29430 , RIbe2aa78_102, RIbe2a910_99);
not \U$29185 ( \29431 , \29430 );
not \U$29186 ( \29432 , \9736 );
or \U$29187 ( \29433 , \29431 , \29432 );
xor \U$29188 ( \29434 , RIbe2b6a8_128, RIbe2a910_99);
nand \U$29189 ( \29435 , \10400 , \29434 );
nand \U$29190 ( \29436 , \29433 , \29435 );
xor \U$29191 ( \29437 , RIbe29b78_70, RIbe2a280_85);
not \U$29192 ( \29438 , \29437 );
not \U$29193 ( \29439 , \13268 );
or \U$29194 ( \29440 , \29438 , \29439 );
xor \U$29195 ( \29441 , RIbe2a280_85, RIbe27b20_1);
nand \U$29196 ( \29442 , \18667 , \29441 );
nand \U$29197 ( \29443 , \29440 , \29442 );
or \U$29198 ( \29444 , \29436 , \29443 );
xor \U$29199 ( \29445 , RIbe29e48_76, RIbe2a4d8_90);
not \U$29200 ( \29446 , \29445 );
not \U$29201 ( \29447 , \16652 );
or \U$29202 ( \29448 , \29446 , \29447 );
xor \U$29203 ( \29449 , RIbe2b2e8_120, RIbe29e48_76);
nand \U$29204 ( \29450 , \4849 , \29449 );
nand \U$29205 ( \29451 , \29448 , \29450 );
nand \U$29206 ( \29452 , \29444 , \29451 );
nand \U$29207 ( \29453 , \29436 , \29443 );
nand \U$29208 ( \29454 , \29452 , \29453 );
not \U$29209 ( \29455 , \29454 );
not \U$29210 ( \29456 , \29455 );
xor \U$29211 ( \29457 , RIbe2b018_114, RIbe29218_50);
not \U$29212 ( \29458 , \29457 );
not \U$29213 ( \29459 , \16811 );
or \U$29214 ( \29460 , \29458 , \29459 );
xor \U$29215 ( \29461 , RIbe2b018_114, RIbe29a10_67);
nand \U$29216 ( \29462 , \18777 , \29461 );
nand \U$29217 ( \29463 , \29460 , \29462 );
not \U$29218 ( \29464 , \29463 );
xor \U$29219 ( \29465 , RIbe2b360_121, RIbe2a028_80);
not \U$29220 ( \29466 , \29465 );
not \U$29221 ( \29467 , \8169 );
or \U$29222 ( \29468 , \29466 , \29467 );
xor \U$29223 ( \29469 , RIbe2a0a0_81, RIbe2a028_80);
nand \U$29224 ( \29470 , \8930 , \29469 );
nand \U$29225 ( \29471 , \29468 , \29470 );
not \U$29226 ( \29472 , \29471 );
or \U$29227 ( \29473 , \29464 , \29472 );
or \U$29228 ( \29474 , \29471 , \29463 );
xor \U$29229 ( \29475 , RIbe2adc0_109, RIbe29c68_72);
not \U$29230 ( \29476 , \29475 );
not \U$29231 ( \29477 , \7513 );
or \U$29232 ( \29478 , \29476 , \29477 );
xor \U$29233 ( \29479 , RIbe2a460_89, RIbe29c68_72);
nand \U$29234 ( \29480 , \4580 , \29479 );
nand \U$29235 ( \29481 , \29478 , \29480 );
nand \U$29236 ( \29482 , \29474 , \29481 );
nand \U$29237 ( \29483 , \29473 , \29482 );
not \U$29238 ( \29484 , \29483 );
and \U$29239 ( \29485 , \29456 , \29484 );
and \U$29240 ( \29486 , \29455 , \29483 );
nor \U$29241 ( \29487 , \29485 , \29486 );
not \U$29242 ( \29488 , \29487 );
not \U$29243 ( \29489 , \29488 );
or \U$29244 ( \29490 , \29429 , \29489 );
nand \U$29245 ( \29491 , \29454 , \29483 );
nand \U$29246 ( \29492 , \29490 , \29491 );
not \U$29247 ( \29493 , RIbe2a3e8_88);
not \U$29248 ( \29494 , RIbe2aa00_101);
and \U$29249 ( \29495 , \29493 , \29494 );
and \U$29250 ( \29496 , RIbe2a3e8_88, RIbe2aa00_101);
nor \U$29251 ( \29497 , \29495 , \29496 );
not \U$29252 ( \29498 , \29497 );
not \U$29253 ( \29499 , \17060 );
or \U$29254 ( \29500 , \29498 , \29499 );
xor \U$29255 ( \29501 , RIbe2aa78_102, RIbe2a3e8_88);
nand \U$29256 ( \29502 , \9268 , \29501 );
nand \U$29257 ( \29503 , \29500 , \29502 );
not \U$29258 ( \29504 , \29503 );
not \U$29259 ( \29505 , \29461 );
not \U$29260 ( \29506 , \20396 );
or \U$29261 ( \29507 , \29505 , \29506 );
nand \U$29262 ( \29508 , \20583 , \25131 );
nand \U$29263 ( \29509 , \29507 , \29508 );
not \U$29264 ( \29510 , \29509 );
and \U$29265 ( \29511 , \29504 , \29510 );
xor \U$29266 ( \29512 , RIbe2b3d8_122, RIbe28390_19);
not \U$29267 ( \29513 , \29512 );
not \U$29268 ( \29514 , \3408 );
or \U$29269 ( \29515 , \29513 , \29514 );
nand \U$29270 ( \29516 , \8654 , \25228 );
nand \U$29271 ( \29517 , \29515 , \29516 );
not \U$29272 ( \29518 , \29517 );
or \U$29273 ( \29519 , RIbe28390_19, RIbe28b10_35);
nand \U$29274 ( \29520 , \29519 , RIbe2ae38_110);
nand \U$29275 ( \29521 , RIbe28390_19, RIbe28b10_35);
and \U$29276 ( \29522 , \29520 , \29521 , RIbe28b88_36);
not \U$29277 ( \29523 , \29522 );
not \U$29278 ( \29524 , \29523 );
and \U$29279 ( \29525 , \29518 , \29524 );
and \U$29280 ( \29526 , \29517 , \29523 );
nor \U$29281 ( \29527 , \29525 , \29526 );
nor \U$29282 ( \29528 , \29511 , \29527 );
and \U$29283 ( \29529 , \29503 , \29509 );
nor \U$29284 ( \29530 , \29528 , \29529 );
xor \U$29285 ( \29531 , RIbe27fd0_11, RIbe2a6b8_94);
not \U$29286 ( \29532 , \29531 );
not \U$29287 ( \29533 , \11366 );
or \U$29288 ( \29534 , \29532 , \29533 );
xor \U$29289 ( \29535 , RIbe27fd0_11, RIbe2b4c8_124);
nand \U$29290 ( \29536 , \2707 , \29535 );
nand \U$29291 ( \29537 , \29534 , \29536 );
xor \U$29292 ( \29538 , RIbe285e8_24, RIbe2a7a8_96);
not \U$29293 ( \29539 , \29538 );
not \U$29294 ( \29540 , \2761 );
or \U$29295 ( \29541 , \29539 , \29540 );
xor \U$29296 ( \29542 , RIbe285e8_24, RIbe2abe0_105);
nand \U$29297 ( \29543 , \2625 , \29542 );
nand \U$29298 ( \29544 , \29541 , \29543 );
or \U$29299 ( \29545 , \29537 , \29544 );
xor \U$29300 ( \29546 , RIbe29998_66, RIbe2b180_117);
not \U$29301 ( \29547 , \29546 );
not \U$29302 ( \29548 , \14852 );
or \U$29303 ( \29549 , \29547 , \29548 );
nand \U$29304 ( \29550 , \14966 , \29314 );
nand \U$29305 ( \29551 , \29549 , \29550 );
nand \U$29306 ( \29552 , \29545 , \29551 );
nand \U$29307 ( \29553 , \29537 , \29544 );
nand \U$29308 ( \29554 , \29552 , \29553 );
xor \U$29309 ( \29555 , RIbe2ac58_106, RIbe27e68_8);
not \U$29310 ( \29556 , \29555 );
not \U$29311 ( \29557 , \2599 );
or \U$29312 ( \29558 , \29556 , \29557 );
nand \U$29313 ( \29559 , \2603 , \29307 );
nand \U$29314 ( \29560 , \29558 , \29559 );
not \U$29315 ( \29561 , RIbe29b00_69);
not \U$29316 ( \29562 , RIbe2aaf0_103);
and \U$29317 ( \29563 , \29561 , \29562 );
and \U$29318 ( \29564 , RIbe29b00_69, RIbe2aaf0_103);
nor \U$29319 ( \29565 , \29563 , \29564 );
not \U$29320 ( \29566 , \29565 );
not \U$29321 ( \29567 , \20574 );
or \U$29322 ( \29568 , \29566 , \29567 );
nand \U$29323 ( \29569 , \29320 , RIbe2ab68_104);
nand \U$29324 ( \29570 , \29568 , \29569 );
or \U$29325 ( \29571 , \29560 , \29570 );
xor \U$29326 ( \29572 , RIbe2a2f8_86, RIbe2a118_82);
not \U$29327 ( \29573 , \29572 );
not \U$29328 ( \29574 , \10792 );
or \U$29329 ( \29575 , \29573 , \29574 );
xor \U$29330 ( \29576 , RIbe2a2f8_86, RIbe2a820_97);
nand \U$29331 ( \29577 , \11094 , \29576 );
nand \U$29332 ( \29578 , \29575 , \29577 );
nand \U$29333 ( \29579 , \29571 , \29578 );
nand \U$29334 ( \29580 , \29560 , \29570 );
nand \U$29335 ( \29581 , \29579 , \29580 );
xor \U$29336 ( \29582 , \29554 , \29581 );
not \U$29337 ( \29583 , RIbe2a3e8_88);
not \U$29338 ( \29584 , RIbe2a898_98);
and \U$29339 ( \29585 , \29583 , \29584 );
and \U$29340 ( \29586 , RIbe2a3e8_88, RIbe2a898_98);
nor \U$29341 ( \29587 , \29585 , \29586 );
not \U$29342 ( \29588 , \29587 );
not \U$29343 ( \29589 , \9263 );
or \U$29344 ( \29590 , \29588 , \29589 );
nand \U$29345 ( \29591 , \9268 , \29497 );
nand \U$29346 ( \29592 , \29590 , \29591 );
not \U$29347 ( \29593 , \29592 );
xor \U$29348 ( \29594 , RIbe28cf0_39, RIbe2b108_116);
not \U$29349 ( \29595 , \29594 );
not \U$29350 ( \29596 , \21852 );
or \U$29351 ( \29597 , \29595 , \29596 );
nand \U$29352 ( \29598 , \13534 , \29347 );
nand \U$29353 ( \29599 , \29597 , \29598 );
not \U$29354 ( \29600 , \29599 );
or \U$29355 ( \29601 , \29593 , \29600 );
or \U$29356 ( \29602 , \29599 , \29592 );
xor \U$29357 ( \29603 , RIbe28390_19, RIbe2aeb0_111);
not \U$29358 ( \29604 , \29603 );
not \U$29359 ( \29605 , \3408 );
or \U$29360 ( \29606 , \29604 , \29605 );
nand \U$29361 ( \29607 , \2777 , \29512 );
nand \U$29362 ( \29608 , \29606 , \29607 );
nand \U$29363 ( \29609 , \29602 , \29608 );
nand \U$29364 ( \29610 , \29601 , \29609 );
and \U$29365 ( \29611 , \29582 , \29610 );
and \U$29366 ( \29612 , \29554 , \29581 );
or \U$29367 ( \29613 , \29611 , \29612 );
xnor \U$29368 ( \29614 , \29530 , \29613 );
xor \U$29369 ( \29615 , \29492 , \29614 );
not \U$29370 ( \29616 , \29615 );
xnor \U$29371 ( \29617 , \29371 , \29390 );
and \U$29372 ( \29618 , \11461 , \29415 );
and \U$29373 ( \29619 , \3249 , \25110 );
nor \U$29374 ( \29620 , \29618 , \29619 );
not \U$29375 ( \29621 , \29620 );
not \U$29376 ( \29622 , \29535 );
not \U$29377 ( \29623 , \3377 );
or \U$29378 ( \29624 , \29622 , \29623 );
nand \U$29379 ( \29625 , \2707 , \25102 );
nand \U$29380 ( \29626 , \29624 , \29625 );
not \U$29381 ( \29627 , \29434 );
not \U$29382 ( \29628 , \11452 );
not \U$29383 ( \29629 , \29628 );
or \U$29384 ( \29630 , \29627 , \29629 );
nand \U$29385 ( \29631 , \9726 , \25271 );
nand \U$29386 ( \29632 , \29630 , \29631 );
xor \U$29387 ( \29633 , \29626 , \29632 );
not \U$29388 ( \29634 , \29633 );
or \U$29389 ( \29635 , \29621 , \29634 );
or \U$29390 ( \29636 , \29633 , \29620 );
nand \U$29391 ( \29637 , \29635 , \29636 );
not \U$29392 ( \29638 , \29637 );
not \U$29393 ( \29639 , \29527 );
xor \U$29394 ( \29640 , \29503 , \29509 );
not \U$29395 ( \29641 , \29640 );
and \U$29396 ( \29642 , \29639 , \29641 );
and \U$29397 ( \29643 , \29527 , \29640 );
nor \U$29398 ( \29644 , \29642 , \29643 );
not \U$29399 ( \29645 , \29644 );
or \U$29400 ( \29646 , \29638 , \29645 );
or \U$29401 ( \29647 , \29644 , \29637 );
nand \U$29402 ( \29648 , \29646 , \29647 );
not \U$29403 ( \29649 , \29648 );
and \U$29404 ( \29650 , RIbe27df0_7, RIbe2b018_114);
nor \U$29405 ( \29651 , RIbe27df0_7, RIbe2b018_114);
nor \U$29406 ( \29652 , \29650 , \29651 );
not \U$29407 ( \29653 , \29652 );
not \U$29408 ( \29654 , \15967 );
or \U$29409 ( \29655 , \29653 , \29654 );
nand \U$29410 ( \29656 , \19371 , \29457 );
nand \U$29411 ( \29657 , \29655 , \29656 );
xor \U$29412 ( \29658 , RIbe28f48_44, RIbe2b4c8_124);
not \U$29413 ( \29659 , \29658 );
not \U$29414 ( \29660 , \9618 );
or \U$29415 ( \29661 , \29659 , \29660 );
nand \U$29416 ( \29662 , \11201 , \29411 );
nand \U$29417 ( \29663 , \29661 , \29662 );
xor \U$29418 ( \29664 , \29657 , \29663 );
xnor \U$29419 ( \29665 , RIbe2ad48_108, RIbe29c68_72);
not \U$29420 ( \29666 , \29665 );
not \U$29421 ( \29667 , \29666 );
not \U$29422 ( \29668 , \8595 );
or \U$29423 ( \29669 , \29667 , \29668 );
nand \U$29424 ( \29670 , \4580 , \29475 );
nand \U$29425 ( \29671 , \29669 , \29670 );
and \U$29426 ( \29672 , \29664 , \29671 );
and \U$29427 ( \29673 , \29657 , \29663 );
or \U$29428 ( \29674 , \29672 , \29673 );
not \U$29429 ( \29675 , \29674 );
nand \U$29430 ( \29676 , RIbe28408_20, RIbe28480_21);
and \U$29431 ( \29677 , \29676 , RIbe28390_19);
or \U$29432 ( \29678 , RIbe28408_20, RIbe28480_21);
nand \U$29433 ( \29679 , \29678 , RIbe2ae38_110);
nand \U$29434 ( \29680 , \29677 , \29679 );
not \U$29435 ( \29681 , \29680 );
xor \U$29436 ( \29682 , RIbe28480_21, RIbe2b3d8_122);
not \U$29437 ( \29683 , \29682 );
not \U$29438 ( \29684 , \2518 );
or \U$29439 ( \29685 , \29683 , \29684 );
xor \U$29440 ( \29686 , RIbe28480_21, RIbe2b450_123);
nand \U$29441 ( \29687 , \3074 , \29686 );
nand \U$29442 ( \29688 , \29685 , \29687 );
nand \U$29443 ( \29689 , \29681 , \29688 );
not \U$29444 ( \29690 , \29689 );
not \U$29445 ( \29691 , RIbe27fd0_11);
not \U$29446 ( \29692 , RIbe2a640_93);
and \U$29447 ( \29693 , \29691 , \29692 );
and \U$29448 ( \29694 , RIbe27fd0_11, RIbe2a640_93);
nor \U$29449 ( \29695 , \29693 , \29694 );
not \U$29450 ( \29696 , \29695 );
not \U$29451 ( \29697 , \9082 );
or \U$29452 ( \29698 , \29696 , \29697 );
nand \U$29453 ( \29699 , \2707 , \29531 );
nand \U$29454 ( \29700 , \29698 , \29699 );
not \U$29455 ( \29701 , \29700 );
not \U$29456 ( \29702 , \29701 );
xor \U$29457 ( \29703 , RIbe29ce0_73, RIbe2a280_85);
not \U$29458 ( \29704 , \29703 );
not \U$29459 ( \29705 , \23353 );
or \U$29460 ( \29706 , \29704 , \29705 );
nand \U$29461 ( \29707 , \10849 , \29437 );
nand \U$29462 ( \29708 , \29706 , \29707 );
not \U$29463 ( \29709 , \29708 );
not \U$29464 ( \29710 , \29709 );
or \U$29465 ( \29711 , \29702 , \29710 );
xor \U$29466 ( \29712 , RIbe2a460_89, RIbe29e48_76);
not \U$29467 ( \29713 , \29712 );
not \U$29468 ( \29714 , \16652 );
or \U$29469 ( \29715 , \29713 , \29714 );
nand \U$29470 ( \29716 , \16655 , \29445 );
nand \U$29471 ( \29717 , \29715 , \29716 );
nand \U$29472 ( \29718 , \29711 , \29717 );
nand \U$29473 ( \29719 , \29708 , \29700 );
nand \U$29474 ( \29720 , \29718 , \29719 );
not \U$29475 ( \29721 , \29720 );
or \U$29476 ( \29722 , \29690 , \29721 );
or \U$29477 ( \29723 , \29720 , \29689 );
nand \U$29478 ( \29724 , \29722 , \29723 );
not \U$29479 ( \29725 , \29724 );
or \U$29480 ( \29726 , \29675 , \29725 );
not \U$29481 ( \29727 , \29689 );
nand \U$29482 ( \29728 , \29727 , \29720 );
nand \U$29483 ( \29729 , \29726 , \29728 );
not \U$29484 ( \29730 , \29729 );
or \U$29485 ( \29731 , \29649 , \29730 );
not \U$29486 ( \29732 , \29644 );
nand \U$29487 ( \29733 , \29732 , \29637 );
nand \U$29488 ( \29734 , \29731 , \29733 );
xnor \U$29489 ( \29735 , \29617 , \29734 );
not \U$29490 ( \29736 , \29735 );
or \U$29491 ( \29737 , \29616 , \29736 );
not \U$29492 ( \29738 , \29617 );
nand \U$29493 ( \29739 , \29738 , \29734 );
nand \U$29494 ( \29740 , \29737 , \29739 );
not \U$29495 ( \29741 , \29740 );
and \U$29496 ( \29742 , \29396 , \29741 );
and \U$29497 ( \29743 , \29740 , \29395 );
nor \U$29498 ( \29744 , \29742 , \29743 );
not \U$29499 ( \29745 , \25100 );
not \U$29500 ( \29746 , \29745 );
not \U$29501 ( \29747 , \25119 );
or \U$29502 ( \29748 , \29746 , \29747 );
or \U$29503 ( \29749 , \25119 , \29745 );
nand \U$29504 ( \29750 , \29748 , \29749 );
not \U$29505 ( \29751 , \29750 );
xor \U$29506 ( \29752 , \25013 , \25027 );
not \U$29507 ( \29753 , \29752 );
not \U$29508 ( \29754 , \29753 );
or \U$29509 ( \29755 , \29751 , \29754 );
or \U$29510 ( \29756 , \29753 , \29750 );
nand \U$29511 ( \29757 , \29755 , \29756 );
not \U$29512 ( \29758 , \29757 );
xnor \U$29513 ( \29759 , \25063 , \25081 );
not \U$29514 ( \29760 , \29759 );
not \U$29515 ( \29761 , \29760 );
or \U$29516 ( \29762 , \29758 , \29761 );
nand \U$29517 ( \29763 , \29752 , \29750 );
nand \U$29518 ( \29764 , \29762 , \29763 );
not \U$29519 ( \29765 , \29764 );
not \U$29520 ( \29766 , \29407 );
not \U$29521 ( \29767 , \16914 );
or \U$29522 ( \29768 , \29766 , \29767 );
nand \U$29523 ( \29769 , \17811 , \25095 );
nand \U$29524 ( \29770 , \29768 , \29769 );
not \U$29525 ( \29771 , \29770 );
not \U$29526 ( \29772 , \29449 );
not \U$29527 ( \29773 , \19978 );
or \U$29528 ( \29774 , \29772 , \29773 );
nand \U$29529 ( \29775 , \4849 , \25144 );
nand \U$29530 ( \29776 , \29774 , \29775 );
not \U$29531 ( \29777 , \29441 );
not \U$29532 ( \29778 , \14382 );
or \U$29533 ( \29779 , \29777 , \29778 );
nand \U$29534 ( \29780 , \14649 , \25138 );
nand \U$29535 ( \29781 , \29779 , \29780 );
xor \U$29536 ( \29782 , \29776 , \29781 );
not \U$29537 ( \29783 , \29782 );
or \U$29538 ( \29784 , \29771 , \29783 );
nand \U$29539 ( \29785 , \29781 , \29776 );
nand \U$29540 ( \29786 , \29784 , \29785 );
not \U$29541 ( \29787 , \29786 );
nor \U$29542 ( \29788 , \29632 , \29626 );
or \U$29543 ( \29789 , \29788 , \29620 );
nand \U$29544 ( \29790 , \29632 , \29626 );
nand \U$29545 ( \29791 , \29789 , \29790 );
not \U$29546 ( \29792 , \29791 );
not \U$29547 ( \29793 , \29469 );
not \U$29548 ( \29794 , \8401 );
or \U$29549 ( \29795 , \29793 , \29794 );
nand \U$29550 ( \29796 , \8172 , \25021 );
nand \U$29551 ( \29797 , \29795 , \29796 );
not \U$29552 ( \29798 , \29797 );
xor \U$29553 ( \29799 , RIbe28480_21, RIbe2a730_95);
not \U$29554 ( \29800 , \29799 );
not \U$29555 ( \29801 , \16953 );
or \U$29556 ( \29802 , \29800 , \29801 );
nand \U$29557 ( \29803 , \16676 , \25015 );
nand \U$29558 ( \29804 , \29802 , \29803 );
not \U$29559 ( \29805 , \29804 );
not \U$29560 ( \29806 , \29542 );
not \U$29561 ( \29807 , \10863 );
or \U$29562 ( \29808 , \29806 , \29807 );
nand \U$29563 ( \29809 , \8270 , \25065 );
nand \U$29564 ( \29810 , \29808 , \29809 );
not \U$29565 ( \29811 , \29810 );
not \U$29566 ( \29812 , \29811 );
or \U$29567 ( \29813 , \29805 , \29812 );
or \U$29568 ( \29814 , \29804 , \29811 );
nand \U$29569 ( \29815 , \29813 , \29814 );
not \U$29570 ( \29816 , \29815 );
or \U$29571 ( \29817 , \29798 , \29816 );
not \U$29572 ( \29818 , \29811 );
nand \U$29573 ( \29819 , \29818 , \29804 );
nand \U$29574 ( \29820 , \29817 , \29819 );
not \U$29575 ( \29821 , \29820 );
not \U$29576 ( \29822 , \29821 );
or \U$29577 ( \29823 , \29792 , \29822 );
or \U$29578 ( \29824 , \29821 , \29791 );
nand \U$29579 ( \29825 , \29823 , \29824 );
not \U$29580 ( \29826 , \29825 );
or \U$29581 ( \29827 , \29787 , \29826 );
not \U$29582 ( \29828 , \29821 );
nand \U$29583 ( \29829 , \29828 , \29791 );
nand \U$29584 ( \29830 , \29827 , \29829 );
not \U$29585 ( \29831 , \29830 );
not \U$29586 ( \29832 , \29501 );
not \U$29587 ( \29833 , \8806 );
or \U$29588 ( \29834 , \29832 , \29833 );
nand \U$29589 ( \29835 , \8794 , \24235 );
nand \U$29590 ( \29836 , \29834 , \29835 );
and \U$29591 ( \29837 , \29517 , \29522 );
xor \U$29592 ( \29838 , \29836 , \29837 );
buf \U$29593 ( \29839 , \29838 );
not \U$29594 ( \29840 , \29576 );
not \U$29595 ( \29841 , \16714 );
or \U$29596 ( \29842 , \29840 , \29841 );
nand \U$29597 ( \29843 , \8705 , \25008 );
nand \U$29598 ( \29844 , \29842 , \29843 );
not \U$29599 ( \29845 , \29844 );
not \U$29600 ( \29846 , \29845 );
xor \U$29601 ( \29847 , RIbe29ce0_73, RIbe2a190_83);
not \U$29602 ( \29848 , \29847 );
not \U$29603 ( \29849 , \15764 );
or \U$29604 ( \29850 , \29848 , \29849 );
nand \U$29605 ( \29851 , \22918 , \25034 );
nand \U$29606 ( \29852 , \29850 , \29851 );
not \U$29607 ( \29853 , \29852 );
not \U$29608 ( \29854 , \29853 );
or \U$29609 ( \29855 , \29846 , \29854 );
not \U$29610 ( \29856 , \29479 );
not \U$29611 ( \29857 , \4578 );
or \U$29612 ( \29858 , \29856 , \29857 );
nand \U$29613 ( \29859 , \7237 , \25049 );
nand \U$29614 ( \29860 , \29858 , \29859 );
nand \U$29615 ( \29861 , \29855 , \29860 );
nand \U$29616 ( \29862 , \29844 , \29852 );
and \U$29617 ( \29863 , \29861 , \29862 );
not \U$29618 ( \29864 , \29863 );
and \U$29619 ( \29865 , \29839 , \29864 );
and \U$29620 ( \29866 , \29836 , \29837 );
nor \U$29621 ( \29867 , \29865 , \29866 );
not \U$29622 ( \29868 , \29867 );
and \U$29623 ( \29869 , \29831 , \29868 );
and \U$29624 ( \29870 , \29830 , \29867 );
nor \U$29625 ( \29871 , \29869 , \29870 );
not \U$29626 ( \29872 , \29871 );
or \U$29627 ( \29873 , \29765 , \29872 );
or \U$29628 ( \29874 , \29764 , \29871 );
nand \U$29629 ( \29875 , \29873 , \29874 );
xor \U$29630 ( \29876 , \25290 , \25297 );
xor \U$29631 ( \29877 , \29876 , \25302 );
not \U$29632 ( \29878 , \29877 );
not \U$29633 ( \29879 , \29492 );
not \U$29634 ( \29880 , \29614 );
or \U$29635 ( \29881 , \29879 , \29880 );
not \U$29636 ( \29882 , \29530 );
nand \U$29637 ( \29883 , \29882 , \29613 );
nand \U$29638 ( \29884 , \29881 , \29883 );
not \U$29639 ( \29885 , \29884 );
not \U$29640 ( \29886 , \29885 );
or \U$29641 ( \29887 , \29878 , \29886 );
not \U$29642 ( \29888 , \29877 );
nand \U$29643 ( \29889 , \29884 , \29888 );
nand \U$29644 ( \29890 , \29887 , \29889 );
not \U$29645 ( \29891 , \29890 );
and \U$29646 ( \29892 , \29875 , \29891 );
not \U$29647 ( \29893 , \29875 );
and \U$29648 ( \29894 , \29893 , \29890 );
nor \U$29649 ( \29895 , \29892 , \29894 );
not \U$29650 ( \29896 , \29895 );
and \U$29651 ( \29897 , \29744 , \29896 );
not \U$29652 ( \29898 , \29744 );
and \U$29653 ( \29899 , \29898 , \29895 );
nor \U$29654 ( \29900 , \29897 , \29899 );
xor \U$29655 ( \29901 , \29729 , \29648 );
not \U$29656 ( \29902 , \29901 );
not \U$29657 ( \29903 , \29409 );
and \U$29658 ( \29904 , \29424 , \29903 );
not \U$29659 ( \29905 , \29424 );
and \U$29660 ( \29906 , \29905 , \29409 );
nor \U$29661 ( \29907 , \29904 , \29906 );
xor \U$29662 ( \29908 , \29481 , \29463 );
not \U$29663 ( \29909 , \29471 );
xor \U$29664 ( \29910 , \29908 , \29909 );
nand \U$29665 ( \29911 , \29907 , \29910 );
not \U$29666 ( \29912 , \29911 );
xor \U$29667 ( \29913 , RIbe27c88_4, RIbe2b018_114);
not \U$29668 ( \29914 , \29913 );
not \U$29669 ( \29915 , \22763 );
or \U$29670 ( \29916 , \29914 , \29915 );
nand \U$29671 ( \29917 , \15953 , \29652 );
nand \U$29672 ( \29918 , \29916 , \29917 );
not \U$29673 ( \29919 , \29918 );
not \U$29674 ( \29920 , \4581 );
not \U$29675 ( \29921 , \29665 );
and \U$29676 ( \29922 , \29920 , \29921 );
xor \U$29677 ( \29923 , RIbe29c68_72, RIbe2b540_125);
and \U$29678 ( \29924 , \8259 , \29923 );
nor \U$29679 ( \29925 , \29922 , \29924 );
nand \U$29680 ( \29926 , \29919 , \29925 );
not \U$29681 ( \29927 , \29926 );
xor \U$29682 ( \29928 , RIbe2adc0_109, RIbe29e48_76);
not \U$29683 ( \29929 , \29928 );
not \U$29684 ( \29930 , \7716 );
or \U$29685 ( \29931 , \29929 , \29930 );
nand \U$29686 ( \29932 , \4850 , \29712 );
nand \U$29687 ( \29933 , \29931 , \29932 );
not \U$29688 ( \29934 , \29933 );
or \U$29689 ( \29935 , \29927 , \29934 );
not \U$29690 ( \29936 , \29925 );
nand \U$29691 ( \29937 , \29936 , \29918 );
nand \U$29692 ( \29938 , \29935 , \29937 );
not \U$29693 ( \29939 , \29938 );
xor \U$29694 ( \29940 , RIbe28390_19, RIbe2ae38_110);
not \U$29695 ( \29941 , \29940 );
not \U$29696 ( \29942 , \2639 );
or \U$29697 ( \29943 , \29941 , \29942 );
nand \U$29698 ( \29944 , \5831 , \29603 );
nand \U$29699 ( \29945 , \29943 , \29944 );
not \U$29700 ( \29946 , \29945 );
not \U$29701 ( \29947 , \29688 );
not \U$29702 ( \29948 , \29680 );
and \U$29703 ( \29949 , \29947 , \29948 );
and \U$29704 ( \29950 , \29688 , \29680 );
nor \U$29705 ( \29951 , \29949 , \29950 );
not \U$29706 ( \29952 , \29951 );
or \U$29707 ( \29953 , \29946 , \29952 );
or \U$29708 ( \29954 , \29951 , \29945 );
nand \U$29709 ( \29955 , \29953 , \29954 );
not \U$29710 ( \29956 , \29955 );
or \U$29711 ( \29957 , \29939 , \29956 );
not \U$29712 ( \29958 , \29951 );
nand \U$29713 ( \29959 , \29958 , \29945 );
nand \U$29714 ( \29960 , \29957 , \29959 );
not \U$29715 ( \29961 , \29960 );
or \U$29716 ( \29962 , \29912 , \29961 );
or \U$29717 ( \29963 , \29907 , \29910 );
nand \U$29718 ( \29964 , \29962 , \29963 );
not \U$29719 ( \29965 , \29964 );
not \U$29720 ( \29966 , \29844 );
not \U$29721 ( \29967 , \29853 );
or \U$29722 ( \29968 , \29966 , \29967 );
nand \U$29723 ( \29969 , \29845 , \29852 );
nand \U$29724 ( \29970 , \29968 , \29969 );
xnor \U$29725 ( \29971 , \29970 , \29860 );
not \U$29726 ( \29972 , \29971 );
not \U$29727 ( \29973 , \29972 );
not \U$29728 ( \29974 , \29686 );
not \U$29729 ( \29975 , \3483 );
or \U$29730 ( \29976 , \29974 , \29975 );
nand \U$29731 ( \29977 , \3074 , \29799 );
nand \U$29732 ( \29978 , \29976 , \29977 );
not \U$29733 ( \29979 , \29978 );
and \U$29734 ( \29980 , \13250 , RIbe2ae38_110);
xor \U$29735 ( \29981 , RIbe29d58_74, RIbe2a190_83);
not \U$29736 ( \29982 , \29981 );
not \U$29737 ( \29983 , \11396 );
or \U$29738 ( \29984 , \29982 , \29983 );
nand \U$29739 ( \29985 , \10695 , \29847 );
nand \U$29740 ( \29986 , \29984 , \29985 );
xor \U$29741 ( \29987 , \29980 , \29986 );
not \U$29742 ( \29988 , \29987 );
or \U$29743 ( \29989 , \29979 , \29988 );
nand \U$29744 ( \29990 , \29986 , \29980 );
nand \U$29745 ( \29991 , \29989 , \29990 );
not \U$29746 ( \29992 , \29991 );
not \U$29747 ( \29993 , \29992 );
or \U$29748 ( \29994 , \29973 , \29993 );
nand \U$29749 ( \29995 , \29971 , \29991 );
nand \U$29750 ( \29996 , \29994 , \29995 );
not \U$29751 ( \29997 , \29312 );
not \U$29752 ( \29998 , \29997 );
not \U$29753 ( \29999 , \29326 );
or \U$29754 ( \30000 , \29998 , \29999 );
or \U$29755 ( \30001 , \29326 , \29997 );
nand \U$29756 ( \30002 , \30000 , \30001 );
not \U$29757 ( \30003 , \30002 );
and \U$29758 ( \30004 , \29996 , \30003 );
not \U$29759 ( \30005 , \29996 );
and \U$29760 ( \30006 , \30005 , \30002 );
nor \U$29761 ( \30007 , \30004 , \30006 );
not \U$29762 ( \30008 , \30007 );
or \U$29763 ( \30009 , \29965 , \30008 );
or \U$29764 ( \30010 , \29964 , \30007 );
nand \U$29765 ( \30011 , \30009 , \30010 );
not \U$29766 ( \30012 , \30011 );
or \U$29767 ( \30013 , \29902 , \30012 );
not \U$29768 ( \30014 , \30007 );
nand \U$29769 ( \30015 , \30014 , \29964 );
nand \U$29770 ( \30016 , \30013 , \30015 );
xor \U$29771 ( \30017 , \29770 , \29782 );
not \U$29772 ( \30018 , \30017 );
xor \U$29773 ( \30019 , \29336 , \29343 );
not \U$29774 ( \30020 , \29352 );
and \U$29775 ( \30021 , \30019 , \30020 );
not \U$29776 ( \30022 , \30019 );
and \U$29777 ( \30023 , \30022 , \29352 );
nor \U$29778 ( \30024 , \30021 , \30023 );
xnor \U$29779 ( \30025 , \29815 , \29797 );
nand \U$29780 ( \30026 , \30024 , \30025 );
not \U$29781 ( \30027 , \30026 );
or \U$29782 ( \30028 , \30018 , \30027 );
not \U$29783 ( \30029 , \30024 );
not \U$29784 ( \30030 , \30025 );
nand \U$29785 ( \30031 , \30029 , \30030 );
nand \U$29786 ( \30032 , \30028 , \30031 );
xor \U$29787 ( \30033 , \29825 , \29786 );
xor \U$29788 ( \30034 , \30032 , \30033 );
not \U$29789 ( \30035 , \29759 );
not \U$29790 ( \30036 , \29757 );
or \U$29791 ( \30037 , \30035 , \30036 );
or \U$29792 ( \30038 , \29757 , \29759 );
nand \U$29793 ( \30039 , \30037 , \30038 );
xor \U$29794 ( \30040 , \30034 , \30039 );
xor \U$29795 ( \30041 , \30016 , \30040 );
xnor \U$29796 ( \30042 , \29735 , \29615 );
and \U$29797 ( \30043 , \30041 , \30042 );
not \U$29798 ( \30044 , \30041 );
not \U$29799 ( \30045 , \30042 );
and \U$29800 ( \30046 , \30044 , \30045 );
or \U$29801 ( \30047 , \30043 , \30046 );
not \U$29802 ( \30048 , \30047 );
xor \U$29803 ( \30049 , \29554 , \29581 );
xor \U$29804 ( \30050 , \30049 , \29610 );
not \U$29805 ( \30051 , \30050 );
not \U$29806 ( \30052 , \29487 );
not \U$29807 ( \30053 , \29428 );
and \U$29808 ( \30054 , \30052 , \30053 );
and \U$29809 ( \30055 , \29487 , \29428 );
nor \U$29810 ( \30056 , \30054 , \30055 );
not \U$29811 ( \30057 , \30056 );
or \U$29812 ( \30058 , \30051 , \30057 );
or \U$29813 ( \30059 , \30056 , \30050 );
nand \U$29814 ( \30060 , \30058 , \30059 );
buf \U$29815 ( \30061 , \30026 );
nand \U$29816 ( \30062 , \30061 , \30031 );
not \U$29817 ( \30063 , \30017 );
and \U$29818 ( \30064 , \30062 , \30063 );
not \U$29819 ( \30065 , \30062 );
and \U$29820 ( \30066 , \30065 , \30017 );
nor \U$29821 ( \30067 , \30064 , \30066 );
xnor \U$29822 ( \30068 , \30060 , \30067 );
not \U$29823 ( \30069 , \30068 );
not \U$29824 ( \30070 , \30069 );
not \U$29825 ( \30071 , \19580 );
xor \U$29826 ( \30072 , RIbe29218_50, RIbe2aaf0_103);
not \U$29827 ( \30073 , \30072 );
not \U$29828 ( \30074 , \30073 );
and \U$29829 ( \30075 , \30071 , \30074 );
xor \U$29830 ( \30076 , RIbe29a10_67, RIbe2aaf0_103);
and \U$29831 ( \30077 , RIbe2ab68_104, \30076 );
nor \U$29832 ( \30078 , \30075 , \30077 );
not \U$29833 ( \30079 , \30078 );
not \U$29834 ( \30080 , \30079 );
xor \U$29835 ( \30081 , RIbe2a2f8_86, RIbe2b360_121);
not \U$29836 ( \30082 , \30081 );
not \U$29837 ( \30083 , \16714 );
or \U$29838 ( \30084 , \30082 , \30083 );
xor \U$29839 ( \30085 , RIbe2a0a0_81, RIbe2a2f8_86);
nand \U$29840 ( \30086 , \8705 , \30085 );
nand \U$29841 ( \30087 , \30084 , \30086 );
not \U$29842 ( \30088 , \30087 );
or \U$29843 ( \30089 , \30080 , \30088 );
not \U$29844 ( \30090 , \30087 );
not \U$29845 ( \30091 , \30090 );
not \U$29846 ( \30092 , \30078 );
or \U$29847 ( \30093 , \30091 , \30092 );
xor \U$29848 ( \30094 , RIbe2a910_99, RIbe2a898_98);
not \U$29849 ( \30095 , \30094 );
not \U$29850 ( \30096 , \9738 );
or \U$29851 ( \30097 , \30095 , \30096 );
xor \U$29852 ( \30098 , RIbe2a910_99, RIbe2aa00_101);
nand \U$29853 ( \30099 , \10400 , \30098 );
nand \U$29854 ( \30100 , \30097 , \30099 );
nand \U$29855 ( \30101 , \30093 , \30100 );
nand \U$29856 ( \30102 , \30089 , \30101 );
not \U$29857 ( \30103 , \30102 );
xor \U$29858 ( \30104 , RIbe285e8_24, RIbe2b450_123);
not \U$29859 ( \30105 , \30104 );
not \U$29860 ( \30106 , \11174 );
or \U$29861 ( \30107 , \30105 , \30106 );
xor \U$29862 ( \30108 , RIbe285e8_24, RIbe2a730_95);
nand \U$29863 ( \30109 , \2758 , \30108 );
nand \U$29864 ( \30110 , \30107 , \30109 );
not \U$29865 ( \30111 , \30110 );
xor \U$29866 ( \30112 , RIbe29d58_74, RIbe2a280_85);
not \U$29867 ( \30113 , \30112 );
not \U$29868 ( \30114 , \27992 );
or \U$29869 ( \30115 , \30113 , \30114 );
nand \U$29870 ( \30116 , \11348 , \29703 );
nand \U$29871 ( \30117 , \30115 , \30116 );
not \U$29872 ( \30118 , \30117 );
or \U$29873 ( \30119 , \30111 , \30118 );
or \U$29874 ( \30120 , \30117 , \30110 );
nand \U$29875 ( \30121 , \2648 , RIbe2ae38_110);
not \U$29876 ( \30122 , \30121 );
nand \U$29877 ( \30123 , \30120 , \30122 );
nand \U$29878 ( \30124 , \30119 , \30123 );
not \U$29879 ( \30125 , \30124 );
or \U$29880 ( \30126 , \30103 , \30125 );
or \U$29881 ( \30127 , \30124 , \30102 );
xor \U$29882 ( \30128 , RIbe28cf0_39, RIbe2b180_117);
not \U$29883 ( \30129 , \30128 );
not \U$29884 ( \30130 , \15353 );
or \U$29885 ( \30131 , \30129 , \30130 );
xor \U$29886 ( \30132 , RIbe298a8_64, RIbe2b180_117);
nand \U$29887 ( \30133 , \16646 , \30132 );
nand \U$29888 ( \30134 , \30131 , \30133 );
xnor \U$29889 ( \30135 , RIbe2a118_82, RIbe2a3e8_88);
or \U$29890 ( \30136 , \11544 , \30135 );
xor \U$29891 ( \30137 , RIbe2a3e8_88, RIbe2a820_97);
nand \U$29892 ( \30138 , \9268 , \30137 );
nand \U$29893 ( \30139 , \30136 , \30138 );
nor \U$29894 ( \30140 , \30134 , \30139 );
xor \U$29895 ( \30141 , RIbe2af28_112, RIbe29998_66);
not \U$29896 ( \30142 , \30141 );
not \U$29897 ( \30143 , \15345 );
or \U$29898 ( \30144 , \30142 , \30143 );
xor \U$29899 ( \30145 , RIbe28d68_40, RIbe2af28_112);
nand \U$29900 ( \30146 , \16917 , \30145 );
nand \U$29901 ( \30147 , \30144 , \30146 );
not \U$29902 ( \30148 , \30147 );
or \U$29903 ( \30149 , \30140 , \30148 );
nand \U$29904 ( \30150 , \30139 , \30134 );
nand \U$29905 ( \30151 , \30149 , \30150 );
nand \U$29906 ( \30152 , \30127 , \30151 );
nand \U$29907 ( \30153 , \30126 , \30152 );
not \U$29908 ( \30154 , \30085 );
not \U$29909 ( \30155 , \16715 );
or \U$29910 ( \30156 , \30154 , \30155 );
nand \U$29911 ( \30157 , \11094 , \29572 );
nand \U$29912 ( \30158 , \30156 , \30157 );
not \U$29913 ( \30159 , \30158 );
not \U$29914 ( \30160 , \30132 );
not \U$29915 ( \30161 , \15353 );
or \U$29916 ( \30162 , \30160 , \30161 );
nand \U$29917 ( \30163 , \16646 , \29546 );
nand \U$29918 ( \30164 , \30162 , \30163 );
not \U$29919 ( \30165 , \30164 );
not \U$29920 ( \30166 , \30108 );
not \U$29921 ( \30167 , \2761 );
or \U$29922 ( \30168 , \30166 , \30167 );
nand \U$29923 ( \30169 , \2758 , \29538 );
nand \U$29924 ( \30170 , \30168 , \30169 );
not \U$29925 ( \30171 , \30170 );
and \U$29926 ( \30172 , \30165 , \30171 );
not \U$29927 ( \30173 , \30165 );
and \U$29928 ( \30174 , \30173 , \30170 );
nor \U$29929 ( \30175 , \30172 , \30174 );
not \U$29930 ( \30176 , \30175 );
or \U$29931 ( \30177 , \30159 , \30176 );
not \U$29932 ( \30178 , \30165 );
nand \U$29933 ( \30179 , \30178 , \30170 );
nand \U$29934 ( \30180 , \30177 , \30179 );
not \U$29935 ( \30181 , \30180 );
not \U$29936 ( \30182 , \30181 );
not \U$29937 ( \30183 , \30137 );
not \U$29938 ( \30184 , \9262 );
or \U$29939 ( \30185 , \30183 , \30184 );
nand \U$29940 ( \30186 , \26573 , \29587 );
nand \U$29941 ( \30187 , \30185 , \30186 );
not \U$29942 ( \30188 , \30187 );
xor \U$29943 ( \30189 , RIbe2a028_80, RIbe2b2e8_120);
not \U$29944 ( \30190 , \30189 );
not \U$29945 ( \30191 , \8168 );
or \U$29946 ( \30192 , \30190 , \30191 );
nand \U$29947 ( \30193 , \8930 , \29465 );
nand \U$29948 ( \30194 , \30192 , \30193 );
not \U$29949 ( \30195 , \30194 );
or \U$29950 ( \30196 , \30188 , \30195 );
or \U$29951 ( \30197 , \30194 , \30187 );
xor \U$29952 ( \30198 , RIbe2b108_116, RIbe27b20_1);
not \U$29953 ( \30199 , \30198 );
not \U$29954 ( \30200 , \14296 );
or \U$29955 ( \30201 , \30199 , \30200 );
nand \U$29956 ( \30202 , \13533 , \29594 );
nand \U$29957 ( \30203 , \30201 , \30202 );
nand \U$29958 ( \30204 , \30197 , \30203 );
nand \U$29959 ( \30205 , \30196 , \30204 );
not \U$29960 ( \30206 , \30205 );
not \U$29961 ( \30207 , \30206 );
not \U$29962 ( \30208 , \30098 );
not \U$29963 ( \30209 , \10987 );
or \U$29964 ( \30210 , \30208 , \30209 );
nand \U$29965 ( \30211 , \11456 , \29430 );
nand \U$29966 ( \30212 , \30210 , \30211 );
not \U$29967 ( \30213 , \30145 );
not \U$29968 ( \30214 , \16913 );
or \U$29969 ( \30215 , \30213 , \30214 );
nand \U$29970 ( \30216 , \17810 , \29401 );
nand \U$29971 ( \30217 , \30215 , \30216 );
nor \U$29972 ( \30218 , \30212 , \30217 );
xor \U$29973 ( \30219 , RIbe2a550_91, RIbe2b6a8_128);
and \U$29974 ( \30220 , \19607 , \30219 );
and \U$29975 ( \30221 , \12004 , \29418 );
nor \U$29976 ( \30222 , \30220 , \30221 );
or \U$29977 ( \30223 , \30218 , \30222 );
nand \U$29978 ( \30224 , \30212 , \30217 );
nand \U$29979 ( \30225 , \30223 , \30224 );
not \U$29980 ( \30226 , \30225 );
or \U$29981 ( \30227 , \30207 , \30226 );
or \U$29982 ( \30228 , \30225 , \30206 );
nand \U$29983 ( \30229 , \30227 , \30228 );
not \U$29984 ( \30230 , \30229 );
or \U$29985 ( \30231 , \30182 , \30230 );
or \U$29986 ( \30232 , \30229 , \30181 );
nand \U$29987 ( \30233 , \30231 , \30232 );
xor \U$29988 ( \30234 , \30153 , \30233 );
not \U$29989 ( \30235 , \30076 );
buf \U$29990 ( \30236 , \28282 );
not \U$29991 ( \30237 , \30236 );
or \U$29992 ( \30238 , \30235 , \30237 );
nand \U$29993 ( \30239 , \29565 , RIbe2ab68_104);
nand \U$29994 ( \30240 , \30238 , \30239 );
xor \U$29995 ( \30241 , RIbe2abe0_105, RIbe27e68_8);
not \U$29996 ( \30242 , \30241 );
not \U$29997 ( \30243 , \2599 );
or \U$29998 ( \30244 , \30242 , \30243 );
nand \U$29999 ( \30245 , \2603 , \29555 );
nand \U$30000 ( \30246 , \30244 , \30245 );
xor \U$30001 ( \30247 , \30240 , \30246 );
not \U$30002 ( \30248 , RIbe29ec0_77);
not \U$30003 ( \30249 , RIbe2a190_83);
and \U$30004 ( \30250 , \30248 , \30249 );
and \U$30005 ( \30251 , RIbe29ec0_77, RIbe2a190_83);
nor \U$30006 ( \30252 , \30250 , \30251 );
not \U$30007 ( \30253 , \30252 );
not \U$30008 ( \30254 , \11396 );
or \U$30009 ( \30255 , \30253 , \30254 );
nand \U$30010 ( \30256 , \11400 , \29981 );
nand \U$30011 ( \30257 , \30255 , \30256 );
not \U$30012 ( \30258 , \30257 );
and \U$30013 ( \30259 , \30247 , \30258 );
not \U$30014 ( \30260 , \30247 );
and \U$30015 ( \30261 , \30260 , \30257 );
nor \U$30016 ( \30262 , \30259 , \30261 );
not \U$30017 ( \30263 , \30262 );
not \U$30018 ( \30264 , \30263 );
not \U$30019 ( \30265 , \29701 );
not \U$30020 ( \30266 , \29708 );
or \U$30021 ( \30267 , \30265 , \30266 );
nand \U$30022 ( \30268 , \29709 , \29700 );
nand \U$30023 ( \30269 , \30267 , \30268 );
xnor \U$30024 ( \30270 , \30269 , \29717 );
not \U$30025 ( \30271 , \30270 );
xor \U$30026 ( \30272 , \30187 , \30203 );
xor \U$30027 ( \30273 , \30272 , \30194 );
not \U$30028 ( \30274 , \30273 );
or \U$30029 ( \30275 , \30271 , \30274 );
or \U$30030 ( \30276 , \30273 , \30270 );
nand \U$30031 ( \30277 , \30275 , \30276 );
not \U$30032 ( \30278 , \30277 );
or \U$30033 ( \30279 , \30264 , \30278 );
not \U$30034 ( \30280 , \30270 );
nand \U$30035 ( \30281 , \30280 , \30273 );
nand \U$30036 ( \30282 , \30279 , \30281 );
and \U$30037 ( \30283 , \30234 , \30282 );
and \U$30038 ( \30284 , \30153 , \30233 );
or \U$30039 ( \30285 , \30283 , \30284 );
not \U$30040 ( \30286 , \30285 );
not \U$30041 ( \30287 , \30286 );
xor \U$30042 ( \30288 , \29674 , \29724 );
not \U$30043 ( \30289 , \30288 );
not \U$30044 ( \30290 , \30175 );
not \U$30045 ( \30291 , \30158 );
not \U$30046 ( \30292 , \30291 );
and \U$30047 ( \30293 , \30290 , \30292 );
and \U$30048 ( \30294 , \30175 , \30291 );
nor \U$30049 ( \30295 , \30293 , \30294 );
not \U$30050 ( \30296 , \30295 );
not \U$30051 ( \30297 , \30296 );
xor \U$30052 ( \30298 , RIbe2a550_91, RIbe2aa78_102);
not \U$30053 ( \30299 , \30298 );
not \U$30054 ( \30300 , \11999 );
or \U$30055 ( \30301 , \30299 , \30300 );
nand \U$30056 ( \30302 , \11484 , \30219 );
nand \U$30057 ( \30303 , \30301 , \30302 );
xor \U$30058 ( \30304 , RIbe28f48_44, RIbe2a6b8_94);
not \U$30059 ( \30305 , \30304 );
not \U$30060 ( \30306 , \23097 );
or \U$30061 ( \30307 , \30305 , \30306 );
nand \U$30062 ( \30308 , \9524 , \29658 );
nand \U$30063 ( \30309 , \30307 , \30308 );
nor \U$30064 ( \30310 , \30303 , \30309 );
not \U$30065 ( \30311 , \30310 );
xor \U$30066 ( \30312 , RIbe2a7a8_96, RIbe27e68_8);
not \U$30067 ( \30313 , \30312 );
not \U$30068 ( \30314 , \4443 );
or \U$30069 ( \30315 , \30313 , \30314 );
nand \U$30070 ( \30316 , \2603 , \30241 );
nand \U$30071 ( \30317 , \30315 , \30316 );
nand \U$30072 ( \30318 , \30311 , \30317 );
nand \U$30073 ( \30319 , \30303 , \30309 );
nand \U$30074 ( \30320 , \30318 , \30319 );
xor \U$30075 ( \30321 , RIbe2a028_80, RIbe2a4d8_90);
not \U$30076 ( \30322 , \30321 );
not \U$30077 ( \30323 , \8168 );
or \U$30078 ( \30324 , \30322 , \30323 );
nand \U$30079 ( \30325 , \8172 , \30189 );
nand \U$30080 ( \30326 , \30324 , \30325 );
not \U$30081 ( \30327 , \30326 );
xor \U$30082 ( \30328 , RIbe2b108_116, RIbe29b78_70);
not \U$30083 ( \30329 , \30328 );
not \U$30084 ( \30330 , \14296 );
or \U$30085 ( \30331 , \30329 , \30330 );
nand \U$30086 ( \30332 , \13533 , \30198 );
nand \U$30087 ( \30333 , \30331 , \30332 );
not \U$30088 ( \30334 , \30333 );
not \U$30089 ( \30335 , \30334 );
or \U$30090 ( \30336 , \30327 , \30335 );
or \U$30091 ( \30337 , \30334 , \30326 );
nand \U$30092 ( \30338 , \30336 , \30337 );
not \U$30093 ( \30339 , \30338 );
not \U$30094 ( \30340 , RIbe29f38_78);
not \U$30095 ( \30341 , RIbe2a190_83);
and \U$30096 ( \30342 , \30340 , \30341 );
and \U$30097 ( \30343 , RIbe29f38_78, RIbe2a190_83);
nor \U$30098 ( \30344 , \30342 , \30343 );
not \U$30099 ( \30345 , \30344 );
not \U$30100 ( \30346 , \10690 );
or \U$30101 ( \30347 , \30345 , \30346 );
nand \U$30102 ( \30348 , \11400 , \30252 );
nand \U$30103 ( \30349 , \30347 , \30348 );
not \U$30104 ( \30350 , \30349 );
or \U$30105 ( \30351 , \30339 , \30350 );
nand \U$30106 ( \30352 , \30326 , \30333 );
nand \U$30107 ( \30353 , \30351 , \30352 );
xor \U$30108 ( \30354 , \30320 , \30353 );
not \U$30109 ( \30355 , \30354 );
or \U$30110 ( \30356 , \30297 , \30355 );
nand \U$30111 ( \30357 , \30318 , \30319 );
nand \U$30112 ( \30358 , \30353 , \30357 );
nand \U$30113 ( \30359 , \30356 , \30358 );
not \U$30114 ( \30360 , \30359 );
or \U$30115 ( \30361 , \30289 , \30360 );
or \U$30116 ( \30362 , \30359 , \30288 );
not \U$30117 ( \30363 , \30218 );
nand \U$30118 ( \30364 , \30363 , \30224 );
xor \U$30119 ( \30365 , \30364 , \30222 );
not \U$30120 ( \30366 , \30365 );
xor \U$30121 ( \30367 , RIbe285e8_24, RIbe2b3d8_122);
not \U$30122 ( \30368 , \30367 );
not \U$30123 ( \30369 , \10863 );
or \U$30124 ( \30370 , \30368 , \30369 );
nand \U$30125 ( \30371 , \2625 , \30104 );
nand \U$30126 ( \30372 , \30370 , \30371 );
or \U$30127 ( \30373 , RIbe285e8_24, RIbe287c8_28);
nand \U$30128 ( \30374 , \30373 , RIbe2ae38_110);
nand \U$30129 ( \30375 , RIbe285e8_24, RIbe287c8_28);
nand \U$30130 ( \30376 , \30374 , \30375 , RIbe28480_21);
not \U$30131 ( \30377 , \30376 );
and \U$30132 ( \30378 , \30372 , \30377 );
not \U$30133 ( \30379 , \30378 );
xor \U$30134 ( \30380 , RIbe28480_21, RIbe2aeb0_111);
not \U$30135 ( \30381 , \30380 );
not \U$30136 ( \30382 , \2518 );
or \U$30137 ( \30383 , \30381 , \30382 );
not \U$30138 ( \30384 , \2526 );
nand \U$30139 ( \30385 , \30384 , \29682 );
nand \U$30140 ( \30386 , \30383 , \30385 );
xor \U$30141 ( \30387 , RIbe27fd0_11, RIbe2ac58_106);
not \U$30142 ( \30388 , \30387 );
not \U$30143 ( \30389 , \10466 );
or \U$30144 ( \30390 , \30388 , \30389 );
nand \U$30145 ( \30391 , \2707 , \29695 );
nand \U$30146 ( \30392 , \30390 , \30391 );
xor \U$30147 ( \30393 , \30386 , \30392 );
not \U$30148 ( \30394 , \30393 );
or \U$30149 ( \30395 , \30379 , \30394 );
nand \U$30150 ( \30396 , \30392 , \30386 );
nand \U$30151 ( \30397 , \30395 , \30396 );
not \U$30152 ( \30398 , \30397 );
not \U$30153 ( \30399 , \30398 );
xor \U$30154 ( \30400 , \29657 , \29663 );
xor \U$30155 ( \30401 , \30400 , \29671 );
not \U$30156 ( \30402 , \30401 );
or \U$30157 ( \30403 , \30399 , \30402 );
or \U$30158 ( \30404 , \30401 , \30398 );
nand \U$30159 ( \30405 , \30403 , \30404 );
not \U$30160 ( \30406 , \30405 );
or \U$30161 ( \30407 , \30366 , \30406 );
nand \U$30162 ( \30408 , \30401 , \30397 );
nand \U$30163 ( \30409 , \30407 , \30408 );
nand \U$30164 ( \30410 , \30362 , \30409 );
nand \U$30165 ( \30411 , \30361 , \30410 );
not \U$30166 ( \30412 , \30411 );
or \U$30167 ( \30413 , \30287 , \30412 );
not \U$30168 ( \30414 , \30285 );
or \U$30169 ( \30415 , \30411 , \30414 );
nand \U$30170 ( \30416 , \30413 , \30415 );
not \U$30171 ( \30417 , \30416 );
or \U$30172 ( \30418 , \30070 , \30417 );
not \U$30173 ( \30419 , \30414 );
nand \U$30174 ( \30420 , \30419 , \30411 );
nand \U$30175 ( \30421 , \30418 , \30420 );
not \U$30176 ( \30422 , \30421 );
xor \U$30177 ( \30423 , \29599 , \29592 );
xor \U$30178 ( \30424 , \30423 , \29608 );
not \U$30179 ( \30425 , \30424 );
xor \U$30180 ( \30426 , \29978 , \29987 );
not \U$30181 ( \30427 , \30426 );
and \U$30182 ( \30428 , \30247 , \30257 );
and \U$30183 ( \30429 , \30240 , \30246 );
nor \U$30184 ( \30430 , \30428 , \30429 );
not \U$30185 ( \30431 , \30430 );
or \U$30186 ( \30432 , \30427 , \30431 );
or \U$30187 ( \30433 , \30430 , \30426 );
nand \U$30188 ( \30434 , \30432 , \30433 );
not \U$30189 ( \30435 , \30434 );
or \U$30190 ( \30436 , \30425 , \30435 );
not \U$30191 ( \30437 , \30430 );
nand \U$30192 ( \30438 , \30437 , \30426 );
nand \U$30193 ( \30439 , \30436 , \30438 );
not \U$30194 ( \30440 , \30180 );
not \U$30195 ( \30441 , \30205 );
or \U$30196 ( \30442 , \30440 , \30441 );
not \U$30197 ( \30443 , \30206 );
not \U$30198 ( \30444 , \30181 );
or \U$30199 ( \30445 , \30443 , \30444 );
nand \U$30200 ( \30446 , \30445 , \30225 );
nand \U$30201 ( \30447 , \30442 , \30446 );
or \U$30202 ( \30448 , \30439 , \30447 );
xor \U$30203 ( \30449 , \29537 , \29544 );
xor \U$30204 ( \30450 , \30449 , \29551 );
xor \U$30205 ( \30451 , \29560 , \29570 );
xor \U$30206 ( \30452 , \30451 , \29578 );
xor \U$30207 ( \30453 , \30450 , \30452 );
xor \U$30208 ( \30454 , \29451 , \29443 );
xor \U$30209 ( \30455 , \30454 , \29436 );
and \U$30210 ( \30456 , \30453 , \30455 );
and \U$30211 ( \30457 , \30450 , \30452 );
or \U$30212 ( \30458 , \30456 , \30457 );
nand \U$30213 ( \30459 , \30448 , \30458 );
nand \U$30214 ( \30460 , \30439 , \30447 );
nand \U$30215 ( \30461 , \30459 , \30460 );
not \U$30216 ( \30462 , \30067 );
not \U$30217 ( \30463 , \30060 );
or \U$30218 ( \30464 , \30462 , \30463 );
not \U$30219 ( \30465 , \30056 );
nand \U$30220 ( \30466 , \30465 , \30050 );
nand \U$30221 ( \30467 , \30464 , \30466 );
xor \U$30222 ( \30468 , \30461 , \30467 );
not \U$30223 ( \30469 , \30468 );
not \U$30224 ( \30470 , \29838 );
not \U$30225 ( \30471 , \29863 );
and \U$30226 ( \30472 , \30470 , \30471 );
and \U$30227 ( \30473 , \29838 , \29863 );
nor \U$30228 ( \30474 , \30472 , \30473 );
not \U$30229 ( \30475 , \30474 );
not \U$30230 ( \30476 , \29991 );
not \U$30231 ( \30477 , \29972 );
or \U$30232 ( \30478 , \30476 , \30477 );
or \U$30233 ( \30479 , \29991 , \29972 );
nand \U$30234 ( \30480 , \30479 , \30002 );
nand \U$30235 ( \30481 , \30478 , \30480 );
not \U$30236 ( \30482 , \30481 );
or \U$30237 ( \30483 , \30475 , \30482 );
or \U$30238 ( \30484 , \30481 , \30474 );
nand \U$30239 ( \30485 , \30483 , \30484 );
buf \U$30240 ( \30486 , \30485 );
xor \U$30241 ( \30487 , \29354 , \29330 );
xnor \U$30242 ( \30488 , \30487 , \29364 );
not \U$30243 ( \30489 , \30488 );
and \U$30244 ( \30490 , \30486 , \30489 );
not \U$30245 ( \30491 , \30486 );
and \U$30246 ( \30492 , \30491 , \30488 );
nor \U$30247 ( \30493 , \30490 , \30492 );
not \U$30248 ( \30494 , \30493 );
and \U$30249 ( \30495 , \30469 , \30494 );
and \U$30250 ( \30496 , \30468 , \30493 );
nor \U$30251 ( \30497 , \30495 , \30496 );
not \U$30252 ( \30498 , \30497 );
or \U$30253 ( \30499 , \30422 , \30498 );
or \U$30254 ( \30500 , \30497 , \30421 );
nand \U$30255 ( \30501 , \30499 , \30500 );
not \U$30256 ( \30502 , \30501 );
or \U$30257 ( \30503 , \30048 , \30502 );
not \U$30258 ( \30504 , \30497 );
nand \U$30259 ( \30505 , \30504 , \30421 );
nand \U$30260 ( \30506 , \30503 , \30505 );
xor \U$30261 ( \30507 , \29900 , \30506 );
not \U$30262 ( \30508 , \25216 );
not \U$30263 ( \30509 , \25214 );
nand \U$30264 ( \30510 , \30509 , \25218 );
not \U$30265 ( \30511 , \30510 );
or \U$30266 ( \30512 , \30508 , \30511 );
or \U$30267 ( \30513 , \30510 , \25216 );
nand \U$30268 ( \30514 , \30512 , \30513 );
not \U$30269 ( \30515 , \30514 );
xor \U$30270 ( \30516 , \25093 , \25158 );
xnor \U$30271 ( \30517 , \30516 , \25124 );
not \U$30272 ( \30518 , \30517 );
not \U$30273 ( \30519 , \30518 );
or \U$30274 ( \30520 , \30515 , \30519 );
not \U$30275 ( \30521 , \30514 );
nand \U$30276 ( \30522 , \30521 , \30517 );
nand \U$30277 ( \30523 , \30520 , \30522 );
not \U$30278 ( \30524 , \25057 );
nand \U$30279 ( \30525 , \30524 , \25089 );
not \U$30280 ( \30526 , \30525 );
not \U$30281 ( \30527 , \25087 );
and \U$30282 ( \30528 , \30526 , \30527 );
and \U$30283 ( \30529 , \30525 , \25087 );
nor \U$30284 ( \30530 , \30528 , \30529 );
not \U$30285 ( \30531 , \30530 );
and \U$30286 ( \30532 , \30523 , \30531 );
not \U$30287 ( \30533 , \30523 );
and \U$30288 ( \30534 , \30533 , \30530 );
nor \U$30289 ( \30535 , \30532 , \30534 );
xor \U$30290 ( \30536 , \30032 , \30033 );
and \U$30291 ( \30537 , \30536 , \30039 );
and \U$30292 ( \30538 , \30032 , \30033 );
or \U$30293 ( \30539 , \30537 , \30538 );
not \U$30294 ( \30540 , \30539 );
not \U$30295 ( \30541 , \30488 );
not \U$30296 ( \30542 , \30485 );
or \U$30297 ( \30543 , \30541 , \30542 );
not \U$30298 ( \30544 , \30474 );
nand \U$30299 ( \30545 , \30544 , \30481 );
nand \U$30300 ( \30546 , \30543 , \30545 );
not \U$30301 ( \30547 , \30546 );
and \U$30302 ( \30548 , \30540 , \30547 );
not \U$30303 ( \30549 , \30540 );
and \U$30304 ( \30550 , \30549 , \30546 );
nor \U$30305 ( \30551 , \30548 , \30550 );
xor \U$30306 ( \30552 , \30535 , \30551 );
not \U$30307 ( \30553 , \30493 );
not \U$30308 ( \30554 , \30553 );
not \U$30309 ( \30555 , \30468 );
or \U$30310 ( \30556 , \30554 , \30555 );
nand \U$30311 ( \30557 , \30467 , \30461 );
nand \U$30312 ( \30558 , \30556 , \30557 );
xnor \U$30313 ( \30559 , \30552 , \30558 );
not \U$30314 ( \30560 , \30045 );
not \U$30315 ( \30561 , \30041 );
or \U$30316 ( \30562 , \30560 , \30561 );
nand \U$30317 ( \30563 , \30040 , \30016 );
nand \U$30318 ( \30564 , \30562 , \30563 );
and \U$30319 ( \30565 , \30559 , \30564 );
not \U$30320 ( \30566 , \30559 );
not \U$30321 ( \30567 , \30564 );
and \U$30322 ( \30568 , \30566 , \30567 );
nor \U$30323 ( \30569 , \30565 , \30568 );
xor \U$30324 ( \30570 , \30507 , \30569 );
not \U$30325 ( \30571 , \29901 );
not \U$30326 ( \30572 , \30571 );
not \U$30327 ( \30573 , \30011 );
or \U$30328 ( \30574 , \30572 , \30573 );
or \U$30329 ( \30575 , \30011 , \30571 );
nand \U$30330 ( \30576 , \30574 , \30575 );
not \U$30331 ( \30577 , \30576 );
xor \U$30332 ( \30578 , \30439 , \30458 );
xnor \U$30333 ( \30579 , \30578 , \30447 );
not \U$30334 ( \30580 , \30579 );
and \U$30335 ( \30581 , \30577 , \30580 );
and \U$30336 ( \30582 , \30576 , \30579 );
nor \U$30337 ( \30583 , \30581 , \30582 );
not \U$30338 ( \30584 , \30583 );
not \U$30339 ( \30585 , \30584 );
xnor \U$30340 ( \30586 , \30434 , \30424 );
not \U$30341 ( \30587 , \30586 );
xor \U$30342 ( \30588 , \30450 , \30452 );
xor \U$30343 ( \30589 , \30588 , \30455 );
not \U$30344 ( \30590 , \30589 );
and \U$30345 ( \30591 , \30587 , \30590 );
and \U$30346 ( \30592 , \30586 , \30589 );
nor \U$30347 ( \30593 , \30591 , \30592 );
not \U$30348 ( \30594 , \30593 );
not \U$30349 ( \30595 , \30594 );
xor \U$30350 ( \30596 , RIbe27b20_1, RIbe2b180_117);
nand \U$30351 ( \30597 , \14849 , \30596 );
or \U$30352 ( \30598 , \30597 , \14845 );
nand \U$30353 ( \30599 , \14845 , \30128 );
nand \U$30354 ( \30600 , \30598 , \30599 );
xor \U$30355 ( \30601 , RIbe28f48_44, RIbe2a640_93);
nand \U$30356 ( \30602 , \3253 , \30601 );
or \U$30357 ( \30603 , \30602 , \3248 );
nand \U$30358 ( \30604 , \3248 , \30304 );
nand \U$30359 ( \30605 , \30603 , \30604 );
xor \U$30360 ( \30606 , \30600 , \30605 );
xor \U$30361 ( \30607 , RIbe27e68_8, RIbe2a730_95);
not \U$30362 ( \30608 , \30607 );
not \U$30363 ( \30609 , \2458 );
or \U$30364 ( \30610 , \30608 , \30609 );
nand \U$30365 ( \30611 , \13306 , \30312 );
nand \U$30366 ( \30612 , \30610 , \30611 );
and \U$30367 ( \30613 , \30606 , \30612 );
and \U$30368 ( \30614 , \30605 , \30600 );
nor \U$30369 ( \30615 , \30613 , \30614 );
not \U$30370 ( \30616 , \30615 );
not \U$30371 ( \30617 , \30616 );
xor \U$30372 ( \30618 , RIbe2abe0_105, RIbe27fd0_11);
and \U$30373 ( \30619 , \30618 , \10466 );
and \U$30374 ( \30620 , \2707 , \30387 );
nor \U$30375 ( \30621 , \30619 , \30620 );
not \U$30376 ( \30622 , \30621 );
not \U$30377 ( \30623 , \30622 );
xor \U$30378 ( \30624 , RIbe2ae38_110, RIbe28480_21);
and \U$30379 ( \30625 , \16953 , \30624 );
not \U$30380 ( \30626 , \30380 );
nor \U$30381 ( \30627 , \30626 , \2670 );
nor \U$30382 ( \30628 , \30625 , \30627 );
not \U$30383 ( \30629 , \30628 );
xor \U$30384 ( \30630 , RIbe27df0_7, RIbe2aaf0_103);
not \U$30385 ( \30631 , \30630 );
not \U$30386 ( \30632 , \18832 );
or \U$30387 ( \30633 , \30631 , \30632 );
nand \U$30388 ( \30634 , \30072 , RIbe2ab68_104);
nand \U$30389 ( \30635 , \30633 , \30634 );
not \U$30390 ( \30636 , \30635 );
or \U$30391 ( \30637 , \30629 , \30636 );
or \U$30392 ( \30638 , \30635 , \30628 );
nand \U$30393 ( \30639 , \30637 , \30638 );
not \U$30394 ( \30640 , \30639 );
or \U$30395 ( \30641 , \30623 , \30640 );
not \U$30396 ( \30642 , \30628 );
nand \U$30397 ( \30643 , \30642 , \30635 );
nand \U$30398 ( \30644 , \30641 , \30643 );
xor \U$30399 ( \30645 , RIbe2a2f8_86, RIbe2b2e8_120);
not \U$30400 ( \30646 , \30645 );
not \U$30401 ( \30647 , \10792 );
or \U$30402 ( \30648 , \30646 , \30647 );
nand \U$30403 ( \30649 , \11094 , \30081 );
nand \U$30404 ( \30650 , \30648 , \30649 );
xor \U$30405 ( \30651 , RIbe29e48_76, RIbe2ad48_108);
not \U$30406 ( \30652 , \30651 );
not \U$30407 ( \30653 , \11039 );
or \U$30408 ( \30654 , \30652 , \30653 );
nand \U$30409 ( \30655 , \7368 , \29928 );
nand \U$30410 ( \30656 , \30654 , \30655 );
xor \U$30411 ( \30657 , \30650 , \30656 );
xor \U$30412 ( \30658 , RIbe2a910_99, RIbe2a820_97);
not \U$30413 ( \30659 , \30658 );
not \U$30414 ( \30660 , \12716 );
or \U$30415 ( \30661 , \30659 , \30660 );
nand \U$30416 ( \30662 , \9726 , \30094 );
nand \U$30417 ( \30663 , \30661 , \30662 );
and \U$30418 ( \30664 , \30657 , \30663 );
and \U$30419 ( \30665 , \30650 , \30656 );
or \U$30420 ( \30666 , \30664 , \30665 );
xor \U$30421 ( \30667 , \30644 , \30666 );
not \U$30422 ( \30668 , \30667 );
or \U$30423 ( \30669 , \30617 , \30668 );
nand \U$30424 ( \30670 , \30666 , \30644 );
nand \U$30425 ( \30671 , \30669 , \30670 );
not \U$30426 ( \30672 , \30671 );
xor \U$30427 ( \30673 , \29955 , \29938 );
not \U$30428 ( \30674 , \30673 );
not \U$30429 ( \30675 , RIbe29ce0_73);
not \U$30430 ( \30676 , RIbe2b108_116);
and \U$30431 ( \30677 , \30675 , \30676 );
and \U$30432 ( \30678 , RIbe29ce0_73, RIbe2b108_116);
nor \U$30433 ( \30679 , \30677 , \30678 );
buf \U$30434 ( \30680 , \30679 );
and \U$30435 ( \30681 , \14297 , \30680 );
not \U$30436 ( \30682 , \30328 );
nor \U$30437 ( \30683 , \30682 , \16876 );
nor \U$30438 ( \30684 , \30681 , \30683 );
not \U$30439 ( \30685 , \30684 );
not \U$30440 ( \30686 , \30685 );
xor \U$30441 ( \30687 , RIbe2aa00_101, RIbe2a550_91);
and \U$30442 ( \30688 , \10432 , \30687 );
and \U$30443 ( \30689 , \11484 , \30298 );
nor \U$30444 ( \30690 , \30688 , \30689 );
not \U$30445 ( \30691 , \30690 );
xor \U$30446 ( \30692 , RIbe2a028_80, RIbe2a460_89);
not \U$30447 ( \30693 , \30692 );
not \U$30448 ( \30694 , \8400 );
or \U$30449 ( \30695 , \30693 , \30694 );
nand \U$30450 ( \30696 , \8930 , \30321 );
nand \U$30451 ( \30697 , \30695 , \30696 );
not \U$30452 ( \30698 , \30697 );
or \U$30453 ( \30699 , \30691 , \30698 );
or \U$30454 ( \30700 , \30697 , \30690 );
nand \U$30455 ( \30701 , \30699 , \30700 );
not \U$30456 ( \30702 , \30701 );
or \U$30457 ( \30703 , \30686 , \30702 );
not \U$30458 ( \30704 , \30690 );
nand \U$30459 ( \30705 , \30704 , \30697 );
nand \U$30460 ( \30706 , \30703 , \30705 );
not \U$30461 ( \30707 , \30706 );
xor \U$30462 ( \30708 , RIbe2b6a8_128, RIbe2a190_83);
not \U$30463 ( \30709 , \30708 );
not \U$30464 ( \30710 , \14730 );
or \U$30465 ( \30711 , \30709 , \30710 );
nand \U$30466 ( \30712 , \13278 , \30344 );
nand \U$30467 ( \30713 , \30711 , \30712 );
not \U$30468 ( \30714 , \30713 );
xor \U$30469 ( \30715 , RIbe29c68_72, RIbe2b4c8_124);
not \U$30470 ( \30716 , \30715 );
not \U$30471 ( \30717 , \14971 );
or \U$30472 ( \30718 , \30716 , \30717 );
nand \U$30473 ( \30719 , \4580 , \29923 );
nand \U$30474 ( \30720 , \30718 , \30719 );
not \U$30475 ( \30721 , \30720 );
xor \U$30476 ( \30722 , RIbe28d68_40, RIbe2b018_114);
not \U$30477 ( \30723 , \19854 );
and \U$30478 ( \30724 , \30722 , \30723 );
and \U$30479 ( \30725 , \21442 , \29913 );
nor \U$30480 ( \30726 , \30724 , \30725 );
not \U$30481 ( \30727 , \30726 );
or \U$30482 ( \30728 , \30721 , \30727 );
or \U$30483 ( \30729 , \30726 , \30720 );
nand \U$30484 ( \30730 , \30728 , \30729 );
not \U$30485 ( \30731 , \30730 );
or \U$30486 ( \30732 , \30714 , \30731 );
not \U$30487 ( \30733 , \30726 );
nand \U$30488 ( \30734 , \30733 , \30720 );
nand \U$30489 ( \30735 , \30732 , \30734 );
xor \U$30490 ( \30736 , RIbe298a8_64, RIbe2af28_112);
not \U$30491 ( \30737 , \30736 );
not \U$30492 ( \30738 , \16913 );
or \U$30493 ( \30739 , \30737 , \30738 );
nand \U$30494 ( \30740 , \17810 , \30141 );
nand \U$30495 ( \30741 , \30739 , \30740 );
not \U$30496 ( \30742 , \30741 );
not \U$30497 ( \30743 , \9095 );
xor \U$30498 ( \30744 , RIbe2a0a0_81, RIbe2a3e8_88);
not \U$30499 ( \30745 , \30744 );
not \U$30500 ( \30746 , \30745 );
and \U$30501 ( \30747 , \30743 , \30746 );
nor \U$30502 ( \30748 , \30135 , \26572 );
nor \U$30503 ( \30749 , \30747 , \30748 );
not \U$30504 ( \30750 , \30749 );
xor \U$30505 ( \30751 , RIbe29ec0_77, RIbe2a280_85);
not \U$30506 ( \30752 , \30751 );
not \U$30507 ( \30753 , \10845 );
or \U$30508 ( \30754 , \30752 , \30753 );
nand \U$30509 ( \30755 , \18667 , \30112 );
nand \U$30510 ( \30756 , \30754 , \30755 );
not \U$30511 ( \30757 , \30756 );
or \U$30512 ( \30758 , \30750 , \30757 );
or \U$30513 ( \30759 , \30756 , \30749 );
nand \U$30514 ( \30760 , \30758 , \30759 );
not \U$30515 ( \30761 , \30760 );
or \U$30516 ( \30762 , \30742 , \30761 );
not \U$30517 ( \30763 , \30749 );
nand \U$30518 ( \30764 , \30763 , \30756 );
nand \U$30519 ( \30765 , \30762 , \30764 );
xor \U$30520 ( \30766 , \30735 , \30765 );
not \U$30521 ( \30767 , \30766 );
or \U$30522 ( \30768 , \30707 , \30767 );
nand \U$30523 ( \30769 , \30735 , \30765 );
nand \U$30524 ( \30770 , \30768 , \30769 );
not \U$30525 ( \30771 , \30770 );
not \U$30526 ( \30772 , \30771 );
or \U$30527 ( \30773 , \30674 , \30772 );
or \U$30528 ( \30774 , \30771 , \30673 );
nand \U$30529 ( \30775 , \30773 , \30774 );
not \U$30530 ( \30776 , \30775 );
or \U$30531 ( \30777 , \30672 , \30776 );
nand \U$30532 ( \30778 , \30770 , \30673 );
nand \U$30533 ( \30779 , \30777 , \30778 );
not \U$30534 ( \30780 , \30779 );
or \U$30535 ( \30781 , \30595 , \30780 );
not \U$30536 ( \30782 , \30586 );
nand \U$30537 ( \30783 , \30782 , \30589 );
nand \U$30538 ( \30784 , \30781 , \30783 );
not \U$30539 ( \30785 , \30784 );
or \U$30540 ( \30786 , \30585 , \30785 );
not \U$30541 ( \30787 , \30579 );
nand \U$30542 ( \30788 , \30787 , \30576 );
nand \U$30543 ( \30789 , \30786 , \30788 );
xor \U$30544 ( \30790 , \30153 , \30233 );
xor \U$30545 ( \30791 , \30790 , \30282 );
not \U$30546 ( \30792 , \30791 );
xor \U$30547 ( \30793 , \30288 , \30359 );
xnor \U$30548 ( \30794 , \30793 , \30409 );
not \U$30549 ( \30795 , \30794 );
or \U$30550 ( \30796 , \30792 , \30795 );
or \U$30551 ( \30797 , \30794 , \30791 );
nand \U$30552 ( \30798 , \30796 , \30797 );
not \U$30553 ( \30799 , \30798 );
and \U$30554 ( \30800 , \30779 , \30594 );
not \U$30555 ( \30801 , \30779 );
and \U$30556 ( \30802 , \30801 , \30593 );
nor \U$30557 ( \30803 , \30800 , \30802 );
not \U$30558 ( \30804 , \30803 );
or \U$30559 ( \30805 , \30799 , \30804 );
not \U$30560 ( \30806 , \30794 );
nand \U$30561 ( \30807 , \30806 , \30791 );
nand \U$30562 ( \30808 , \30805 , \30807 );
not \U$30563 ( \30809 , \30808 );
xor \U$30564 ( \30810 , \30405 , \30365 );
not \U$30565 ( \30811 , \30810 );
xor \U$30566 ( \30812 , \30262 , \30277 );
xor \U$30567 ( \30813 , \30124 , \30102 );
xor \U$30568 ( \30814 , \30813 , \30151 );
xnor \U$30569 ( \30815 , \30812 , \30814 );
not \U$30570 ( \30816 , \30815 );
or \U$30571 ( \30817 , \30811 , \30816 );
nand \U$30572 ( \30818 , \30277 , \30262 );
not \U$30573 ( \30819 , \30818 );
not \U$30574 ( \30820 , \30277 );
nand \U$30575 ( \30821 , \30820 , \30263 );
not \U$30576 ( \30822 , \30821 );
or \U$30577 ( \30823 , \30819 , \30822 );
nand \U$30578 ( \30824 , \30823 , \30814 );
nand \U$30579 ( \30825 , \30817 , \30824 );
not \U$30580 ( \30826 , \30825 );
not \U$30581 ( \30827 , \30295 );
not \U$30582 ( \30828 , \30354 );
or \U$30583 ( \30829 , \30827 , \30828 );
or \U$30584 ( \30830 , \30354 , \30295 );
nand \U$30585 ( \30831 , \30829 , \30830 );
not \U$30586 ( \30832 , \30310 );
nand \U$30587 ( \30833 , \30832 , \30319 );
not \U$30588 ( \30834 , \30833 );
not \U$30589 ( \30835 , \30317 );
and \U$30590 ( \30836 , \30834 , \30835 );
and \U$30591 ( \30837 , \30833 , \30317 );
nor \U$30592 ( \30838 , \30836 , \30837 );
not \U$30593 ( \30839 , \30838 );
not \U$30594 ( \30840 , \30839 );
xor \U$30595 ( \30841 , \30121 , \30110 );
xor \U$30596 ( \30842 , \30841 , \30117 );
not \U$30597 ( \30843 , \30842 );
not \U$30598 ( \30844 , \30843 );
or \U$30599 ( \30845 , \30840 , \30844 );
not \U$30600 ( \30846 , \30842 );
not \U$30601 ( \30847 , \30838 );
or \U$30602 ( \30848 , \30846 , \30847 );
not \U$30603 ( \30849 , \30140 );
nand \U$30604 ( \30850 , \30849 , \30150 );
and \U$30605 ( \30851 , \30850 , \30148 );
not \U$30606 ( \30852 , \30850 );
and \U$30607 ( \30853 , \30852 , \30147 );
nor \U$30608 ( \30854 , \30851 , \30853 );
nand \U$30609 ( \30855 , \30848 , \30854 );
nand \U$30610 ( \30856 , \30845 , \30855 );
nand \U$30611 ( \30857 , \30831 , \30856 );
not \U$30612 ( \30858 , \30079 );
not \U$30613 ( \30859 , \30090 );
or \U$30614 ( \30860 , \30858 , \30859 );
nand \U$30615 ( \30861 , \30087 , \30078 );
nand \U$30616 ( \30862 , \30860 , \30861 );
xnor \U$30617 ( \30863 , \30862 , \30100 );
not \U$30618 ( \30864 , \30863 );
not \U$30619 ( \30865 , \30864 );
not \U$30620 ( \30866 , \30349 );
and \U$30621 ( \30867 , \30338 , \30866 );
not \U$30622 ( \30868 , \30338 );
and \U$30623 ( \30869 , \30868 , \30349 );
nor \U$30624 ( \30870 , \30867 , \30869 );
not \U$30625 ( \30871 , \30870 );
not \U$30626 ( \30872 , \30871 );
or \U$30627 ( \30873 , \30865 , \30872 );
not \U$30628 ( \30874 , \30870 );
not \U$30629 ( \30875 , \30863 );
or \U$30630 ( \30876 , \30874 , \30875 );
not \U$30631 ( \30877 , \29925 );
xor \U$30632 ( \30878 , \29918 , \29933 );
not \U$30633 ( \30879 , \30878 );
or \U$30634 ( \30880 , \30877 , \30879 );
or \U$30635 ( \30881 , \30878 , \29925 );
nand \U$30636 ( \30882 , \30880 , \30881 );
nand \U$30637 ( \30883 , \30876 , \30882 );
nand \U$30638 ( \30884 , \30873 , \30883 );
nand \U$30639 ( \30885 , \30831 , \30884 );
nand \U$30640 ( \30886 , \30856 , \30884 );
and \U$30641 ( \30887 , \30857 , \30885 , \30886 );
nand \U$30642 ( \30888 , \29963 , \29911 );
not \U$30643 ( \30889 , \30888 );
not \U$30644 ( \30890 , \29960 );
and \U$30645 ( \30891 , \30889 , \30890 );
and \U$30646 ( \30892 , \30888 , \29960 );
nor \U$30647 ( \30893 , \30891 , \30892 );
and \U$30648 ( \30894 , \30887 , \30893 );
not \U$30649 ( \30895 , \30887 );
not \U$30650 ( \30896 , \30893 );
and \U$30651 ( \30897 , \30895 , \30896 );
nor \U$30652 ( \30898 , \30894 , \30897 );
not \U$30653 ( \30899 , \30898 );
or \U$30654 ( \30900 , \30826 , \30899 );
not \U$30655 ( \30901 , \30887 );
nand \U$30656 ( \30902 , \30901 , \30896 );
nand \U$30657 ( \30903 , \30900 , \30902 );
not \U$30658 ( \30904 , \30903 );
not \U$30659 ( \30905 , \30068 );
not \U$30660 ( \30906 , \30416 );
or \U$30661 ( \30907 , \30905 , \30906 );
or \U$30662 ( \30908 , \30416 , \30068 );
nand \U$30663 ( \30909 , \30907 , \30908 );
not \U$30664 ( \30910 , \30909 );
not \U$30665 ( \30911 , \30910 );
or \U$30666 ( \30912 , \30904 , \30911 );
not \U$30667 ( \30913 , \30903 );
nand \U$30668 ( \30914 , \30913 , \30909 );
nand \U$30669 ( \30915 , \30912 , \30914 );
not \U$30670 ( \30916 , \30915 );
or \U$30671 ( \30917 , \30809 , \30916 );
nand \U$30672 ( \30918 , \30909 , \30903 );
nand \U$30673 ( \30919 , \30917 , \30918 );
xor \U$30674 ( \30920 , \30789 , \30919 );
xnor \U$30675 ( \30921 , \30501 , \30047 );
not \U$30676 ( \30922 , \30921 );
and \U$30677 ( \30923 , \30920 , \30922 );
and \U$30678 ( \30924 , \30789 , \30919 );
nor \U$30679 ( \30925 , \30923 , \30924 );
nand \U$30680 ( \30926 , \30570 , \30925 );
not \U$30681 ( \30927 , \30920 );
not \U$30682 ( \30928 , \30921 );
and \U$30683 ( \30929 , \30927 , \30928 );
and \U$30684 ( \30930 , \30920 , \30921 );
nor \U$30685 ( \30931 , \30929 , \30930 );
not \U$30686 ( \30932 , \30583 );
not \U$30687 ( \30933 , \30784 );
and \U$30688 ( \30934 , \30932 , \30933 );
and \U$30689 ( \30935 , \30784 , \30583 );
nor \U$30690 ( \30936 , \30934 , \30935 );
not \U$30691 ( \30937 , \30798 );
not \U$30692 ( \30938 , \30937 );
not \U$30693 ( \30939 , \30803 );
or \U$30694 ( \30940 , \30938 , \30939 );
or \U$30695 ( \30941 , \30803 , \30937 );
nand \U$30696 ( \30942 , \30940 , \30941 );
not \U$30697 ( \30943 , \30942 );
not \U$30698 ( \30944 , \30775 );
not \U$30699 ( \30945 , \30671 );
not \U$30700 ( \30946 , \30945 );
and \U$30701 ( \30947 , \30944 , \30946 );
and \U$30702 ( \30948 , \30775 , \30945 );
nor \U$30703 ( \30949 , \30947 , \30948 );
not \U$30704 ( \30950 , \30949 );
not \U$30705 ( \30951 , \30950 );
xor \U$30706 ( \30952 , RIbe29998_66, RIbe2b018_114);
not \U$30707 ( \30953 , \30952 );
not \U$30708 ( \30954 , \22763 );
or \U$30709 ( \30955 , \30953 , \30954 );
nand \U$30710 ( \30956 , \19371 , \30722 );
nand \U$30711 ( \30957 , \30955 , \30956 );
not \U$30712 ( \30958 , \30957 );
xor \U$30713 ( \30959 , RIbe29c68_72, RIbe2a6b8_94);
not \U$30714 ( \30960 , \30959 );
not \U$30715 ( \30961 , \7513 );
or \U$30716 ( \30962 , \30960 , \30961 );
nand \U$30717 ( \30963 , \4580 , \30715 );
nand \U$30718 ( \30964 , \30962 , \30963 );
not \U$30719 ( \30965 , \30964 );
xor \U$30720 ( \30966 , RIbe2a550_91, RIbe2a898_98);
not \U$30721 ( \30967 , \30966 );
not \U$30722 ( \30968 , \10433 );
or \U$30723 ( \30969 , \30967 , \30968 );
nand \U$30724 ( \30970 , \11485 , \30687 );
nand \U$30725 ( \30971 , \30969 , \30970 );
not \U$30726 ( \30972 , \30971 );
not \U$30727 ( \30973 , \30972 );
or \U$30728 ( \30974 , \30965 , \30973 );
or \U$30729 ( \30975 , \30972 , \30964 );
nand \U$30730 ( \30976 , \30974 , \30975 );
not \U$30731 ( \30977 , \30976 );
or \U$30732 ( \30978 , \30958 , \30977 );
nand \U$30733 ( \30979 , \30971 , \30964 );
nand \U$30734 ( \30980 , \30978 , \30979 );
not \U$30735 ( \30981 , \30980 );
xor \U$30736 ( \30982 , RIbe2a910_99, RIbe2a118_82);
not \U$30737 ( \30983 , \30982 );
not \U$30738 ( \30984 , \11453 );
or \U$30739 ( \30985 , \30983 , \30984 );
nand \U$30740 ( \30986 , \11456 , \30658 );
nand \U$30741 ( \30987 , \30985 , \30986 );
not \U$30742 ( \30988 , \30987 );
xor \U$30743 ( \30989 , RIbe27c88_4, RIbe2aaf0_103);
not \U$30744 ( \30990 , \30989 );
not \U$30745 ( \30991 , \18832 );
or \U$30746 ( \30992 , \30990 , \30991 );
nand \U$30747 ( \30993 , \30630 , RIbe2ab68_104);
nand \U$30748 ( \30994 , \30992 , \30993 );
not \U$30749 ( \30995 , \30994 );
xor \U$30750 ( \30996 , RIbe2a2f8_86, RIbe2a4d8_90);
not \U$30751 ( \30997 , \30996 );
not \U$30752 ( \30998 , \14826 );
or \U$30753 ( \30999 , \30997 , \30998 );
nand \U$30754 ( \31000 , \18963 , \30645 );
nand \U$30755 ( \31001 , \30999 , \31000 );
not \U$30756 ( \31002 , \31001 );
not \U$30757 ( \31003 , \31002 );
or \U$30758 ( \31004 , \30995 , \31003 );
not \U$30759 ( \31005 , \30994 );
nand \U$30760 ( \31006 , \31005 , \31001 );
nand \U$30761 ( \31007 , \31004 , \31006 );
not \U$30762 ( \31008 , \31007 );
or \U$30763 ( \31009 , \30988 , \31008 );
not \U$30764 ( \31010 , \31002 );
nand \U$30765 ( \31011 , \31010 , \30994 );
nand \U$30766 ( \31012 , \31009 , \31011 );
not \U$30767 ( \31013 , \31012 );
xor \U$30768 ( \31014 , RIbe2b450_123, RIbe27e68_8);
not \U$30769 ( \31015 , \31014 );
not \U$30770 ( \31016 , \2458 );
or \U$30771 ( \31017 , \31015 , \31016 );
nand \U$30772 ( \31018 , \2603 , \30607 );
nand \U$30773 ( \31019 , \31017 , \31018 );
not \U$30774 ( \31020 , \31019 );
nand \U$30775 ( \31021 , \16676 , RIbe2ae38_110);
not \U$30776 ( \31022 , \31021 );
xor \U$30777 ( \31023 , RIbe29d58_74, RIbe2b108_116);
not \U$30778 ( \31024 , \31023 );
not \U$30779 ( \31025 , \13527 );
or \U$30780 ( \31026 , \31024 , \31025 );
nand \U$30781 ( \31027 , \13533 , \30679 );
nand \U$30782 ( \31028 , \31026 , \31027 );
not \U$30783 ( \31029 , \31028 );
or \U$30784 ( \31030 , \31022 , \31029 );
or \U$30785 ( \31031 , \31028 , \31021 );
nand \U$30786 ( \31032 , \31030 , \31031 );
not \U$30787 ( \31033 , \31032 );
or \U$30788 ( \31034 , \31020 , \31033 );
not \U$30789 ( \31035 , \31021 );
nand \U$30790 ( \31036 , \31035 , \31028 );
nand \U$30791 ( \31037 , \31034 , \31036 );
not \U$30792 ( \31038 , \31037 );
not \U$30793 ( \31039 , \31038 );
or \U$30794 ( \31040 , \31013 , \31039 );
or \U$30795 ( \31041 , \31038 , \31012 );
nand \U$30796 ( \31042 , \31040 , \31041 );
not \U$30797 ( \31043 , \31042 );
or \U$30798 ( \31044 , \30981 , \31043 );
not \U$30799 ( \31045 , \31038 );
nand \U$30800 ( \31046 , \31045 , \31012 );
nand \U$30801 ( \31047 , \31044 , \31046 );
not \U$30802 ( \31048 , \31047 );
xor \U$30803 ( \31049 , \30378 , \30393 );
not \U$30804 ( \31050 , \31049 );
xor \U$30805 ( \31051 , RIbe2adc0_109, RIbe2a028_80);
not \U$30806 ( \31052 , \31051 );
not \U$30807 ( \31053 , \14513 );
or \U$30808 ( \31054 , \31052 , \31053 );
nand \U$30809 ( \31055 , \8172 , \30692 );
nand \U$30810 ( \31056 , \31054 , \31055 );
xor \U$30811 ( \31057 , RIbe2a3e8_88, RIbe2b360_121);
not \U$30812 ( \31058 , \31057 );
not \U$30813 ( \31059 , \9262 );
or \U$30814 ( \31060 , \31058 , \31059 );
nand \U$30815 ( \31061 , \9089 , \30744 );
nand \U$30816 ( \31062 , \31060 , \31061 );
or \U$30817 ( \31063 , \31056 , \31062 );
xor \U$30818 ( \31064 , RIbe29e48_76, RIbe2b540_125);
not \U$30819 ( \31065 , \31064 );
not \U$30820 ( \31066 , \4842 );
or \U$30821 ( \31067 , \31065 , \31066 );
nand \U$30822 ( \31068 , \4849 , \30651 );
nand \U$30823 ( \31069 , \31067 , \31068 );
nand \U$30824 ( \31070 , \31063 , \31069 );
nand \U$30825 ( \31071 , \31056 , \31062 );
nand \U$30826 ( \31072 , \31070 , \31071 );
not \U$30827 ( \31073 , \31072 );
xor \U$30828 ( \31074 , RIbe285e8_24, RIbe2aeb0_111);
not \U$30829 ( \31075 , \31074 );
not \U$30830 ( \31076 , \10863 );
or \U$30831 ( \31077 , \31075 , \31076 );
nand \U$30832 ( \31078 , \2758 , \30367 );
nand \U$30833 ( \31079 , \31077 , \31078 );
not \U$30834 ( \31080 , \31079 );
xor \U$30835 ( \31081 , RIbe2af28_112, RIbe28cf0_39);
not \U$30836 ( \31082 , \31081 );
not \U$30837 ( \31083 , \14423 );
or \U$30838 ( \31084 , \31082 , \31083 );
nand \U$30839 ( \31085 , \17809 , \30736 );
nand \U$30840 ( \31086 , \31084 , \31085 );
not \U$30841 ( \31087 , \31086 );
or \U$30842 ( \31088 , \31080 , \31087 );
or \U$30843 ( \31089 , \31086 , \31079 );
xor \U$30844 ( \31090 , RIbe28f48_44, RIbe2ac58_106);
not \U$30845 ( \31091 , \31090 );
not \U$30846 ( \31092 , \23097 );
or \U$30847 ( \31093 , \31091 , \31092 );
nand \U$30848 ( \31094 , \9524 , \30601 );
nand \U$30849 ( \31095 , \31093 , \31094 );
nand \U$30850 ( \31096 , \31089 , \31095 );
nand \U$30851 ( \31097 , \31088 , \31096 );
not \U$30852 ( \31098 , \31097 );
and \U$30853 ( \31099 , \30372 , \30376 );
not \U$30854 ( \31100 , \30372 );
and \U$30855 ( \31101 , \31100 , \30377 );
nor \U$30856 ( \31102 , \31099 , \31101 );
not \U$30857 ( \31103 , \31102 );
or \U$30858 ( \31104 , \31098 , \31103 );
or \U$30859 ( \31105 , \31102 , \31097 );
nand \U$30860 ( \31106 , \31104 , \31105 );
not \U$30861 ( \31107 , \31106 );
or \U$30862 ( \31108 , \31073 , \31107 );
not \U$30863 ( \31109 , \31102 );
nand \U$30864 ( \31110 , \31109 , \31097 );
nand \U$30865 ( \31111 , \31108 , \31110 );
not \U$30866 ( \31112 , \31111 );
not \U$30867 ( \31113 , \31112 );
or \U$30868 ( \31114 , \31050 , \31113 );
or \U$30869 ( \31115 , \31112 , \31049 );
nand \U$30870 ( \31116 , \31114 , \31115 );
not \U$30871 ( \31117 , \31116 );
or \U$30872 ( \31118 , \31048 , \31117 );
not \U$30873 ( \31119 , \31112 );
nand \U$30874 ( \31120 , \31119 , \31049 );
nand \U$30875 ( \31121 , \31118 , \31120 );
not \U$30876 ( \31122 , \31121 );
xor \U$30877 ( \31123 , \30706 , \30766 );
not \U$30878 ( \31124 , \31123 );
not \U$30879 ( \31125 , \30612 );
not \U$30880 ( \31126 , \30606 );
not \U$30881 ( \31127 , \31126 );
or \U$30882 ( \31128 , \31125 , \31127 );
not \U$30883 ( \31129 , \30612 );
nand \U$30884 ( \31130 , \31129 , \30606 );
nand \U$30885 ( \31131 , \31128 , \31130 );
not \U$30886 ( \31132 , \31131 );
not \U$30887 ( \31133 , \30639 );
not \U$30888 ( \31134 , \30621 );
and \U$30889 ( \31135 , \31133 , \31134 );
and \U$30890 ( \31136 , \30639 , \30621 );
nor \U$30891 ( \31137 , \31135 , \31136 );
nand \U$30892 ( \31138 , \31132 , \31137 );
not \U$30893 ( \31139 , \31138 );
xor \U$30894 ( \31140 , \30730 , \30713 );
not \U$30895 ( \31141 , \31140 );
or \U$30896 ( \31142 , \31139 , \31141 );
not \U$30897 ( \31143 , \31137 );
nand \U$30898 ( \31144 , \31131 , \31143 );
nand \U$30899 ( \31145 , \31142 , \31144 );
not \U$30900 ( \31146 , \31145 );
not \U$30901 ( \31147 , \30684 );
not \U$30902 ( \31148 , \30701 );
or \U$30903 ( \31149 , \31147 , \31148 );
or \U$30904 ( \31150 , \30701 , \30684 );
nand \U$30905 ( \31151 , \31149 , \31150 );
not \U$30906 ( \31152 , \30741 );
not \U$30907 ( \31153 , \30760 );
not \U$30908 ( \31154 , \31153 );
or \U$30909 ( \31155 , \31152 , \31154 );
not \U$30910 ( \31156 , \30741 );
nand \U$30911 ( \31157 , \31156 , \30760 );
nand \U$30912 ( \31158 , \31155 , \31157 );
or \U$30913 ( \31159 , \31151 , \31158 );
xor \U$30914 ( \31160 , RIbe2aa78_102, RIbe2a190_83);
not \U$30915 ( \31161 , \31160 );
not \U$30916 ( \31162 , \10690 );
or \U$30917 ( \31163 , \31161 , \31162 );
nand \U$30918 ( \31164 , \15693 , \30708 );
nand \U$30919 ( \31165 , \31163 , \31164 );
not \U$30920 ( \31166 , \31165 );
and \U$30921 ( \31167 , \2707 , \30618 );
xor \U$30922 ( \31168 , RIbe27fd0_11, RIbe2a7a8_96);
not \U$30923 ( \31169 , \31168 );
nor \U$30924 ( \31170 , \31169 , \9081 );
nor \U$30925 ( \31171 , \31167 , \31170 );
not \U$30926 ( \31172 , \31171 );
xor \U$30927 ( \31173 , RIbe29f38_78, RIbe2a280_85);
not \U$30928 ( \31174 , \31173 );
not \U$30929 ( \31175 , \27992 );
or \U$30930 ( \31176 , \31174 , \31175 );
nand \U$30931 ( \31177 , \18667 , \30751 );
nand \U$30932 ( \31178 , \31176 , \31177 );
not \U$30933 ( \31179 , \31178 );
or \U$30934 ( \31180 , \31172 , \31179 );
or \U$30935 ( \31181 , \31178 , \31171 );
nand \U$30936 ( \31182 , \31180 , \31181 );
not \U$30937 ( \31183 , \31182 );
or \U$30938 ( \31184 , \31166 , \31183 );
not \U$30939 ( \31185 , \31171 );
nand \U$30940 ( \31186 , \31185 , \31178 );
nand \U$30941 ( \31187 , \31184 , \31186 );
nand \U$30942 ( \31188 , \31159 , \31187 );
nand \U$30943 ( \31189 , \31151 , \31158 );
nand \U$30944 ( \31190 , \31188 , \31189 );
not \U$30945 ( \31191 , \31190 );
not \U$30946 ( \31192 , \31191 );
or \U$30947 ( \31193 , \31146 , \31192 );
or \U$30948 ( \31194 , \31191 , \31145 );
nand \U$30949 ( \31195 , \31193 , \31194 );
not \U$30950 ( \31196 , \31195 );
or \U$30951 ( \31197 , \31124 , \31196 );
not \U$30952 ( \31198 , \31191 );
nand \U$30953 ( \31199 , \31198 , \31145 );
nand \U$30954 ( \31200 , \31197 , \31199 );
not \U$30955 ( \31201 , \31200 );
not \U$30956 ( \31202 , \31201 );
or \U$30957 ( \31203 , \31122 , \31202 );
not \U$30958 ( \31204 , \31121 );
nand \U$30959 ( \31205 , \31204 , \31200 );
nand \U$30960 ( \31206 , \31203 , \31205 );
not \U$30961 ( \31207 , \31206 );
or \U$30962 ( \31208 , \30951 , \31207 );
nand \U$30963 ( \31209 , \31200 , \31121 );
nand \U$30964 ( \31210 , \31208 , \31209 );
not \U$30965 ( \31211 , \31210 );
xnor \U$30966 ( \31212 , \30825 , \30898 );
not \U$30967 ( \31213 , \31212 );
or \U$30968 ( \31214 , \31211 , \31213 );
or \U$30969 ( \31215 , \31212 , \31210 );
nand \U$30970 ( \31216 , \31214 , \31215 );
not \U$30971 ( \31217 , \31216 );
or \U$30972 ( \31218 , \30943 , \31217 );
not \U$30973 ( \31219 , \31212 );
nand \U$30974 ( \31220 , \31219 , \31210 );
nand \U$30975 ( \31221 , \31218 , \31220 );
not \U$30976 ( \31222 , \31221 );
xor \U$30977 ( \31223 , \30936 , \31222 );
not \U$30978 ( \31224 , \30808 );
and \U$30979 ( \31225 , \30915 , \31224 );
not \U$30980 ( \31226 , \30915 );
and \U$30981 ( \31227 , \31226 , \30808 );
nor \U$30982 ( \31228 , \31225 , \31227 );
and \U$30983 ( \31229 , \31223 , \31228 );
and \U$30984 ( \31230 , \30936 , \31222 );
or \U$30985 ( \31231 , \31229 , \31230 );
nand \U$30986 ( \31232 , \30931 , \31231 );
and \U$30987 ( \31233 , \31206 , \30950 );
not \U$30988 ( \31234 , \31206 );
and \U$30989 ( \31235 , \31234 , \30949 );
nor \U$30990 ( \31236 , \31233 , \31235 );
and \U$30991 ( \31237 , \30854 , \30838 );
not \U$30992 ( \31238 , \30854 );
and \U$30993 ( \31239 , \31238 , \30839 );
or \U$30994 ( \31240 , \31237 , \31239 );
and \U$30995 ( \31241 , \31240 , \30842 );
not \U$30996 ( \31242 , \31240 );
and \U$30997 ( \31243 , \31242 , \30843 );
nor \U$30998 ( \31244 , \31241 , \31243 );
not \U$30999 ( \31245 , \31244 );
not \U$31000 ( \31246 , \30870 );
not \U$31001 ( \31247 , \30864 );
or \U$31002 ( \31248 , \31246 , \31247 );
nand \U$31003 ( \31249 , \30863 , \30871 );
nand \U$31004 ( \31250 , \31248 , \31249 );
not \U$31005 ( \31251 , \30882 );
and \U$31006 ( \31252 , \31250 , \31251 );
not \U$31007 ( \31253 , \31250 );
and \U$31008 ( \31254 , \31253 , \30882 );
nor \U$31009 ( \31255 , \31252 , \31254 );
not \U$31010 ( \31256 , \31255 );
not \U$31011 ( \31257 , \31256 );
not \U$31012 ( \31258 , \30615 );
not \U$31013 ( \31259 , \30667 );
or \U$31014 ( \31260 , \31258 , \31259 );
or \U$31015 ( \31261 , \30667 , \30615 );
nand \U$31016 ( \31262 , \31260 , \31261 );
not \U$31017 ( \31263 , \31262 );
not \U$31018 ( \31264 , \31263 );
or \U$31019 ( \31265 , \31257 , \31264 );
nand \U$31020 ( \31266 , \31262 , \31255 );
nand \U$31021 ( \31267 , \31265 , \31266 );
not \U$31022 ( \31268 , \31267 );
or \U$31023 ( \31269 , \31245 , \31268 );
or \U$31024 ( \31270 , \31267 , \31244 );
nand \U$31025 ( \31271 , \31269 , \31270 );
not \U$31026 ( \31272 , \31271 );
xnor \U$31027 ( \31273 , \31123 , \31195 );
not \U$31028 ( \31274 , \31273 );
buf \U$31029 ( \31275 , \31158 );
xor \U$31030 ( \31276 , \31151 , \31275 );
xor \U$31031 ( \31277 , \31276 , \31187 );
not \U$31032 ( \31278 , \31277 );
buf \U$31033 ( \31279 , \31072 );
xor \U$31034 ( \31280 , \31106 , \31279 );
not \U$31035 ( \31281 , \31280 );
xor \U$31036 ( \31282 , \31131 , \31143 );
xnor \U$31037 ( \31283 , \31282 , \31140 );
not \U$31038 ( \31284 , \31283 );
or \U$31039 ( \31285 , \31281 , \31284 );
or \U$31040 ( \31286 , \31283 , \31280 );
nand \U$31041 ( \31287 , \31285 , \31286 );
not \U$31042 ( \31288 , \31287 );
or \U$31043 ( \31289 , \31278 , \31288 );
not \U$31044 ( \31290 , \31283 );
nand \U$31045 ( \31291 , \31290 , \31280 );
nand \U$31046 ( \31292 , \31289 , \31291 );
not \U$31047 ( \31293 , \31292 );
or \U$31048 ( \31294 , \31274 , \31293 );
or \U$31049 ( \31295 , \31292 , \31273 );
nand \U$31050 ( \31296 , \31294 , \31295 );
not \U$31051 ( \31297 , \31296 );
or \U$31052 ( \31298 , \31272 , \31297 );
not \U$31053 ( \31299 , \31273 );
nand \U$31054 ( \31300 , \31299 , \31292 );
nand \U$31055 ( \31301 , \31298 , \31300 );
xor \U$31056 ( \31302 , \31236 , \31301 );
xor \U$31057 ( \31303 , \30650 , \30656 );
xor \U$31058 ( \31304 , \31303 , \30663 );
not \U$31059 ( \31305 , \31304 );
xor \U$31060 ( \31306 , RIbe29b78_70, RIbe2b180_117);
not \U$31061 ( \31307 , \31306 );
not \U$31062 ( \31308 , \14852 );
or \U$31063 ( \31309 , \31307 , \31308 );
nand \U$31064 ( \31310 , \21759 , \30596 );
nand \U$31065 ( \31311 , \31309 , \31310 );
xor \U$31066 ( \31312 , RIbe2b3d8_122, RIbe27e68_8);
not \U$31067 ( \31313 , \31312 );
not \U$31068 ( \31314 , \2457 );
or \U$31069 ( \31315 , \31313 , \31314 );
nand \U$31070 ( \31316 , \2463 , \31014 );
nand \U$31071 ( \31317 , \31315 , \31316 );
or \U$31072 ( \31318 , RIbe27e68_8, RIbe28660_25);
nand \U$31073 ( \31319 , \31318 , RIbe2ae38_110);
nand \U$31074 ( \31320 , RIbe27e68_8, RIbe28660_25);
nand \U$31075 ( \31321 , \31319 , \31320 , RIbe285e8_24);
not \U$31076 ( \31322 , \31321 );
and \U$31077 ( \31323 , \31317 , \31322 );
xor \U$31078 ( \31324 , \31311 , \31323 );
xor \U$31079 ( \31325 , RIbe285e8_24, RIbe2ae38_110);
not \U$31080 ( \31326 , \31325 );
not \U$31081 ( \31327 , \10863 );
or \U$31082 ( \31328 , \31326 , \31327 );
nand \U$31083 ( \31329 , \8270 , \31074 );
nand \U$31084 ( \31330 , \31328 , \31329 );
xor \U$31085 ( \31331 , RIbe2a3e8_88, RIbe2b2e8_120);
not \U$31086 ( \31332 , \31331 );
not \U$31087 ( \31333 , \8805 );
or \U$31088 ( \31334 , \31332 , \31333 );
nand \U$31089 ( \31335 , \9089 , \31057 );
nand \U$31090 ( \31336 , \31334 , \31335 );
nor \U$31091 ( \31337 , \31330 , \31336 );
xor \U$31092 ( \31338 , RIbe27b20_1, RIbe2af28_112);
and \U$31093 ( \31339 , \31338 , \16913 );
and \U$31094 ( \31340 , \17810 , \31081 );
nor \U$31095 ( \31341 , \31339 , \31340 );
or \U$31096 ( \31342 , \31337 , \31341 );
nand \U$31097 ( \31343 , \31330 , \31336 );
nand \U$31098 ( \31344 , \31342 , \31343 );
and \U$31099 ( \31345 , \31324 , \31344 );
and \U$31100 ( \31346 , \31311 , \31323 );
nor \U$31101 ( \31347 , \31345 , \31346 );
not \U$31102 ( \31348 , \31347 );
and \U$31103 ( \31349 , \31305 , \31348 );
and \U$31104 ( \31350 , \31347 , \31304 );
nor \U$31105 ( \31351 , \31349 , \31350 );
not \U$31106 ( \31352 , \31351 );
not \U$31107 ( \31353 , \31352 );
xor \U$31108 ( \31354 , RIbe2aa00_101, RIbe2a190_83);
not \U$31109 ( \31355 , \31354 );
not \U$31110 ( \31356 , \15690 );
or \U$31111 ( \31357 , \31355 , \31356 );
not \U$31112 ( \31358 , \11971 );
nand \U$31113 ( \31359 , \31358 , \31160 );
nand \U$31114 ( \31360 , \31357 , \31359 );
not \U$31115 ( \31361 , \31360 );
xor \U$31116 ( \31362 , RIbe2a730_95, RIbe27fd0_11);
not \U$31117 ( \31363 , \31362 );
not \U$31118 ( \31364 , \9825 );
or \U$31119 ( \31365 , \31363 , \31364 );
nand \U$31120 ( \31366 , \2707 , \31168 );
nand \U$31121 ( \31367 , \31365 , \31366 );
xor \U$31122 ( \31368 , RIbe2a640_93, RIbe29c68_72);
not \U$31123 ( \31369 , \31368 );
not \U$31124 ( \31370 , \4578 );
or \U$31125 ( \31371 , \31369 , \31370 );
nand \U$31126 ( \31372 , \7237 , \30959 );
nand \U$31127 ( \31373 , \31371 , \31372 );
xor \U$31128 ( \31374 , \31367 , \31373 );
not \U$31129 ( \31375 , \31374 );
or \U$31130 ( \31376 , \31361 , \31375 );
nand \U$31131 ( \31377 , \31373 , \31367 );
nand \U$31132 ( \31378 , \31376 , \31377 );
not \U$31133 ( \31379 , \31378 );
xor \U$31134 ( \31380 , RIbe2ad48_108, RIbe2a028_80);
not \U$31135 ( \31381 , \31380 );
not \U$31136 ( \31382 , \8168 );
or \U$31137 ( \31383 , \31381 , \31382 );
nand \U$31138 ( \31384 , \8172 , \31051 );
nand \U$31139 ( \31385 , \31383 , \31384 );
xor \U$31140 ( \31386 , RIbe2a910_99, RIbe2a0a0_81);
not \U$31141 ( \31387 , \31386 );
not \U$31142 ( \31388 , \9736 );
or \U$31143 ( \31389 , \31387 , \31388 );
nand \U$31144 ( \31390 , \10400 , \30982 );
nand \U$31145 ( \31391 , \31389 , \31390 );
xor \U$31146 ( \31392 , \31385 , \31391 );
xor \U$31147 ( \31393 , RIbe2b4c8_124, RIbe29e48_76);
not \U$31148 ( \31394 , \31393 );
not \U$31149 ( \31395 , \7716 );
or \U$31150 ( \31396 , \31394 , \31395 );
nand \U$31151 ( \31397 , \7368 , \31064 );
nand \U$31152 ( \31398 , \31396 , \31397 );
and \U$31153 ( \31399 , \31392 , \31398 );
and \U$31154 ( \31400 , \31385 , \31391 );
or \U$31155 ( \31401 , \31399 , \31400 );
xor \U$31156 ( \31402 , RIbe298a8_64, RIbe2b018_114);
not \U$31157 ( \31403 , \31402 );
not \U$31158 ( \31404 , \30723 );
or \U$31159 ( \31405 , \31403 , \31404 );
nand \U$31160 ( \31406 , \21442 , \30952 );
nand \U$31161 ( \31407 , \31405 , \31406 );
xor \U$31162 ( \31408 , RIbe29ec0_77, RIbe2b108_116);
not \U$31163 ( \31409 , \31408 );
not \U$31164 ( \31410 , \14296 );
or \U$31165 ( \31411 , \31409 , \31410 );
nand \U$31166 ( \31412 , \13533 , \31023 );
nand \U$31167 ( \31413 , \31411 , \31412 );
or \U$31168 ( \31414 , \31407 , \31413 );
xor \U$31169 ( \31415 , RIbe2a820_97, RIbe2a550_91);
not \U$31170 ( \31416 , \31415 );
not \U$31171 ( \31417 , \10433 );
or \U$31172 ( \31418 , \31416 , \31417 );
nand \U$31173 ( \31419 , \15995 , \30966 );
nand \U$31174 ( \31420 , \31418 , \31419 );
nand \U$31175 ( \31421 , \31414 , \31420 );
nand \U$31176 ( \31422 , \31413 , \31407 );
nand \U$31177 ( \31423 , \31421 , \31422 );
and \U$31178 ( \31424 , \31401 , \31423 );
not \U$31179 ( \31425 , \31401 );
not \U$31180 ( \31426 , \31423 );
and \U$31181 ( \31427 , \31425 , \31426 );
nor \U$31182 ( \31428 , \31424 , \31427 );
not \U$31183 ( \31429 , \31428 );
or \U$31184 ( \31430 , \31379 , \31429 );
not \U$31185 ( \31431 , \31426 );
nand \U$31186 ( \31432 , \31431 , \31401 );
nand \U$31187 ( \31433 , \31430 , \31432 );
not \U$31188 ( \31434 , \31433 );
or \U$31189 ( \31435 , \31353 , \31434 );
not \U$31190 ( \31436 , \31347 );
nand \U$31191 ( \31437 , \31436 , \31304 );
nand \U$31192 ( \31438 , \31435 , \31437 );
not \U$31193 ( \31439 , \31438 );
xor \U$31194 ( \31440 , \30980 , \31042 );
not \U$31195 ( \31441 , \31440 );
xor \U$31196 ( \31442 , \31086 , \31095 );
xor \U$31197 ( \31443 , \31442 , \31079 );
not \U$31198 ( \31444 , \31443 );
not \U$31199 ( \31445 , \31165 );
not \U$31200 ( \31446 , \31182 );
not \U$31201 ( \31447 , \31446 );
or \U$31202 ( \31448 , \31445 , \31447 );
not \U$31203 ( \31449 , \31165 );
nand \U$31204 ( \31450 , \31449 , \31182 );
nand \U$31205 ( \31451 , \31448 , \31450 );
not \U$31206 ( \31452 , \31451 );
not \U$31207 ( \31453 , \31007 );
not \U$31208 ( \31454 , \30987 );
not \U$31209 ( \31455 , \31454 );
and \U$31210 ( \31456 , \31453 , \31455 );
and \U$31211 ( \31457 , \31007 , \31454 );
nor \U$31212 ( \31458 , \31456 , \31457 );
not \U$31213 ( \31459 , \31458 );
or \U$31214 ( \31460 , \31452 , \31459 );
or \U$31215 ( \31461 , \31458 , \31451 );
nand \U$31216 ( \31462 , \31460 , \31461 );
not \U$31217 ( \31463 , \31462 );
or \U$31218 ( \31464 , \31444 , \31463 );
not \U$31219 ( \31465 , \31458 );
nand \U$31220 ( \31466 , \31465 , \31451 );
nand \U$31221 ( \31467 , \31464 , \31466 );
not \U$31222 ( \31468 , \31467 );
nand \U$31223 ( \31469 , \31441 , \31468 );
not \U$31224 ( \31470 , \31469 );
xor \U$31225 ( \31471 , \30976 , \30957 );
not \U$31226 ( \31472 , \31471 );
xor \U$31227 ( \31473 , \31019 , \31032 );
xor \U$31228 ( \31474 , RIbe2a2f8_86, RIbe2a460_89);
not \U$31229 ( \31475 , \31474 );
not \U$31230 ( \31476 , \8989 );
or \U$31231 ( \31477 , \31475 , \31476 );
nand \U$31232 ( \31478 , \8706 , \30996 );
nand \U$31233 ( \31479 , \31477 , \31478 );
not \U$31234 ( \31480 , \31479 );
xor \U$31235 ( \31481 , RIbe2a280_85, RIbe2b6a8_128);
not \U$31236 ( \31482 , \31481 );
not \U$31237 ( \31483 , \10845 );
or \U$31238 ( \31484 , \31482 , \31483 );
nand \U$31239 ( \31485 , \11348 , \31173 );
nand \U$31240 ( \31486 , \31484 , \31485 );
xor \U$31241 ( \31487 , RIbe28d68_40, RIbe2aaf0_103);
not \U$31242 ( \31488 , \31487 );
not \U$31243 ( \31489 , \18832 );
or \U$31244 ( \31490 , \31488 , \31489 );
nand \U$31245 ( \31491 , \30989 , RIbe2ab68_104);
nand \U$31246 ( \31492 , \31490 , \31491 );
xor \U$31247 ( \31493 , \31486 , \31492 );
not \U$31248 ( \31494 , \31493 );
or \U$31249 ( \31495 , \31480 , \31494 );
nand \U$31250 ( \31496 , \31486 , \31492 );
nand \U$31251 ( \31497 , \31495 , \31496 );
and \U$31252 ( \31498 , \31473 , \31497 );
not \U$31253 ( \31499 , \31473 );
not \U$31254 ( \31500 , \31497 );
and \U$31255 ( \31501 , \31499 , \31500 );
nor \U$31256 ( \31502 , \31498 , \31501 );
not \U$31257 ( \31503 , \31502 );
or \U$31258 ( \31504 , \31472 , \31503 );
nand \U$31259 ( \31505 , \31473 , \31497 );
nand \U$31260 ( \31506 , \31504 , \31505 );
not \U$31261 ( \31507 , \31506 );
or \U$31262 ( \31508 , \31470 , \31507 );
nand \U$31263 ( \31509 , \31440 , \31467 );
nand \U$31264 ( \31510 , \31508 , \31509 );
and \U$31265 ( \31511 , \31439 , \31510 );
not \U$31266 ( \31512 , \31439 );
not \U$31267 ( \31513 , \31510 );
and \U$31268 ( \31514 , \31512 , \31513 );
nor \U$31269 ( \31515 , \31511 , \31514 );
not \U$31270 ( \31516 , \31116 );
not \U$31271 ( \31517 , \31516 );
not \U$31272 ( \31518 , \31047 );
and \U$31273 ( \31519 , \31517 , \31518 );
and \U$31274 ( \31520 , \31516 , \31047 );
nor \U$31275 ( \31521 , \31519 , \31520 );
or \U$31276 ( \31522 , \31515 , \31521 );
or \U$31277 ( \31523 , \31513 , \31439 );
nand \U$31278 ( \31524 , \31522 , \31523 );
and \U$31279 ( \31525 , \31302 , \31524 );
and \U$31280 ( \31526 , \31236 , \31301 );
or \U$31281 ( \31527 , \31525 , \31526 );
not \U$31282 ( \31528 , \31527 );
xor \U$31283 ( \31529 , \30856 , \30884 );
xor \U$31284 ( \31530 , \31529 , \30831 );
xor \U$31285 ( \31531 , \30815 , \30810 );
xor \U$31286 ( \31532 , \31530 , \31531 );
not \U$31287 ( \31533 , \31244 );
not \U$31288 ( \31534 , \31533 );
not \U$31289 ( \31535 , \31267 );
or \U$31290 ( \31536 , \31534 , \31535 );
nand \U$31291 ( \31537 , \31262 , \31256 );
nand \U$31292 ( \31538 , \31536 , \31537 );
and \U$31293 ( \31539 , \31532 , \31538 );
and \U$31294 ( \31540 , \31530 , \31531 );
or \U$31295 ( \31541 , \31539 , \31540 );
not \U$31296 ( \31542 , \31541 );
and \U$31297 ( \31543 , \31528 , \31542 );
not \U$31298 ( \31544 , \31528 );
and \U$31299 ( \31545 , \31544 , \31541 );
nor \U$31300 ( \31546 , \31543 , \31545 );
buf \U$31301 ( \31547 , \31216 );
buf \U$31302 ( \31548 , \30942 );
and \U$31303 ( \31549 , \31547 , \31548 );
not \U$31304 ( \31550 , \31547 );
not \U$31305 ( \31551 , \30942 );
and \U$31306 ( \31552 , \31550 , \31551 );
nor \U$31307 ( \31553 , \31549 , \31552 );
not \U$31308 ( \31554 , \31553 );
and \U$31309 ( \31555 , \31546 , \31554 );
not \U$31310 ( \31556 , \31546 );
and \U$31311 ( \31557 , \31556 , \31553 );
nor \U$31312 ( \31558 , \31555 , \31557 );
xor \U$31313 ( \31559 , \31236 , \31301 );
xor \U$31314 ( \31560 , \31559 , \31524 );
not \U$31315 ( \31561 , \31560 );
not \U$31316 ( \31562 , \31561 );
xor \U$31317 ( \31563 , \31530 , \31531 );
xor \U$31318 ( \31564 , \31563 , \31538 );
not \U$31319 ( \31565 , \31564 );
not \U$31320 ( \31566 , \31277 );
not \U$31321 ( \31567 , \31566 );
not \U$31322 ( \31568 , \31287 );
or \U$31323 ( \31569 , \31567 , \31568 );
or \U$31324 ( \31570 , \31287 , \31566 );
nand \U$31325 ( \31571 , \31569 , \31570 );
not \U$31326 ( \31572 , \31571 );
not \U$31327 ( \31573 , \31341 );
not \U$31328 ( \31574 , \31337 );
nand \U$31329 ( \31575 , \31574 , \31343 );
not \U$31330 ( \31576 , \31575 );
or \U$31331 ( \31577 , \31573 , \31576 );
or \U$31332 ( \31578 , \31575 , \31341 );
nand \U$31333 ( \31579 , \31577 , \31578 );
xor \U$31334 ( \31580 , \31407 , \31413 );
not \U$31335 ( \31581 , \31420 );
and \U$31336 ( \31582 , \31580 , \31581 );
not \U$31337 ( \31583 , \31580 );
and \U$31338 ( \31584 , \31583 , \31420 );
nor \U$31339 ( \31585 , \31582 , \31584 );
and \U$31340 ( \31586 , \31579 , \31585 );
xor \U$31341 ( \31587 , \31367 , \31373 );
xnor \U$31342 ( \31588 , \31587 , \31360 );
or \U$31343 ( \31589 , \31586 , \31588 );
or \U$31344 ( \31590 , \31585 , \31579 );
nand \U$31345 ( \31591 , \31589 , \31590 );
not \U$31346 ( \31592 , \31591 );
not \U$31347 ( \31593 , \31592 );
xnor \U$31348 ( \31594 , \31462 , \31443 );
not \U$31349 ( \31595 , \31594 );
or \U$31350 ( \31596 , \31593 , \31595 );
not \U$31351 ( \31597 , \31471 );
not \U$31352 ( \31598 , \31597 );
buf \U$31353 ( \31599 , \31502 );
not \U$31354 ( \31600 , \31599 );
or \U$31355 ( \31601 , \31598 , \31600 );
or \U$31356 ( \31602 , \31599 , \31597 );
nand \U$31357 ( \31603 , \31601 , \31602 );
nand \U$31358 ( \31604 , \31596 , \31603 );
not \U$31359 ( \31605 , \31594 );
nand \U$31360 ( \31606 , \31605 , \31591 );
nand \U$31361 ( \31607 , \31604 , \31606 );
not \U$31362 ( \31608 , \31607 );
xor \U$31363 ( \31609 , \31506 , \31440 );
not \U$31364 ( \31610 , \31609 );
not \U$31365 ( \31611 , \31468 );
and \U$31366 ( \31612 , \31610 , \31611 );
and \U$31367 ( \31613 , \31609 , \31468 );
nor \U$31368 ( \31614 , \31612 , \31613 );
not \U$31369 ( \31615 , \31614 );
or \U$31370 ( \31616 , \31608 , \31615 );
or \U$31371 ( \31617 , \31614 , \31607 );
nand \U$31372 ( \31618 , \31616 , \31617 );
not \U$31373 ( \31619 , \31618 );
or \U$31374 ( \31620 , \31572 , \31619 );
not \U$31375 ( \31621 , \31614 );
nand \U$31376 ( \31622 , \31621 , \31607 );
nand \U$31377 ( \31623 , \31620 , \31622 );
not \U$31378 ( \31624 , \31623 );
not \U$31379 ( \31625 , \31378 );
and \U$31380 ( \31626 , \31428 , \31625 );
not \U$31381 ( \31627 , \31428 );
and \U$31382 ( \31628 , \31627 , \31378 );
nor \U$31383 ( \31629 , \31626 , \31628 );
not \U$31384 ( \31630 , \31629 );
not \U$31385 ( \31631 , \31630 );
nand \U$31386 ( \31632 , \8270 , RIbe2ae38_110);
not \U$31387 ( \31633 , \31632 );
not \U$31388 ( \31634 , \31633 );
not \U$31389 ( \31635 , \2717 );
xor \U$31390 ( \31636 , RIbe27fd0_11, RIbe2b450_123);
not \U$31391 ( \31637 , \31636 );
not \U$31392 ( \31638 , \31637 );
and \U$31393 ( \31639 , \31635 , \31638 );
and \U$31394 ( \31640 , \7709 , \31362 );
nor \U$31395 ( \31641 , \31639 , \31640 );
not \U$31396 ( \31642 , \31641 );
not \U$31397 ( \31643 , \31642 );
or \U$31398 ( \31644 , \31634 , \31643 );
not \U$31399 ( \31645 , \31641 );
not \U$31400 ( \31646 , \31632 );
or \U$31401 ( \31647 , \31645 , \31646 );
and \U$31402 ( \31648 , RIbe29d58_74, RIbe2b180_117);
nor \U$31403 ( \31649 , RIbe29d58_74, RIbe2b180_117);
nor \U$31404 ( \31650 , \31648 , \31649 );
not \U$31405 ( \31651 , \31650 );
not \U$31406 ( \31652 , \14852 );
or \U$31407 ( \31653 , \31651 , \31652 );
xor \U$31408 ( \31654 , RIbe2b180_117, RIbe29ce0_73);
nand \U$31409 ( \31655 , \14845 , \31654 );
nand \U$31410 ( \31656 , \31653 , \31655 );
nand \U$31411 ( \31657 , \31647 , \31656 );
nand \U$31412 ( \31658 , \31644 , \31657 );
not \U$31413 ( \31659 , \31658 );
xor \U$31414 ( \31660 , RIbe29998_66, RIbe2aaf0_103);
not \U$31415 ( \31661 , \31660 );
not \U$31416 ( \31662 , \28282 );
or \U$31417 ( \31663 , \31661 , \31662 );
nand \U$31418 ( \31664 , \31487 , RIbe2ab68_104);
nand \U$31419 ( \31665 , \31663 , \31664 );
not \U$31420 ( \31666 , \31665 );
xor \U$31421 ( \31667 , RIbe2b108_116, RIbe29f38_78);
not \U$31422 ( \31668 , \31667 );
not \U$31423 ( \31669 , \25617 );
or \U$31424 ( \31670 , \31668 , \31669 );
nand \U$31425 ( \31671 , \16898 , \31408 );
nand \U$31426 ( \31672 , \31670 , \31671 );
not \U$31427 ( \31673 , \31672 );
or \U$31428 ( \31674 , \31666 , \31673 );
or \U$31429 ( \31675 , \31672 , \31665 );
xor \U$31430 ( \31676 , RIbe28f48_44, RIbe2a7a8_96);
not \U$31431 ( \31677 , \31676 );
not \U$31432 ( \31678 , \8221 );
or \U$31433 ( \31679 , \31677 , \31678 );
xor \U$31434 ( \31680 , RIbe2abe0_105, RIbe28f48_44);
nand \U$31435 ( \31681 , \3249 , \31680 );
nand \U$31436 ( \31682 , \31679 , \31681 );
nand \U$31437 ( \31683 , \31675 , \31682 );
nand \U$31438 ( \31684 , \31674 , \31683 );
not \U$31439 ( \31685 , \31684 );
or \U$31440 ( \31686 , \31659 , \31685 );
or \U$31441 ( \31687 , \31684 , \31658 );
xor \U$31442 ( \31688 , RIbe2b360_121, RIbe2a910_99);
not \U$31443 ( \31689 , \31688 );
not \U$31444 ( \31690 , \9738 );
or \U$31445 ( \31691 , \31689 , \31690 );
nand \U$31446 ( \31692 , \9726 , \31386 );
nand \U$31447 ( \31693 , \31691 , \31692 );
not \U$31448 ( \31694 , \31693 );
xor \U$31449 ( \31695 , RIbe2a3e8_88, RIbe2a4d8_90);
not \U$31450 ( \31696 , \31695 );
not \U$31451 ( \31697 , \8806 );
or \U$31452 ( \31698 , \31696 , \31697 );
nand \U$31453 ( \31699 , \8794 , \31331 );
nand \U$31454 ( \31700 , \31698 , \31699 );
not \U$31455 ( \31701 , \31700 );
not \U$31456 ( \31702 , \31701 );
xor \U$31457 ( \31703 , RIbe2a028_80, RIbe2b540_125);
not \U$31458 ( \31704 , \31703 );
not \U$31459 ( \31705 , \8400 );
or \U$31460 ( \31706 , \31704 , \31705 );
nand \U$31461 ( \31707 , \8172 , \31380 );
nand \U$31462 ( \31708 , \31706 , \31707 );
not \U$31463 ( \31709 , \31708 );
or \U$31464 ( \31710 , \31702 , \31709 );
or \U$31465 ( \31711 , \31708 , \31701 );
nand \U$31466 ( \31712 , \31710 , \31711 );
not \U$31467 ( \31713 , \31712 );
or \U$31468 ( \31714 , \31694 , \31713 );
nand \U$31469 ( \31715 , \31708 , \31700 );
nand \U$31470 ( \31716 , \31714 , \31715 );
nand \U$31471 ( \31717 , \31687 , \31716 );
nand \U$31472 ( \31718 , \31686 , \31717 );
not \U$31473 ( \31719 , \31718 );
xor \U$31474 ( \31720 , RIbe2a898_98, RIbe2a190_83);
not \U$31475 ( \31721 , \31720 );
not \U$31476 ( \31722 , \10831 );
or \U$31477 ( \31723 , \31721 , \31722 );
nand \U$31478 ( \31724 , \10834 , \31354 );
nand \U$31479 ( \31725 , \31723 , \31724 );
not \U$31480 ( \31726 , \31725 );
xor \U$31481 ( \31727 , RIbe28cf0_39, RIbe2b018_114);
not \U$31482 ( \31728 , \31727 );
not \U$31483 ( \31729 , \30723 );
or \U$31484 ( \31730 , \31728 , \31729 );
nand \U$31485 ( \31731 , \15952 , \31402 );
nand \U$31486 ( \31732 , \31730 , \31731 );
not \U$31487 ( \31733 , \31732 );
or \U$31488 ( \31734 , \31726 , \31733 );
or \U$31489 ( \31735 , \31725 , \31732 );
xor \U$31490 ( \31736 , RIbe2af28_112, RIbe29b78_70);
not \U$31491 ( \31737 , \31736 );
not \U$31492 ( \31738 , \16913 );
or \U$31493 ( \31739 , \31737 , \31738 );
nand \U$31494 ( \31740 , \17810 , \31338 );
nand \U$31495 ( \31741 , \31739 , \31740 );
nand \U$31496 ( \31742 , \31735 , \31741 );
nand \U$31497 ( \31743 , \31734 , \31742 );
not \U$31498 ( \31744 , \31743 );
xor \U$31499 ( \31745 , RIbe2aa78_102, RIbe2a280_85);
not \U$31500 ( \31746 , \31745 );
not \U$31501 ( \31747 , \23353 );
or \U$31502 ( \31748 , \31746 , \31747 );
nand \U$31503 ( \31749 , \18667 , \31481 );
nand \U$31504 ( \31750 , \31748 , \31749 );
xor \U$31505 ( \31751 , RIbe2a118_82, RIbe2a550_91);
not \U$31506 ( \31752 , \31751 );
not \U$31507 ( \31753 , \10433 );
or \U$31508 ( \31754 , \31752 , \31753 );
nand \U$31509 ( \31755 , \11484 , \31415 );
nand \U$31510 ( \31756 , \31754 , \31755 );
nand \U$31511 ( \31757 , \31750 , \31756 );
not \U$31512 ( \31758 , \31757 );
xor \U$31513 ( \31759 , RIbe2a6b8_94, RIbe29e48_76);
not \U$31514 ( \31760 , \31759 );
not \U$31515 ( \31761 , \11039 );
or \U$31516 ( \31762 , \31760 , \31761 );
nand \U$31517 ( \31763 , \8245 , \31393 );
nand \U$31518 ( \31764 , \31762 , \31763 );
not \U$31519 ( \31765 , \31764 );
nor \U$31520 ( \31766 , \31750 , \31756 );
nor \U$31521 ( \31767 , \31765 , \31766 );
nor \U$31522 ( \31768 , \31758 , \31767 );
nand \U$31523 ( \31769 , \31744 , \31768 );
not \U$31524 ( \31770 , \31769 );
xor \U$31525 ( \31771 , RIbe2ac58_106, RIbe29c68_72);
not \U$31526 ( \31772 , \31771 );
not \U$31527 ( \31773 , \8259 );
or \U$31528 ( \31774 , \31772 , \31773 );
nand \U$31529 ( \31775 , \4580 , \31368 );
nand \U$31530 ( \31776 , \31774 , \31775 );
not \U$31531 ( \31777 , \31776 );
xor \U$31532 ( \31778 , RIbe2aeb0_111, RIbe27e68_8);
not \U$31533 ( \31779 , \31778 );
not \U$31534 ( \31780 , \2458 );
or \U$31535 ( \31781 , \31779 , \31780 );
nand \U$31536 ( \31782 , \2463 , \31312 );
nand \U$31537 ( \31783 , \31781 , \31782 );
xor \U$31538 ( \31784 , RIbe2a2f8_86, RIbe2adc0_109);
not \U$31539 ( \31785 , \31784 );
not \U$31540 ( \31786 , \8697 );
or \U$31541 ( \31787 , \31785 , \31786 );
nand \U$31542 ( \31788 , \11094 , \31474 );
nand \U$31543 ( \31789 , \31787 , \31788 );
and \U$31544 ( \31790 , \31783 , \31789 );
not \U$31545 ( \31791 , \31783 );
not \U$31546 ( \31792 , \31789 );
and \U$31547 ( \31793 , \31791 , \31792 );
nor \U$31548 ( \31794 , \31790 , \31793 );
not \U$31549 ( \31795 , \31794 );
or \U$31550 ( \31796 , \31777 , \31795 );
not \U$31551 ( \31797 , \31792 );
nand \U$31552 ( \31798 , \31797 , \31783 );
nand \U$31553 ( \31799 , \31796 , \31798 );
not \U$31554 ( \31800 , \31799 );
or \U$31555 ( \31801 , \31770 , \31800 );
not \U$31556 ( \31802 , \31768 );
nand \U$31557 ( \31803 , \31802 , \31743 );
nand \U$31558 ( \31804 , \31801 , \31803 );
not \U$31559 ( \31805 , \31804 );
not \U$31560 ( \31806 , \31805 );
or \U$31561 ( \31807 , \31719 , \31806 );
or \U$31562 ( \31808 , \31805 , \31718 );
nand \U$31563 ( \31809 , \31807 , \31808 );
not \U$31564 ( \31810 , \31809 );
or \U$31565 ( \31811 , \31631 , \31810 );
not \U$31566 ( \31812 , \31805 );
nand \U$31567 ( \31813 , \31812 , \31718 );
nand \U$31568 ( \31814 , \31811 , \31813 );
not \U$31569 ( \31815 , \31814 );
xnor \U$31570 ( \31816 , \31324 , \31344 );
not \U$31571 ( \31817 , \31816 );
not \U$31572 ( \31818 , \31817 );
not \U$31573 ( \31819 , \31680 );
not \U$31574 ( \31820 , \12721 );
or \U$31575 ( \31821 , \31819 , \31820 );
nand \U$31576 ( \31822 , \9524 , \31090 );
nand \U$31577 ( \31823 , \31821 , \31822 );
not \U$31578 ( \31824 , \31654 );
not \U$31579 ( \31825 , \15353 );
or \U$31580 ( \31826 , \31824 , \31825 );
nand \U$31581 ( \31827 , \16646 , \31306 );
nand \U$31582 ( \31828 , \31826 , \31827 );
nor \U$31583 ( \31829 , \31823 , \31828 );
and \U$31584 ( \31830 , \31317 , \31322 );
not \U$31585 ( \31831 , \31317 );
and \U$31586 ( \31832 , \31831 , \31321 );
or \U$31587 ( \31833 , \31830 , \31832 );
or \U$31588 ( \31834 , \31829 , \31833 );
nand \U$31589 ( \31835 , \31828 , \31823 );
nand \U$31590 ( \31836 , \31834 , \31835 );
not \U$31591 ( \31837 , \31836 );
not \U$31592 ( \31838 , \31069 );
not \U$31593 ( \31839 , \31062 );
not \U$31594 ( \31840 , \31839 );
or \U$31595 ( \31841 , \31838 , \31840 );
or \U$31596 ( \31842 , \31069 , \31839 );
nand \U$31597 ( \31843 , \31841 , \31842 );
not \U$31598 ( \31844 , \31056 );
and \U$31599 ( \31845 , \31843 , \31844 );
not \U$31600 ( \31846 , \31843 );
and \U$31601 ( \31847 , \31846 , \31056 );
nor \U$31602 ( \31848 , \31845 , \31847 );
not \U$31603 ( \31849 , \31848 );
or \U$31604 ( \31850 , \31837 , \31849 );
or \U$31605 ( \31851 , \31836 , \31848 );
nand \U$31606 ( \31852 , \31850 , \31851 );
not \U$31607 ( \31853 , \31852 );
or \U$31608 ( \31854 , \31818 , \31853 );
not \U$31609 ( \31855 , \31848 );
nand \U$31610 ( \31856 , \31855 , \31836 );
nand \U$31611 ( \31857 , \31854 , \31856 );
not \U$31612 ( \31858 , \31351 );
not \U$31613 ( \31859 , \31433 );
or \U$31614 ( \31860 , \31858 , \31859 );
or \U$31615 ( \31861 , \31433 , \31351 );
nand \U$31616 ( \31862 , \31860 , \31861 );
xor \U$31617 ( \31863 , \31857 , \31862 );
not \U$31618 ( \31864 , \31863 );
or \U$31619 ( \31865 , \31815 , \31864 );
nand \U$31620 ( \31866 , \31862 , \31857 );
nand \U$31621 ( \31867 , \31865 , \31866 );
not \U$31622 ( \31868 , \31867 );
xor \U$31623 ( \31869 , \31438 , \31521 );
xor \U$31624 ( \31870 , \31869 , \31513 );
not \U$31625 ( \31871 , \31870 );
not \U$31626 ( \31872 , \31871 );
or \U$31627 ( \31873 , \31868 , \31872 );
not \U$31628 ( \31874 , \31867 );
nand \U$31629 ( \31875 , \31874 , \31870 );
nand \U$31630 ( \31876 , \31873 , \31875 );
not \U$31631 ( \31877 , \31876 );
or \U$31632 ( \31878 , \31624 , \31877 );
nand \U$31633 ( \31879 , \31870 , \31867 );
nand \U$31634 ( \31880 , \31878 , \31879 );
not \U$31635 ( \31881 , \31880 );
not \U$31636 ( \31882 , \31881 );
or \U$31637 ( \31883 , \31565 , \31882 );
or \U$31638 ( \31884 , \31881 , \31564 );
nand \U$31639 ( \31885 , \31883 , \31884 );
not \U$31640 ( \31886 , \31885 );
or \U$31641 ( \31887 , \31562 , \31886 );
not \U$31642 ( \31888 , \31564 );
nand \U$31643 ( \31889 , \31888 , \31881 );
nand \U$31644 ( \31890 , \31887 , \31889 );
nand \U$31645 ( \31891 , \31558 , \31890 );
xor \U$31646 ( \31892 , \30936 , \31222 );
xor \U$31647 ( \31893 , \31892 , \31228 );
not \U$31648 ( \31894 , \31542 );
not \U$31649 ( \31895 , \31528 );
or \U$31650 ( \31896 , \31894 , \31895 );
nand \U$31651 ( \31897 , \31896 , \31553 );
nand \U$31652 ( \31898 , \31527 , \31541 );
nand \U$31653 ( \31899 , \31897 , \31898 );
not \U$31654 ( \31900 , \31899 );
nand \U$31655 ( \31901 , \31893 , \31900 );
and \U$31656 ( \31902 , \30926 , \31232 , \31891 , \31901 );
not \U$31657 ( \31903 , \31902 );
xor \U$31658 ( \31904 , \31725 , \31732 );
xor \U$31659 ( \31905 , \31741 , \31904 );
and \U$31660 ( \31906 , \31712 , \31693 );
not \U$31661 ( \31907 , \31712 );
not \U$31662 ( \31908 , \31693 );
and \U$31663 ( \31909 , \31907 , \31908 );
nor \U$31664 ( \31910 , \31906 , \31909 );
xor \U$31665 ( \31911 , \31905 , \31910 );
xor \U$31666 ( \31912 , \31776 , \31794 );
xor \U$31667 ( \31913 , \31911 , \31912 );
xor \U$31668 ( \31914 , \31665 , \31672 );
xnor \U$31669 ( \31915 , \31914 , \31682 );
not \U$31670 ( \31916 , \31915 );
not \U$31671 ( \31917 , \31916 );
not \U$31672 ( \31918 , \31766 );
nand \U$31673 ( \31919 , \31918 , \31757 );
buf \U$31674 ( \31920 , \31764 );
and \U$31675 ( \31921 , \31919 , \31920 );
not \U$31676 ( \31922 , \31919 );
not \U$31677 ( \31923 , \31920 );
and \U$31678 ( \31924 , \31922 , \31923 );
nor \U$31679 ( \31925 , \31921 , \31924 );
not \U$31680 ( \31926 , \31925 );
not \U$31681 ( \31927 , \31926 );
or \U$31682 ( \31928 , \31917 , \31927 );
nand \U$31683 ( \31929 , \31925 , \31915 );
nand \U$31684 ( \31930 , \31928 , \31929 );
xor \U$31685 ( \31931 , \31633 , \31642 );
xnor \U$31686 ( \31932 , \31931 , \31656 );
not \U$31687 ( \31933 , \31932 );
and \U$31688 ( \31934 , \31930 , \31933 );
not \U$31689 ( \31935 , \31930 );
and \U$31690 ( \31936 , \31935 , \31932 );
nor \U$31691 ( \31937 , \31934 , \31936 );
and \U$31692 ( \31938 , \31913 , \31937 );
not \U$31693 ( \31939 , \31913 );
not \U$31694 ( \31940 , \31937 );
and \U$31695 ( \31941 , \31939 , \31940 );
or \U$31696 ( \31942 , \31938 , \31941 );
buf \U$31697 ( \31943 , \10690 );
not \U$31698 ( \31944 , \31943 );
xor \U$31699 ( \31945 , RIbe2a820_97, RIbe2a190_83);
not \U$31700 ( \31946 , \31945 );
or \U$31701 ( \31947 , \31944 , \31946 );
buf \U$31702 ( \31948 , \10696 );
nand \U$31703 ( \31949 , \31948 , \31720 );
nand \U$31704 ( \31950 , \31947 , \31949 );
not \U$31705 ( \31951 , \2451 );
nand \U$31706 ( \31952 , \31951 , RIbe2ae38_110);
nand \U$31707 ( \31953 , RIbe27f58_10, RIbe27fd0_11);
and \U$31708 ( \31954 , \31952 , \31953 , RIbe27e68_8);
xor \U$31709 ( \31955 , RIbe27fd0_11, RIbe2b3d8_122);
not \U$31710 ( \31956 , \31955 );
not \U$31711 ( \31957 , \3377 );
or \U$31712 ( \31958 , \31956 , \31957 );
nand \U$31713 ( \31959 , \2707 , \31636 );
nand \U$31714 ( \31960 , \31958 , \31959 );
xor \U$31715 ( \31961 , \31954 , \31960 );
xor \U$31716 ( \31962 , \31950 , \31961 );
xor \U$31717 ( \31963 , RIbe2a190_83, RIbe2a118_82);
not \U$31718 ( \31964 , \31963 );
not \U$31719 ( \31965 , \25032 );
or \U$31720 ( \31966 , \31964 , \31965 );
nand \U$31721 ( \31967 , \15693 , \31945 );
nand \U$31722 ( \31968 , \31966 , \31967 );
xor \U$31723 ( \31969 , RIbe2b360_121, RIbe2a550_91);
not \U$31724 ( \31970 , \31969 );
not \U$31725 ( \31971 , \19607 );
or \U$31726 ( \31972 , \31970 , \31971 );
not \U$31727 ( \31973 , RIbe2a0a0_81);
not \U$31728 ( \31974 , RIbe2a550_91);
and \U$31729 ( \31975 , \31973 , \31974 );
and \U$31730 ( \31976 , RIbe2a0a0_81, RIbe2a550_91);
nor \U$31731 ( \31977 , \31975 , \31976 );
nand \U$31732 ( \31978 , \11228 , \31977 );
nand \U$31733 ( \31979 , \31972 , \31978 );
xor \U$31734 ( \31980 , \31968 , \31979 );
and \U$31735 ( \31981 , RIbe29e48_76, RIbe2ac58_106);
nor \U$31736 ( \31982 , RIbe29e48_76, RIbe2ac58_106);
nor \U$31737 ( \31983 , \31981 , \31982 );
not \U$31738 ( \31984 , \31983 );
not \U$31739 ( \31985 , \7372 );
or \U$31740 ( \31986 , \31984 , \31985 );
xor \U$31741 ( \31987 , RIbe29e48_76, RIbe2a640_93);
nand \U$31742 ( \31988 , \7368 , \31987 );
nand \U$31743 ( \31989 , \31986 , \31988 );
and \U$31744 ( \31990 , \31980 , \31989 );
and \U$31745 ( \31991 , \31968 , \31979 );
or \U$31746 ( \31992 , \31990 , \31991 );
xor \U$31747 ( \31993 , \31962 , \31992 );
not \U$31748 ( \31994 , \31993 );
xor \U$31749 ( \31995 , RIbe28f48_44, RIbe2b3d8_122);
not \U$31750 ( \31996 , \31995 );
not \U$31751 ( \31997 , \11461 );
or \U$31752 ( \31998 , \31996 , \31997 );
xor \U$31753 ( \31999 , RIbe28f48_44, RIbe2b450_123);
nand \U$31754 ( \32000 , \3249 , \31999 );
nand \U$31755 ( \32001 , \31998 , \32000 );
or \U$31756 ( \32002 , RIbe28ed0_43, RIbe28f48_44);
nand \U$31757 ( \32003 , \32002 , RIbe2ae38_110);
nand \U$31758 ( \32004 , RIbe28ed0_43, RIbe28f48_44);
and \U$31759 ( \32005 , \32003 , \32004 , RIbe27fd0_11);
nand \U$31760 ( \32006 , \32001 , \32005 );
not \U$31761 ( \32007 , \32006 );
not \U$31762 ( \32008 , \32007 );
xor \U$31763 ( \32009 , RIbe2a6b8_94, RIbe2a028_80);
not \U$31764 ( \32010 , \32009 );
not \U$31765 ( \32011 , \22849 );
or \U$31766 ( \32012 , \32010 , \32011 );
xor \U$31767 ( \32013 , RIbe2a028_80, RIbe2b4c8_124);
nand \U$31768 ( \32014 , \8172 , \32013 );
nand \U$31769 ( \32015 , \32012 , \32014 );
not \U$31770 ( \32016 , \32015 );
xor \U$31771 ( \32017 , RIbe2a898_98, RIbe2a280_85);
and \U$31772 ( \32018 , \20237 , \32017 );
xor \U$31773 ( \32019 , RIbe2aa00_101, RIbe2a280_85);
and \U$31774 ( \32020 , \10849 , \32019 );
nor \U$31775 ( \32021 , \32018 , \32020 );
not \U$31776 ( \32022 , \32021 );
or \U$31777 ( \32023 , \32016 , \32022 );
or \U$31778 ( \32024 , \32015 , \32021 );
nand \U$31779 ( \32025 , \32023 , \32024 );
not \U$31780 ( \32026 , \32025 );
or \U$31781 ( \32027 , \32008 , \32026 );
not \U$31782 ( \32028 , \32021 );
nand \U$31783 ( \32029 , \32028 , \32015 );
nand \U$31784 ( \32030 , \32027 , \32029 );
not \U$31785 ( \32031 , \32030 );
not \U$31786 ( \32032 , \32031 );
xor \U$31787 ( \32033 , RIbe2a460_89, RIbe2a910_99);
not \U$31788 ( \32034 , \32033 );
not \U$31789 ( \32035 , \9737 );
or \U$31790 ( \32036 , \32034 , \32035 );
xor \U$31791 ( \32037 , RIbe2a4d8_90, RIbe2a910_99);
nand \U$31792 ( \32038 , \9726 , \32037 );
nand \U$31793 ( \32039 , \32036 , \32038 );
not \U$31794 ( \32040 , \32039 );
xor \U$31795 ( \32041 , RIbe29ce0_73, RIbe2b018_114);
not \U$31796 ( \32042 , \32041 );
not \U$31797 ( \32043 , \30723 );
or \U$31798 ( \32044 , \32042 , \32043 );
xor \U$31799 ( \32045 , RIbe29b78_70, RIbe2b018_114);
nand \U$31800 ( \32046 , \18777 , \32045 );
nand \U$31801 ( \32047 , \32044 , \32046 );
not \U$31802 ( \32048 , \32047 );
nand \U$31803 ( \32049 , \32040 , \32048 );
xor \U$31804 ( \32050 , RIbe2b6a8_128, RIbe2b180_117);
not \U$31805 ( \32051 , \32050 );
not \U$31806 ( \32052 , \15353 );
or \U$31807 ( \32053 , \32051 , \32052 );
xor \U$31808 ( \32054 , RIbe29f38_78, RIbe2b180_117);
nand \U$31809 ( \32055 , \21759 , \32054 );
nand \U$31810 ( \32056 , \32053 , \32055 );
and \U$31811 ( \32057 , \32049 , \32056 );
nor \U$31812 ( \32058 , \32040 , \32048 );
nor \U$31813 ( \32059 , \32057 , \32058 );
not \U$31814 ( \32060 , \32059 );
not \U$31815 ( \32061 , \32060 );
xor \U$31816 ( \32062 , RIbe2a640_93, RIbe2a028_80);
not \U$31817 ( \32063 , \32062 );
not \U$31818 ( \32064 , \8400 );
or \U$31819 ( \32065 , \32063 , \32064 );
nand \U$31820 ( \32066 , \8172 , \32009 );
nand \U$31821 ( \32067 , \32065 , \32066 );
xor \U$31822 ( \32068 , RIbe2a820_97, RIbe2a280_85);
not \U$31823 ( \32069 , \32068 );
not \U$31824 ( \32070 , \27992 );
or \U$31825 ( \32071 , \32069 , \32070 );
nand \U$31826 ( \32072 , \18667 , \32017 );
nand \U$31827 ( \32073 , \32071 , \32072 );
nor \U$31828 ( \32074 , \32067 , \32073 );
not \U$31829 ( \32075 , \32074 );
xor \U$31830 ( \32076 , RIbe2a550_91, RIbe2b2e8_120);
not \U$31831 ( \32077 , \32076 );
not \U$31832 ( \32078 , \18635 );
or \U$31833 ( \32079 , \32077 , \32078 );
not \U$31834 ( \32080 , \23307 );
nand \U$31835 ( \32081 , \32080 , \31969 );
nand \U$31836 ( \32082 , \32079 , \32081 );
and \U$31837 ( \32083 , \32075 , \32082 );
nand \U$31838 ( \32084 , \32067 , \32073 );
not \U$31839 ( \32085 , \32084 );
nor \U$31840 ( \32086 , \32083 , \32085 );
not \U$31841 ( \32087 , \32086 );
not \U$31842 ( \32088 , \32087 );
or \U$31843 ( \32089 , \32061 , \32088 );
not \U$31844 ( \32090 , \32059 );
not \U$31845 ( \32091 , \32086 );
or \U$31846 ( \32092 , \32090 , \32091 );
xor \U$31847 ( \32093 , RIbe2b108_116, RIbe2aa00_101);
not \U$31848 ( \32094 , \32093 );
not \U$31849 ( \32095 , \14297 );
or \U$31850 ( \32096 , \32094 , \32095 );
not \U$31851 ( \32097 , RIbe2aa78_102);
not \U$31852 ( \32098 , RIbe2b108_116);
and \U$31853 ( \32099 , \32097 , \32098 );
and \U$31854 ( \32100 , RIbe2aa78_102, RIbe2b108_116);
nor \U$31855 ( \32101 , \32099 , \32100 );
nand \U$31856 ( \32102 , \16875 , \32101 );
nand \U$31857 ( \32103 , \32096 , \32102 );
not \U$31858 ( \32104 , \32103 );
xor \U$31859 ( \32105 , RIbe29c68_72, RIbe2a730_95);
not \U$31860 ( \32106 , \32105 );
not \U$31861 ( \32107 , \8594 );
or \U$31862 ( \32108 , \32106 , \32107 );
xor \U$31863 ( \32109 , RIbe29c68_72, RIbe2a7a8_96);
nand \U$31864 ( \32110 , \4580 , \32109 );
nand \U$31865 ( \32111 , \32108 , \32110 );
xor \U$31866 ( \32112 , RIbe27b20_1, RIbe2aaf0_103);
not \U$31867 ( \32113 , \32112 );
not \U$31868 ( \32114 , \28282 );
or \U$31869 ( \32115 , \32113 , \32114 );
xor \U$31870 ( \32116 , RIbe28cf0_39, RIbe2aaf0_103);
nand \U$31871 ( \32117 , \32116 , RIbe2ab68_104);
nand \U$31872 ( \32118 , \32115 , \32117 );
xor \U$31873 ( \32119 , \32111 , \32118 );
not \U$31874 ( \32120 , \32119 );
or \U$31875 ( \32121 , \32104 , \32120 );
nand \U$31876 ( \32122 , \32111 , \32118 );
nand \U$31877 ( \32123 , \32121 , \32122 );
nand \U$31878 ( \32124 , \32092 , \32123 );
nand \U$31879 ( \32125 , \32089 , \32124 );
not \U$31880 ( \32126 , \32125 );
or \U$31881 ( \32127 , \32032 , \32126 );
or \U$31882 ( \32128 , \32125 , \32031 );
nand \U$31883 ( \32129 , \32127 , \32128 );
not \U$31884 ( \32130 , \32129 );
or \U$31885 ( \32131 , \31994 , \32130 );
not \U$31886 ( \32132 , \32031 );
nand \U$31887 ( \32133 , \32132 , \32125 );
nand \U$31888 ( \32134 , \32131 , \32133 );
xor \U$31889 ( \32135 , \31942 , \32134 );
not \U$31890 ( \32136 , \32135 );
xor \U$31891 ( \32137 , RIbe27b20_1, RIbe2b018_114);
not \U$31892 ( \32138 , \32137 );
not \U$31893 ( \32139 , \15967 );
or \U$31894 ( \32140 , \32138 , \32139 );
nand \U$31895 ( \32141 , \15953 , \31727 );
nand \U$31896 ( \32142 , \32140 , \32141 );
not \U$31897 ( \32143 , RIbe29ce0_73);
not \U$31898 ( \32144 , RIbe2af28_112);
and \U$31899 ( \32145 , \32143 , \32144 );
and \U$31900 ( \32146 , RIbe29ce0_73, RIbe2af28_112);
nor \U$31901 ( \32147 , \32145 , \32146 );
and \U$31902 ( \32148 , \16913 , \32147 );
and \U$31903 ( \32149 , \16917 , \31736 );
nor \U$31904 ( \32150 , \32148 , \32149 );
not \U$31905 ( \32151 , \32150 );
xor \U$31906 ( \32152 , \32142 , \32151 );
xor \U$31907 ( \32153 , RIbe29c68_72, RIbe2abe0_105);
not \U$31908 ( \32154 , \32153 );
not \U$31909 ( \32155 , \8595 );
or \U$31910 ( \32156 , \32154 , \32155 );
nand \U$31911 ( \32157 , \7642 , \31771 );
nand \U$31912 ( \32158 , \32156 , \32157 );
xor \U$31913 ( \32159 , \32152 , \32158 );
xor \U$31914 ( \32160 , RIbe2aeb0_111, RIbe27fd0_11);
not \U$31915 ( \32161 , \32160 );
not \U$31916 ( \32162 , \11366 );
or \U$31917 ( \32163 , \32161 , \32162 );
nand \U$31918 ( \32164 , \2707 , \31955 );
nand \U$31919 ( \32165 , \32163 , \32164 );
not \U$31920 ( \32166 , \32165 );
xor \U$31921 ( \32167 , RIbe2b540_125, RIbe2a2f8_86);
not \U$31922 ( \32168 , \32167 );
not \U$31923 ( \32169 , \16714 );
or \U$31924 ( \32170 , \32168 , \32169 );
xor \U$31925 ( \32171 , RIbe2ad48_108, RIbe2a2f8_86);
nand \U$31926 ( \32172 , \8705 , \32171 );
nand \U$31927 ( \32173 , \32170 , \32172 );
xor \U$31928 ( \32174 , RIbe2a3e8_88, RIbe2adc0_109);
not \U$31929 ( \32175 , \32174 );
not \U$31930 ( \32176 , \8806 );
or \U$31931 ( \32177 , \32175 , \32176 );
xor \U$31932 ( \32178 , RIbe2a3e8_88, RIbe2a460_89);
nand \U$31933 ( \32179 , \8794 , \32178 );
nand \U$31934 ( \32180 , \32177 , \32179 );
and \U$31935 ( \32181 , \32173 , \32180 );
not \U$31936 ( \32182 , \32173 );
not \U$31937 ( \32183 , \32180 );
and \U$31938 ( \32184 , \32182 , \32183 );
nor \U$31939 ( \32185 , \32181 , \32184 );
not \U$31940 ( \32186 , \32185 );
or \U$31941 ( \32187 , \32166 , \32186 );
not \U$31942 ( \32188 , \32183 );
nand \U$31943 ( \32189 , \32188 , \32173 );
nand \U$31944 ( \32190 , \32187 , \32189 );
not \U$31945 ( \32191 , \32190 );
and \U$31946 ( \32192 , \32159 , \32191 );
not \U$31947 ( \32193 , \32159 );
and \U$31948 ( \32194 , \32193 , \32190 );
or \U$31949 ( \32195 , \32192 , \32194 );
not \U$31950 ( \32196 , \31987 );
not \U$31951 ( \32197 , \16652 );
or \U$31952 ( \32198 , \32196 , \32197 );
nand \U$31953 ( \32199 , \4850 , \31759 );
nand \U$31954 ( \32200 , \32198 , \32199 );
xor \U$31955 ( \32201 , RIbe29ec0_77, RIbe2b180_117);
not \U$31956 ( \32202 , \32201 );
not \U$31957 ( \32203 , \15353 );
or \U$31958 ( \32204 , \32202 , \32203 );
nand \U$31959 ( \32205 , \21759 , \31650 );
nand \U$31960 ( \32206 , \32204 , \32205 );
xor \U$31961 ( \32207 , \32200 , \32206 );
not \U$31962 ( \32208 , \31977 );
not \U$31963 ( \32209 , \12000 );
or \U$31964 ( \32210 , \32208 , \32209 );
nand \U$31965 ( \32211 , \15995 , \31751 );
nand \U$31966 ( \32212 , \32210 , \32211 );
xnor \U$31967 ( \32213 , \32207 , \32212 );
and \U$31968 ( \32214 , \32195 , \32213 );
not \U$31969 ( \32215 , \32195 );
not \U$31970 ( \32216 , \32213 );
and \U$31971 ( \32217 , \32215 , \32216 );
nor \U$31972 ( \32218 , \32214 , \32217 );
not \U$31973 ( \32219 , \32218 );
not \U$31974 ( \32220 , \32219 );
xor \U$31975 ( \32221 , RIbe29d58_74, RIbe2b018_114);
not \U$31976 ( \32222 , \32221 );
not \U$31977 ( \32223 , \20396 );
or \U$31978 ( \32224 , \32222 , \32223 );
nand \U$31979 ( \32225 , \19371 , \32041 );
nand \U$31980 ( \32226 , \32224 , \32225 );
not \U$31981 ( \32227 , \32226 );
xor \U$31982 ( \32228 , RIbe29c68_72, RIbe2b450_123);
not \U$31983 ( \32229 , \32228 );
not \U$31984 ( \32230 , \7513 );
or \U$31985 ( \32231 , \32229 , \32230 );
nand \U$31986 ( \32232 , \7237 , \32105 );
nand \U$31987 ( \32233 , \32231 , \32232 );
nand \U$31988 ( \32234 , \4897 , RIbe2ae38_110);
not \U$31989 ( \32235 , \32234 );
and \U$31990 ( \32236 , \32233 , \32235 );
not \U$31991 ( \32237 , \32233 );
and \U$31992 ( \32238 , \32237 , \32234 );
nor \U$31993 ( \32239 , \32236 , \32238 );
not \U$31994 ( \32240 , \32239 );
or \U$31995 ( \32241 , \32227 , \32240 );
nand \U$31996 ( \32242 , \32233 , \32235 );
nand \U$31997 ( \32243 , \32241 , \32242 );
not \U$31998 ( \32244 , \32243 );
xor \U$31999 ( \32245 , RIbe2a2f8_86, RIbe2a6b8_94);
not \U$32000 ( \32246 , \32245 );
not \U$32001 ( \32247 , \14827 );
or \U$32002 ( \32248 , \32246 , \32247 );
xor \U$32003 ( \32249 , RIbe2a2f8_86, RIbe2b4c8_124);
nand \U$32004 ( \32250 , \8705 , \32249 );
nand \U$32005 ( \32251 , \32248 , \32250 );
not \U$32006 ( \32252 , \32251 );
xor \U$32007 ( \32253 , RIbe2a898_98, RIbe2b108_116);
not \U$32008 ( \32254 , \32253 );
not \U$32009 ( \32255 , \13529 );
or \U$32010 ( \32256 , \32254 , \32255 );
nand \U$32011 ( \32257 , \16875 , \32093 );
nand \U$32012 ( \32258 , \32256 , \32257 );
not \U$32013 ( \32259 , \32258 );
or \U$32014 ( \32260 , \32252 , \32259 );
or \U$32015 ( \32261 , \32258 , \32251 );
xor \U$32016 ( \32262 , RIbe2a7a8_96, RIbe29e48_76);
not \U$32017 ( \32263 , \32262 );
not \U$32018 ( \32264 , \7716 );
or \U$32019 ( \32265 , \32263 , \32264 );
xor \U$32020 ( \32266 , RIbe2abe0_105, RIbe29e48_76);
nand \U$32021 ( \32267 , \7368 , \32266 );
nand \U$32022 ( \32268 , \32265 , \32267 );
nand \U$32023 ( \32269 , \32261 , \32268 );
nand \U$32024 ( \32270 , \32260 , \32269 );
not \U$32025 ( \32271 , \32005 );
not \U$32026 ( \32272 , \32001 );
not \U$32027 ( \32273 , \32272 );
or \U$32028 ( \32274 , \32271 , \32273 );
or \U$32029 ( \32275 , \32272 , \32005 );
nand \U$32030 ( \32276 , \32274 , \32275 );
xor \U$32031 ( \32277 , \32270 , \32276 );
not \U$32032 ( \32278 , \32277 );
or \U$32033 ( \32279 , \32244 , \32278 );
nand \U$32034 ( \32280 , \32276 , \32270 );
nand \U$32035 ( \32281 , \32279 , \32280 );
not \U$32036 ( \32282 , \32281 );
and \U$32037 ( \32283 , \21852 , \32101 );
xor \U$32038 ( \32284 , RIbe2b6a8_128, RIbe2b108_116);
and \U$32039 ( \32285 , \13534 , \32284 );
nor \U$32040 ( \32286 , \32283 , \32285 );
not \U$32041 ( \32287 , \32286 );
and \U$32042 ( \32288 , \4574 , \32109 );
not \U$32043 ( \32289 , \32288 );
not \U$32044 ( \32290 , \4581 );
or \U$32045 ( \32291 , \32289 , \32290 );
nand \U$32046 ( \32292 , \4580 , \32153 );
nand \U$32047 ( \32293 , \32291 , \32292 );
not \U$32048 ( \32294 , \32054 );
not \U$32049 ( \32295 , \14852 );
or \U$32050 ( \32296 , \32294 , \32295 );
nand \U$32051 ( \32297 , \16646 , \32201 );
nand \U$32052 ( \32298 , \32296 , \32297 );
xor \U$32053 ( \32299 , \32293 , \32298 );
not \U$32054 ( \32300 , \32299 );
or \U$32055 ( \32301 , \32287 , \32300 );
or \U$32056 ( \32302 , \32299 , \32286 );
nand \U$32057 ( \32303 , \32301 , \32302 );
not \U$32058 ( \32304 , \32303 );
not \U$32059 ( \32305 , \32025 );
not \U$32060 ( \32306 , \32006 );
and \U$32061 ( \32307 , \32305 , \32306 );
and \U$32062 ( \32308 , \32025 , \32006 );
nor \U$32063 ( \32309 , \32307 , \32308 );
not \U$32064 ( \32310 , \32309 );
or \U$32065 ( \32311 , \32304 , \32310 );
or \U$32066 ( \32312 , \32309 , \32303 );
nand \U$32067 ( \32313 , \32311 , \32312 );
not \U$32068 ( \32314 , \32313 );
or \U$32069 ( \32315 , \32282 , \32314 );
not \U$32070 ( \32316 , \32309 );
nand \U$32071 ( \32317 , \32316 , \32303 );
nand \U$32072 ( \32318 , \32315 , \32317 );
not \U$32073 ( \32319 , \32013 );
not \U$32074 ( \32320 , \8169 );
or \U$32075 ( \32321 , \32319 , \32320 );
nand \U$32076 ( \32322 , \9065 , \31703 );
nand \U$32077 ( \32323 , \32321 , \32322 );
not \U$32078 ( \32324 , \32323 );
not \U$32079 ( \32325 , \32324 );
not \U$32080 ( \32326 , \32171 );
not \U$32081 ( \32327 , \8697 );
or \U$32082 ( \32328 , \32326 , \32327 );
not \U$32083 ( \32329 , \9378 );
nand \U$32084 ( \32330 , \32329 , \31784 );
nand \U$32085 ( \32331 , \32328 , \32330 );
xor \U$32086 ( \32332 , RIbe2ae38_110, RIbe27e68_8);
not \U$32087 ( \32333 , \32332 );
not \U$32088 ( \32334 , \2599 );
or \U$32089 ( \32335 , \32333 , \32334 );
nand \U$32090 ( \32336 , \2464 , \31778 );
nand \U$32091 ( \32337 , \32335 , \32336 );
xor \U$32092 ( \32338 , \32331 , \32337 );
not \U$32093 ( \32339 , \32338 );
or \U$32094 ( \32340 , \32325 , \32339 );
or \U$32095 ( \32341 , \32338 , \32324 );
nand \U$32096 ( \32342 , \32340 , \32341 );
not \U$32097 ( \32343 , \32342 );
not \U$32098 ( \32344 , \32178 );
not \U$32099 ( \32345 , \9096 );
or \U$32100 ( \32346 , \32344 , \32345 );
nand \U$32101 ( \32347 , \8793 , \31695 );
nand \U$32102 ( \32348 , \32346 , \32347 );
not \U$32103 ( \32349 , \32348 );
not \U$32104 ( \32350 , \32349 );
xor \U$32105 ( \32351 , RIbe298a8_64, RIbe2aaf0_103);
not \U$32106 ( \32352 , \32351 );
not \U$32107 ( \32353 , \18832 );
or \U$32108 ( \32354 , \32352 , \32353 );
nand \U$32109 ( \32355 , \31660 , RIbe2ab68_104);
nand \U$32110 ( \32356 , \32354 , \32355 );
not \U$32111 ( \32357 , \32356 );
and \U$32112 ( \32358 , \32350 , \32357 );
and \U$32113 ( \32359 , \32349 , \32356 );
nor \U$32114 ( \32360 , \32358 , \32359 );
xor \U$32115 ( \32361 , RIbe2b2e8_120, RIbe2a910_99);
not \U$32116 ( \32362 , \32361 );
not \U$32117 ( \32363 , \10987 );
or \U$32118 ( \32364 , \32362 , \32363 );
nand \U$32119 ( \32365 , \10401 , \31688 );
nand \U$32120 ( \32366 , \32364 , \32365 );
xor \U$32121 ( \32367 , \32360 , \32366 );
not \U$32122 ( \32368 , \32367 );
xor \U$32123 ( \32369 , RIbe28f48_44, RIbe2a730_95);
not \U$32124 ( \32370 , \32369 );
not \U$32125 ( \32371 , \9618 );
or \U$32126 ( \32372 , \32370 , \32371 );
nand \U$32127 ( \32373 , \9524 , \31676 );
nand \U$32128 ( \32374 , \32372 , \32373 );
not \U$32129 ( \32375 , \32019 );
not \U$32130 ( \32376 , \27992 );
or \U$32131 ( \32377 , \32375 , \32376 );
nand \U$32132 ( \32378 , \14649 , \31745 );
nand \U$32133 ( \32379 , \32377 , \32378 );
xor \U$32134 ( \32380 , \32374 , \32379 );
not \U$32135 ( \32381 , \32284 );
not \U$32136 ( \32382 , \14297 );
or \U$32137 ( \32383 , \32381 , \32382 );
nand \U$32138 ( \32384 , \23015 , \31667 );
nand \U$32139 ( \32385 , \32383 , \32384 );
xor \U$32140 ( \32386 , \32380 , \32385 );
not \U$32141 ( \32387 , \32386 );
or \U$32142 ( \32388 , \32368 , \32387 );
or \U$32143 ( \32389 , \32386 , \32367 );
nand \U$32144 ( \32390 , \32388 , \32389 );
not \U$32145 ( \32391 , \32390 );
not \U$32146 ( \32392 , \32391 );
or \U$32147 ( \32393 , \32343 , \32392 );
not \U$32148 ( \32394 , \32342 );
nand \U$32149 ( \32395 , \32394 , \32390 );
nand \U$32150 ( \32396 , \32393 , \32395 );
xor \U$32151 ( \32397 , \32318 , \32396 );
not \U$32152 ( \32398 , \32397 );
or \U$32153 ( \32399 , \32220 , \32398 );
nand \U$32154 ( \32400 , \32318 , \32396 );
nand \U$32155 ( \32401 , \32399 , \32400 );
not \U$32156 ( \32402 , \32401 );
not \U$32157 ( \32403 , \32402 );
or \U$32158 ( \32404 , \32136 , \32403 );
not \U$32159 ( \32405 , \32135 );
nand \U$32160 ( \32406 , \32405 , \32401 );
nand \U$32161 ( \32407 , \32404 , \32406 );
not \U$32162 ( \32408 , \32407 );
not \U$32163 ( \32409 , \32185 );
not \U$32164 ( \32410 , \32165 );
not \U$32165 ( \32411 , \32410 );
and \U$32166 ( \32412 , \32409 , \32411 );
and \U$32167 ( \32413 , \32185 , \32410 );
nor \U$32168 ( \32414 , \32412 , \32413 );
not \U$32169 ( \32415 , \32414 );
not \U$32170 ( \32416 , \32045 );
not \U$32171 ( \32417 , \16811 );
or \U$32172 ( \32418 , \32416 , \32417 );
nand \U$32173 ( \32419 , \18777 , \32137 );
nand \U$32174 ( \32420 , \32418 , \32419 );
xor \U$32175 ( \32421 , RIbe29d58_74, RIbe2af28_112);
not \U$32176 ( \32422 , \32421 );
not \U$32177 ( \32423 , \16913 );
or \U$32178 ( \32424 , \32422 , \32423 );
nand \U$32179 ( \32425 , \16917 , \32147 );
nand \U$32180 ( \32426 , \32424 , \32425 );
xor \U$32181 ( \32427 , \32420 , \32426 );
not \U$32182 ( \32428 , \32037 );
not \U$32183 ( \32429 , \11453 );
or \U$32184 ( \32430 , \32428 , \32429 );
nand \U$32185 ( \32431 , \11456 , \32361 );
nand \U$32186 ( \32432 , \32430 , \32431 );
xnor \U$32187 ( \32433 , \32427 , \32432 );
not \U$32188 ( \32434 , \32433 );
or \U$32189 ( \32435 , \32415 , \32434 );
xor \U$32190 ( \32436 , \31968 , \31979 );
xor \U$32191 ( \32437 , \32436 , \31989 );
nand \U$32192 ( \32438 , \32435 , \32437 );
not \U$32193 ( \32439 , \32414 );
not \U$32194 ( \32440 , \32433 );
nand \U$32195 ( \32441 , \32439 , \32440 );
nand \U$32196 ( \32442 , \32438 , \32441 );
not \U$32197 ( \32443 , \32442 );
xor \U$32198 ( \32444 , RIbe2ae38_110, RIbe27fd0_11);
not \U$32199 ( \32445 , \32444 );
not \U$32200 ( \32446 , \4893 );
or \U$32201 ( \32447 , \32445 , \32446 );
nand \U$32202 ( \32448 , \7709 , \32160 );
nand \U$32203 ( \32449 , \32447 , \32448 );
not \U$32204 ( \32450 , \32449 );
xor \U$32205 ( \32451 , RIbe2af28_112, RIbe29ec0_77);
not \U$32206 ( \32452 , \32451 );
not \U$32207 ( \32453 , \15345 );
or \U$32208 ( \32454 , \32452 , \32453 );
nand \U$32209 ( \32455 , \16917 , \32421 );
nand \U$32210 ( \32456 , \32454 , \32455 );
not \U$32211 ( \32457 , \32456 );
or \U$32212 ( \32458 , \32450 , \32457 );
or \U$32213 ( \32459 , \32456 , \32449 );
not \U$32214 ( \32460 , \32249 );
not \U$32215 ( \32461 , \9375 );
or \U$32216 ( \32462 , \32460 , \32461 );
nand \U$32217 ( \32463 , \11094 , \32167 );
nand \U$32218 ( \32464 , \32462 , \32463 );
nand \U$32219 ( \32465 , \32459 , \32464 );
nand \U$32220 ( \32466 , \32458 , \32465 );
and \U$32221 ( \32467 , \2463 , RIbe2ae38_110);
not \U$32222 ( \32468 , \32467 );
not \U$32223 ( \32469 , \32116 );
not \U$32224 ( \32470 , \23169 );
or \U$32225 ( \32471 , \32469 , \32470 );
nand \U$32226 ( \32472 , \32351 , RIbe2ab68_104);
nand \U$32227 ( \32473 , \32471 , \32472 );
not \U$32228 ( \32474 , \32473 );
not \U$32229 ( \32475 , \32474 );
or \U$32230 ( \32476 , \32468 , \32475 );
or \U$32231 ( \32477 , \32474 , \32467 );
nand \U$32232 ( \32478 , \32476 , \32477 );
not \U$32233 ( \32479 , \31999 );
not \U$32234 ( \32480 , \3256 );
or \U$32235 ( \32481 , \32479 , \32480 );
nand \U$32236 ( \32482 , \4181 , \32369 );
nand \U$32237 ( \32483 , \32481 , \32482 );
xor \U$32238 ( \32484 , \32478 , \32483 );
or \U$32239 ( \32485 , \32466 , \32484 );
not \U$32240 ( \32486 , \32266 );
not \U$32241 ( \32487 , \7716 );
or \U$32242 ( \32488 , \32486 , \32487 );
nand \U$32243 ( \32489 , \4851 , \31983 );
nand \U$32244 ( \32490 , \32488 , \32489 );
xor \U$32245 ( \32491 , RIbe2a3e8_88, RIbe2ad48_108);
not \U$32246 ( \32492 , \32491 );
or \U$32247 ( \32493 , \11544 , \32492 );
nand \U$32248 ( \32494 , \10476 , \32174 );
nand \U$32249 ( \32495 , \32493 , \32494 );
nor \U$32250 ( \32496 , \32490 , \32495 );
xor \U$32251 ( \32497 , RIbe2a0a0_81, RIbe2a190_83);
not \U$32252 ( \32498 , \32497 );
not \U$32253 ( \32499 , \15690 );
or \U$32254 ( \32500 , \32498 , \32499 );
nand \U$32255 ( \32501 , \15693 , \31963 );
nand \U$32256 ( \32502 , \32500 , \32501 );
not \U$32257 ( \32503 , \32502 );
or \U$32258 ( \32504 , \32496 , \32503 );
nand \U$32259 ( \32505 , \32490 , \32495 );
nand \U$32260 ( \32506 , \32504 , \32505 );
and \U$32261 ( \32507 , \32485 , \32506 );
and \U$32262 ( \32508 , \32466 , \32484 );
nor \U$32263 ( \32509 , \32507 , \32508 );
not \U$32264 ( \32510 , \32509 );
or \U$32265 ( \32511 , \32443 , \32510 );
or \U$32266 ( \32512 , \32442 , \32509 );
nand \U$32267 ( \32513 , \32511 , \32512 );
buf \U$32268 ( \32514 , \32513 );
not \U$32269 ( \32515 , \32286 );
not \U$32270 ( \32516 , \32515 );
not \U$32271 ( \32517 , \32299 );
or \U$32272 ( \32518 , \32516 , \32517 );
nand \U$32273 ( \32519 , \32298 , \32293 );
nand \U$32274 ( \32520 , \32518 , \32519 );
not \U$32275 ( \32521 , \32483 );
not \U$32276 ( \32522 , \32478 );
or \U$32277 ( \32523 , \32521 , \32522 );
nand \U$32278 ( \32524 , \32473 , \32467 );
nand \U$32279 ( \32525 , \32523 , \32524 );
not \U$32280 ( \32526 , \32525 );
not \U$32281 ( \32527 , \32526 );
not \U$32282 ( \32528 , \32426 );
not \U$32283 ( \32529 , \32420 );
nand \U$32284 ( \32530 , \32528 , \32529 );
not \U$32285 ( \32531 , \32530 );
not \U$32286 ( \32532 , \32432 );
or \U$32287 ( \32533 , \32531 , \32532 );
not \U$32288 ( \32534 , \32529 );
nand \U$32289 ( \32535 , \32534 , \32426 );
nand \U$32290 ( \32536 , \32533 , \32535 );
not \U$32291 ( \32537 , \32536 );
or \U$32292 ( \32538 , \32527 , \32537 );
or \U$32293 ( \32539 , \32536 , \32526 );
nand \U$32294 ( \32540 , \32538 , \32539 );
xor \U$32295 ( \32541 , \32520 , \32540 );
and \U$32296 ( \32542 , \32514 , \32541 );
not \U$32297 ( \32543 , \32514 );
not \U$32298 ( \32544 , \32541 );
and \U$32299 ( \32545 , \32543 , \32544 );
nor \U$32300 ( \32546 , \32542 , \32545 );
not \U$32301 ( \32547 , \32546 );
not \U$32302 ( \32548 , \31993 );
not \U$32303 ( \32549 , \32548 );
not \U$32304 ( \32550 , \32129 );
or \U$32305 ( \32551 , \32549 , \32550 );
or \U$32306 ( \32552 , \32129 , \32548 );
nand \U$32307 ( \32553 , \32551 , \32552 );
not \U$32308 ( \32554 , \32553 );
xor \U$32309 ( \32555 , \32484 , \32466 );
xor \U$32310 ( \32556 , \32555 , \32506 );
not \U$32311 ( \32557 , \32556 );
xor \U$32312 ( \32558 , RIbe2a118_82, RIbe2a280_85);
not \U$32313 ( \32559 , \32558 );
not \U$32314 ( \32560 , \14383 );
or \U$32315 ( \32561 , \32559 , \32560 );
nand \U$32316 ( \32562 , \11348 , \32068 );
nand \U$32317 ( \32563 , \32561 , \32562 );
not \U$32318 ( \32564 , \32563 );
xor \U$32319 ( \32565 , RIbe2b540_125, RIbe2a3e8_88);
not \U$32320 ( \32566 , \32565 );
not \U$32321 ( \32567 , \9263 );
or \U$32322 ( \32568 , \32566 , \32567 );
nand \U$32323 ( \32569 , \10476 , \32491 );
nand \U$32324 ( \32570 , \32568 , \32569 );
xor \U$32325 ( \32571 , RIbe2a910_99, RIbe2adc0_109);
not \U$32326 ( \32572 , \32571 );
not \U$32327 ( \32573 , \9737 );
or \U$32328 ( \32574 , \32572 , \32573 );
nand \U$32329 ( \32575 , \10400 , \32033 );
nand \U$32330 ( \32576 , \32574 , \32575 );
xor \U$32331 ( \32577 , \32570 , \32576 );
not \U$32332 ( \32578 , \32577 );
or \U$32333 ( \32579 , \32564 , \32578 );
nand \U$32334 ( \32580 , \32576 , \32570 );
nand \U$32335 ( \32581 , \32579 , \32580 );
not \U$32336 ( \32582 , \32581 );
xor \U$32337 ( \32583 , RIbe2a190_83, RIbe2b360_121);
not \U$32338 ( \32584 , \32583 );
not \U$32339 ( \32585 , \23387 );
or \U$32340 ( \32586 , \32584 , \32585 );
nand \U$32341 ( \32587 , \10834 , \32497 );
nand \U$32342 ( \32588 , \32586 , \32587 );
not \U$32343 ( \32589 , \32588 );
xor \U$32344 ( \32590 , RIbe2a028_80, RIbe2ac58_106);
not \U$32345 ( \32591 , \32590 );
not \U$32346 ( \32592 , \10674 );
or \U$32347 ( \32593 , \32591 , \32592 );
nand \U$32348 ( \32594 , \8172 , \32062 );
nand \U$32349 ( \32595 , \32593 , \32594 );
not \U$32350 ( \32596 , \32595 );
or \U$32351 ( \32597 , \32589 , \32596 );
or \U$32352 ( \32598 , \32595 , \32588 );
xor \U$32353 ( \32599 , RIbe28f48_44, RIbe2aeb0_111);
not \U$32354 ( \32600 , \32599 );
not \U$32355 ( \32601 , \8221 );
or \U$32356 ( \32602 , \32600 , \32601 );
nand \U$32357 ( \32603 , \3249 , \31995 );
nand \U$32358 ( \32604 , \32602 , \32603 );
nand \U$32359 ( \32605 , \32598 , \32604 );
nand \U$32360 ( \32606 , \32597 , \32605 );
not \U$32361 ( \32607 , \32606 );
xor \U$32362 ( \32608 , RIbe29b78_70, RIbe2aaf0_103);
not \U$32363 ( \32609 , \32608 );
not \U$32364 ( \32610 , \28282 );
or \U$32365 ( \32611 , \32609 , \32610 );
nand \U$32366 ( \32612 , \32112 , RIbe2ab68_104);
nand \U$32367 ( \32613 , \32611 , \32612 );
xor \U$32368 ( \32614 , RIbe2a4d8_90, RIbe2a550_91);
not \U$32369 ( \32615 , \32614 );
not \U$32370 ( \32616 , \26415 );
or \U$32371 ( \32617 , \32615 , \32616 );
nand \U$32372 ( \32618 , \11227 , \32076 );
nand \U$32373 ( \32619 , \32617 , \32618 );
xor \U$32374 ( \32620 , \32613 , \32619 );
and \U$32375 ( \32621 , RIbe29f38_78, RIbe2af28_112);
nor \U$32376 ( \32622 , RIbe29f38_78, RIbe2af28_112);
nor \U$32377 ( \32623 , \32621 , \32622 );
not \U$32378 ( \32624 , \32623 );
not \U$32379 ( \32625 , \15345 );
or \U$32380 ( \32626 , \32624 , \32625 );
nand \U$32381 ( \32627 , \19721 , \32451 );
nand \U$32382 ( \32628 , \32626 , \32627 );
and \U$32383 ( \32629 , \32620 , \32628 );
and \U$32384 ( \32630 , \32613 , \32619 );
nor \U$32385 ( \32631 , \32629 , \32630 );
not \U$32386 ( \32632 , \32631 );
or \U$32387 ( \32633 , \32607 , \32632 );
or \U$32388 ( \32634 , \32631 , \32606 );
nand \U$32389 ( \32635 , \32633 , \32634 );
not \U$32390 ( \32636 , \32635 );
or \U$32391 ( \32637 , \32582 , \32636 );
not \U$32392 ( \32638 , \32631 );
nand \U$32393 ( \32639 , \32638 , \32606 );
nand \U$32394 ( \32640 , \32637 , \32639 );
not \U$32395 ( \32641 , \32074 );
nand \U$32396 ( \32642 , \32641 , \32084 );
not \U$32397 ( \32643 , \32082 );
and \U$32398 ( \32644 , \32642 , \32643 );
not \U$32399 ( \32645 , \32642 );
and \U$32400 ( \32646 , \32645 , \32082 );
nor \U$32401 ( \32647 , \32644 , \32646 );
xor \U$32402 ( \32648 , \32047 , \32040 );
xnor \U$32403 ( \32649 , \32648 , \32056 );
nor \U$32404 ( \32650 , \32647 , \32649 );
xnor \U$32405 ( \32651 , \32119 , \32103 );
or \U$32406 ( \32652 , \32650 , \32651 );
nand \U$32407 ( \32653 , \32647 , \32649 );
nand \U$32408 ( \32654 , \32652 , \32653 );
and \U$32409 ( \32655 , \32640 , \32654 );
not \U$32410 ( \32656 , \32640 );
not \U$32411 ( \32657 , \32654 );
and \U$32412 ( \32658 , \32656 , \32657 );
nor \U$32413 ( \32659 , \32655 , \32658 );
not \U$32414 ( \32660 , \32659 );
or \U$32415 ( \32661 , \32557 , \32660 );
not \U$32416 ( \32662 , \32657 );
nand \U$32417 ( \32663 , \32662 , \32640 );
nand \U$32418 ( \32664 , \32661 , \32663 );
not \U$32419 ( \32665 , \32664 );
not \U$32420 ( \32666 , \32665 );
or \U$32421 ( \32667 , \32554 , \32666 );
not \U$32422 ( \32668 , \32664 );
or \U$32423 ( \32669 , \32668 , \32553 );
nand \U$32424 ( \32670 , \32667 , \32669 );
not \U$32425 ( \32671 , \32670 );
or \U$32426 ( \32672 , \32547 , \32671 );
not \U$32427 ( \32673 , \32668 );
nand \U$32428 ( \32674 , \32673 , \32553 );
nand \U$32429 ( \32675 , \32672 , \32674 );
not \U$32430 ( \32676 , \32675 );
not \U$32431 ( \32677 , \32676 );
and \U$32432 ( \32678 , \32408 , \32677 );
and \U$32433 ( \32679 , \32407 , \32676 );
nor \U$32434 ( \32680 , \32678 , \32679 );
not \U$32435 ( \32681 , \32680 );
not \U$32436 ( \32682 , \32681 );
not \U$32437 ( \32683 , \16646 );
not \U$32438 ( \32684 , RIbe2aa78_102);
not \U$32439 ( \32685 , RIbe2b180_117);
and \U$32440 ( \32686 , \32684 , \32685 );
and \U$32441 ( \32687 , RIbe2aa78_102, RIbe2b180_117);
nor \U$32442 ( \32688 , \32686 , \32687 );
not \U$32443 ( \32689 , \32688 );
or \U$32444 ( \32690 , \32683 , \32689 );
xnor \U$32445 ( \32691 , RIbe2b180_117, RIbe2aa00_101);
not \U$32446 ( \32692 , \32691 );
nand \U$32447 ( \32693 , \32692 , \14852 );
nand \U$32448 ( \32694 , \32690 , \32693 );
not \U$32449 ( \32695 , RIbe2a2f8_86);
not \U$32450 ( \32696 , RIbe2a640_93);
and \U$32451 ( \32697 , \32695 , \32696 );
and \U$32452 ( \32698 , RIbe2a2f8_86, RIbe2a640_93);
nor \U$32453 ( \32699 , \32697 , \32698 );
not \U$32454 ( \32700 , \32699 );
not \U$32455 ( \32701 , \10446 );
or \U$32456 ( \32702 , \32700 , \32701 );
nand \U$32457 ( \32703 , \8706 , \32245 );
nand \U$32458 ( \32704 , \32702 , \32703 );
nor \U$32459 ( \32705 , \32694 , \32704 );
xor \U$32460 ( \32706 , RIbe2b3d8_122, RIbe29c68_72);
not \U$32461 ( \32707 , \32706 );
not \U$32462 ( \32708 , \8595 );
or \U$32463 ( \32709 , \32707 , \32708 );
nand \U$32464 ( \32710 , \4580 , \32228 );
nand \U$32465 ( \32711 , \32709 , \32710 );
or \U$32466 ( \32712 , RIbe29bf0_71, RIbe29c68_72);
nand \U$32467 ( \32713 , \32712 , RIbe2ae38_110);
nand \U$32468 ( \32714 , RIbe29bf0_71, RIbe29c68_72);
and \U$32469 ( \32715 , \32713 , \32714 , RIbe28f48_44);
or \U$32470 ( \32716 , \32711 , \32715 );
nand \U$32471 ( \32717 , \32711 , \32715 );
nand \U$32472 ( \32718 , \32716 , \32717 );
or \U$32473 ( \32719 , \32705 , \32718 );
nand \U$32474 ( \32720 , \32694 , \32704 );
nand \U$32475 ( \32721 , \32719 , \32720 );
not \U$32476 ( \32722 , \32721 );
not \U$32477 ( \32723 , \32628 );
xor \U$32478 ( \32724 , \32620 , \32723 );
not \U$32479 ( \32725 , \32724 );
xnor \U$32480 ( \32726 , \32604 , \32588 );
not \U$32481 ( \32727 , \32595 );
and \U$32482 ( \32728 , \32726 , \32727 );
not \U$32483 ( \32729 , \32726 );
and \U$32484 ( \32730 , \32729 , \32595 );
nor \U$32485 ( \32731 , \32728 , \32730 );
not \U$32486 ( \32732 , \32731 );
or \U$32487 ( \32733 , \32725 , \32732 );
or \U$32488 ( \32734 , \32731 , \32724 );
nand \U$32489 ( \32735 , \32733 , \32734 );
not \U$32490 ( \32736 , \32735 );
or \U$32491 ( \32737 , \32722 , \32736 );
not \U$32492 ( \32738 , \32724 );
nand \U$32493 ( \32739 , \32738 , \32731 );
nand \U$32494 ( \32740 , \32737 , \32739 );
xnor \U$32495 ( \32741 , \32649 , \32647 );
and \U$32496 ( \32742 , \32741 , \32651 );
not \U$32497 ( \32743 , \32741 );
not \U$32498 ( \32744 , \32651 );
and \U$32499 ( \32745 , \32743 , \32744 );
nor \U$32500 ( \32746 , \32742 , \32745 );
xor \U$32501 ( \32747 , \32740 , \32746 );
xor \U$32502 ( \32748 , \32577 , \32563 );
not \U$32503 ( \32749 , \32748 );
not \U$32504 ( \32750 , \32226 );
and \U$32505 ( \32751 , \32239 , \32750 );
not \U$32506 ( \32752 , \32239 );
and \U$32507 ( \32753 , \32752 , \32226 );
nor \U$32508 ( \32754 , \32751 , \32753 );
not \U$32509 ( \32755 , \32754 );
xor \U$32510 ( \32756 , \32251 , \32258 );
and \U$32511 ( \32757 , \32756 , \32268 );
not \U$32512 ( \32758 , \32756 );
not \U$32513 ( \32759 , \32268 );
and \U$32514 ( \32760 , \32758 , \32759 );
nor \U$32515 ( \32761 , \32757 , \32760 );
not \U$32516 ( \32762 , \32761 );
and \U$32517 ( \32763 , \32755 , \32762 );
and \U$32518 ( \32764 , \32754 , \32761 );
nor \U$32519 ( \32765 , \32763 , \32764 );
not \U$32520 ( \32766 , \32765 );
not \U$32521 ( \32767 , \32766 );
or \U$32522 ( \32768 , \32749 , \32767 );
not \U$32523 ( \32769 , \32754 );
nand \U$32524 ( \32770 , \32769 , \32761 );
nand \U$32525 ( \32771 , \32768 , \32770 );
and \U$32526 ( \32772 , \32747 , \32771 );
and \U$32527 ( \32773 , \32740 , \32746 );
or \U$32528 ( \32774 , \32772 , \32773 );
not \U$32529 ( \32775 , \32774 );
xor \U$32530 ( \32776 , RIbe2af28_112, RIbe2b6a8_128);
not \U$32531 ( \32777 , \32776 );
not \U$32532 ( \32778 , \18649 );
or \U$32533 ( \32779 , \32777 , \32778 );
nand \U$32534 ( \32780 , \19721 , \32623 );
nand \U$32535 ( \32781 , \32779 , \32780 );
not \U$32536 ( \32782 , \32781 );
xor \U$32537 ( \32783 , RIbe2b2e8_120, RIbe2a190_83);
not \U$32538 ( \32784 , \32783 );
not \U$32539 ( \32785 , \14730 );
or \U$32540 ( \32786 , \32784 , \32785 );
nand \U$32541 ( \32787 , \13278 , \32583 );
nand \U$32542 ( \32788 , \32786 , \32787 );
xor \U$32543 ( \32789 , RIbe28f48_44, RIbe2ae38_110);
not \U$32544 ( \32790 , \32789 );
not \U$32545 ( \32791 , \9618 );
or \U$32546 ( \32792 , \32790 , \32791 );
nand \U$32547 ( \32793 , \11201 , \32599 );
nand \U$32548 ( \32794 , \32792 , \32793 );
xor \U$32549 ( \32795 , \32788 , \32794 );
not \U$32550 ( \32796 , \32795 );
or \U$32551 ( \32797 , \32782 , \32796 );
nand \U$32552 ( \32798 , \32794 , \32788 );
nand \U$32553 ( \32799 , \32797 , \32798 );
not \U$32554 ( \32800 , \32799 );
xor \U$32555 ( \32801 , RIbe2a3e8_88, RIbe2b4c8_124);
not \U$32556 ( \32802 , \32801 );
not \U$32557 ( \32803 , \12590 );
or \U$32558 ( \32804 , \32802 , \32803 );
nand \U$32559 ( \32805 , \8794 , \32565 );
nand \U$32560 ( \32806 , \32804 , \32805 );
not \U$32561 ( \32807 , \32806 );
xor \U$32562 ( \32808 , RIbe2a028_80, RIbe2abe0_105);
not \U$32563 ( \32809 , \32808 );
not \U$32564 ( \32810 , \8168 );
or \U$32565 ( \32811 , \32809 , \32810 );
nand \U$32566 ( \32812 , \8930 , \32590 );
nand \U$32567 ( \32813 , \32811 , \32812 );
xor \U$32568 ( \32814 , RIbe2a910_99, RIbe2ad48_108);
not \U$32569 ( \32815 , \32814 );
not \U$32570 ( \32816 , \9736 );
or \U$32571 ( \32817 , \32815 , \32816 );
nand \U$32572 ( \32818 , \10400 , \32571 );
nand \U$32573 ( \32819 , \32817 , \32818 );
and \U$32574 ( \32820 , \32813 , \32819 );
not \U$32575 ( \32821 , \32813 );
not \U$32576 ( \32822 , \32819 );
and \U$32577 ( \32823 , \32821 , \32822 );
nor \U$32578 ( \32824 , \32820 , \32823 );
not \U$32579 ( \32825 , \32824 );
or \U$32580 ( \32826 , \32807 , \32825 );
not \U$32581 ( \32827 , \32822 );
nand \U$32582 ( \32828 , \32827 , \32813 );
nand \U$32583 ( \32829 , \32826 , \32828 );
xor \U$32584 ( \32830 , RIbe2a730_95, RIbe29e48_76);
not \U$32585 ( \32831 , \32830 );
not \U$32586 ( \32832 , \4843 );
or \U$32587 ( \32833 , \32831 , \32832 );
nand \U$32588 ( \32834 , \4851 , \32262 );
nand \U$32589 ( \32835 , \32833 , \32834 );
not \U$32590 ( \32836 , \32835 );
xor \U$32591 ( \32837 , RIbe2a0a0_81, RIbe2a280_85);
not \U$32592 ( \32838 , \32837 );
not \U$32593 ( \32839 , \10845 );
or \U$32594 ( \32840 , \32838 , \32839 );
nand \U$32595 ( \32841 , \18667 , \32558 );
nand \U$32596 ( \32842 , \32840 , \32841 );
not \U$32597 ( \32843 , \32842 );
not \U$32598 ( \32844 , \32843 );
xor \U$32599 ( \32845 , RIbe2b108_116, RIbe2a820_97);
not \U$32600 ( \32846 , \32845 );
not \U$32601 ( \32847 , \14296 );
or \U$32602 ( \32848 , \32846 , \32847 );
nand \U$32603 ( \32849 , \16875 , \32253 );
nand \U$32604 ( \32850 , \32848 , \32849 );
not \U$32605 ( \32851 , \32850 );
or \U$32606 ( \32852 , \32844 , \32851 );
or \U$32607 ( \32853 , \32850 , \32843 );
nand \U$32608 ( \32854 , \32852 , \32853 );
not \U$32609 ( \32855 , \32854 );
or \U$32610 ( \32856 , \32836 , \32855 );
nand \U$32611 ( \32857 , \32850 , \32842 );
nand \U$32612 ( \32858 , \32856 , \32857 );
xor \U$32613 ( \32859 , \32829 , \32858 );
not \U$32614 ( \32860 , \32859 );
or \U$32615 ( \32861 , \32800 , \32860 );
nand \U$32616 ( \32862 , \32858 , \32829 );
nand \U$32617 ( \32863 , \32861 , \32862 );
xor \U$32618 ( \32864 , \32277 , \32243 );
nor \U$32619 ( \32865 , \32863 , \32864 );
xnor \U$32620 ( \32866 , \32635 , \32581 );
or \U$32621 ( \32867 , \32865 , \32866 );
nand \U$32622 ( \32868 , \32863 , \32864 );
nand \U$32623 ( \32869 , \32867 , \32868 );
buf \U$32624 ( \32870 , \32313 );
buf \U$32625 ( \32871 , \32281 );
xor \U$32626 ( \32872 , \32870 , \32871 );
xor \U$32627 ( \32873 , \32869 , \32872 );
not \U$32628 ( \32874 , \32873 );
or \U$32629 ( \32875 , \32775 , \32874 );
nand \U$32630 ( \32876 , \32869 , \32872 );
nand \U$32631 ( \32877 , \32875 , \32876 );
not \U$32632 ( \32878 , \32877 );
xnor \U$32633 ( \32879 , \32218 , \32397 );
not \U$32634 ( \32880 , \32879 );
xor \U$32635 ( \32881 , \32414 , \32437 );
xnor \U$32636 ( \32882 , \32881 , \32440 );
not \U$32637 ( \32883 , \32882 );
xor \U$32638 ( \32884 , \32060 , \32087 );
xnor \U$32639 ( \32885 , \32884 , \32123 );
not \U$32640 ( \32886 , \32885 );
not \U$32641 ( \32887 , \32886 );
not \U$32642 ( \32888 , \32496 );
nand \U$32643 ( \32889 , \32888 , \32505 );
and \U$32644 ( \32890 , \32889 , \32502 );
not \U$32645 ( \32891 , \32889 );
and \U$32646 ( \32892 , \32891 , \32503 );
nor \U$32647 ( \32893 , \32890 , \32892 );
xor \U$32648 ( \32894 , \32449 , \32464 );
xnor \U$32649 ( \32895 , \32894 , \32456 );
nand \U$32650 ( \32896 , \32893 , \32895 );
not \U$32651 ( \32897 , \32896 );
not \U$32652 ( \32898 , \32717 );
not \U$32653 ( \32899 , \32898 );
buf \U$32654 ( \32900 , \14852 );
and \U$32655 ( \32901 , \32900 , \32688 );
and \U$32656 ( \32902 , \14966 , \32050 );
nor \U$32657 ( \32903 , \32901 , \32902 );
not \U$32658 ( \32904 , \32903 );
xor \U$32659 ( \32905 , RIbe29ce0_73, RIbe2aaf0_103);
not \U$32660 ( \32906 , \32905 );
not \U$32661 ( \32907 , \19581 );
or \U$32662 ( \32908 , \32906 , \32907 );
nand \U$32663 ( \32909 , \32608 , RIbe2ab68_104);
nand \U$32664 ( \32910 , \32908 , \32909 );
not \U$32665 ( \32911 , \32910 );
xor \U$32666 ( \32912 , RIbe29ec0_77, RIbe2b018_114);
not \U$32667 ( \32913 , \32912 );
not \U$32668 ( \32914 , \16811 );
or \U$32669 ( \32915 , \32913 , \32914 );
nand \U$32670 ( \32916 , \15953 , \32221 );
nand \U$32671 ( \32917 , \32915 , \32916 );
buf \U$32672 ( \32918 , \32917 );
not \U$32673 ( \32919 , \32918 );
or \U$32674 ( \32920 , \32911 , \32919 );
not \U$32675 ( \32921 , \32917 );
not \U$32676 ( \32922 , \32910 );
nand \U$32677 ( \32923 , \32921 , \32922 );
xor \U$32678 ( \32924 , RIbe2a550_91, RIbe2a460_89);
not \U$32679 ( \32925 , \32924 );
not \U$32680 ( \32926 , \10433 );
or \U$32681 ( \32927 , \32925 , \32926 );
nand \U$32682 ( \32928 , \14612 , \32614 );
nand \U$32683 ( \32929 , \32927 , \32928 );
nand \U$32684 ( \32930 , \32923 , \32929 );
nand \U$32685 ( \32931 , \32920 , \32930 );
not \U$32686 ( \32932 , \32931 );
or \U$32687 ( \32933 , \32904 , \32932 );
or \U$32688 ( \32934 , \32903 , \32931 );
nand \U$32689 ( \32935 , \32933 , \32934 );
not \U$32690 ( \32936 , \32935 );
or \U$32691 ( \32937 , \32899 , \32936 );
not \U$32692 ( \32938 , \32903 );
nand \U$32693 ( \32939 , \32938 , \32931 );
nand \U$32694 ( \32940 , \32937 , \32939 );
not \U$32695 ( \32941 , \32940 );
or \U$32696 ( \32942 , \32897 , \32941 );
not \U$32697 ( \32943 , \32893 );
not \U$32698 ( \32944 , \32895 );
nand \U$32699 ( \32945 , \32943 , \32944 );
nand \U$32700 ( \32946 , \32942 , \32945 );
not \U$32701 ( \32947 , \32946 );
not \U$32702 ( \32948 , \32947 );
or \U$32703 ( \32949 , \32887 , \32948 );
nand \U$32704 ( \32950 , \32946 , \32885 );
nand \U$32705 ( \32951 , \32949 , \32950 );
not \U$32706 ( \32952 , \32951 );
or \U$32707 ( \32953 , \32883 , \32952 );
nand \U$32708 ( \32954 , \32946 , \32886 );
nand \U$32709 ( \32955 , \32953 , \32954 );
not \U$32710 ( \32956 , \32955 );
not \U$32711 ( \32957 , \32956 );
and \U$32712 ( \32958 , \32880 , \32957 );
and \U$32713 ( \32959 , \32879 , \32956 );
nor \U$32714 ( \32960 , \32958 , \32959 );
not \U$32715 ( \32961 , \32960 );
not \U$32716 ( \32962 , \32961 );
or \U$32717 ( \32963 , \32878 , \32962 );
not \U$32718 ( \32964 , \32956 );
nand \U$32719 ( \32965 , \32964 , \32879 );
nand \U$32720 ( \32966 , \32963 , \32965 );
not \U$32721 ( \32967 , \32966 );
not \U$32722 ( \32968 , \31992 );
not \U$32723 ( \32969 , \31962 );
or \U$32724 ( \32970 , \32968 , \32969 );
nand \U$32725 ( \32971 , \31961 , \31950 );
nand \U$32726 ( \32972 , \32970 , \32971 );
not \U$32727 ( \32973 , \32525 );
not \U$32728 ( \32974 , \32536 );
or \U$32729 ( \32975 , \32973 , \32974 );
nand \U$32730 ( \32976 , \32540 , \32520 );
nand \U$32731 ( \32977 , \32975 , \32976 );
xor \U$32732 ( \32978 , \32972 , \32977 );
xor \U$32733 ( \32979 , \32374 , \32379 );
and \U$32734 ( \32980 , \32979 , \32385 );
and \U$32735 ( \32981 , \32374 , \32379 );
or \U$32736 ( \32982 , \32980 , \32981 );
not \U$32737 ( \32983 , \32323 );
not \U$32738 ( \32984 , \32337 );
or \U$32739 ( \32985 , \32983 , \32984 );
or \U$32740 ( \32986 , \32337 , \32323 );
nand \U$32741 ( \32987 , \32986 , \32331 );
nand \U$32742 ( \32988 , \32985 , \32987 );
xor \U$32743 ( \32989 , \32982 , \32988 );
not \U$32744 ( \32990 , \32348 );
not \U$32745 ( \32991 , \32356 );
or \U$32746 ( \32992 , \32990 , \32991 );
not \U$32747 ( \32993 , \32366 );
or \U$32748 ( \32994 , \32360 , \32993 );
nand \U$32749 ( \32995 , \32992 , \32994 );
buf \U$32750 ( \32996 , \32995 );
xor \U$32751 ( \32997 , \32989 , \32996 );
xor \U$32752 ( \32998 , \32978 , \32997 );
not \U$32753 ( \32999 , \32541 );
not \U$32754 ( \33000 , \32513 );
or \U$32755 ( \33001 , \32999 , \33000 );
not \U$32756 ( \33002 , \32509 );
nand \U$32757 ( \33003 , \33002 , \32442 );
nand \U$32758 ( \33004 , \33001 , \33003 );
nor \U$32759 ( \33005 , \32998 , \33004 );
not \U$32760 ( \33006 , \33005 );
nand \U$32761 ( \33007 , \32998 , \33004 );
nand \U$32762 ( \33008 , \33006 , \33007 );
not \U$32763 ( \33009 , \33008 );
not \U$32764 ( \33010 , \32342 );
not \U$32765 ( \33011 , \32390 );
or \U$32766 ( \33012 , \33010 , \33011 );
not \U$32767 ( \33013 , \32367 );
nand \U$32768 ( \33014 , \33013 , \32386 );
nand \U$32769 ( \33015 , \33012 , \33014 );
nand \U$32770 ( \33016 , \31960 , \31954 );
not \U$32771 ( \33017 , \32206 );
not \U$32772 ( \33018 , \32212 );
or \U$32773 ( \33019 , \33017 , \33018 );
or \U$32774 ( \33020 , \32212 , \32206 );
nand \U$32775 ( \33021 , \33020 , \32200 );
nand \U$32776 ( \33022 , \33019 , \33021 );
xor \U$32777 ( \33023 , \33016 , \33022 );
not \U$32778 ( \33024 , \32142 );
nand \U$32779 ( \33025 , \33024 , \32150 );
not \U$32780 ( \33026 , \33025 );
not \U$32781 ( \33027 , \32158 );
or \U$32782 ( \33028 , \33026 , \33027 );
nand \U$32783 ( \33029 , \32151 , \32142 );
nand \U$32784 ( \33030 , \33028 , \33029 );
not \U$32785 ( \33031 , \33030 );
xnor \U$32786 ( \33032 , \33023 , \33031 );
not \U$32787 ( \33033 , \33032 );
not \U$32788 ( \33034 , \33033 );
not \U$32789 ( \33035 , \32190 );
not \U$32790 ( \33036 , \32216 );
or \U$32791 ( \33037 , \33035 , \33036 );
not \U$32792 ( \33038 , \32213 );
not \U$32793 ( \33039 , \32191 );
or \U$32794 ( \33040 , \33038 , \33039 );
nand \U$32795 ( \33041 , \33040 , \32159 );
nand \U$32796 ( \33042 , \33037 , \33041 );
not \U$32797 ( \33043 , \33042 );
not \U$32798 ( \33044 , \33043 );
or \U$32799 ( \33045 , \33034 , \33044 );
or \U$32800 ( \33046 , \33043 , \33033 );
nand \U$32801 ( \33047 , \33045 , \33046 );
xnor \U$32802 ( \33048 , \33015 , \33047 );
not \U$32803 ( \33049 , \33048 );
not \U$32804 ( \33050 , \33049 );
and \U$32805 ( \33051 , \33009 , \33050 );
and \U$32806 ( \33052 , \33049 , \33008 );
nor \U$32807 ( \33053 , \33051 , \33052 );
nand \U$32808 ( \33054 , \32967 , \33053 );
not \U$32809 ( \33055 , \33054 );
or \U$32810 ( \33056 , \32682 , \33055 );
not \U$32811 ( \33057 , \33053 );
nand \U$32812 ( \33058 , \33057 , \32966 );
nand \U$32813 ( \33059 , \33056 , \33058 );
not \U$32814 ( \33060 , \33042 );
not \U$32815 ( \33061 , \33033 );
or \U$32816 ( \33062 , \33060 , \33061 );
not \U$32817 ( \33063 , \33032 );
not \U$32818 ( \33064 , \33043 );
or \U$32819 ( \33065 , \33063 , \33064 );
nand \U$32820 ( \33066 , \33065 , \33015 );
nand \U$32821 ( \33067 , \33062 , \33066 );
xor \U$32822 ( \33068 , \32972 , \32977 );
and \U$32823 ( \33069 , \33068 , \32997 );
and \U$32824 ( \33070 , \32972 , \32977 );
or \U$32825 ( \33071 , \33069 , \33070 );
and \U$32826 ( \33072 , \33067 , \33071 );
not \U$32827 ( \33073 , \33067 );
not \U$32828 ( \33074 , \33071 );
and \U$32829 ( \33075 , \33073 , \33074 );
nor \U$32830 ( \33076 , \33072 , \33075 );
xor \U$32831 ( \33077 , \31658 , \31684 );
xor \U$32832 ( \33078 , \33077 , \31716 );
not \U$32833 ( \33079 , \31933 );
not \U$32834 ( \33080 , \31916 );
or \U$32835 ( \33081 , \33079 , \33080 );
not \U$32836 ( \33082 , \31932 );
not \U$32837 ( \33083 , \31915 );
or \U$32838 ( \33084 , \33082 , \33083 );
nand \U$32839 ( \33085 , \33084 , \31926 );
nand \U$32840 ( \33086 , \33081 , \33085 );
not \U$32841 ( \33087 , \33086 );
xor \U$32842 ( \33088 , \31743 , \31768 );
xor \U$32843 ( \33089 , \33088 , \31799 );
not \U$32844 ( \33090 , \33089 );
or \U$32845 ( \33091 , \33087 , \33090 );
or \U$32846 ( \33092 , \33089 , \33086 );
nand \U$32847 ( \33093 , \33091 , \33092 );
xor \U$32848 ( \33094 , \33078 , \33093 );
not \U$32849 ( \33095 , \33094 );
and \U$32850 ( \33096 , \33076 , \33095 );
not \U$32851 ( \33097 , \33076 );
and \U$32852 ( \33098 , \33097 , \33094 );
nor \U$32853 ( \33099 , \33096 , \33098 );
not \U$32854 ( \33100 , \33099 );
not \U$32855 ( \33101 , \31829 );
nand \U$32856 ( \33102 , \33101 , \31835 );
not \U$32857 ( \33103 , \31833 );
and \U$32858 ( \33104 , \33102 , \33103 );
not \U$32859 ( \33105 , \33102 );
and \U$32860 ( \33106 , \33105 , \31833 );
nor \U$32861 ( \33107 , \33104 , \33106 );
xnor \U$32862 ( \33108 , \31479 , \31493 );
not \U$32863 ( \33109 , \33108 );
xor \U$32864 ( \33110 , \31385 , \31391 );
xor \U$32865 ( \33111 , \33110 , \31398 );
not \U$32866 ( \33112 , \33111 );
or \U$32867 ( \33113 , \33109 , \33112 );
or \U$32868 ( \33114 , \33111 , \33108 );
nand \U$32869 ( \33115 , \33113 , \33114 );
buf \U$32870 ( \33116 , \33115 );
xor \U$32871 ( \33117 , \33107 , \33116 );
not \U$32872 ( \33118 , \31579 );
not \U$32873 ( \33119 , \31585 );
or \U$32874 ( \33120 , \33118 , \33119 );
or \U$32875 ( \33121 , \31585 , \31579 );
nand \U$32876 ( \33122 , \33120 , \33121 );
not \U$32877 ( \33123 , \33122 );
not \U$32878 ( \33124 , \31588 );
and \U$32879 ( \33125 , \33123 , \33124 );
and \U$32880 ( \33126 , \33122 , \31588 );
nor \U$32881 ( \33127 , \33125 , \33126 );
xnor \U$32882 ( \33128 , \33117 , \33127 );
xor \U$32883 ( \33129 , \31905 , \31910 );
and \U$32884 ( \33130 , \33129 , \31912 );
and \U$32885 ( \33131 , \31905 , \31910 );
or \U$32886 ( \33132 , \33130 , \33131 );
not \U$32887 ( \33133 , \33132 );
not \U$32888 ( \33134 , \33133 );
or \U$32889 ( \33135 , \32988 , \32995 );
nand \U$32890 ( \33136 , \33135 , \32982 );
nand \U$32891 ( \33137 , \32988 , \32995 );
and \U$32892 ( \33138 , \33136 , \33137 );
not \U$32893 ( \33139 , \33016 );
not \U$32894 ( \33140 , \33031 );
or \U$32895 ( \33141 , \33139 , \33140 );
nand \U$32896 ( \33142 , \33141 , \33022 );
not \U$32897 ( \33143 , \33016 );
nand \U$32898 ( \33144 , \33143 , \33030 );
nand \U$32899 ( \33145 , \33142 , \33144 );
not \U$32900 ( \33146 , \33145 );
and \U$32901 ( \33147 , \33138 , \33146 );
not \U$32902 ( \33148 , \33138 );
and \U$32903 ( \33149 , \33148 , \33145 );
nor \U$32904 ( \33150 , \33147 , \33149 );
not \U$32905 ( \33151 , \33150 );
or \U$32906 ( \33152 , \33134 , \33151 );
or \U$32907 ( \33153 , \33150 , \33133 );
nand \U$32908 ( \33154 , \33152 , \33153 );
and \U$32909 ( \33155 , \33128 , \33154 );
not \U$32910 ( \33156 , \33128 );
not \U$32911 ( \33157 , \33154 );
and \U$32912 ( \33158 , \33156 , \33157 );
nor \U$32913 ( \33159 , \33155 , \33158 );
not \U$32914 ( \33160 , \32134 );
not \U$32915 ( \33161 , \31942 );
or \U$32916 ( \33162 , \33160 , \33161 );
nand \U$32917 ( \33163 , \31913 , \31940 );
nand \U$32918 ( \33164 , \33162 , \33163 );
xor \U$32919 ( \33165 , \33159 , \33164 );
not \U$32920 ( \33166 , \33165 );
or \U$32921 ( \33167 , \33048 , \33005 );
nand \U$32922 ( \33168 , \33167 , \33007 );
not \U$32923 ( \33169 , \33168 );
not \U$32924 ( \33170 , \33169 );
and \U$32925 ( \33171 , \33166 , \33170 );
and \U$32926 ( \33172 , \33165 , \33169 );
nor \U$32927 ( \33173 , \33171 , \33172 );
xor \U$32928 ( \33174 , \33100 , \33173 );
not \U$32929 ( \33175 , \32675 );
not \U$32930 ( \33176 , \32407 );
or \U$32931 ( \33177 , \33175 , \33176 );
nand \U$32932 ( \33178 , \32401 , \32135 );
nand \U$32933 ( \33179 , \33177 , \33178 );
buf \U$32934 ( \33180 , \33179 );
xnor \U$32935 ( \33181 , \33174 , \33180 );
nand \U$32936 ( \33182 , \33059 , \33181 );
buf \U$32937 ( \33183 , \32659 );
buf \U$32938 ( \33184 , \32556 );
not \U$32939 ( \33185 , \33184 );
and \U$32940 ( \33186 , \33183 , \33185 );
not \U$32941 ( \33187 , \33183 );
and \U$32942 ( \33188 , \33187 , \33184 );
nor \U$32943 ( \33189 , \33186 , \33188 );
not \U$32944 ( \33190 , \33189 );
and \U$32945 ( \33191 , \32951 , \32882 );
not \U$32946 ( \33192 , \32951 );
not \U$32947 ( \33193 , \32882 );
and \U$32948 ( \33194 , \33192 , \33193 );
nor \U$32949 ( \33195 , \33191 , \33194 );
not \U$32950 ( \33196 , \33195 );
or \U$32951 ( \33197 , \33190 , \33196 );
or \U$32952 ( \33198 , \33195 , \33189 );
nand \U$32953 ( \33199 , \33197 , \33198 );
xor \U$32954 ( \33200 , \32873 , \32774 );
and \U$32955 ( \33201 , \33199 , \33200 );
not \U$32956 ( \33202 , \33195 );
nor \U$32957 ( \33203 , \33202 , \33189 );
nor \U$32958 ( \33204 , \33201 , \33203 );
not \U$32959 ( \33205 , \33204 );
not \U$32960 ( \33206 , \33205 );
not \U$32961 ( \33207 , \32877 );
not \U$32962 ( \33208 , \33207 );
not \U$32963 ( \33209 , \32961 );
or \U$32964 ( \33210 , \33208 , \33209 );
nand \U$32965 ( \33211 , \32960 , \32877 );
nand \U$32966 ( \33212 , \33210 , \33211 );
xor \U$32967 ( \33213 , \32670 , \32546 );
or \U$32968 ( \33214 , \33212 , \33213 );
not \U$32969 ( \33215 , \33214 );
or \U$32970 ( \33216 , \33206 , \33215 );
nand \U$32971 ( \33217 , \33212 , \33213 );
nand \U$32972 ( \33218 , \33216 , \33217 );
xor \U$32973 ( \33219 , \33053 , \32680 );
xor \U$32974 ( \33220 , \33219 , \32966 );
nand \U$32975 ( \33221 , \33218 , \33220 );
nand \U$32976 ( \33222 , \33182 , \33221 );
not \U$32977 ( \33223 , \33222 );
not \U$32978 ( \33224 , \33223 );
nor \U$32979 ( \33225 , \33218 , \33220 );
xor \U$32980 ( \33226 , \33213 , \33204 );
xnor \U$32981 ( \33227 , \33226 , \33212 );
not \U$32982 ( \33228 , \33200 );
xor \U$32983 ( \33229 , \33199 , \33228 );
not \U$32984 ( \33230 , \33229 );
not \U$32985 ( \33231 , \33230 );
xnor \U$32986 ( \33232 , \32735 , \32721 );
not \U$32987 ( \33233 , \33232 );
not \U$32988 ( \33234 , \33233 );
xor \U$32989 ( \33235 , \32781 , \32795 );
xor \U$32990 ( \33236 , \32806 , \32824 );
nor \U$32991 ( \33237 , \33235 , \33236 );
xnor \U$32992 ( \33238 , \32854 , \32835 );
or \U$32993 ( \33239 , \33237 , \33238 );
nand \U$32994 ( \33240 , \33235 , \33236 );
nand \U$32995 ( \33241 , \33239 , \33240 );
not \U$32996 ( \33242 , \33241 );
not \U$32997 ( \33243 , \32799 );
and \U$32998 ( \33244 , \32859 , \33243 );
not \U$32999 ( \33245 , \32859 );
and \U$33000 ( \33246 , \33245 , \32799 );
nor \U$33001 ( \33247 , \33244 , \33246 );
not \U$33002 ( \33248 , \33247 );
or \U$33003 ( \33249 , \33242 , \33248 );
or \U$33004 ( \33250 , \33241 , \33247 );
nand \U$33005 ( \33251 , \33249 , \33250 );
not \U$33006 ( \33252 , \33251 );
or \U$33007 ( \33253 , \33234 , \33252 );
not \U$33008 ( \33254 , \33247 );
nand \U$33009 ( \33255 , \33254 , \33241 );
nand \U$33010 ( \33256 , \33253 , \33255 );
not \U$33011 ( \33257 , \33256 );
xor \U$33012 ( \33258 , \32944 , \32893 );
xnor \U$33013 ( \33259 , \33258 , \32940 );
xor \U$33014 ( \33260 , RIbe2b450_123, RIbe29e48_76);
and \U$33015 ( \33261 , \4843 , \33260 );
and \U$33016 ( \33262 , \4851 , \32830 );
nor \U$33017 ( \33263 , \33261 , \33262 );
not \U$33018 ( \33264 , \33263 );
not \U$33019 ( \33265 , \33264 );
not \U$33020 ( \33266 , \24871 );
nand \U$33021 ( \33267 , \33266 , \9524 );
not \U$33022 ( \33268 , \33267 );
xor \U$33023 ( \33269 , RIbe2a4d8_90, RIbe2a190_83);
not \U$33024 ( \33270 , \33269 );
not \U$33025 ( \33271 , \10690 );
or \U$33026 ( \33272 , \33270 , \33271 );
nand \U$33027 ( \33273 , \10695 , \32783 );
nand \U$33028 ( \33274 , \33272 , \33273 );
not \U$33029 ( \33275 , \33274 );
or \U$33030 ( \33276 , \33268 , \33275 );
or \U$33031 ( \33277 , \33274 , \33267 );
nand \U$33032 ( \33278 , \33276 , \33277 );
not \U$33033 ( \33279 , \33278 );
or \U$33034 ( \33280 , \33265 , \33279 );
not \U$33035 ( \33281 , \33267 );
nand \U$33036 ( \33282 , \33281 , \33274 );
nand \U$33037 ( \33283 , \33280 , \33282 );
not \U$33038 ( \33284 , RIbe2a2f8_86);
not \U$33039 ( \33285 , RIbe2ac58_106);
and \U$33040 ( \33286 , \33284 , \33285 );
and \U$33041 ( \33287 , RIbe2a2f8_86, RIbe2ac58_106);
nor \U$33042 ( \33288 , \33286 , \33287 );
not \U$33043 ( \33289 , \33288 );
not \U$33044 ( \33290 , \10446 );
or \U$33045 ( \33291 , \33289 , \33290 );
nand \U$33046 ( \33292 , \9379 , \32699 );
nand \U$33047 ( \33293 , \33291 , \33292 );
not \U$33048 ( \33294 , \33293 );
xor \U$33049 ( \33295 , RIbe2b108_116, RIbe2a118_82);
not \U$33050 ( \33296 , \33295 );
not \U$33051 ( \33297 , \14296 );
or \U$33052 ( \33298 , \33296 , \33297 );
nand \U$33053 ( \33299 , \13533 , \32845 );
nand \U$33054 ( \33300 , \33298 , \33299 );
not \U$33055 ( \33301 , \33300 );
xor \U$33056 ( \33302 , RIbe2a910_99, RIbe2b540_125);
not \U$33057 ( \33303 , \33302 );
not \U$33058 ( \33304 , \9736 );
or \U$33059 ( \33305 , \33303 , \33304 );
nand \U$33060 ( \33306 , \10400 , \32814 );
nand \U$33061 ( \33307 , \33305 , \33306 );
not \U$33062 ( \33308 , \33307 );
not \U$33063 ( \33309 , \33308 );
or \U$33064 ( \33310 , \33301 , \33309 );
not \U$33065 ( \33311 , \33300 );
nand \U$33066 ( \33312 , \33311 , \33307 );
nand \U$33067 ( \33313 , \33310 , \33312 );
not \U$33068 ( \33314 , \33313 );
or \U$33069 ( \33315 , \33294 , \33314 );
nand \U$33070 ( \33316 , \33300 , \33307 );
nand \U$33071 ( \33317 , \33315 , \33316 );
xor \U$33072 ( \33318 , \33283 , \33317 );
and \U$33073 ( \33319 , \7642 , \32706 );
not \U$33074 ( \33320 , \8595 );
xnor \U$33075 ( \33321 , RIbe2aeb0_111, RIbe29c68_72);
nor \U$33076 ( \33322 , \33320 , \33321 );
nor \U$33077 ( \33323 , \33319 , \33322 );
not \U$33078 ( \33324 , \33323 );
not \U$33079 ( \33325 , \33324 );
xor \U$33080 ( \33326 , RIbe2adc0_109, RIbe2a550_91);
not \U$33081 ( \33327 , \33326 );
not \U$33082 ( \33328 , \10433 );
or \U$33083 ( \33329 , \33327 , \33328 );
nand \U$33084 ( \33330 , \23306 , \32924 );
nand \U$33085 ( \33331 , \33329 , \33330 );
xor \U$33086 ( \33332 , RIbe2a280_85, RIbe2b360_121);
not \U$33087 ( \33333 , \33332 );
not \U$33088 ( \33334 , \14942 );
or \U$33089 ( \33335 , \33333 , \33334 );
nand \U$33090 ( \33336 , \11348 , \32837 );
nand \U$33091 ( \33337 , \33335 , \33336 );
xor \U$33092 ( \33338 , \33331 , \33337 );
not \U$33093 ( \33339 , \33338 );
or \U$33094 ( \33340 , \33325 , \33339 );
nand \U$33095 ( \33341 , \33337 , \33331 );
nand \U$33096 ( \33342 , \33340 , \33341 );
and \U$33097 ( \33343 , \33318 , \33342 );
and \U$33098 ( \33344 , \33283 , \33317 );
or \U$33099 ( \33345 , \33343 , \33344 );
not \U$33100 ( \33346 , \33345 );
and \U$33101 ( \33347 , \32935 , \32717 );
not \U$33102 ( \33348 , \32935 );
and \U$33103 ( \33349 , \33348 , \32898 );
nor \U$33104 ( \33350 , \33347 , \33349 );
not \U$33105 ( \33351 , \33350 );
xor \U$33106 ( \33352 , RIbe29d58_74, RIbe2aaf0_103);
not \U$33107 ( \33353 , \33352 );
not \U$33108 ( \33354 , \19581 );
or \U$33109 ( \33355 , \33353 , \33354 );
nand \U$33110 ( \33356 , \32905 , RIbe2ab68_104);
nand \U$33111 ( \33357 , \33355 , \33356 );
xor \U$33112 ( \33358 , RIbe2af28_112, RIbe2aa78_102);
not \U$33113 ( \33359 , \33358 );
not \U$33114 ( \33360 , \16913 );
or \U$33115 ( \33361 , \33359 , \33360 );
nand \U$33116 ( \33362 , \17810 , \32776 );
nand \U$33117 ( \33363 , \33361 , \33362 );
xor \U$33118 ( \33364 , \33357 , \33363 );
not \U$33119 ( \33365 , \32912 );
not \U$33120 ( \33366 , \15953 );
or \U$33121 ( \33367 , \33365 , \33366 );
not \U$33122 ( \33368 , \20396 );
xor \U$33123 ( \33369 , RIbe2b018_114, RIbe29f38_78);
not \U$33124 ( \33370 , \33369 );
or \U$33125 ( \33371 , \33368 , \33370 );
nand \U$33126 ( \33372 , \33367 , \33371 );
and \U$33127 ( \33373 , \33364 , \33372 );
and \U$33128 ( \33374 , \33357 , \33363 );
or \U$33129 ( \33375 , \33373 , \33374 );
buf \U$33130 ( \33376 , \32918 );
not \U$33131 ( \33377 , \33376 );
not \U$33132 ( \33378 , \32929 );
not \U$33133 ( \33379 , \32922 );
and \U$33134 ( \33380 , \33378 , \33379 );
and \U$33135 ( \33381 , \32929 , \32922 );
nor \U$33136 ( \33382 , \33380 , \33381 );
not \U$33137 ( \33383 , \33382 );
or \U$33138 ( \33384 , \33377 , \33383 );
or \U$33139 ( \33385 , \33382 , \33376 );
nand \U$33140 ( \33386 , \33384 , \33385 );
xor \U$33141 ( \33387 , \33375 , \33386 );
xor \U$33142 ( \33388 , RIbe2a898_98, RIbe2b180_117);
nand \U$33143 ( \33389 , \33388 , \14849 );
and \U$33144 ( \33390 , \25254 , \33389 );
not \U$33145 ( \33391 , \25254 );
and \U$33146 ( \33392 , \33391 , \32691 );
or \U$33147 ( \33393 , \33390 , \33392 );
not \U$33148 ( \33394 , \33393 );
not \U$33149 ( \33395 , \33394 );
xor \U$33150 ( \33396 , RIbe2a7a8_96, RIbe2a028_80);
not \U$33151 ( \33397 , \33396 );
not \U$33152 ( \33398 , \8401 );
or \U$33153 ( \33399 , \33397 , \33398 );
nand \U$33154 ( \33400 , \9065 , \32808 );
nand \U$33155 ( \33401 , \33399 , \33400 );
not \U$33156 ( \33402 , \33401 );
or \U$33157 ( \33403 , \33395 , \33402 );
not \U$33158 ( \33404 , \33393 );
not \U$33159 ( \33405 , \33401 );
or \U$33160 ( \33406 , \33404 , \33405 );
or \U$33161 ( \33407 , \33401 , \33393 );
nand \U$33162 ( \33408 , \33406 , \33407 );
xor \U$33163 ( \33409 , RIbe2a3e8_88, RIbe2a6b8_94);
not \U$33164 ( \33410 , \33409 );
not \U$33165 ( \33411 , \9263 );
or \U$33166 ( \33412 , \33410 , \33411 );
nand \U$33167 ( \33413 , \11541 , \32801 );
nand \U$33168 ( \33414 , \33412 , \33413 );
nand \U$33169 ( \33415 , \33408 , \33414 );
nand \U$33170 ( \33416 , \33403 , \33415 );
and \U$33171 ( \33417 , \33387 , \33416 );
and \U$33172 ( \33418 , \33375 , \33386 );
or \U$33173 ( \33419 , \33417 , \33418 );
not \U$33174 ( \33420 , \33419 );
or \U$33175 ( \33421 , \33351 , \33420 );
or \U$33176 ( \33422 , \33419 , \33350 );
nand \U$33177 ( \33423 , \33421 , \33422 );
not \U$33178 ( \33424 , \33423 );
or \U$33179 ( \33425 , \33346 , \33424 );
not \U$33180 ( \33426 , \33350 );
nand \U$33181 ( \33427 , \33426 , \33419 );
nand \U$33182 ( \33428 , \33425 , \33427 );
xor \U$33183 ( \33429 , \33259 , \33428 );
not \U$33184 ( \33430 , \33429 );
or \U$33185 ( \33431 , \33257 , \33430 );
nand \U$33186 ( \33432 , \33428 , \33259 );
nand \U$33187 ( \33433 , \33431 , \33432 );
xor \U$33188 ( \33434 , \32740 , \32746 );
xor \U$33189 ( \33435 , \33434 , \32771 );
not \U$33190 ( \33436 , \33435 );
xnor \U$33191 ( \33437 , \32748 , \32765 );
not \U$33192 ( \33438 , \33437 );
xor \U$33193 ( \33439 , RIbe2a460_89, RIbe2a190_83);
not \U$33194 ( \33440 , \33439 );
not \U$33195 ( \33441 , \15690 );
or \U$33196 ( \33442 , \33440 , \33441 );
nand \U$33197 ( \33443 , \11400 , \33269 );
nand \U$33198 ( \33444 , \33442 , \33443 );
xor \U$33199 ( \33445 , RIbe2b2e8_120, RIbe2a280_85);
not \U$33200 ( \33446 , \33445 );
not \U$33201 ( \33447 , \20237 );
or \U$33202 ( \33448 , \33446 , \33447 );
nand \U$33203 ( \33449 , \11348 , \33332 );
nand \U$33204 ( \33450 , \33448 , \33449 );
or \U$33205 ( \33451 , \33444 , \33450 );
xor \U$33206 ( \33452 , RIbe29c68_72, RIbe2ae38_110);
not \U$33207 ( \33453 , \33452 );
not \U$33208 ( \33454 , \8259 );
or \U$33209 ( \33455 , \33453 , \33454 );
not \U$33210 ( \33456 , \33321 );
nand \U$33211 ( \33457 , \33456 , \4580 );
nand \U$33212 ( \33458 , \33455 , \33457 );
nand \U$33213 ( \33459 , \33451 , \33458 );
nand \U$33214 ( \33460 , \33450 , \33444 );
nand \U$33215 ( \33461 , \33459 , \33460 );
not \U$33216 ( \33462 , \33461 );
nand \U$33217 ( \33463 , RIbe29dd0_75, RIbe29e48_76);
or \U$33218 ( \33464 , RIbe29dd0_75, RIbe29e48_76);
nand \U$33219 ( \33465 , \33464 , RIbe2ae38_110);
nand \U$33220 ( \33466 , \33463 , RIbe29c68_72, \33465 );
not \U$33221 ( \33467 , \33466 );
xor \U$33222 ( \33468 , RIbe29e48_76, RIbe2b3d8_122);
not \U$33223 ( \33469 , \33468 );
not \U$33224 ( \33470 , \19978 );
or \U$33225 ( \33471 , \33469 , \33470 );
nand \U$33226 ( \33472 , \16655 , \33260 );
nand \U$33227 ( \33473 , \33471 , \33472 );
nand \U$33228 ( \33474 , \33467 , \33473 );
not \U$33229 ( \33475 , \33474 );
xor \U$33230 ( \33476 , RIbe2a2f8_86, RIbe2abe0_105);
not \U$33231 ( \33477 , \33476 );
not \U$33232 ( \33478 , \10792 );
or \U$33233 ( \33479 , \33477 , \33478 );
nand \U$33234 ( \33480 , \8706 , \33288 );
nand \U$33235 ( \33481 , \33479 , \33480 );
not \U$33236 ( \33482 , \33481 );
xor \U$33237 ( \33483 , RIbe2ad48_108, RIbe2a550_91);
not \U$33238 ( \33484 , \33483 );
not \U$33239 ( \33485 , \10433 );
or \U$33240 ( \33486 , \33484 , \33485 );
nand \U$33241 ( \33487 , \15995 , \33326 );
nand \U$33242 ( \33488 , \33486 , \33487 );
not \U$33243 ( \33489 , \33488 );
or \U$33244 ( \33490 , \33482 , \33489 );
or \U$33245 ( \33491 , \33488 , \33481 );
xor \U$33246 ( \33492 , RIbe2b108_116, RIbe2a0a0_81);
not \U$33247 ( \33493 , \33492 );
not \U$33248 ( \33494 , \14297 );
or \U$33249 ( \33495 , \33493 , \33494 );
nand \U$33250 ( \33496 , \13534 , \33295 );
nand \U$33251 ( \33497 , \33495 , \33496 );
nand \U$33252 ( \33498 , \33491 , \33497 );
nand \U$33253 ( \33499 , \33490 , \33498 );
not \U$33254 ( \33500 , \33499 );
or \U$33255 ( \33501 , \33475 , \33500 );
or \U$33256 ( \33502 , \33499 , \33474 );
nand \U$33257 ( \33503 , \33501 , \33502 );
not \U$33258 ( \33504 , \33503 );
or \U$33259 ( \33505 , \33462 , \33504 );
not \U$33260 ( \33506 , \33474 );
nand \U$33261 ( \33507 , \33506 , \33499 );
nand \U$33262 ( \33508 , \33505 , \33507 );
not \U$33263 ( \33509 , \33508 );
not \U$33264 ( \33510 , \32720 );
nor \U$33265 ( \33511 , \33510 , \32705 );
xor \U$33266 ( \33512 , \33511 , \32718 );
not \U$33267 ( \33513 , \33512 );
xor \U$33268 ( \33514 , \33313 , \33293 );
not \U$33269 ( \33515 , \33514 );
not \U$33270 ( \33516 , \33278 );
not \U$33271 ( \33517 , \33263 );
and \U$33272 ( \33518 , \33516 , \33517 );
and \U$33273 ( \33519 , \33278 , \33263 );
nor \U$33274 ( \33520 , \33518 , \33519 );
nand \U$33275 ( \33521 , \33515 , \33520 );
not \U$33276 ( \33522 , \33521 );
xor \U$33277 ( \33523 , \33357 , \33363 );
xor \U$33278 ( \33524 , \33523 , \33372 );
not \U$33279 ( \33525 , \33524 );
or \U$33280 ( \33526 , \33522 , \33525 );
buf \U$33281 ( \33527 , \33514 );
not \U$33282 ( \33528 , \33520 );
nand \U$33283 ( \33529 , \33527 , \33528 );
nand \U$33284 ( \33530 , \33526 , \33529 );
not \U$33285 ( \33531 , \33530 );
or \U$33286 ( \33532 , \33513 , \33531 );
or \U$33287 ( \33533 , \33530 , \33512 );
nand \U$33288 ( \33534 , \33532 , \33533 );
not \U$33289 ( \33535 , \33534 );
or \U$33290 ( \33536 , \33509 , \33535 );
not \U$33291 ( \33537 , \33512 );
nand \U$33292 ( \33538 , \33537 , \33530 );
nand \U$33293 ( \33539 , \33536 , \33538 );
not \U$33294 ( \33540 , \33539 );
or \U$33295 ( \33541 , \33438 , \33540 );
or \U$33296 ( \33542 , \33539 , \33437 );
not \U$33297 ( \33543 , \33338 );
not \U$33298 ( \33544 , \33323 );
and \U$33299 ( \33545 , \33543 , \33544 );
and \U$33300 ( \33546 , \33338 , \33323 );
nor \U$33301 ( \33547 , \33545 , \33546 );
not \U$33302 ( \33548 , \33547 );
not \U$33303 ( \33549 , \33548 );
xor \U$33304 ( \33550 , RIbe2a910_99, RIbe2b4c8_124);
not \U$33305 ( \33551 , \33550 );
not \U$33306 ( \33552 , \9737 );
or \U$33307 ( \33553 , \33551 , \33552 );
nand \U$33308 ( \33554 , \10400 , \33302 );
nand \U$33309 ( \33555 , \33553 , \33554 );
xor \U$33310 ( \33556 , RIbe2a028_80, RIbe2a730_95);
not \U$33311 ( \33557 , \33556 );
not \U$33312 ( \33558 , \22849 );
or \U$33313 ( \33559 , \33557 , \33558 );
nand \U$33314 ( \33560 , \8930 , \33396 );
nand \U$33315 ( \33561 , \33559 , \33560 );
nor \U$33316 ( \33562 , \33555 , \33561 );
xor \U$33317 ( \33563 , RIbe2b180_117, RIbe2a820_97);
not \U$33318 ( \33564 , \33563 );
not \U$33319 ( \33565 , \15353 );
or \U$33320 ( \33566 , \33564 , \33565 );
nand \U$33321 ( \33567 , \14966 , \33388 );
nand \U$33322 ( \33568 , \33566 , \33567 );
not \U$33323 ( \33569 , \33568 );
or \U$33324 ( \33570 , \33562 , \33569 );
nand \U$33325 ( \33571 , \33555 , \33561 );
nand \U$33326 ( \33572 , \33570 , \33571 );
not \U$33327 ( \33573 , \33572 );
xor \U$33328 ( \33574 , RIbe2af28_112, RIbe2aa00_101);
not \U$33329 ( \33575 , \33574 );
not \U$33330 ( \33576 , \16913 );
or \U$33331 ( \33577 , \33575 , \33576 );
nand \U$33332 ( \33578 , \19721 , \33358 );
nand \U$33333 ( \33579 , \33577 , \33578 );
not \U$33334 ( \33580 , \33579 );
xor \U$33335 ( \33581 , RIbe29ec0_77, RIbe2aaf0_103);
not \U$33336 ( \33582 , \33581 );
not \U$33337 ( \33583 , \20574 );
or \U$33338 ( \33584 , \33582 , \33583 );
nand \U$33339 ( \33585 , \33352 , RIbe2ab68_104);
nand \U$33340 ( \33586 , \33584 , \33585 );
not \U$33341 ( \33587 , \33586 );
xor \U$33342 ( \33588 , RIbe2a3e8_88, RIbe2a640_93);
not \U$33343 ( \33589 , \33588 );
not \U$33344 ( \33590 , \9096 );
or \U$33345 ( \33591 , \33589 , \33590 );
nand \U$33346 ( \33592 , \8793 , \33409 );
nand \U$33347 ( \33593 , \33591 , \33592 );
not \U$33348 ( \33594 , \33593 );
not \U$33349 ( \33595 , \33594 );
or \U$33350 ( \33596 , \33587 , \33595 );
or \U$33351 ( \33597 , \33594 , \33586 );
nand \U$33352 ( \33598 , \33596 , \33597 );
not \U$33353 ( \33599 , \33598 );
or \U$33354 ( \33600 , \33580 , \33599 );
nand \U$33355 ( \33601 , \33593 , \33586 );
nand \U$33356 ( \33602 , \33600 , \33601 );
not \U$33357 ( \33603 , \33602 );
not \U$33358 ( \33604 , \33603 );
or \U$33359 ( \33605 , \33573 , \33604 );
not \U$33360 ( \33606 , \33572 );
nand \U$33361 ( \33607 , \33606 , \33602 );
nand \U$33362 ( \33608 , \33605 , \33607 );
not \U$33363 ( \33609 , \33608 );
or \U$33364 ( \33610 , \33549 , \33609 );
nand \U$33365 ( \33611 , \33572 , \33602 );
nand \U$33366 ( \33612 , \33610 , \33611 );
xor \U$33367 ( \33613 , \33375 , \33386 );
xor \U$33368 ( \33614 , \33613 , \33416 );
or \U$33369 ( \33615 , \33612 , \33614 );
xor \U$33370 ( \33616 , \33283 , \33317 );
xor \U$33371 ( \33617 , \33616 , \33342 );
nand \U$33372 ( \33618 , \33615 , \33617 );
nand \U$33373 ( \33619 , \33612 , \33614 );
nand \U$33374 ( \33620 , \33618 , \33619 );
nand \U$33375 ( \33621 , \33542 , \33620 );
nand \U$33376 ( \33622 , \33541 , \33621 );
xor \U$33377 ( \33623 , \32864 , \32866 );
xor \U$33378 ( \33624 , \33623 , \32863 );
not \U$33379 ( \33625 , \33624 );
and \U$33380 ( \33626 , \33622 , \33625 );
not \U$33381 ( \33627 , \33622 );
and \U$33382 ( \33628 , \33627 , \33624 );
nor \U$33383 ( \33629 , \33626 , \33628 );
not \U$33384 ( \33630 , \33629 );
or \U$33385 ( \33631 , \33436 , \33630 );
nand \U$33386 ( \33632 , \33622 , \33625 );
nand \U$33387 ( \33633 , \33631 , \33632 );
xor \U$33388 ( \33634 , \33433 , \33633 );
not \U$33389 ( \33635 , \33634 );
or \U$33390 ( \33636 , \33231 , \33635 );
nand \U$33391 ( \33637 , \33633 , \33433 );
nand \U$33392 ( \33638 , \33636 , \33637 );
nor \U$33393 ( \33639 , \33227 , \33638 );
nor \U$33394 ( \33640 , \33225 , \33639 );
nand \U$33395 ( \33641 , \33227 , \33638 );
not \U$33396 ( \33642 , \33229 );
not \U$33397 ( \33643 , \33634 );
or \U$33398 ( \33644 , \33642 , \33643 );
not \U$33399 ( \33645 , \33229 );
not \U$33400 ( \33646 , \33634 );
nand \U$33401 ( \33647 , \33645 , \33646 );
nand \U$33402 ( \33648 , \33644 , \33647 );
xor \U$33403 ( \33649 , \33450 , \33444 );
xnor \U$33404 ( \33650 , \33649 , \33458 );
not \U$33405 ( \33651 , \33650 );
not \U$33406 ( \33652 , \33651 );
xor \U$33407 ( \33653 , \33598 , \33579 );
not \U$33408 ( \33654 , \33653 );
not \U$33409 ( \33655 , \33562 );
nand \U$33410 ( \33656 , \33655 , \33571 );
and \U$33411 ( \33657 , \33656 , \33568 );
not \U$33412 ( \33658 , \33656 );
and \U$33413 ( \33659 , \33658 , \33569 );
nor \U$33414 ( \33660 , \33657 , \33659 );
not \U$33415 ( \33661 , \33660 );
or \U$33416 ( \33662 , \33654 , \33661 );
or \U$33417 ( \33663 , \33660 , \33653 );
nand \U$33418 ( \33664 , \33662 , \33663 );
not \U$33419 ( \33665 , \33664 );
or \U$33420 ( \33666 , \33652 , \33665 );
not \U$33421 ( \33667 , \33660 );
nand \U$33422 ( \33668 , \33667 , \33653 );
nand \U$33423 ( \33669 , \33666 , \33668 );
not \U$33424 ( \33670 , \33669 );
not \U$33425 ( \33671 , \33461 );
xor \U$33426 ( \33672 , \33503 , \33671 );
not \U$33427 ( \33673 , \33672 );
and \U$33428 ( \33674 , \33608 , \33548 );
not \U$33429 ( \33675 , \33608 );
and \U$33430 ( \33676 , \33675 , \33547 );
nor \U$33431 ( \33677 , \33674 , \33676 );
not \U$33432 ( \33678 , \33677 );
or \U$33433 ( \33679 , \33673 , \33678 );
or \U$33434 ( \33680 , \33677 , \33672 );
nand \U$33435 ( \33681 , \33679 , \33680 );
not \U$33436 ( \33682 , \33681 );
or \U$33437 ( \33683 , \33670 , \33682 );
not \U$33438 ( \33684 , \33672 );
nand \U$33439 ( \33685 , \33684 , \33677 );
nand \U$33440 ( \33686 , \33683 , \33685 );
not \U$33441 ( \33687 , \33686 );
not \U$33442 ( \33688 , \33235 );
not \U$33443 ( \33689 , \33688 );
not \U$33444 ( \33690 , \33236 );
not \U$33445 ( \33691 , \33238 );
or \U$33446 ( \33692 , \33690 , \33691 );
or \U$33447 ( \33693 , \33238 , \33236 );
nand \U$33448 ( \33694 , \33692 , \33693 );
not \U$33449 ( \33695 , \33694 );
or \U$33450 ( \33696 , \33689 , \33695 );
or \U$33451 ( \33697 , \33694 , \33688 );
nand \U$33452 ( \33698 , \33696 , \33697 );
not \U$33453 ( \33699 , \33698 );
xor \U$33454 ( \33700 , RIbe2af28_112, RIbe2a898_98);
not \U$33455 ( \33701 , \33700 );
not \U$33456 ( \33702 , \15345 );
or \U$33457 ( \33703 , \33701 , \33702 );
nand \U$33458 ( \33704 , \17810 , \33574 );
nand \U$33459 ( \33705 , \33703 , \33704 );
not \U$33460 ( \33706 , \33705 );
xor \U$33461 ( \33707 , RIbe2b540_125, RIbe2a550_91);
not \U$33462 ( \33708 , \33707 );
not \U$33463 ( \33709 , \12000 );
or \U$33464 ( \33710 , \33708 , \33709 );
nand \U$33465 ( \33711 , \12004 , \33483 );
nand \U$33466 ( \33712 , \33710 , \33711 );
not \U$33467 ( \33713 , \33712 );
or \U$33468 ( \33714 , \33706 , \33713 );
or \U$33469 ( \33715 , \33712 , \33705 );
not \U$33470 ( \33716 , RIbe2a118_82);
not \U$33471 ( \33717 , RIbe2b180_117);
and \U$33472 ( \33718 , \33716 , \33717 );
and \U$33473 ( \33719 , RIbe2a118_82, RIbe2b180_117);
nor \U$33474 ( \33720 , \33718 , \33719 );
not \U$33475 ( \33721 , \33720 );
not \U$33476 ( \33722 , \15353 );
or \U$33477 ( \33723 , \33721 , \33722 );
nand \U$33478 ( \33724 , \14966 , \33563 );
nand \U$33479 ( \33725 , \33723 , \33724 );
nand \U$33480 ( \33726 , \33715 , \33725 );
nand \U$33481 ( \33727 , \33714 , \33726 );
not \U$33482 ( \33728 , \33727 );
not \U$33483 ( \33729 , \33728 );
not \U$33484 ( \33730 , RIbe2a6b8_94);
not \U$33485 ( \33731 , RIbe2a910_99);
and \U$33486 ( \33732 , \33730 , \33731 );
and \U$33487 ( \33733 , RIbe2a6b8_94, RIbe2a910_99);
nor \U$33488 ( \33734 , \33732 , \33733 );
not \U$33489 ( \33735 , \33734 );
not \U$33490 ( \33736 , \11453 );
or \U$33491 ( \33737 , \33735 , \33736 );
nand \U$33492 ( \33738 , \10401 , \33550 );
nand \U$33493 ( \33739 , \33737 , \33738 );
xor \U$33494 ( \33740 , RIbe2aa78_102, RIbe2b018_114);
not \U$33495 ( \33741 , \33740 );
not \U$33496 ( \33742 , \15967 );
or \U$33497 ( \33743 , \33741 , \33742 );
xor \U$33498 ( \33744 , RIbe2b018_114, RIbe2b6a8_128);
nand \U$33499 ( \33745 , \19371 , \33744 );
nand \U$33500 ( \33746 , \33743 , \33745 );
nor \U$33501 ( \33747 , \33739 , \33746 );
xor \U$33502 ( \33748 , RIbe2a4d8_90, RIbe2a280_85);
and \U$33503 ( \33749 , \20237 , \33748 );
and \U$33504 ( \33750 , \11348 , \33445 );
nor \U$33505 ( \33751 , \33749 , \33750 );
or \U$33506 ( \33752 , \33747 , \33751 );
nand \U$33507 ( \33753 , \33739 , \33746 );
nand \U$33508 ( \33754 , \33752 , \33753 );
not \U$33509 ( \33755 , \33754 );
not \U$33510 ( \33756 , \33755 );
or \U$33511 ( \33757 , \33729 , \33756 );
xor \U$33512 ( \33758 , RIbe2a7a8_96, RIbe2a2f8_86);
not \U$33513 ( \33759 , \33758 );
not \U$33514 ( \33760 , \9375 );
or \U$33515 ( \33761 , \33759 , \33760 );
nand \U$33516 ( \33762 , \8706 , \33476 );
nand \U$33517 ( \33763 , \33761 , \33762 );
not \U$33518 ( \33764 , \33763 );
xor \U$33519 ( \33765 , RIbe29e48_76, RIbe2aeb0_111);
not \U$33520 ( \33766 , \33765 );
not \U$33521 ( \33767 , \16652 );
or \U$33522 ( \33768 , \33766 , \33767 );
nand \U$33523 ( \33769 , \7368 , \33468 );
nand \U$33524 ( \33770 , \33768 , \33769 );
xor \U$33525 ( \33771 , RIbe2a3e8_88, RIbe2ac58_106);
not \U$33526 ( \33772 , \33771 );
not \U$33527 ( \33773 , \9263 );
or \U$33528 ( \33774 , \33772 , \33773 );
nand \U$33529 ( \33775 , \10476 , \33588 );
nand \U$33530 ( \33776 , \33774 , \33775 );
xor \U$33531 ( \33777 , \33770 , \33776 );
not \U$33532 ( \33778 , \33777 );
or \U$33533 ( \33779 , \33764 , \33778 );
nand \U$33534 ( \33780 , \33770 , \33776 );
nand \U$33535 ( \33781 , \33779 , \33780 );
nand \U$33536 ( \33782 , \33757 , \33781 );
nand \U$33537 ( \33783 , \33754 , \33727 );
nand \U$33538 ( \33784 , \33782 , \33783 );
not \U$33539 ( \33785 , \33784 );
not \U$33540 ( \33786 , \33414 );
not \U$33541 ( \33787 , \33786 );
not \U$33542 ( \33788 , \33408 );
or \U$33543 ( \33789 , \33787 , \33788 );
or \U$33544 ( \33790 , \33408 , \33786 );
nand \U$33545 ( \33791 , \33789 , \33790 );
not \U$33546 ( \33792 , \33744 );
not \U$33547 ( \33793 , \16812 );
or \U$33548 ( \33794 , \33792 , \33793 );
nand \U$33549 ( \33795 , \20583 , \33369 );
nand \U$33550 ( \33796 , \33794 , \33795 );
not \U$33551 ( \33797 , \33796 );
not \U$33552 ( \33798 , \33473 );
not \U$33553 ( \33799 , \33466 );
and \U$33554 ( \33800 , \33798 , \33799 );
and \U$33555 ( \33801 , \33473 , \33466 );
nor \U$33556 ( \33802 , \33800 , \33801 );
not \U$33557 ( \33803 , \33802 );
or \U$33558 ( \33804 , \33797 , \33803 );
or \U$33559 ( \33805 , \33802 , \33796 );
nand \U$33560 ( \33806 , \33804 , \33805 );
not \U$33561 ( \33807 , \33806 );
xor \U$33562 ( \33808 , RIbe2b450_123, RIbe2a028_80);
not \U$33563 ( \33809 , \33808 );
not \U$33564 ( \33810 , \8400 );
or \U$33565 ( \33811 , \33809 , \33810 );
nand \U$33566 ( \33812 , \8172 , \33556 );
nand \U$33567 ( \33813 , \33811 , \33812 );
nand \U$33568 ( \33814 , \4580 , RIbe2ae38_110);
nor \U$33569 ( \33815 , \33813 , \33814 );
not \U$33570 ( \33816 , \33815 );
nand \U$33571 ( \33817 , \33813 , \33814 );
nand \U$33572 ( \33818 , \33816 , \33817 );
not \U$33573 ( \33819 , \33818 );
xor \U$33574 ( \33820 , RIbe2a190_83, RIbe2adc0_109);
not \U$33575 ( \33821 , \33820 );
not \U$33576 ( \33822 , \31943 );
or \U$33577 ( \33823 , \33821 , \33822 );
nand \U$33578 ( \33824 , \31948 , \33439 );
nand \U$33579 ( \33825 , \33823 , \33824 );
not \U$33580 ( \33826 , \33825 );
or \U$33581 ( \33827 , \33819 , \33826 );
not \U$33582 ( \33828 , \33814 );
nand \U$33583 ( \33829 , \33828 , \33813 );
nand \U$33584 ( \33830 , \33827 , \33829 );
not \U$33585 ( \33831 , \33830 );
or \U$33586 ( \33832 , \33807 , \33831 );
not \U$33587 ( \33833 , \33802 );
nand \U$33588 ( \33834 , \33833 , \33796 );
nand \U$33589 ( \33835 , \33832 , \33834 );
and \U$33590 ( \33836 , \33791 , \33835 );
not \U$33591 ( \33837 , \33791 );
not \U$33592 ( \33838 , \33835 );
and \U$33593 ( \33839 , \33837 , \33838 );
nor \U$33594 ( \33840 , \33836 , \33839 );
not \U$33595 ( \33841 , \33840 );
or \U$33596 ( \33842 , \33785 , \33841 );
not \U$33597 ( \33843 , \33838 );
nand \U$33598 ( \33844 , \33843 , \33791 );
nand \U$33599 ( \33845 , \33842 , \33844 );
not \U$33600 ( \33846 , \33845 );
not \U$33601 ( \33847 , \33846 );
or \U$33602 ( \33848 , \33699 , \33847 );
or \U$33603 ( \33849 , \33846 , \33698 );
nand \U$33604 ( \33850 , \33848 , \33849 );
not \U$33605 ( \33851 , \33850 );
or \U$33606 ( \33852 , \33687 , \33851 );
not \U$33607 ( \33853 , \33846 );
nand \U$33608 ( \33854 , \33853 , \33698 );
nand \U$33609 ( \33855 , \33852 , \33854 );
not \U$33610 ( \33856 , \33855 );
xor \U$33611 ( \33857 , \33423 , \33345 );
not \U$33612 ( \33858 , \33857 );
not \U$33613 ( \33859 , \33858 );
not \U$33614 ( \33860 , \33251 );
not \U$33615 ( \33861 , \33232 );
and \U$33616 ( \33862 , \33860 , \33861 );
and \U$33617 ( \33863 , \33251 , \33232 );
nor \U$33618 ( \33864 , \33862 , \33863 );
not \U$33619 ( \33865 , \33864 );
not \U$33620 ( \33866 , \33865 );
or \U$33621 ( \33867 , \33859 , \33866 );
nand \U$33622 ( \33868 , \33864 , \33857 );
nand \U$33623 ( \33869 , \33867 , \33868 );
not \U$33624 ( \33870 , \33869 );
or \U$33625 ( \33871 , \33856 , \33870 );
not \U$33626 ( \33872 , \33858 );
nand \U$33627 ( \33873 , \33872 , \33865 );
nand \U$33628 ( \33874 , \33871 , \33873 );
xor \U$33629 ( \33875 , \33256 , \33429 );
or \U$33630 ( \33876 , \33874 , \33875 );
xor \U$33631 ( \33877 , \33629 , \33435 );
nand \U$33632 ( \33878 , \33876 , \33877 );
nand \U$33633 ( \33879 , \33874 , \33875 );
nand \U$33634 ( \33880 , \33878 , \33879 );
nand \U$33635 ( \33881 , \33648 , \33880 );
nand \U$33636 ( \33882 , \33641 , \33881 );
nand \U$33637 ( \33883 , \33640 , \33882 );
not \U$33638 ( \33884 , \33883 );
or \U$33639 ( \33885 , \33224 , \33884 );
nor \U$33640 ( \33886 , \33059 , \33181 );
not \U$33641 ( \33887 , \33886 );
nand \U$33642 ( \33888 , \33885 , \33887 );
not \U$33643 ( \33889 , \31885 );
not \U$33644 ( \33890 , \31560 );
and \U$33645 ( \33891 , \33889 , \33890 );
and \U$33646 ( \33892 , \31885 , \31560 );
nor \U$33647 ( \33893 , \33891 , \33892 );
not \U$33648 ( \33894 , \33893 );
buf \U$33649 ( \33895 , \31296 );
not \U$33650 ( \33896 , \31271 );
and \U$33651 ( \33897 , \33895 , \33896 );
not \U$33652 ( \33898 , \33895 );
and \U$33653 ( \33899 , \33898 , \31271 );
nor \U$33654 ( \33900 , \33897 , \33899 );
not \U$33655 ( \33901 , \33900 );
xor \U$33656 ( \33902 , \31571 , \31618 );
not \U$33657 ( \33903 , \33902 );
not \U$33658 ( \33904 , \33107 );
not \U$33659 ( \33905 , \33904 );
not \U$33660 ( \33906 , \33115 );
or \U$33661 ( \33907 , \33905 , \33906 );
not \U$33662 ( \33908 , \33108 );
nand \U$33663 ( \33909 , \33908 , \33111 );
nand \U$33664 ( \33910 , \33907 , \33909 );
not \U$33665 ( \33911 , \33910 );
not \U$33666 ( \33912 , \33911 );
xnor \U$33667 ( \33913 , \31816 , \31852 );
not \U$33668 ( \33914 , \33913 );
and \U$33669 ( \33915 , \33912 , \33914 );
not \U$33670 ( \33916 , \33910 );
and \U$33671 ( \33917 , \33916 , \33913 );
nor \U$33672 ( \33918 , \33915 , \33917 );
not \U$33673 ( \33919 , \33918 );
not \U$33674 ( \33920 , \33919 );
and \U$33675 ( \33921 , \31809 , \31629 );
not \U$33676 ( \33922 , \31809 );
and \U$33677 ( \33923 , \33922 , \31630 );
or \U$33678 ( \33924 , \33921 , \33923 );
not \U$33679 ( \33925 , \33924 );
or \U$33680 ( \33926 , \33920 , \33925 );
nand \U$33681 ( \33927 , \33910 , \33913 );
nand \U$33682 ( \33928 , \33926 , \33927 );
not \U$33683 ( \33929 , \33928 );
not \U$33684 ( \33930 , \31814 );
not \U$33685 ( \33931 , \33930 );
not \U$33686 ( \33932 , \31863 );
or \U$33687 ( \33933 , \33931 , \33932 );
or \U$33688 ( \33934 , \31863 , \33930 );
nand \U$33689 ( \33935 , \33933 , \33934 );
not \U$33690 ( \33936 , \33935 );
not \U$33691 ( \33937 , \33936 );
or \U$33692 ( \33938 , \33929 , \33937 );
not \U$33693 ( \33939 , \33928 );
nand \U$33694 ( \33940 , \33939 , \33935 );
nand \U$33695 ( \33941 , \33938 , \33940 );
not \U$33696 ( \33942 , \33941 );
or \U$33697 ( \33943 , \33903 , \33942 );
nand \U$33698 ( \33944 , \33935 , \33928 );
nand \U$33699 ( \33945 , \33943 , \33944 );
buf \U$33700 ( \33946 , \33945 );
not \U$33701 ( \33947 , \33946 );
not \U$33702 ( \33948 , \33947 );
or \U$33703 ( \33949 , \33901 , \33948 );
not \U$33704 ( \33950 , \31623 );
and \U$33705 ( \33951 , \31876 , \33950 );
not \U$33706 ( \33952 , \31876 );
and \U$33707 ( \33953 , \33952 , \31623 );
nor \U$33708 ( \33954 , \33951 , \33953 );
not \U$33709 ( \33955 , \33954 );
nand \U$33710 ( \33956 , \33949 , \33955 );
not \U$33711 ( \33957 , \33900 );
nand \U$33712 ( \33958 , \33957 , \33946 );
nand \U$33713 ( \33959 , \33956 , \33958 );
not \U$33714 ( \33960 , \33959 );
nand \U$33715 ( \33961 , \33894 , \33960 );
xor \U$33716 ( \33962 , \33900 , \33945 );
xnor \U$33717 ( \33963 , \33962 , \33954 );
not \U$33718 ( \33964 , \33094 );
not \U$33719 ( \33965 , \33076 );
or \U$33720 ( \33966 , \33964 , \33965 );
not \U$33721 ( \33967 , \33074 );
nand \U$33722 ( \33968 , \33967 , \33067 );
nand \U$33723 ( \33969 , \33966 , \33968 );
not \U$33724 ( \33970 , \33969 );
not \U$33725 ( \33971 , \33918 );
not \U$33726 ( \33972 , \33924 );
and \U$33727 ( \33973 , \33971 , \33972 );
and \U$33728 ( \33974 , \33924 , \33918 );
nor \U$33729 ( \33975 , \33973 , \33974 );
not \U$33730 ( \33976 , \33154 );
not \U$33731 ( \33977 , \33128 );
or \U$33732 ( \33978 , \33976 , \33977 );
nand \U$33733 ( \33979 , \33116 , \33107 );
not \U$33734 ( \33980 , \33979 );
not \U$33735 ( \33981 , \33116 );
nand \U$33736 ( \33982 , \33981 , \33904 );
not \U$33737 ( \33983 , \33982 );
or \U$33738 ( \33984 , \33980 , \33983 );
nand \U$33739 ( \33985 , \33984 , \33127 );
nand \U$33740 ( \33986 , \33978 , \33985 );
not \U$33741 ( \33987 , \33986 );
and \U$33742 ( \33988 , \33975 , \33987 );
not \U$33743 ( \33989 , \33975 );
and \U$33744 ( \33990 , \33989 , \33986 );
nor \U$33745 ( \33991 , \33988 , \33990 );
not \U$33746 ( \33992 , \33991 );
or \U$33747 ( \33993 , \33970 , \33992 );
not \U$33748 ( \33994 , \33975 );
nand \U$33749 ( \33995 , \33994 , \33986 );
nand \U$33750 ( \33996 , \33993 , \33995 );
and \U$33751 ( \33997 , \31603 , \31592 );
not \U$33752 ( \33998 , \31603 );
and \U$33753 ( \33999 , \33998 , \31591 );
nor \U$33754 ( \34000 , \33997 , \33999 );
xor \U$33755 ( \34001 , \34000 , \31605 );
not \U$33756 ( \34002 , \34001 );
not \U$33757 ( \34003 , \34002 );
not \U$33758 ( \34004 , \33132 );
not \U$33759 ( \34005 , \33150 );
or \U$33760 ( \34006 , \34004 , \34005 );
not \U$33761 ( \34007 , \33138 );
nand \U$33762 ( \34008 , \34007 , \33145 );
nand \U$33763 ( \34009 , \34006 , \34008 );
not \U$33764 ( \34010 , \33078 );
not \U$33765 ( \34011 , \33093 );
or \U$33766 ( \34012 , \34010 , \34011 );
not \U$33767 ( \34013 , \33089 );
nand \U$33768 ( \34014 , \34013 , \33086 );
nand \U$33769 ( \34015 , \34012 , \34014 );
xor \U$33770 ( \34016 , \34009 , \34015 );
not \U$33771 ( \34017 , \34016 );
or \U$33772 ( \34018 , \34003 , \34017 );
nand \U$33773 ( \34019 , \34015 , \34009 );
nand \U$33774 ( \34020 , \34018 , \34019 );
or \U$33775 ( \34021 , \33996 , \34020 );
and \U$33776 ( \34022 , \33941 , \33902 );
not \U$33777 ( \34023 , \33941 );
not \U$33778 ( \34024 , \33902 );
and \U$33779 ( \34025 , \34023 , \34024 );
nor \U$33780 ( \34026 , \34022 , \34025 );
nand \U$33781 ( \34027 , \34021 , \34026 );
nand \U$33782 ( \34028 , \33996 , \34020 );
and \U$33783 ( \34029 , \34027 , \34028 );
nand \U$33784 ( \34030 , \33963 , \34029 );
xor \U$33785 ( \34031 , \34020 , \33996 );
xnor \U$33786 ( \34032 , \34031 , \34026 );
not \U$33787 ( \34033 , \33969 );
and \U$33788 ( \34034 , \33991 , \34033 );
not \U$33789 ( \34035 , \33991 );
and \U$33790 ( \34036 , \34035 , \33969 );
nor \U$33791 ( \34037 , \34034 , \34036 );
or \U$33792 ( \34038 , \33168 , \33164 );
nand \U$33793 ( \34039 , \34038 , \33159 );
nand \U$33794 ( \34040 , \33168 , \33164 );
nand \U$33795 ( \34041 , \34039 , \34040 );
not \U$33796 ( \34042 , \34041 );
nand \U$33797 ( \34043 , \34037 , \34042 );
not \U$33798 ( \34044 , \34016 );
not \U$33799 ( \34045 , \34001 );
and \U$33800 ( \34046 , \34044 , \34045 );
and \U$33801 ( \34047 , \34016 , \34001 );
nor \U$33802 ( \34048 , \34046 , \34047 );
not \U$33803 ( \34049 , \34048 );
and \U$33804 ( \34050 , \34043 , \34049 );
nor \U$33805 ( \34051 , \34037 , \34042 );
nor \U$33806 ( \34052 , \34050 , \34051 );
nand \U$33807 ( \34053 , \34032 , \34052 );
not \U$33808 ( \34054 , \34049 );
not \U$33809 ( \34055 , \34042 );
or \U$33810 ( \34056 , \34054 , \34055 );
nand \U$33811 ( \34057 , \34048 , \34041 );
nand \U$33812 ( \34058 , \34056 , \34057 );
not \U$33813 ( \34059 , \34037 );
and \U$33814 ( \34060 , \34058 , \34059 );
not \U$33815 ( \34061 , \34058 );
and \U$33816 ( \34062 , \34061 , \34037 );
nor \U$33817 ( \34063 , \34060 , \34062 );
not \U$33818 ( \34064 , \34063 );
not \U$33819 ( \34065 , \33173 );
not \U$33820 ( \34066 , \33099 );
not \U$33821 ( \34067 , \33179 );
or \U$33822 ( \34068 , \34066 , \34067 );
or \U$33823 ( \34069 , \33179 , \33099 );
nand \U$33824 ( \34070 , \34068 , \34069 );
nand \U$33825 ( \34071 , \34065 , \34070 );
nand \U$33826 ( \34072 , \33180 , \33100 );
nand \U$33827 ( \34073 , \34064 , \34071 , \34072 );
and \U$33828 ( \34074 , \34030 , \34053 , \34073 );
nand \U$33829 ( \34075 , \33961 , \34074 );
or \U$33830 ( \34076 , \33888 , \34075 );
not \U$33831 ( \34077 , \34072 );
not \U$33832 ( \34078 , \34071 );
or \U$33833 ( \34079 , \34077 , \34078 );
nand \U$33834 ( \34080 , \34079 , \34063 );
not \U$33835 ( \34081 , \34080 );
nand \U$33836 ( \34082 , \34081 , \34053 );
not \U$33837 ( \34083 , \34032 );
not \U$33838 ( \34084 , \34052 );
nand \U$33839 ( \34085 , \34083 , \34084 );
nand \U$33840 ( \34086 , \34082 , \34085 );
nand \U$33841 ( \34087 , \34086 , \34030 );
nand \U$33842 ( \34088 , \33893 , \33959 );
or \U$33843 ( \34089 , \33963 , \34029 );
nand \U$33844 ( \34090 , \34087 , \34088 , \34089 );
nand \U$33845 ( \34091 , \34090 , \33961 );
nand \U$33846 ( \34092 , \34076 , \34091 );
not \U$33847 ( \34093 , \34092 );
or \U$33848 ( \34094 , \31903 , \34093 );
buf \U$33849 ( \34095 , \31232 );
not \U$33850 ( \34096 , \34095 );
nor \U$33851 ( \34097 , \31558 , \31890 );
nand \U$33852 ( \34098 , \34097 , \31901 );
not \U$33853 ( \34099 , \30931 );
not \U$33854 ( \34100 , \31231 );
nand \U$33855 ( \34101 , \34099 , \34100 );
not \U$33856 ( \34102 , \31893 );
nand \U$33857 ( \34103 , \34102 , \31899 );
nand \U$33858 ( \34104 , \34098 , \34101 , \34103 );
not \U$33859 ( \34105 , \34104 );
or \U$33860 ( \34106 , \34096 , \34105 );
or \U$33861 ( \34107 , \30570 , \30925 );
nand \U$33862 ( \34108 , \34106 , \34107 );
buf \U$33863 ( \34109 , \30926 );
nand \U$33864 ( \34110 , \34108 , \34109 );
nand \U$33865 ( \34111 , \34094 , \34110 );
buf \U$33866 ( \34112 , \25194 );
xor \U$33867 ( \34113 , \25202 , \25188 );
xor \U$33868 ( \34114 , \34112 , \34113 );
not \U$33869 ( \34115 , \34114 );
not \U$33870 ( \34116 , \29890 );
not \U$33871 ( \34117 , \29875 );
or \U$33872 ( \34118 , \34116 , \34117 );
nand \U$33873 ( \34119 , \29884 , \29877 );
nand \U$33874 ( \34120 , \34118 , \34119 );
not \U$33875 ( \34121 , \34120 );
not \U$33876 ( \34122 , \34121 );
or \U$33877 ( \34123 , \34115 , \34122 );
not \U$33878 ( \34124 , \34120 );
or \U$33879 ( \34125 , \34124 , \34114 );
nand \U$33880 ( \34126 , \34123 , \34125 );
and \U$33881 ( \34127 , \24417 , \24404 );
not \U$33882 ( \34128 , \24417 );
and \U$33883 ( \34129 , \34128 , \24418 );
nor \U$33884 ( \34130 , \34127 , \34129 );
xnor \U$33885 ( \34131 , \34130 , \24415 );
not \U$33886 ( \34132 , \25005 );
not \U$33887 ( \34133 , \25166 );
or \U$33888 ( \34134 , \34132 , \34133 );
or \U$33889 ( \34135 , \25166 , \25005 );
nand \U$33890 ( \34136 , \34134 , \34135 );
xor \U$33891 ( \34137 , \34131 , \34136 );
not \U$33892 ( \34138 , \29867 );
not \U$33893 ( \34139 , \34138 );
not \U$33894 ( \34140 , \29830 );
or \U$33895 ( \34141 , \34139 , \34140 );
not \U$33896 ( \34142 , \29764 );
or \U$33897 ( \34143 , \29871 , \34142 );
nand \U$33898 ( \34144 , \34141 , \34143 );
xor \U$33899 ( \34145 , \34137 , \34144 );
xor \U$33900 ( \34146 , \34126 , \34145 );
not \U$33901 ( \34147 , \30564 );
not \U$33902 ( \34148 , \30559 );
or \U$33903 ( \34149 , \34147 , \34148 );
and \U$33904 ( \34150 , \30551 , \30535 );
not \U$33905 ( \34151 , \30551 );
not \U$33906 ( \34152 , \30535 );
and \U$33907 ( \34153 , \34151 , \34152 );
or \U$33908 ( \34154 , \34150 , \34153 );
nand \U$33909 ( \34155 , \34154 , \30558 );
nand \U$33910 ( \34156 , \34149 , \34155 );
xor \U$33911 ( \34157 , \34146 , \34156 );
not \U$33912 ( \34158 , \30514 );
not \U$33913 ( \34159 , \30517 );
or \U$33914 ( \34160 , \34158 , \34159 );
nand \U$33915 ( \34161 , \34160 , \30530 );
nand \U$33916 ( \34162 , \30518 , \30521 );
nand \U$33917 ( \34163 , \34161 , \34162 );
not \U$33918 ( \34164 , \34163 );
not \U$33919 ( \34165 , \34164 );
nor \U$33920 ( \34166 , \29368 , \29394 );
or \U$33921 ( \34167 , \34166 , \29366 );
nand \U$33922 ( \34168 , \29368 , \29394 );
nand \U$33923 ( \34169 , \34167 , \34168 );
not \U$33924 ( \34170 , \34169 );
or \U$33925 ( \34171 , \34165 , \34170 );
or \U$33926 ( \34172 , \34169 , \34164 );
nand \U$33927 ( \34173 , \34171 , \34172 );
not \U$33928 ( \34174 , \34173 );
xnor \U$33929 ( \34175 , \25219 , \25305 );
not \U$33930 ( \34176 , \34175 );
and \U$33931 ( \34177 , \34174 , \34176 );
and \U$33932 ( \34178 , \34175 , \34173 );
nor \U$33933 ( \34179 , \34177 , \34178 );
not \U$33934 ( \34180 , \34179 );
not \U$33935 ( \34181 , \34152 );
not \U$33936 ( \34182 , \30551 );
or \U$33937 ( \34183 , \34181 , \34182 );
not \U$33938 ( \34184 , \30540 );
nand \U$33939 ( \34185 , \34184 , \30546 );
nand \U$33940 ( \34186 , \34183 , \34185 );
not \U$33941 ( \34187 , \34186 );
or \U$33942 ( \34188 , \34180 , \34187 );
or \U$33943 ( \34189 , \34186 , \34179 );
nand \U$33944 ( \34190 , \34188 , \34189 );
buf \U$33945 ( \34191 , \34190 );
or \U$33946 ( \34192 , \29744 , \29895 );
not \U$33947 ( \34193 , \29395 );
nand \U$33948 ( \34194 , \34193 , \29740 );
nand \U$33949 ( \34195 , \34192 , \34194 );
not \U$33950 ( \34196 , \34195 );
and \U$33951 ( \34197 , \34191 , \34196 );
not \U$33952 ( \34198 , \34191 );
and \U$33953 ( \34199 , \34198 , \34195 );
nor \U$33954 ( \34200 , \34197 , \34199 );
not \U$33955 ( \34201 , \34200 );
and \U$33956 ( \34202 , \34157 , \34201 );
and \U$33957 ( \34203 , \34146 , \34156 );
nor \U$33958 ( \34204 , \34202 , \34203 );
not \U$33959 ( \34205 , \34195 );
not \U$33960 ( \34206 , \34190 );
or \U$33961 ( \34207 , \34205 , \34206 );
not \U$33962 ( \34208 , \34179 );
nand \U$33963 ( \34209 , \34208 , \34186 );
nand \U$33964 ( \34210 , \34207 , \34209 );
not \U$33965 ( \34211 , \34210 );
xor \U$33966 ( \34212 , \25172 , \25003 );
xnor \U$33967 ( \34213 , \34212 , \25171 );
not \U$33968 ( \34214 , \34213 );
xor \U$33969 ( \34215 , \23903 , \23900 );
xnor \U$33970 ( \34216 , \34215 , \23980 );
not \U$33971 ( \34217 , \34216 );
xor \U$33972 ( \34218 , \34131 , \34136 );
and \U$33973 ( \34219 , \34218 , \34144 );
and \U$33974 ( \34220 , \34131 , \34136 );
or \U$33975 ( \34221 , \34219 , \34220 );
not \U$33976 ( \34222 , \34221 );
or \U$33977 ( \34223 , \34217 , \34222 );
or \U$33978 ( \34224 , \34221 , \34216 );
nand \U$33979 ( \34225 , \34223 , \34224 );
not \U$33980 ( \34226 , \34225 );
and \U$33981 ( \34227 , \34214 , \34226 );
and \U$33982 ( \34228 , \34225 , \34213 );
nor \U$33983 ( \34229 , \34227 , \34228 );
not \U$33984 ( \34230 , \34229 );
and \U$33985 ( \34231 , \34211 , \34230 );
and \U$33986 ( \34232 , \34210 , \34229 );
nor \U$33987 ( \34233 , \34231 , \34232 );
not \U$33988 ( \34234 , \34145 );
not \U$33989 ( \34235 , \34126 );
or \U$33990 ( \34236 , \34234 , \34235 );
not \U$33991 ( \34237 , \34124 );
nand \U$33992 ( \34238 , \34237 , \34114 );
nand \U$33993 ( \34239 , \34236 , \34238 );
not \U$33994 ( \34240 , \25204 );
and \U$33995 ( \34241 , \25309 , \34240 );
not \U$33996 ( \34242 , \25309 );
and \U$33997 ( \34243 , \34242 , \25204 );
nor \U$33998 ( \34244 , \34241 , \34243 );
buf \U$33999 ( \34245 , \25206 );
xor \U$34000 ( \34246 , \34244 , \34245 );
not \U$34001 ( \34247 , \34246 );
not \U$34002 ( \34248 , \34247 );
not \U$34003 ( \34249 , \34175 );
not \U$34004 ( \34250 , \34249 );
not \U$34005 ( \34251 , \34173 );
or \U$34006 ( \34252 , \34250 , \34251 );
not \U$34007 ( \34253 , \34164 );
nand \U$34008 ( \34254 , \34253 , \34169 );
nand \U$34009 ( \34255 , \34252 , \34254 );
not \U$34010 ( \34256 , \34255 );
not \U$34011 ( \34257 , \34256 );
or \U$34012 ( \34258 , \34248 , \34257 );
nand \U$34013 ( \34259 , \34246 , \34255 );
nand \U$34014 ( \34260 , \34258 , \34259 );
xor \U$34015 ( \34261 , \34239 , \34260 );
xor \U$34016 ( \34262 , \34233 , \34261 );
nand \U$34017 ( \34263 , \34204 , \34262 );
not \U$34018 ( \34264 , \34213 );
not \U$34019 ( \34265 , \34264 );
not \U$34020 ( \34266 , \34225 );
or \U$34021 ( \34267 , \34265 , \34266 );
not \U$34022 ( \34268 , \34216 );
nand \U$34023 ( \34269 , \34268 , \34221 );
nand \U$34024 ( \34270 , \34267 , \34269 );
not \U$34025 ( \34271 , \34239 );
not \U$34026 ( \34272 , \34260 );
or \U$34027 ( \34273 , \34271 , \34272 );
nand \U$34028 ( \34274 , \34255 , \34247 );
nand \U$34029 ( \34275 , \34273 , \34274 );
xor \U$34030 ( \34276 , \34270 , \34275 );
xor \U$34031 ( \34277 , \25368 , \25375 );
xor \U$34032 ( \34278 , \34276 , \34277 );
not \U$34033 ( \34279 , \34261 );
not \U$34034 ( \34280 , \34233 );
not \U$34035 ( \34281 , \34280 );
or \U$34036 ( \34282 , \34279 , \34281 );
not \U$34037 ( \34283 , \34229 );
nand \U$34038 ( \34284 , \34283 , \34210 );
nand \U$34039 ( \34285 , \34282 , \34284 );
nor \U$34040 ( \34286 , \34278 , \34285 );
xor \U$34041 ( \34287 , \34270 , \34275 );
and \U$34042 ( \34288 , \34287 , \34277 );
and \U$34043 ( \34289 , \34270 , \34275 );
or \U$34044 ( \34290 , \34288 , \34289 );
xor \U$34045 ( \34291 , \25355 , \25380 );
xor \U$34046 ( \34292 , \34291 , \25382 );
nor \U$34047 ( \34293 , \34290 , \34292 );
nor \U$34048 ( \34294 , \34286 , \34293 );
xor \U$34049 ( \34295 , \34157 , \34200 );
not \U$34050 ( \34296 , \29900 );
xor \U$34051 ( \34297 , \34296 , \30506 );
and \U$34052 ( \34298 , \34297 , \30569 );
and \U$34053 ( \34299 , \34296 , \30506 );
nor \U$34054 ( \34300 , \34298 , \34299 );
nand \U$34055 ( \34301 , \34295 , \34300 );
and \U$34056 ( \34302 , \34263 , \34294 , \34301 );
nand \U$34057 ( \34303 , \34111 , \34302 );
nor \U$34058 ( \34304 , \33648 , \33880 );
nor \U$34059 ( \34305 , \33886 , \34304 );
and \U$34060 ( \34306 , \33961 , \34074 , \33640 , \34305 );
and \U$34061 ( \34307 , \34306 , \31902 );
and \U$34062 ( \34308 , \34263 , \34301 );
not \U$34063 ( \34309 , \17059 );
xnor \U$34064 ( \34310 , RIbe2a3e8_88, RIbe2a7a8_96);
not \U$34065 ( \34311 , \34310 );
and \U$34066 ( \34312 , \34309 , \34311 );
xor \U$34067 ( \34313 , RIbe2a3e8_88, RIbe2abe0_105);
and \U$34068 ( \34314 , \11541 , \34313 );
nor \U$34069 ( \34315 , \34312 , \34314 );
not \U$34070 ( \34316 , \34315 );
not \U$34071 ( \34317 , \34316 );
xor \U$34072 ( \34318 , RIbe2a910_99, RIbe2ac58_106);
not \U$34073 ( \34319 , \34318 );
not \U$34074 ( \34320 , \9737 );
or \U$34075 ( \34321 , \34319 , \34320 );
xor \U$34076 ( \34322 , RIbe2a640_93, RIbe2a910_99);
nand \U$34077 ( \34323 , \10400 , \34322 );
nand \U$34078 ( \34324 , \34321 , \34323 );
not \U$34079 ( \34325 , \34324 );
not \U$34080 ( \34326 , \34325 );
xor \U$34081 ( \34327 , RIbe2a028_80, RIbe2aeb0_111);
not \U$34082 ( \34328 , \34327 );
not \U$34083 ( \34329 , \8400 );
or \U$34084 ( \34330 , \34328 , \34329 );
xor \U$34085 ( \34331 , RIbe2a028_80, RIbe2b3d8_122);
nand \U$34086 ( \34332 , \8930 , \34331 );
nand \U$34087 ( \34333 , \34330 , \34332 );
not \U$34088 ( \34334 , \34333 );
or \U$34089 ( \34335 , \34326 , \34334 );
not \U$34090 ( \34336 , \34324 );
or \U$34091 ( \34337 , \34333 , \34336 );
nand \U$34092 ( \34338 , \34335 , \34337 );
not \U$34093 ( \34339 , \34338 );
or \U$34094 ( \34340 , \34317 , \34339 );
nand \U$34095 ( \34341 , \34333 , \34324 );
nand \U$34096 ( \34342 , \34340 , \34341 );
not \U$34097 ( \34343 , \34342 );
not \U$34098 ( \34344 , \34331 );
not \U$34099 ( \34345 , \8169 );
or \U$34100 ( \34346 , \34344 , \34345 );
nand \U$34101 ( \34347 , \9065 , \33808 );
nand \U$34102 ( \34348 , \34346 , \34347 );
not \U$34103 ( \34349 , \34348 );
or \U$34104 ( \34350 , RIbe2a028_80, RIbe29fb0_79);
nand \U$34105 ( \34351 , \34350 , RIbe2ae38_110);
nand \U$34106 ( \34352 , RIbe29fb0_79, RIbe2a028_80);
nand \U$34107 ( \34353 , \34351 , \34352 , RIbe29e48_76);
not \U$34108 ( \34354 , \34353 );
and \U$34109 ( \34355 , \34349 , \34354 );
and \U$34110 ( \34356 , \34348 , \34353 );
nor \U$34111 ( \34357 , \34355 , \34356 );
not \U$34112 ( \34358 , \34357 );
and \U$34113 ( \34359 , RIbe2a190_83, RIbe2b540_125);
nor \U$34114 ( \34360 , RIbe2a190_83, RIbe2b540_125);
nor \U$34115 ( \34361 , \34359 , \34360 );
not \U$34116 ( \34362 , \34361 );
not \U$34117 ( \34363 , \10690 );
or \U$34118 ( \34364 , \34362 , \34363 );
xor \U$34119 ( \34365 , RIbe2a190_83, RIbe2ad48_108);
nand \U$34120 ( \34366 , \13278 , \34365 );
nand \U$34121 ( \34367 , \34364 , \34366 );
not \U$34122 ( \34368 , \34367 );
not \U$34123 ( \34369 , \34368 );
xor \U$34124 ( \34370 , RIbe2af28_112, RIbe2a118_82);
not \U$34125 ( \34371 , \34370 );
not \U$34126 ( \34372 , \15345 );
or \U$34127 ( \34373 , \34371 , \34372 );
not \U$34128 ( \34374 , \14414 );
xor \U$34129 ( \34375 , RIbe2af28_112, RIbe2a820_97);
nand \U$34130 ( \34376 , \34374 , \34375 );
nand \U$34131 ( \34377 , \34373 , \34376 );
not \U$34132 ( \34378 , \34377 );
not \U$34133 ( \34379 , \34378 );
or \U$34134 ( \34380 , \34369 , \34379 );
xor \U$34135 ( \34381 , RIbe2adc0_109, RIbe2a280_85);
not \U$34136 ( \34382 , \34381 );
not \U$34137 ( \34383 , \20237 );
or \U$34138 ( \34384 , \34382 , \34383 );
xor \U$34139 ( \34385 , RIbe2a460_89, RIbe2a280_85);
nand \U$34140 ( \34386 , \11348 , \34385 );
nand \U$34141 ( \34387 , \34384 , \34386 );
nand \U$34142 ( \34388 , \34380 , \34387 );
nand \U$34143 ( \34389 , \34367 , \34377 );
nand \U$34144 ( \34390 , \34388 , \34389 );
not \U$34145 ( \34391 , \34390 );
or \U$34146 ( \34392 , \34358 , \34391 );
or \U$34147 ( \34393 , \34390 , \34357 );
nand \U$34148 ( \34394 , \34392 , \34393 );
not \U$34149 ( \34395 , \34394 );
or \U$34150 ( \34396 , \34343 , \34395 );
not \U$34151 ( \34397 , \34357 );
nand \U$34152 ( \34398 , \34397 , \34390 );
nand \U$34153 ( \34399 , \34396 , \34398 );
not \U$34154 ( \34400 , \34399 );
not \U$34155 ( \34401 , \34385 );
not \U$34156 ( \34402 , \24028 );
or \U$34157 ( \34403 , \34401 , \34402 );
nand \U$34158 ( \34404 , \11348 , \33748 );
nand \U$34159 ( \34405 , \34403 , \34404 );
not \U$34160 ( \34406 , \34405 );
xor \U$34161 ( \34407 , RIbe2b2e8_120, RIbe2b108_116);
not \U$34162 ( \34408 , \34407 );
not \U$34163 ( \34409 , \25618 );
or \U$34164 ( \34410 , \34408 , \34409 );
xor \U$34165 ( \34411 , RIbe2b108_116, RIbe2b360_121);
nand \U$34166 ( \34412 , \13534 , \34411 );
nand \U$34167 ( \34413 , \34410 , \34412 );
not \U$34168 ( \34414 , \34413 );
not \U$34169 ( \34415 , \34414 );
or \U$34170 ( \34416 , \34406 , \34415 );
not \U$34171 ( \34417 , \34405 );
nand \U$34172 ( \34418 , \34417 , \34413 );
nand \U$34173 ( \34419 , \34416 , \34418 );
not \U$34174 ( \34420 , \34322 );
not \U$34175 ( \34421 , \10987 );
or \U$34176 ( \34422 , \34420 , \34421 );
nand \U$34177 ( \34423 , \11456 , \33734 );
nand \U$34178 ( \34424 , \34422 , \34423 );
and \U$34179 ( \34425 , \34419 , \34424 );
not \U$34180 ( \34426 , \34419 );
not \U$34181 ( \34427 , \34424 );
and \U$34182 ( \34428 , \34426 , \34427 );
nor \U$34183 ( \34429 , \34425 , \34428 );
not \U$34184 ( \34430 , \34429 );
xor \U$34185 ( \34431 , RIbe2aa78_102, RIbe2aaf0_103);
not \U$34186 ( \34432 , \34431 );
not \U$34187 ( \34433 , \20574 );
or \U$34188 ( \34434 , \34432 , \34433 );
xor \U$34189 ( \34435 , RIbe2aaf0_103, RIbe2b6a8_128);
nand \U$34190 ( \34436 , \34435 , RIbe2ab68_104);
nand \U$34191 ( \34437 , \34434 , \34436 );
not \U$34192 ( \34438 , \34437 );
xor \U$34193 ( \34439 , RIbe2b108_116, RIbe2a4d8_90);
not \U$34194 ( \34440 , \34439 );
not \U$34195 ( \34441 , \14297 );
or \U$34196 ( \34442 , \34440 , \34441 );
nand \U$34197 ( \34443 , \16898 , \34407 );
nand \U$34198 ( \34444 , \34442 , \34443 );
not \U$34199 ( \34445 , \34444 );
or \U$34200 ( \34446 , \34438 , \34445 );
or \U$34201 ( \34447 , \34444 , \34437 );
xor \U$34202 ( \34448 , RIbe2a6b8_94, RIbe2a550_91);
not \U$34203 ( \34449 , \34448 );
not \U$34204 ( \34450 , \10433 );
or \U$34205 ( \34451 , \34449 , \34450 );
xor \U$34206 ( \34452 , RIbe2a550_91, RIbe2b4c8_124);
nand \U$34207 ( \34453 , \15995 , \34452 );
nand \U$34208 ( \34454 , \34451 , \34453 );
nand \U$34209 ( \34455 , \34447 , \34454 );
nand \U$34210 ( \34456 , \34446 , \34455 );
not \U$34211 ( \34457 , RIbe2a898_98);
not \U$34212 ( \34458 , RIbe2b018_114);
and \U$34213 ( \34459 , \34457 , \34458 );
and \U$34214 ( \34460 , RIbe2a898_98, RIbe2b018_114);
nor \U$34215 ( \34461 , \34459 , \34460 );
not \U$34216 ( \34462 , \34461 );
not \U$34217 ( \34463 , \16812 );
or \U$34218 ( \34464 , \34462 , \34463 );
xor \U$34219 ( \34465 , RIbe2b018_114, RIbe2aa00_101);
nand \U$34220 ( \34466 , \20583 , \34465 );
nand \U$34221 ( \34467 , \34464 , \34466 );
not \U$34222 ( \34468 , \34467 );
xor \U$34223 ( \34469 , RIbe2a2f8_86, RIbe2b450_123);
not \U$34224 ( \34470 , \34469 );
not \U$34225 ( \34471 , \9374 );
or \U$34226 ( \34472 , \34470 , \34471 );
xor \U$34227 ( \34473 , RIbe2a2f8_86, RIbe2a730_95);
nand \U$34228 ( \34474 , \8705 , \34473 );
nand \U$34229 ( \34475 , \34472 , \34474 );
not \U$34230 ( \34476 , \34475 );
not \U$34231 ( \34477 , \34476 );
nand \U$34232 ( \34478 , \4849 , RIbe2ae38_110);
not \U$34233 ( \34479 , \34478 );
not \U$34234 ( \34480 , \34479 );
or \U$34235 ( \34481 , \34477 , \34480 );
nand \U$34236 ( \34482 , \34475 , \34478 );
nand \U$34237 ( \34483 , \34481 , \34482 );
not \U$34238 ( \34484 , \34483 );
or \U$34239 ( \34485 , \34468 , \34484 );
nand \U$34240 ( \34486 , \34479 , \34475 );
nand \U$34241 ( \34487 , \34485 , \34486 );
xor \U$34242 ( \34488 , \34456 , \34487 );
not \U$34243 ( \34489 , \34488 );
or \U$34244 ( \34490 , \34430 , \34489 );
nand \U$34245 ( \34491 , \34487 , \34456 );
nand \U$34246 ( \34492 , \34490 , \34491 );
not \U$34247 ( \34493 , \34492 );
nand \U$34248 ( \34494 , \34400 , \34493 );
nand \U$34249 ( \34495 , \34399 , \34492 );
nand \U$34250 ( \34496 , \34494 , \34495 );
not \U$34251 ( \34497 , \34375 );
not \U$34252 ( \34498 , \16913 );
or \U$34253 ( \34499 , \34497 , \34498 );
nand \U$34254 ( \34500 , \14413 , \33700 );
nand \U$34255 ( \34501 , \34499 , \34500 );
xor \U$34256 ( \34502 , RIbe2a0a0_81, RIbe2b180_117);
not \U$34257 ( \34503 , \34502 );
not \U$34258 ( \34504 , \14852 );
or \U$34259 ( \34505 , \34503 , \34504 );
nand \U$34260 ( \34506 , \16646 , \33720 );
nand \U$34261 ( \34507 , \34505 , \34506 );
xor \U$34262 ( \34508 , \34501 , \34507 );
not \U$34263 ( \34509 , \34473 );
not \U$34264 ( \34510 , \8989 );
or \U$34265 ( \34511 , \34509 , \34510 );
nand \U$34266 ( \34512 , \11094 , \33758 );
nand \U$34267 ( \34513 , \34511 , \34512 );
xor \U$34268 ( \34514 , \34508 , \34513 );
not \U$34269 ( \34515 , \34514 );
xor \U$34270 ( \34516 , RIbe29e48_76, RIbe2ae38_110);
not \U$34271 ( \34517 , \34516 );
not \U$34272 ( \34518 , \9252 );
or \U$34273 ( \34519 , \34517 , \34518 );
nand \U$34274 ( \34520 , \4851 , \33765 );
nand \U$34275 ( \34521 , \34519 , \34520 );
not \U$34276 ( \34522 , \34521 );
not \U$34277 ( \34523 , \34522 );
not \U$34278 ( \34524 , \34313 );
not \U$34279 ( \34525 , \8806 );
or \U$34280 ( \34526 , \34524 , \34525 );
nand \U$34281 ( \34527 , \10476 , \33771 );
nand \U$34282 ( \34528 , \34526 , \34527 );
not \U$34283 ( \34529 , \34365 );
not \U$34284 ( \34530 , \17563 );
or \U$34285 ( \34531 , \34529 , \34530 );
nand \U$34286 ( \34532 , \13278 , \33820 );
nand \U$34287 ( \34533 , \34531 , \34532 );
not \U$34288 ( \34534 , \34533 );
xnor \U$34289 ( \34535 , \34528 , \34534 );
not \U$34290 ( \34536 , \34535 );
or \U$34291 ( \34537 , \34523 , \34536 );
or \U$34292 ( \34538 , \34535 , \34522 );
nand \U$34293 ( \34539 , \34537 , \34538 );
not \U$34294 ( \34540 , \34539 );
not \U$34295 ( \34541 , \34452 );
not \U$34296 ( \34542 , \12000 );
or \U$34297 ( \34543 , \34541 , \34542 );
nand \U$34298 ( \34544 , \11485 , \33707 );
nand \U$34299 ( \34545 , \34543 , \34544 );
xor \U$34300 ( \34546 , RIbe2aaf0_103, RIbe29f38_78);
not \U$34301 ( \34547 , \34546 );
not \U$34302 ( \34548 , RIbe2ab68_104);
or \U$34303 ( \34549 , \34547 , \34548 );
buf \U$34304 ( \34550 , \19580 );
not \U$34305 ( \34551 , \34435 );
or \U$34306 ( \34552 , \34550 , \34551 );
nand \U$34307 ( \34553 , \34549 , \34552 );
nor \U$34308 ( \34554 , \34545 , \34553 );
not \U$34309 ( \34555 , \34554 );
nand \U$34310 ( \34556 , \34545 , \34553 );
nand \U$34311 ( \34557 , \34555 , \34556 );
not \U$34312 ( \34558 , \17571 );
not \U$34313 ( \34559 , \34558 );
not \U$34314 ( \34560 , \34465 );
not \U$34315 ( \34561 , \34560 );
and \U$34316 ( \34562 , \34559 , \34561 );
buf \U$34317 ( \34563 , \15953 );
and \U$34318 ( \34564 , \34563 , \33740 );
nor \U$34319 ( \34565 , \34562 , \34564 );
not \U$34320 ( \34566 , \34565 );
and \U$34321 ( \34567 , \34557 , \34566 );
not \U$34322 ( \34568 , \34557 );
and \U$34323 ( \34569 , \34568 , \34565 );
nor \U$34324 ( \34570 , \34567 , \34569 );
not \U$34325 ( \34571 , \34570 );
or \U$34326 ( \34572 , \34540 , \34571 );
or \U$34327 ( \34573 , \34570 , \34539 );
nand \U$34328 ( \34574 , \34572 , \34573 );
not \U$34329 ( \34575 , \34574 );
or \U$34330 ( \34576 , \34515 , \34575 );
not \U$34331 ( \34577 , \34570 );
nand \U$34332 ( \34578 , \34577 , \34539 );
nand \U$34333 ( \34579 , \34576 , \34578 );
buf \U$34334 ( \34580 , \34579 );
xor \U$34335 ( \34581 , \34496 , \34580 );
not \U$34336 ( \34582 , \34581 );
xnor \U$34337 ( \34583 , \34488 , \34429 );
not \U$34338 ( \34584 , \34583 );
not \U$34339 ( \34585 , \34584 );
xor \U$34340 ( \34586 , RIbe2b180_117, RIbe2b360_121);
not \U$34341 ( \34587 , \34586 );
not \U$34342 ( \34588 , \14853 );
not \U$34343 ( \34589 , \34588 );
or \U$34344 ( \34590 , \34587 , \34589 );
nand \U$34345 ( \34591 , \14966 , \34502 );
nand \U$34346 ( \34592 , \34590 , \34591 );
xor \U$34347 ( \34593 , RIbe2b3d8_122, RIbe2a2f8_86);
not \U$34348 ( \34594 , \34593 );
not \U$34349 ( \34595 , \8989 );
or \U$34350 ( \34596 , \34594 , \34595 );
nand \U$34351 ( \34597 , \9379 , \34469 );
nand \U$34352 ( \34598 , \34596 , \34597 );
not \U$34353 ( \34599 , \8162 );
nand \U$34354 ( \34600 , \34599 , RIbe2ae38_110);
nand \U$34355 ( \34601 , RIbe2a2f8_86, RIbe2acd0_107);
and \U$34356 ( \34602 , \34601 , RIbe2a028_80);
and \U$34357 ( \34603 , \34600 , \34602 );
and \U$34358 ( \34604 , \34598 , \34603 );
xor \U$34359 ( \34605 , \34592 , \34604 );
xor \U$34360 ( \34606 , RIbe2aa00_101, RIbe2aaf0_103);
not \U$34361 ( \34607 , \34606 );
not \U$34362 ( \34608 , \19580 );
not \U$34363 ( \34609 , \34608 );
or \U$34364 ( \34610 , \34607 , \34609 );
nand \U$34365 ( \34611 , \34431 , RIbe2ab68_104);
nand \U$34366 ( \34612 , \34610 , \34611 );
not \U$34367 ( \34613 , \34612 );
xor \U$34368 ( \34614 , RIbe2a3e8_88, RIbe2a730_95);
not \U$34369 ( \34615 , \34614 );
not \U$34370 ( \34616 , \9263 );
or \U$34371 ( \34617 , \34615 , \34616 );
not \U$34372 ( \34618 , \34310 );
nand \U$34373 ( \34619 , \34618 , \9268 );
nand \U$34374 ( \34620 , \34617 , \34619 );
not \U$34375 ( \34621 , \34620 );
or \U$34376 ( \34622 , \34613 , \34621 );
not \U$34377 ( \34623 , \34612 );
not \U$34378 ( \34624 , \34623 );
not \U$34379 ( \34625 , \34620 );
not \U$34380 ( \34626 , \34625 );
or \U$34381 ( \34627 , \34624 , \34626 );
xor \U$34382 ( \34628 , RIbe2a0a0_81, RIbe2af28_112);
not \U$34383 ( \34629 , \34628 );
not \U$34384 ( \34630 , \15345 );
or \U$34385 ( \34631 , \34629 , \34630 );
nand \U$34386 ( \34632 , \17811 , \34370 );
nand \U$34387 ( \34633 , \34631 , \34632 );
nand \U$34388 ( \34634 , \34627 , \34633 );
nand \U$34389 ( \34635 , \34622 , \34634 );
and \U$34390 ( \34636 , \34605 , \34635 );
and \U$34391 ( \34637 , \34592 , \34604 );
nor \U$34392 ( \34638 , \34636 , \34637 );
not \U$34393 ( \34639 , \34638 );
xor \U$34394 ( \34640 , RIbe2ad48_108, RIbe2a280_85);
not \U$34395 ( \34641 , \34640 );
not \U$34396 ( \34642 , \24028 );
or \U$34397 ( \34643 , \34641 , \34642 );
nand \U$34398 ( \34644 , \11348 , \34381 );
nand \U$34399 ( \34645 , \34643 , \34644 );
xor \U$34400 ( \34646 , RIbe2b108_116, RIbe2a460_89);
not \U$34401 ( \34647 , \34646 );
not \U$34402 ( \34648 , \25617 );
or \U$34403 ( \34649 , \34647 , \34648 );
nand \U$34404 ( \34650 , \23015 , \34439 );
nand \U$34405 ( \34651 , \34649 , \34650 );
nor \U$34406 ( \34652 , \34645 , \34651 );
and \U$34407 ( \34653 , \31948 , \34361 );
and \U$34408 ( \34654 , RIbe2a190_83, RIbe2b4c8_124);
nor \U$34409 ( \34655 , RIbe2a190_83, RIbe2b4c8_124);
nor \U$34410 ( \34656 , \34654 , \34655 );
not \U$34411 ( \34657 , \34656 );
not \U$34412 ( \34658 , \10690 );
nor \U$34413 ( \34659 , \34657 , \34658 );
nor \U$34414 ( \34660 , \34653 , \34659 );
or \U$34415 ( \34661 , \34652 , \34660 );
nand \U$34416 ( \34662 , \34645 , \34651 );
nand \U$34417 ( \34663 , \34661 , \34662 );
not \U$34418 ( \34664 , \34663 );
not \U$34419 ( \34665 , \34664 );
xor \U$34420 ( \34666 , \34437 , \34454 );
xnor \U$34421 ( \34667 , \34666 , \34444 );
not \U$34422 ( \34668 , \34667 );
or \U$34423 ( \34669 , \34665 , \34668 );
not \U$34424 ( \34670 , RIbe2a820_97);
not \U$34425 ( \34671 , RIbe2b018_114);
and \U$34426 ( \34672 , \34670 , \34671 );
and \U$34427 ( \34673 , RIbe2a820_97, RIbe2b018_114);
nor \U$34428 ( \34674 , \34672 , \34673 );
not \U$34429 ( \34675 , \34674 );
not \U$34430 ( \34676 , \17571 );
or \U$34431 ( \34677 , \34675 , \34676 );
nand \U$34432 ( \34678 , \20583 , \34461 );
nand \U$34433 ( \34679 , \34677 , \34678 );
not \U$34434 ( \34680 , \34679 );
xor \U$34435 ( \34681 , RIbe2a028_80, RIbe2ae38_110);
not \U$34436 ( \34682 , \34681 );
not \U$34437 ( \34683 , \9530 );
or \U$34438 ( \34684 , \34682 , \34683 );
nand \U$34439 ( \34685 , \8930 , \34327 );
nand \U$34440 ( \34686 , \34684 , \34685 );
not \U$34441 ( \34687 , \34686 );
or \U$34442 ( \34688 , \34680 , \34687 );
xor \U$34443 ( \34689 , RIbe2a910_99, RIbe2abe0_105);
and \U$34444 ( \34690 , \34689 , \10987 );
and \U$34445 ( \34691 , \10401 , \34318 );
nor \U$34446 ( \34692 , \34690 , \34691 );
nand \U$34447 ( \34693 , \34688 , \34692 );
not \U$34448 ( \34694 , \34686 );
not \U$34449 ( \34695 , \34679 );
nand \U$34450 ( \34696 , \34694 , \34695 );
nand \U$34451 ( \34697 , \34693 , \34696 );
not \U$34452 ( \34698 , \34697 );
nand \U$34453 ( \34699 , \34669 , \34698 );
not \U$34454 ( \34700 , \34667 );
nand \U$34455 ( \34701 , \34700 , \34663 );
nand \U$34456 ( \34702 , \34699 , \34701 );
not \U$34457 ( \34703 , \34702 );
or \U$34458 ( \34704 , \34639 , \34703 );
or \U$34459 ( \34705 , \34702 , \34638 );
nand \U$34460 ( \34706 , \34704 , \34705 );
not \U$34461 ( \34707 , \34706 );
or \U$34462 ( \34708 , \34585 , \34707 );
not \U$34463 ( \34709 , \34638 );
nand \U$34464 ( \34710 , \34709 , \34702 );
nand \U$34465 ( \34711 , \34708 , \34710 );
not \U$34466 ( \34712 , \34711 );
xor \U$34467 ( \34713 , \34514 , \34574 );
not \U$34468 ( \34714 , \34713 );
not \U$34469 ( \34715 , \34394 );
not \U$34470 ( \34716 , \34342 );
not \U$34471 ( \34717 , \34716 );
and \U$34472 ( \34718 , \34715 , \34717 );
and \U$34473 ( \34719 , \34394 , \34716 );
nor \U$34474 ( \34720 , \34718 , \34719 );
not \U$34475 ( \34721 , \34720 );
xor \U$34476 ( \34722 , \34368 , \34387 );
xnor \U$34477 ( \34723 , \34722 , \34377 );
not \U$34478 ( \34724 , \34723 );
not \U$34479 ( \34725 , \34338 );
not \U$34480 ( \34726 , \34315 );
and \U$34481 ( \34727 , \34725 , \34726 );
and \U$34482 ( \34728 , \34338 , \34315 );
nor \U$34483 ( \34729 , \34727 , \34728 );
not \U$34484 ( \34730 , \34483 );
not \U$34485 ( \34731 , \34467 );
not \U$34486 ( \34732 , \34731 );
and \U$34487 ( \34733 , \34730 , \34732 );
and \U$34488 ( \34734 , \34483 , \34731 );
nor \U$34489 ( \34735 , \34733 , \34734 );
and \U$34490 ( \34736 , \34729 , \34735 );
not \U$34491 ( \34737 , \34729 );
not \U$34492 ( \34738 , \34735 );
and \U$34493 ( \34739 , \34737 , \34738 );
nor \U$34494 ( \34740 , \34736 , \34739 );
not \U$34495 ( \34741 , \34740 );
or \U$34496 ( \34742 , \34724 , \34741 );
or \U$34497 ( \34743 , \34735 , \34729 );
nand \U$34498 ( \34744 , \34742 , \34743 );
not \U$34499 ( \34745 , \34744 );
or \U$34500 ( \34746 , \34721 , \34745 );
or \U$34501 ( \34747 , \34744 , \34720 );
nand \U$34502 ( \34748 , \34746 , \34747 );
not \U$34503 ( \34749 , \34748 );
or \U$34504 ( \34750 , \34714 , \34749 );
not \U$34505 ( \34751 , \34720 );
nand \U$34506 ( \34752 , \34751 , \34744 );
nand \U$34507 ( \34753 , \34750 , \34752 );
not \U$34508 ( \34754 , \34753 );
not \U$34509 ( \34755 , \34754 );
or \U$34510 ( \34756 , \34712 , \34755 );
not \U$34511 ( \34757 , \34711 );
nand \U$34512 ( \34758 , \34757 , \34753 );
nand \U$34513 ( \34759 , \34756 , \34758 );
not \U$34514 ( \34760 , \34759 );
or \U$34515 ( \34761 , \34582 , \34760 );
or \U$34516 ( \34762 , \34759 , \34581 );
nand \U$34517 ( \34763 , \34761 , \34762 );
xor \U$34518 ( \34764 , \33725 , \33712 );
xor \U$34519 ( \34765 , \34764 , \33705 );
not \U$34520 ( \34766 , \34765 );
not \U$34521 ( \34767 , \34766 );
or \U$34522 ( \34768 , \34554 , \34565 );
nand \U$34523 ( \34769 , \34768 , \34556 );
not \U$34524 ( \34770 , \34769 );
xor \U$34525 ( \34771 , \33818 , \33825 );
not \U$34526 ( \34772 , \34771 );
not \U$34527 ( \34773 , \34772 );
or \U$34528 ( \34774 , \34770 , \34773 );
not \U$34529 ( \34775 , \34769 );
nand \U$34530 ( \34776 , \34775 , \34771 );
nand \U$34531 ( \34777 , \34774 , \34776 );
not \U$34532 ( \34778 , \34777 );
or \U$34533 ( \34779 , \34767 , \34778 );
or \U$34534 ( \34780 , \34777 , \34766 );
nand \U$34535 ( \34781 , \34779 , \34780 );
and \U$34536 ( \34782 , \33777 , \33763 );
not \U$34537 ( \34783 , \33777 );
not \U$34538 ( \34784 , \33763 );
and \U$34539 ( \34785 , \34783 , \34784 );
nor \U$34540 ( \34786 , \34782 , \34785 );
not \U$34541 ( \34787 , \33747 );
nand \U$34542 ( \34788 , \34787 , \33753 );
not \U$34543 ( \34789 , \34788 );
not \U$34544 ( \34790 , \33751 );
and \U$34545 ( \34791 , \34789 , \34790 );
and \U$34546 ( \34792 , \34788 , \33751 );
nor \U$34547 ( \34793 , \34791 , \34792 );
xor \U$34548 ( \34794 , \34786 , \34793 );
not \U$34549 ( \34795 , \34546 );
or \U$34550 ( \34796 , \34550 , \34795 );
not \U$34551 ( \34797 , \33581 );
or \U$34552 ( \34798 , \18830 , \34797 );
nand \U$34553 ( \34799 , \34796 , \34798 );
not \U$34554 ( \34800 , \34411 );
not \U$34555 ( \34801 , \13543 );
or \U$34556 ( \34802 , \34800 , \34801 );
nand \U$34557 ( \34803 , \13534 , \33492 );
nand \U$34558 ( \34804 , \34802 , \34803 );
xor \U$34559 ( \34805 , \34799 , \34804 );
not \U$34560 ( \34806 , \34348 );
nor \U$34561 ( \34807 , \34806 , \34353 );
xor \U$34562 ( \34808 , \34805 , \34807 );
xor \U$34563 ( \34809 , \34794 , \34808 );
not \U$34564 ( \34810 , \34533 );
not \U$34565 ( \34811 , \34528 );
or \U$34566 ( \34812 , \34810 , \34811 );
not \U$34567 ( \34813 , \34528 );
nand \U$34568 ( \34814 , \34813 , \34534 );
nand \U$34569 ( \34815 , \34814 , \34521 );
nand \U$34570 ( \34816 , \34812 , \34815 );
not \U$34571 ( \34817 , \34513 );
not \U$34572 ( \34818 , \34501 );
or \U$34573 ( \34819 , \34817 , \34818 );
or \U$34574 ( \34820 , \34501 , \34513 );
nand \U$34575 ( \34821 , \34820 , \34507 );
nand \U$34576 ( \34822 , \34819 , \34821 );
not \U$34577 ( \34823 , \34822 );
and \U$34578 ( \34824 , \34816 , \34823 );
not \U$34579 ( \34825 , \34816 );
and \U$34580 ( \34826 , \34825 , \34822 );
or \U$34581 ( \34827 , \34824 , \34826 );
not \U$34582 ( \34828 , \34424 );
not \U$34583 ( \34829 , \34405 );
or \U$34584 ( \34830 , \34828 , \34829 );
or \U$34585 ( \34831 , \34405 , \34424 );
nand \U$34586 ( \34832 , \34831 , \34413 );
nand \U$34587 ( \34833 , \34830 , \34832 );
and \U$34588 ( \34834 , \34827 , \34833 );
not \U$34589 ( \34835 , \34827 );
not \U$34590 ( \34836 , \34833 );
and \U$34591 ( \34837 , \34835 , \34836 );
nor \U$34592 ( \34838 , \34834 , \34837 );
not \U$34593 ( \34839 , \34838 );
and \U$34594 ( \34840 , \34809 , \34839 );
not \U$34595 ( \34841 , \34809 );
and \U$34596 ( \34842 , \34841 , \34838 );
nor \U$34597 ( \34843 , \34840 , \34842 );
xor \U$34598 ( \34844 , \34781 , \34843 );
not \U$34599 ( \34845 , \34844 );
or \U$34600 ( \34846 , \34763 , \34845 );
and \U$34601 ( \34847 , RIbe2af28_112, RIbe2b360_121);
not \U$34602 ( \34848 , RIbe2af28_112);
and \U$34603 ( \34849 , \34848 , \26908 );
nor \U$34604 ( \34850 , \34847 , \34849 );
not \U$34605 ( \34851 , \34850 );
not \U$34606 ( \34852 , \16914 );
or \U$34607 ( \34853 , \34851 , \34852 );
nand \U$34608 ( \34854 , \15348 , \34628 );
nand \U$34609 ( \34855 , \34853 , \34854 );
not \U$34610 ( \34856 , \34855 );
xor \U$34611 ( \34857 , RIbe2b180_117, RIbe2a4d8_90);
not \U$34612 ( \34858 , \34857 );
not \U$34613 ( \34859 , \15353 );
or \U$34614 ( \34860 , \34858 , \34859 );
xor \U$34615 ( \34861 , RIbe2b180_117, RIbe2b2e8_120);
nand \U$34616 ( \34862 , \16646 , \34861 );
nand \U$34617 ( \34863 , \34860 , \34862 );
not \U$34618 ( \34864 , \34863 );
xor \U$34619 ( \34865 , RIbe2a6b8_94, RIbe2a190_83);
not \U$34620 ( \34866 , \34865 );
not \U$34621 ( \34867 , \17563 );
or \U$34622 ( \34868 , \34866 , \34867 );
nand \U$34623 ( \34869 , \13278 , \34656 );
nand \U$34624 ( \34870 , \34868 , \34869 );
not \U$34625 ( \34871 , \34870 );
not \U$34626 ( \34872 , \34871 );
or \U$34627 ( \34873 , \34864 , \34872 );
or \U$34628 ( \34874 , \34871 , \34863 );
nand \U$34629 ( \34875 , \34873 , \34874 );
not \U$34630 ( \34876 , \34875 );
or \U$34631 ( \34877 , \34856 , \34876 );
nand \U$34632 ( \34878 , \34870 , \34863 );
nand \U$34633 ( \34879 , \34877 , \34878 );
xor \U$34634 ( \34880 , RIbe2a910_99, RIbe2a7a8_96);
not \U$34635 ( \34881 , \34880 );
not \U$34636 ( \34882 , \12715 );
or \U$34637 ( \34883 , \34881 , \34882 );
nand \U$34638 ( \34884 , \10400 , \34689 );
nand \U$34639 ( \34885 , \34883 , \34884 );
xor \U$34640 ( \34886 , RIbe2aeb0_111, RIbe2a2f8_86);
not \U$34641 ( \34887 , \34886 );
not \U$34642 ( \34888 , \9374 );
or \U$34643 ( \34889 , \34887 , \34888 );
nand \U$34644 ( \34890 , \8705 , \34593 );
nand \U$34645 ( \34891 , \34889 , \34890 );
nor \U$34646 ( \34892 , \34885 , \34891 );
xor \U$34647 ( \34893 , RIbe2ac58_106, RIbe2a550_91);
and \U$34648 ( \34894 , \10434 , \34893 );
xnor \U$34649 ( \34895 , RIbe2a640_93, RIbe2a550_91);
nor \U$34650 ( \34896 , \23307 , \34895 );
nor \U$34651 ( \34897 , \34894 , \34896 );
or \U$34652 ( \34898 , \34892 , \34897 );
nand \U$34653 ( \34899 , \34885 , \34891 );
nand \U$34654 ( \34900 , \34898 , \34899 );
not \U$34655 ( \34901 , \34900 );
not \U$34656 ( \34902 , RIbe2a118_82);
not \U$34657 ( \34903 , RIbe2b018_114);
and \U$34658 ( \34904 , \34902 , \34903 );
and \U$34659 ( \34905 , RIbe2a118_82, RIbe2b018_114);
nor \U$34660 ( \34906 , \34904 , \34905 );
not \U$34661 ( \34907 , \34906 );
not \U$34662 ( \34908 , \22763 );
or \U$34663 ( \34909 , \34907 , \34908 );
nand \U$34664 ( \34910 , \20583 , \34674 );
nand \U$34665 ( \34911 , \34909 , \34910 );
not \U$34666 ( \34912 , \34911 );
xor \U$34667 ( \34913 , RIbe2a3e8_88, RIbe2b450_123);
not \U$34668 ( \34914 , \34913 );
not \U$34669 ( \34915 , \8806 );
or \U$34670 ( \34916 , \34914 , \34915 );
nand \U$34671 ( \34917 , \8794 , \34614 );
nand \U$34672 ( \34918 , \34916 , \34917 );
nand \U$34673 ( \34919 , \8172 , RIbe2ae38_110);
not \U$34674 ( \34920 , \34919 );
and \U$34675 ( \34921 , \34918 , \34920 );
not \U$34676 ( \34922 , \34918 );
and \U$34677 ( \34923 , \34922 , \34919 );
nor \U$34678 ( \34924 , \34921 , \34923 );
not \U$34679 ( \34925 , \34924 );
or \U$34680 ( \34926 , \34912 , \34925 );
nand \U$34681 ( \34927 , \34918 , \34920 );
nand \U$34682 ( \34928 , \34926 , \34927 );
not \U$34683 ( \34929 , \34928 );
not \U$34684 ( \34930 , \34929 );
or \U$34685 ( \34931 , \34901 , \34930 );
or \U$34686 ( \34932 , \34900 , \34929 );
nand \U$34687 ( \34933 , \34931 , \34932 );
and \U$34688 ( \34934 , \34879 , \34933 );
and \U$34689 ( \34935 , \34928 , \34900 );
nor \U$34690 ( \34936 , \34934 , \34935 );
not \U$34691 ( \34937 , \34603 );
and \U$34692 ( \34938 , \34598 , \34937 );
not \U$34693 ( \34939 , \34598 );
and \U$34694 ( \34940 , \34939 , \34603 );
nor \U$34695 ( \34941 , \34938 , \34940 );
not \U$34696 ( \34942 , \34941 );
not \U$34697 ( \34943 , \34942 );
not \U$34698 ( \34944 , \34861 );
not \U$34699 ( \34945 , \14852 );
or \U$34700 ( \34946 , \34944 , \34945 );
nand \U$34701 ( \34947 , \14966 , \34586 );
nand \U$34702 ( \34948 , \34946 , \34947 );
not \U$34703 ( \34949 , \34948 );
not \U$34704 ( \34950 , \34895 );
not \U$34705 ( \34951 , \34950 );
not \U$34706 ( \34952 , \22975 );
or \U$34707 ( \34953 , \34951 , \34952 );
nand \U$34708 ( \34954 , \11228 , \34448 );
nand \U$34709 ( \34955 , \34953 , \34954 );
not \U$34710 ( \34956 , \34955 );
not \U$34711 ( \34957 , \34956 );
or \U$34712 ( \34958 , \34949 , \34957 );
or \U$34713 ( \34959 , \34948 , \34956 );
nand \U$34714 ( \34960 , \34958 , \34959 );
not \U$34715 ( \34961 , \34960 );
or \U$34716 ( \34962 , \34943 , \34961 );
nand \U$34717 ( \34963 , \34955 , \34948 );
nand \U$34718 ( \34964 , \34962 , \34963 );
not \U$34719 ( \34965 , \34964 );
not \U$34720 ( \34966 , \34965 );
xor \U$34721 ( \34967 , \34605 , \34635 );
not \U$34722 ( \34968 , \34967 );
and \U$34723 ( \34969 , \34966 , \34968 );
and \U$34724 ( \34970 , \34965 , \34967 );
nor \U$34725 ( \34971 , \34969 , \34970 );
or \U$34726 ( \34972 , \34936 , \34971 );
nand \U$34727 ( \34973 , \34964 , \34967 );
nand \U$34728 ( \34974 , \34972 , \34973 );
not \U$34729 ( \34975 , \34583 );
not \U$34730 ( \34976 , \34706 );
or \U$34731 ( \34977 , \34975 , \34976 );
or \U$34732 ( \34978 , \34706 , \34583 );
nand \U$34733 ( \34979 , \34977 , \34978 );
xor \U$34734 ( \34980 , \34974 , \34979 );
not \U$34735 ( \34981 , \34633 );
not \U$34736 ( \34982 , \34612 );
not \U$34737 ( \34983 , \34625 );
or \U$34738 ( \34984 , \34982 , \34983 );
or \U$34739 ( \34985 , \34625 , \34612 );
nand \U$34740 ( \34986 , \34984 , \34985 );
not \U$34741 ( \34987 , \34986 );
or \U$34742 ( \34988 , \34981 , \34987 );
or \U$34743 ( \34989 , \34986 , \34633 );
nand \U$34744 ( \34990 , \34988 , \34989 );
not \U$34745 ( \34991 , \34990 );
not \U$34746 ( \34992 , \34991 );
xor \U$34747 ( \34993 , RIbe2a898_98, RIbe2aaf0_103);
not \U$34748 ( \34994 , \34993 );
not \U$34749 ( \34995 , \34608 );
or \U$34750 ( \34996 , \34994 , \34995 );
nand \U$34751 ( \34997 , \34606 , RIbe2ab68_104);
nand \U$34752 ( \34998 , \34996 , \34997 );
xor \U$34753 ( \34999 , RIbe2b108_116, RIbe2adc0_109);
not \U$34754 ( \35000 , \34999 );
not \U$34755 ( \35001 , \25617 );
or \U$34756 ( \35002 , \35000 , \35001 );
nand \U$34757 ( \35003 , \13534 , \34646 );
nand \U$34758 ( \35004 , \35002 , \35003 );
xor \U$34759 ( \35005 , \34998 , \35004 );
not \U$34760 ( \35006 , RIbe2a280_85);
not \U$34761 ( \35007 , RIbe2b540_125);
and \U$34762 ( \35008 , \35006 , \35007 );
and \U$34763 ( \35009 , RIbe2a280_85, RIbe2b540_125);
nor \U$34764 ( \35010 , \35008 , \35009 );
and \U$34765 ( \35011 , \23047 , \35010 );
not \U$34766 ( \35012 , \34640 );
nor \U$34767 ( \35013 , \35012 , \10848 );
nor \U$34768 ( \35014 , \35011 , \35013 );
not \U$34769 ( \35015 , \35014 );
and \U$34770 ( \35016 , \35005 , \35015 );
and \U$34771 ( \35017 , \34998 , \35004 );
nor \U$34772 ( \35018 , \35016 , \35017 );
not \U$34773 ( \35019 , \35018 );
not \U$34774 ( \35020 , \35019 );
or \U$34775 ( \35021 , \34992 , \35020 );
not \U$34776 ( \35022 , \34990 );
not \U$34777 ( \35023 , \35018 );
or \U$34778 ( \35024 , \35022 , \35023 );
not \U$34779 ( \35025 , \34652 );
nand \U$34780 ( \35026 , \35025 , \34662 );
xor \U$34781 ( \35027 , \35026 , \34660 );
nand \U$34782 ( \35028 , \35024 , \35027 );
nand \U$34783 ( \35029 , \35021 , \35028 );
buf \U$34784 ( \35030 , \34667 );
not \U$34785 ( \35031 , \35030 );
not \U$34786 ( \35032 , \34663 );
not \U$34787 ( \35033 , \35032 );
not \U$34788 ( \35034 , \34698 );
or \U$34789 ( \35035 , \35033 , \35034 );
or \U$34790 ( \35036 , \35032 , \34698 );
nand \U$34791 ( \35037 , \35035 , \35036 );
not \U$34792 ( \35038 , \35037 );
or \U$34793 ( \35039 , \35031 , \35038 );
or \U$34794 ( \35040 , \35037 , \35030 );
nand \U$34795 ( \35041 , \35039 , \35040 );
xor \U$34796 ( \35042 , \35029 , \35041 );
xor \U$34797 ( \35043 , \34740 , \34723 );
and \U$34798 ( \35044 , \35042 , \35043 );
and \U$34799 ( \35045 , \35029 , \35041 );
or \U$34800 ( \35046 , \35044 , \35045 );
and \U$34801 ( \35047 , \34980 , \35046 );
and \U$34802 ( \35048 , \34974 , \34979 );
or \U$34803 ( \35049 , \35047 , \35048 );
nand \U$34804 ( \35050 , \34846 , \35049 );
nand \U$34805 ( \35051 , \34763 , \34845 );
nand \U$34806 ( \35052 , \35050 , \35051 );
xnor \U$34807 ( \35053 , \33830 , \33806 );
not \U$34808 ( \35054 , \35053 );
not \U$34809 ( \35055 , \35054 );
xor \U$34810 ( \35056 , \34799 , \34804 );
and \U$34811 ( \35057 , \35056 , \34807 );
and \U$34812 ( \35058 , \34799 , \34804 );
or \U$34813 ( \35059 , \35057 , \35058 );
not \U$34814 ( \35060 , \35059 );
xor \U$34815 ( \35061 , \33497 , \33481 );
xnor \U$34816 ( \35062 , \35061 , \33488 );
not \U$34817 ( \35063 , \35062 );
and \U$34818 ( \35064 , \35060 , \35063 );
and \U$34819 ( \35065 , \35059 , \35062 );
nor \U$34820 ( \35066 , \35064 , \35065 );
not \U$34821 ( \35067 , \35066 );
or \U$34822 ( \35068 , \35055 , \35067 );
or \U$34823 ( \35069 , \35066 , \35054 );
nand \U$34824 ( \35070 , \35068 , \35069 );
not \U$34825 ( \35071 , \33664 );
not \U$34826 ( \35072 , \33650 );
and \U$34827 ( \35073 , \35071 , \35072 );
and \U$34828 ( \35074 , \33664 , \33650 );
nor \U$34829 ( \35075 , \35073 , \35074 );
xor \U$34830 ( \35076 , \34786 , \34793 );
and \U$34831 ( \35077 , \35076 , \34808 );
and \U$34832 ( \35078 , \34786 , \34793 );
or \U$34833 ( \35079 , \35077 , \35078 );
not \U$34834 ( \35080 , \35079 );
and \U$34835 ( \35081 , \35075 , \35080 );
not \U$34836 ( \35082 , \35075 );
and \U$34837 ( \35083 , \35082 , \35079 );
nor \U$34838 ( \35084 , \35081 , \35083 );
buf \U$34839 ( \35085 , \35084 );
xor \U$34840 ( \35086 , \35070 , \35085 );
nand \U$34841 ( \35087 , \34494 , \34579 );
nand \U$34842 ( \35088 , \35087 , \34495 );
not \U$34843 ( \35089 , \35088 );
or \U$34844 ( \35090 , \34781 , \34838 );
nand \U$34845 ( \35091 , \35090 , \34809 );
nand \U$34846 ( \35092 , \34781 , \34838 );
nand \U$34847 ( \35093 , \35091 , \35092 );
not \U$34848 ( \35094 , \35093 );
not \U$34849 ( \35095 , \35094 );
or \U$34850 ( \35096 , \35089 , \35095 );
not \U$34851 ( \35097 , \35088 );
nand \U$34852 ( \35098 , \35097 , \35093 );
nand \U$34853 ( \35099 , \35096 , \35098 );
not \U$34854 ( \35100 , \34823 );
not \U$34855 ( \35101 , \34816 );
not \U$34856 ( \35102 , \35101 );
or \U$34857 ( \35103 , \35100 , \35102 );
nand \U$34858 ( \35104 , \35103 , \34833 );
nand \U$34859 ( \35105 , \34816 , \34822 );
nand \U$34860 ( \35106 , \35104 , \35105 );
not \U$34861 ( \35107 , \35106 );
xor \U$34862 ( \35108 , \33754 , \33728 );
xor \U$34863 ( \35109 , \35108 , \33781 );
xor \U$34864 ( \35110 , \35107 , \35109 );
not \U$34865 ( \35111 , \34765 );
not \U$34866 ( \35112 , \34777 );
or \U$34867 ( \35113 , \35111 , \35112 );
nand \U$34868 ( \35114 , \34771 , \34769 );
nand \U$34869 ( \35115 , \35113 , \35114 );
xnor \U$34870 ( \35116 , \35110 , \35115 );
and \U$34871 ( \35117 , \35099 , \35116 );
not \U$34872 ( \35118 , \35099 );
not \U$34873 ( \35119 , \35116 );
and \U$34874 ( \35120 , \35118 , \35119 );
nor \U$34875 ( \35121 , \35117 , \35120 );
xor \U$34876 ( \35122 , \35086 , \35121 );
not \U$34877 ( \35123 , \34581 );
nand \U$34878 ( \35124 , \35123 , \34759 );
nand \U$34879 ( \35125 , \34753 , \34711 );
nand \U$34880 ( \35126 , \35124 , \35125 );
xnor \U$34881 ( \35127 , \35122 , \35126 );
nor \U$34882 ( \35128 , \35052 , \35127 );
not \U$34883 ( \35129 , \34844 );
not \U$34884 ( \35130 , \35049 );
or \U$34885 ( \35131 , \35129 , \35130 );
or \U$34886 ( \35132 , \35049 , \34844 );
nand \U$34887 ( \35133 , \35131 , \35132 );
not \U$34888 ( \35134 , \35133 );
not \U$34889 ( \35135 , \34763 );
or \U$34890 ( \35136 , \35134 , \35135 );
or \U$34891 ( \35137 , \34763 , \35133 );
nand \U$34892 ( \35138 , \35136 , \35137 );
xor \U$34893 ( \35139 , \34748 , \34713 );
xor \U$34894 ( \35140 , \34974 , \34979 );
xor \U$34895 ( \35141 , \35140 , \35046 );
xor \U$34896 ( \35142 , \35139 , \35141 );
not \U$34897 ( \35143 , \34971 );
and \U$34898 ( \35144 , \34936 , \35143 );
not \U$34899 ( \35145 , \34936 );
and \U$34900 ( \35146 , \35145 , \34971 );
nor \U$34901 ( \35147 , \35144 , \35146 );
not \U$34902 ( \35148 , \35147 );
not \U$34903 ( \35149 , \35148 );
not \U$34904 ( \35150 , \34991 );
not \U$34905 ( \35151 , \35018 );
or \U$34906 ( \35152 , \35150 , \35151 );
nand \U$34907 ( \35153 , \35019 , \34990 );
nand \U$34908 ( \35154 , \35152 , \35153 );
xor \U$34909 ( \35155 , \35154 , \35027 );
not \U$34910 ( \35156 , \35155 );
not \U$34911 ( \35157 , \34875 );
not \U$34912 ( \35158 , \34855 );
not \U$34913 ( \35159 , \35158 );
and \U$34914 ( \35160 , \35157 , \35159 );
and \U$34915 ( \35161 , \34875 , \35158 );
nor \U$34916 ( \35162 , \35160 , \35161 );
and \U$34917 ( \35163 , RIbe2a730_95, RIbe2a910_99);
nor \U$34918 ( \35164 , RIbe2a730_95, RIbe2a910_99);
nor \U$34919 ( \35165 , \35163 , \35164 );
not \U$34920 ( \35166 , \35165 );
not \U$34921 ( \35167 , \13325 );
or \U$34922 ( \35168 , \35166 , \35167 );
nand \U$34923 ( \35169 , \10401 , \34880 );
nand \U$34924 ( \35170 , \35168 , \35169 );
not \U$34925 ( \35171 , \35170 );
xor \U$34926 ( \35172 , RIbe2b108_116, RIbe2ad48_108);
not \U$34927 ( \35173 , \35172 );
not \U$34928 ( \35174 , \14297 );
or \U$34929 ( \35175 , \35173 , \35174 );
nand \U$34930 ( \35176 , \13534 , \34999 );
nand \U$34931 ( \35177 , \35175 , \35176 );
not \U$34932 ( \35178 , \19580 );
xor \U$34933 ( \35179 , RIbe2a820_97, RIbe2aaf0_103);
and \U$34934 ( \35180 , \35178 , \35179 );
and \U$34935 ( \35181 , RIbe2ab68_104, \34993 );
nor \U$34936 ( \35182 , \35180 , \35181 );
nor \U$34937 ( \35183 , \35177 , \35182 );
not \U$34938 ( \35184 , \35183 );
nand \U$34939 ( \35185 , \35177 , \35182 );
nand \U$34940 ( \35186 , \35184 , \35185 );
not \U$34941 ( \35187 , \35186 );
or \U$34942 ( \35188 , \35171 , \35187 );
not \U$34943 ( \35189 , \35182 );
nand \U$34944 ( \35190 , \35189 , \35177 );
nand \U$34945 ( \35191 , \35188 , \35190 );
not \U$34946 ( \35192 , \35191 );
nand \U$34947 ( \35193 , \35162 , \35192 );
not \U$34948 ( \35194 , \34892 );
nand \U$34949 ( \35195 , \35194 , \34899 );
not \U$34950 ( \35196 , \34897 );
and \U$34951 ( \35197 , \35195 , \35196 );
not \U$34952 ( \35198 , \35195 );
and \U$34953 ( \35199 , \35198 , \34897 );
nor \U$34954 ( \35200 , \35197 , \35199 );
not \U$34955 ( \35201 , \35200 );
and \U$34956 ( \35202 , \35193 , \35201 );
nor \U$34957 ( \35203 , \35192 , \35162 );
nor \U$34958 ( \35204 , \35202 , \35203 );
not \U$34959 ( \35205 , \35204 );
not \U$34960 ( \35206 , \34879 );
not \U$34961 ( \35207 , \34933 );
not \U$34962 ( \35208 , \35207 );
or \U$34963 ( \35209 , \35206 , \35208 );
not \U$34964 ( \35210 , \34879 );
nand \U$34965 ( \35211 , \35210 , \34933 );
nand \U$34966 ( \35212 , \35209 , \35211 );
not \U$34967 ( \35213 , \35212 );
or \U$34968 ( \35214 , \35205 , \35213 );
or \U$34969 ( \35215 , \35212 , \35204 );
nand \U$34970 ( \35216 , \35214 , \35215 );
not \U$34971 ( \35217 , \35216 );
or \U$34972 ( \35218 , \35156 , \35217 );
not \U$34973 ( \35219 , \35204 );
nand \U$34974 ( \35220 , \35219 , \35212 );
nand \U$34975 ( \35221 , \35218 , \35220 );
not \U$34976 ( \35222 , \35221 );
not \U$34977 ( \35223 , \34686 );
not \U$34978 ( \35224 , \34692 );
or \U$34979 ( \35225 , \35223 , \35224 );
or \U$34980 ( \35226 , \34692 , \34686 );
nand \U$34981 ( \35227 , \35225 , \35226 );
xor \U$34982 ( \35228 , \35227 , \34695 );
not \U$34983 ( \35229 , \35228 );
not \U$34984 ( \35230 , \34942 );
not \U$34985 ( \35231 , \34960 );
not \U$34986 ( \35232 , \35231 );
or \U$34987 ( \35233 , \35230 , \35232 );
nand \U$34988 ( \35234 , \34960 , \34941 );
nand \U$34989 ( \35235 , \35233 , \35234 );
not \U$34990 ( \35236 , \35235 );
or \U$34991 ( \35237 , \35229 , \35236 );
or \U$34992 ( \35238 , \35235 , \35228 );
nand \U$34993 ( \35239 , \35237 , \35238 );
not \U$34994 ( \35240 , \35239 );
xor \U$34995 ( \35241 , RIbe2a2f8_86, RIbe2ae38_110);
not \U$34996 ( \35242 , \35241 );
not \U$34997 ( \35243 , \16715 );
or \U$34998 ( \35244 , \35242 , \35243 );
nand \U$34999 ( \35245 , \8706 , \34886 );
nand \U$35000 ( \35246 , \35244 , \35245 );
not \U$35001 ( \35247 , RIbe2a0a0_81);
not \U$35002 ( \35248 , RIbe2b018_114);
and \U$35003 ( \35249 , \35247 , \35248 );
and \U$35004 ( \35250 , RIbe2a0a0_81, RIbe2b018_114);
nor \U$35005 ( \35251 , \35249 , \35250 );
not \U$35006 ( \35252 , \35251 );
not \U$35007 ( \35253 , \17571 );
or \U$35008 ( \35254 , \35252 , \35253 );
nand \U$35009 ( \35255 , \34563 , \34906 );
nand \U$35010 ( \35256 , \35254 , \35255 );
xor \U$35011 ( \35257 , \35246 , \35256 );
not \U$35012 ( \35258 , \34893 );
not \U$35013 ( \35259 , \11228 );
or \U$35014 ( \35260 , \35258 , \35259 );
xnor \U$35015 ( \35261 , RIbe2abe0_105, RIbe2a550_91);
or \U$35016 ( \35262 , \15539 , \35261 );
nand \U$35017 ( \35263 , \35260 , \35262 );
and \U$35018 ( \35264 , \35257 , \35263 );
and \U$35019 ( \35265 , \35246 , \35256 );
or \U$35020 ( \35266 , \35264 , \35265 );
not \U$35021 ( \35267 , \35266 );
or \U$35022 ( \35268 , RIbe2a370_87, RIbe2a3e8_88);
nand \U$35023 ( \35269 , \35268 , RIbe2ae38_110);
nand \U$35024 ( \35270 , RIbe2a370_87, RIbe2a3e8_88);
and \U$35025 ( \35271 , \35269 , \35270 , RIbe2a2f8_86);
not \U$35026 ( \35272 , \8806 );
xor \U$35027 ( \35273 , RIbe2b3d8_122, RIbe2a3e8_88);
not \U$35028 ( \35274 , \35273 );
or \U$35029 ( \35275 , \35272 , \35274 );
nand \U$35030 ( \35276 , \11541 , \34913 );
nand \U$35031 ( \35277 , \35275 , \35276 );
and \U$35032 ( \35278 , \35271 , \35277 );
not \U$35033 ( \35279 , \35278 );
not \U$35034 ( \35280 , \15693 );
not \U$35035 ( \35281 , \34865 );
or \U$35036 ( \35282 , \35280 , \35281 );
not \U$35037 ( \35283 , \11973 );
and \U$35038 ( \35284 , RIbe2a190_83, RIbe2a640_93);
nor \U$35039 ( \35285 , RIbe2a190_83, RIbe2a640_93);
nor \U$35040 ( \35286 , \35284 , \35285 );
nand \U$35041 ( \35287 , \35283 , \35286 );
nand \U$35042 ( \35288 , \35282 , \35287 );
not \U$35043 ( \35289 , \35288 );
xor \U$35044 ( \35290 , RIbe2b180_117, RIbe2a460_89);
not \U$35045 ( \35291 , \35290 );
not \U$35046 ( \35292 , \14852 );
or \U$35047 ( \35293 , \35291 , \35292 );
nand \U$35048 ( \35294 , \16646 , \34857 );
nand \U$35049 ( \35295 , \35293 , \35294 );
xor \U$35050 ( \35296 , RIbe2a280_85, RIbe2b4c8_124);
not \U$35051 ( \35297 , \35296 );
not \U$35052 ( \35298 , \14942 );
or \U$35053 ( \35299 , \35297 , \35298 );
nand \U$35054 ( \35300 , \14649 , \35010 );
nand \U$35055 ( \35301 , \35299 , \35300 );
xor \U$35056 ( \35302 , \35295 , \35301 );
not \U$35057 ( \35303 , \35302 );
or \U$35058 ( \35304 , \35289 , \35303 );
nand \U$35059 ( \35305 , \35301 , \35295 );
nand \U$35060 ( \35306 , \35304 , \35305 );
not \U$35061 ( \35307 , \35306 );
not \U$35062 ( \35308 , \35307 );
or \U$35063 ( \35309 , \35279 , \35308 );
not \U$35064 ( \35310 , \35278 );
nand \U$35065 ( \35311 , \35310 , \35306 );
nand \U$35066 ( \35312 , \35309 , \35311 );
not \U$35067 ( \35313 , \35312 );
or \U$35068 ( \35314 , \35267 , \35313 );
nand \U$35069 ( \35315 , \35306 , \35278 );
nand \U$35070 ( \35316 , \35314 , \35315 );
not \U$35071 ( \35317 , \35316 );
or \U$35072 ( \35318 , \35240 , \35317 );
not \U$35073 ( \35319 , \35228 );
nand \U$35074 ( \35320 , \35319 , \35235 );
nand \U$35075 ( \35321 , \35318 , \35320 );
not \U$35076 ( \35322 , \35321 );
and \U$35077 ( \35323 , \35222 , \35322 );
not \U$35078 ( \35324 , \35222 );
and \U$35079 ( \35325 , \35324 , \35321 );
nor \U$35080 ( \35326 , \35323 , \35325 );
not \U$35081 ( \35327 , \35326 );
or \U$35082 ( \35328 , \35149 , \35327 );
nand \U$35083 ( \35329 , \35221 , \35321 );
nand \U$35084 ( \35330 , \35328 , \35329 );
and \U$35085 ( \35331 , \35142 , \35330 );
and \U$35086 ( \35332 , \35139 , \35141 );
or \U$35087 ( \35333 , \35331 , \35332 );
not \U$35088 ( \35334 , \35333 );
nand \U$35089 ( \35335 , \35138 , \35334 );
not \U$35090 ( \35336 , \35335 );
nor \U$35091 ( \35337 , \35128 , \35336 );
xor \U$35092 ( \35338 , \35029 , \35041 );
xor \U$35093 ( \35339 , \35338 , \35043 );
buf \U$35094 ( \35340 , \35216 );
and \U$35095 ( \35341 , \35340 , \35155 );
not \U$35096 ( \35342 , \35340 );
not \U$35097 ( \35343 , \35155 );
and \U$35098 ( \35344 , \35342 , \35343 );
nor \U$35099 ( \35345 , \35341 , \35344 );
not \U$35100 ( \35346 , \35345 );
buf \U$35101 ( \35347 , \34924 );
not \U$35102 ( \35348 , \34911 );
and \U$35103 ( \35349 , \35347 , \35348 );
not \U$35104 ( \35350 , \35347 );
and \U$35105 ( \35351 , \35350 , \34911 );
nor \U$35106 ( \35352 , \35349 , \35351 );
and \U$35107 ( \35353 , \35005 , \35014 );
not \U$35108 ( \35354 , \35005 );
and \U$35109 ( \35355 , \35354 , \35015 );
nor \U$35110 ( \35356 , \35353 , \35355 );
not \U$35111 ( \35357 , \35356 );
and \U$35112 ( \35358 , \35352 , \35357 );
not \U$35113 ( \35359 , \35352 );
and \U$35114 ( \35360 , \35359 , \35356 );
nor \U$35115 ( \35361 , \35358 , \35360 );
not \U$35116 ( \35362 , \35361 );
not \U$35117 ( \35363 , \35362 );
xor \U$35118 ( \35364 , RIbe2af28_112, RIbe2b2e8_120);
not \U$35119 ( \35365 , \35364 );
buf \U$35120 ( \35366 , \16913 );
not \U$35121 ( \35367 , \35366 );
or \U$35122 ( \35368 , \35365 , \35367 );
nand \U$35123 ( \35369 , \15348 , \34850 );
nand \U$35124 ( \35370 , \35368 , \35369 );
xor \U$35125 ( \35371 , \35271 , \35277 );
xor \U$35126 ( \35372 , \35370 , \35371 );
xor \U$35127 ( \35373 , RIbe2b450_123, RIbe2a910_99);
not \U$35128 ( \35374 , \35373 );
not \U$35129 ( \35375 , \15395 );
or \U$35130 ( \35376 , \35374 , \35375 );
nand \U$35131 ( \35377 , \10401 , \35165 );
nand \U$35132 ( \35378 , \35376 , \35377 );
not \U$35133 ( \35379 , \35378 );
xor \U$35134 ( \35380 , RIbe2b180_117, RIbe2adc0_109);
not \U$35135 ( \35381 , \35380 );
not \U$35136 ( \35382 , \14852 );
or \U$35137 ( \35383 , \35381 , \35382 );
nand \U$35138 ( \35384 , \21759 , \35290 );
nand \U$35139 ( \35385 , \35383 , \35384 );
not \U$35140 ( \35386 , \35385 );
nand \U$35141 ( \35387 , \9379 , RIbe2ae38_110);
not \U$35142 ( \35388 , \35387 );
and \U$35143 ( \35389 , \35386 , \35388 );
and \U$35144 ( \35390 , \35385 , \35387 );
nor \U$35145 ( \35391 , \35389 , \35390 );
not \U$35146 ( \35392 , \35391 );
not \U$35147 ( \35393 , \35392 );
or \U$35148 ( \35394 , \35379 , \35393 );
not \U$35149 ( \35395 , \35387 );
nand \U$35150 ( \35396 , \35395 , \35385 );
nand \U$35151 ( \35397 , \35394 , \35396 );
and \U$35152 ( \35398 , \35372 , \35397 );
and \U$35153 ( \35399 , \35370 , \35371 );
or \U$35154 ( \35400 , \35398 , \35399 );
not \U$35155 ( \35401 , \35400 );
or \U$35156 ( \35402 , \35363 , \35401 );
not \U$35157 ( \35403 , \35352 );
nand \U$35158 ( \35404 , \35403 , \35357 );
nand \U$35159 ( \35405 , \35402 , \35404 );
not \U$35160 ( \35406 , \35239 );
not \U$35161 ( \35407 , \35316 );
not \U$35162 ( \35408 , \35407 );
or \U$35163 ( \35409 , \35406 , \35408 );
or \U$35164 ( \35410 , \35407 , \35239 );
nand \U$35165 ( \35411 , \35409 , \35410 );
xor \U$35166 ( \35412 , \35405 , \35411 );
not \U$35167 ( \35413 , \35412 );
or \U$35168 ( \35414 , \35346 , \35413 );
nand \U$35169 ( \35415 , \35411 , \35405 );
nand \U$35170 ( \35416 , \35414 , \35415 );
xor \U$35171 ( \35417 , \35339 , \35416 );
not \U$35172 ( \35418 , \35147 );
not \U$35173 ( \35419 , \35326 );
or \U$35174 ( \35420 , \35418 , \35419 );
or \U$35175 ( \35421 , \35326 , \35147 );
nand \U$35176 ( \35422 , \35420 , \35421 );
xor \U$35177 ( \35423 , \35417 , \35422 );
not \U$35178 ( \35424 , \35423 );
and \U$35179 ( \35425 , \35412 , \35345 );
not \U$35180 ( \35426 , \35412 );
not \U$35181 ( \35427 , \35345 );
and \U$35182 ( \35428 , \35426 , \35427 );
nor \U$35183 ( \35429 , \35425 , \35428 );
not \U$35184 ( \35430 , \35429 );
not \U$35185 ( \35431 , \35430 );
xor \U$35186 ( \35432 , \35302 , \35288 );
not \U$35187 ( \35433 , \15693 );
not \U$35188 ( \35434 , \35286 );
or \U$35189 ( \35435 , \35433 , \35434 );
xnor \U$35190 ( \35436 , RIbe2ac58_106, RIbe2a190_83);
or \U$35191 ( \35437 , \34658 , \35436 );
nand \U$35192 ( \35438 , \35435 , \35437 );
not \U$35193 ( \35439 , \35438 );
not \U$35194 ( \35440 , \8794 );
not \U$35195 ( \35441 , \35273 );
or \U$35196 ( \35442 , \35440 , \35441 );
xor \U$35197 ( \35443 , RIbe2aeb0_111, RIbe2a3e8_88);
not \U$35198 ( \35444 , \35443 );
or \U$35199 ( \35445 , \11544 , \35444 );
nand \U$35200 ( \35446 , \35442 , \35445 );
not \U$35201 ( \35447 , \35446 );
or \U$35202 ( \35448 , \35439 , \35447 );
or \U$35203 ( \35449 , \35446 , \35438 );
xor \U$35204 ( \35450 , RIbe2a7a8_96, RIbe2a550_91);
not \U$35205 ( \35451 , \35450 );
not \U$35206 ( \35452 , \10434 );
or \U$35207 ( \35453 , \35451 , \35452 );
not \U$35208 ( \35454 , \35261 );
nand \U$35209 ( \35455 , \35454 , \12004 );
nand \U$35210 ( \35456 , \35453 , \35455 );
nand \U$35211 ( \35457 , \35449 , \35456 );
nand \U$35212 ( \35458 , \35448 , \35457 );
or \U$35213 ( \35459 , \35432 , \35458 );
xor \U$35214 ( \35460 , RIbe2b018_114, RIbe2b360_121);
not \U$35215 ( \35461 , \35460 );
not \U$35216 ( \35462 , \17571 );
or \U$35217 ( \35463 , \35461 , \35462 );
nand \U$35218 ( \35464 , \34563 , \35251 );
nand \U$35219 ( \35465 , \35463 , \35464 );
not \U$35220 ( \35466 , \35465 );
not \U$35221 ( \35467 , \19580 );
xnor \U$35222 ( \35468 , RIbe2a118_82, RIbe2aaf0_103);
not \U$35223 ( \35469 , \35468 );
and \U$35224 ( \35470 , \35467 , \35469 );
and \U$35225 ( \35471 , RIbe2ab68_104, \35179 );
nor \U$35226 ( \35472 , \35470 , \35471 );
not \U$35227 ( \35473 , \35472 );
xor \U$35228 ( \35474 , RIbe2a280_85, RIbe2a6b8_94);
not \U$35229 ( \35475 , \35474 );
not \U$35230 ( \35476 , \14942 );
or \U$35231 ( \35477 , \35475 , \35476 );
nand \U$35232 ( \35478 , \11348 , \35296 );
nand \U$35233 ( \35479 , \35477 , \35478 );
not \U$35234 ( \35480 , \35479 );
or \U$35235 ( \35481 , \35473 , \35480 );
or \U$35236 ( \35482 , \35479 , \35472 );
nand \U$35237 ( \35483 , \35481 , \35482 );
not \U$35238 ( \35484 , \35483 );
or \U$35239 ( \35485 , \35466 , \35484 );
not \U$35240 ( \35486 , \35472 );
nand \U$35241 ( \35487 , \35486 , \35479 );
nand \U$35242 ( \35488 , \35485 , \35487 );
nand \U$35243 ( \35489 , \35459 , \35488 );
nand \U$35244 ( \35490 , \35432 , \35458 );
and \U$35245 ( \35491 , \35489 , \35490 );
not \U$35246 ( \35492 , \35491 );
not \U$35247 ( \35493 , \35492 );
xor \U$35248 ( \35494 , \35246 , \35256 );
xor \U$35249 ( \35495 , \35494 , \35263 );
not \U$35250 ( \35496 , \35495 );
nand \U$35251 ( \35497 , RIbe2a910_99, RIbe2ae38_110);
and \U$35252 ( \35498 , \35497 , RIbe2a3e8_88);
or \U$35253 ( \35499 , RIbe2a910_99, RIbe2ae38_110);
nand \U$35254 ( \35500 , \35499 , RIbe2b5b8_126);
nand \U$35255 ( \35501 , \35498 , \35500 );
not \U$35256 ( \35502 , \35501 );
xor \U$35257 ( \35503 , RIbe2a910_99, RIbe2b3d8_122);
not \U$35258 ( \35504 , \35503 );
not \U$35259 ( \35505 , \12716 );
or \U$35260 ( \35506 , \35504 , \35505 );
nand \U$35261 ( \35507 , \11456 , \35373 );
nand \U$35262 ( \35508 , \35506 , \35507 );
nand \U$35263 ( \35509 , \35502 , \35508 );
xor \U$35264 ( \35510 , RIbe2a4d8_90, RIbe2af28_112);
not \U$35265 ( \35511 , \35510 );
not \U$35266 ( \35512 , \16913 );
or \U$35267 ( \35513 , \35511 , \35512 );
nand \U$35268 ( \35514 , \16917 , \35364 );
nand \U$35269 ( \35515 , \35513 , \35514 );
xor \U$35270 ( \35516 , RIbe2b540_125, RIbe2b108_116);
not \U$35271 ( \35517 , \35516 );
not \U$35272 ( \35518 , \25618 );
or \U$35273 ( \35519 , \35517 , \35518 );
nand \U$35274 ( \35520 , \23015 , \35172 );
nand \U$35275 ( \35521 , \35519 , \35520 );
nor \U$35276 ( \35522 , \35515 , \35521 );
or \U$35277 ( \35523 , \35509 , \35522 );
nand \U$35278 ( \35524 , \35521 , \35515 );
nand \U$35279 ( \35525 , \35523 , \35524 );
not \U$35280 ( \35526 , \35525 );
not \U$35281 ( \35527 , \35170 );
and \U$35282 ( \35528 , \35186 , \35527 );
not \U$35283 ( \35529 , \35186 );
and \U$35284 ( \35530 , \35529 , \35170 );
nor \U$35285 ( \35531 , \35528 , \35530 );
not \U$35286 ( \35532 , \35531 );
or \U$35287 ( \35533 , \35526 , \35532 );
or \U$35288 ( \35534 , \35525 , \35531 );
nand \U$35289 ( \35535 , \35533 , \35534 );
not \U$35290 ( \35536 , \35535 );
or \U$35291 ( \35537 , \35496 , \35536 );
not \U$35292 ( \35538 , \35531 );
nand \U$35293 ( \35539 , \35538 , \35525 );
nand \U$35294 ( \35540 , \35537 , \35539 );
not \U$35295 ( \35541 , \35540 );
not \U$35296 ( \35542 , \35266 );
and \U$35297 ( \35543 , \35312 , \35542 );
not \U$35298 ( \35544 , \35312 );
and \U$35299 ( \35545 , \35544 , \35266 );
nor \U$35300 ( \35546 , \35543 , \35545 );
not \U$35301 ( \35547 , \35546 );
or \U$35302 ( \35548 , \35541 , \35547 );
or \U$35303 ( \35549 , \35540 , \35546 );
nand \U$35304 ( \35550 , \35548 , \35549 );
not \U$35305 ( \35551 , \35550 );
or \U$35306 ( \35552 , \35493 , \35551 );
not \U$35307 ( \35553 , \35546 );
nand \U$35308 ( \35554 , \35553 , \35540 );
nand \U$35309 ( \35555 , \35552 , \35554 );
not \U$35310 ( \35556 , \35555 );
not \U$35311 ( \35557 , \35556 );
or \U$35312 ( \35558 , \35431 , \35557 );
not \U$35313 ( \35559 , \35555 );
not \U$35314 ( \35560 , \35429 );
or \U$35315 ( \35561 , \35559 , \35560 );
xor \U$35316 ( \35562 , RIbe2a730_95, RIbe2a550_91);
not \U$35317 ( \35563 , \35562 );
not \U$35318 ( \35564 , \10434 );
or \U$35319 ( \35565 , \35563 , \35564 );
nand \U$35320 ( \35566 , \10440 , \35450 );
nand \U$35321 ( \35567 , \35565 , \35566 );
xnor \U$35322 ( \35568 , RIbe2a0a0_81, RIbe2aaf0_103);
or \U$35323 ( \35569 , \19580 , \35568 );
or \U$35324 ( \35570 , \18830 , \35468 );
nand \U$35325 ( \35571 , \35569 , \35570 );
nor \U$35326 ( \35572 , \35567 , \35571 );
xor \U$35327 ( \35573 , RIbe2a640_93, RIbe2a280_85);
and \U$35328 ( \35574 , \24029 , \35573 );
and \U$35329 ( \35575 , \11348 , \35474 );
nor \U$35330 ( \35576 , \35574 , \35575 );
or \U$35331 ( \35577 , \35572 , \35576 );
nand \U$35332 ( \35578 , \35567 , \35571 );
nand \U$35333 ( \35579 , \35577 , \35578 );
not \U$35334 ( \35580 , \35579 );
xor \U$35335 ( \35581 , RIbe2b108_116, RIbe2b4c8_124);
not \U$35336 ( \35582 , \35581 );
not \U$35337 ( \35583 , \14297 );
or \U$35338 ( \35584 , \35582 , \35583 );
nand \U$35339 ( \35585 , \13534 , \35516 );
nand \U$35340 ( \35586 , \35584 , \35585 );
not \U$35341 ( \35587 , \35586 );
xor \U$35342 ( \35588 , RIbe2b018_114, RIbe2b2e8_120);
not \U$35343 ( \35589 , \35588 );
not \U$35344 ( \35590 , \16811 );
or \U$35345 ( \35591 , \35589 , \35590 );
nand \U$35346 ( \35592 , \15953 , \35460 );
nand \U$35347 ( \35593 , \35591 , \35592 );
not \U$35348 ( \35594 , \35593 );
not \U$35349 ( \35595 , \35594 );
xor \U$35350 ( \35596 , RIbe2af28_112, RIbe2a460_89);
not \U$35351 ( \35597 , \35596 );
not \U$35352 ( \35598 , \14423 );
or \U$35353 ( \35599 , \35597 , \35598 );
nand \U$35354 ( \35600 , \17810 , \35510 );
nand \U$35355 ( \35601 , \35599 , \35600 );
not \U$35356 ( \35602 , \35601 );
or \U$35357 ( \35603 , \35595 , \35602 );
or \U$35358 ( \35604 , \35601 , \35594 );
nand \U$35359 ( \35605 , \35603 , \35604 );
not \U$35360 ( \35606 , \35605 );
or \U$35361 ( \35607 , \35587 , \35606 );
nand \U$35362 ( \35608 , \35601 , \35593 );
nand \U$35363 ( \35609 , \35607 , \35608 );
not \U$35364 ( \35610 , \35609 );
or \U$35365 ( \35611 , \35580 , \35610 );
or \U$35366 ( \35612 , \35609 , \35579 );
xor \U$35367 ( \35613 , RIbe2ad48_108, RIbe2b180_117);
not \U$35368 ( \35614 , \35613 );
not \U$35369 ( \35615 , \32900 );
or \U$35370 ( \35616 , \35614 , \35615 );
nand \U$35371 ( \35617 , \21759 , \35380 );
nand \U$35372 ( \35618 , \35616 , \35617 );
xor \U$35373 ( \35619 , RIbe2a3e8_88, RIbe2ae38_110);
not \U$35374 ( \35620 , \35619 );
not \U$35375 ( \35621 , \15475 );
or \U$35376 ( \35622 , \35620 , \35621 );
nand \U$35377 ( \35623 , \10476 , \35443 );
nand \U$35378 ( \35624 , \35622 , \35623 );
nor \U$35379 ( \35625 , \35618 , \35624 );
xor \U$35380 ( \35626 , RIbe2abe0_105, RIbe2a190_83);
not \U$35381 ( \35627 , \35626 );
not \U$35382 ( \35628 , \15690 );
or \U$35383 ( \35629 , \35627 , \35628 );
not \U$35384 ( \35630 , \35436 );
nand \U$35385 ( \35631 , \35630 , \11400 );
nand \U$35386 ( \35632 , \35629 , \35631 );
not \U$35387 ( \35633 , \35632 );
or \U$35388 ( \35634 , \35625 , \35633 );
nand \U$35389 ( \35635 , \35618 , \35624 );
nand \U$35390 ( \35636 , \35634 , \35635 );
nand \U$35391 ( \35637 , \35612 , \35636 );
nand \U$35392 ( \35638 , \35611 , \35637 );
xor \U$35393 ( \35639 , \35370 , \35371 );
xor \U$35394 ( \35640 , \35639 , \35397 );
xor \U$35395 ( \35641 , \35638 , \35640 );
xor \U$35396 ( \35642 , \35458 , \35488 );
xor \U$35397 ( \35643 , \35642 , \35432 );
and \U$35398 ( \35644 , \35641 , \35643 );
and \U$35399 ( \35645 , \35638 , \35640 );
or \U$35400 ( \35646 , \35644 , \35645 );
not \U$35401 ( \35647 , \35646 );
not \U$35402 ( \35648 , \35201 );
not \U$35403 ( \35649 , \35192 );
or \U$35404 ( \35650 , \35648 , \35649 );
nand \U$35405 ( \35651 , \35200 , \35191 );
nand \U$35406 ( \35652 , \35650 , \35651 );
xor \U$35407 ( \35653 , \35652 , \35162 );
not \U$35408 ( \35654 , \35653 );
not \U$35409 ( \35655 , \35361 );
not \U$35410 ( \35656 , \35400 );
or \U$35411 ( \35657 , \35655 , \35656 );
or \U$35412 ( \35658 , \35400 , \35361 );
nand \U$35413 ( \35659 , \35657 , \35658 );
not \U$35414 ( \35660 , \35659 );
or \U$35415 ( \35661 , \35654 , \35660 );
or \U$35416 ( \35662 , \35659 , \35653 );
nand \U$35417 ( \35663 , \35661 , \35662 );
not \U$35418 ( \35664 , \35663 );
or \U$35419 ( \35665 , \35647 , \35664 );
not \U$35420 ( \35666 , \35653 );
nand \U$35421 ( \35667 , \35666 , \35659 );
nand \U$35422 ( \35668 , \35665 , \35667 );
not \U$35423 ( \35669 , \35668 );
nand \U$35424 ( \35670 , \35561 , \35669 );
nand \U$35425 ( \35671 , \35558 , \35670 );
nand \U$35426 ( \35672 , \35424 , \35671 );
xor \U$35427 ( \35673 , \35139 , \35141 );
xor \U$35428 ( \35674 , \35673 , \35330 );
xor \U$35429 ( \35675 , \35339 , \35416 );
and \U$35430 ( \35676 , \35675 , \35422 );
and \U$35431 ( \35677 , \35339 , \35416 );
or \U$35432 ( \35678 , \35676 , \35677 );
nor \U$35433 ( \35679 , \35674 , \35678 );
not \U$35434 ( \35680 , \35679 );
nand \U$35435 ( \35681 , \35337 , \35672 , \35680 );
not \U$35436 ( \35682 , \35086 );
nand \U$35437 ( \35683 , \35682 , \35121 );
not \U$35438 ( \35684 , \35683 );
not \U$35439 ( \35685 , \35126 );
or \U$35440 ( \35686 , \35684 , \35685 );
not \U$35441 ( \35687 , \35121 );
nand \U$35442 ( \35688 , \35687 , \35086 );
nand \U$35443 ( \35689 , \35686 , \35688 );
not \U$35444 ( \35690 , \35689 );
xnor \U$35445 ( \35691 , \33840 , \33784 );
not \U$35446 ( \35692 , \33669 );
not \U$35447 ( \35693 , \33681 );
not \U$35448 ( \35694 , \35693 );
or \U$35449 ( \35695 , \35692 , \35694 );
not \U$35450 ( \35696 , \33669 );
nand \U$35451 ( \35697 , \35696 , \33681 );
nand \U$35452 ( \35698 , \35695 , \35697 );
xor \U$35453 ( \35699 , \35691 , \35698 );
not \U$35454 ( \35700 , \35070 );
not \U$35455 ( \35701 , \35084 );
or \U$35456 ( \35702 , \35700 , \35701 );
not \U$35457 ( \35703 , \35075 );
nand \U$35458 ( \35704 , \35703 , \35079 );
nand \U$35459 ( \35705 , \35702 , \35704 );
xor \U$35460 ( \35706 , \35699 , \35705 );
not \U$35461 ( \35707 , \35706 );
not \U$35462 ( \35708 , \35707 );
not \U$35463 ( \35709 , \35093 );
not \U$35464 ( \35710 , \35119 );
or \U$35465 ( \35711 , \35709 , \35710 );
not \U$35466 ( \35712 , \35116 );
not \U$35467 ( \35713 , \35094 );
or \U$35468 ( \35714 , \35712 , \35713 );
nand \U$35469 ( \35715 , \35714 , \35088 );
nand \U$35470 ( \35716 , \35711 , \35715 );
not \U$35471 ( \35717 , \35716 );
or \U$35472 ( \35718 , \35066 , \35053 );
not \U$35473 ( \35719 , \35062 );
nand \U$35474 ( \35720 , \35719 , \35059 );
nand \U$35475 ( \35721 , \35718 , \35720 );
not \U$35476 ( \35722 , \35721 );
nand \U$35477 ( \35723 , \33521 , \33529 );
not \U$35478 ( \35724 , \33524 );
xnor \U$35479 ( \35725 , \35723 , \35724 );
not \U$35480 ( \35726 , \35725 );
and \U$35481 ( \35727 , \35722 , \35726 );
and \U$35482 ( \35728 , \35721 , \35725 );
nor \U$35483 ( \35729 , \35727 , \35728 );
or \U$35484 ( \35730 , \35115 , \35106 );
not \U$35485 ( \35731 , \35109 );
nand \U$35486 ( \35732 , \35730 , \35731 );
nand \U$35487 ( \35733 , \35115 , \35106 );
nand \U$35488 ( \35734 , \35732 , \35733 );
xnor \U$35489 ( \35735 , \35729 , \35734 );
not \U$35490 ( \35736 , \35735 );
and \U$35491 ( \35737 , \35717 , \35736 );
not \U$35492 ( \35738 , \35717 );
and \U$35493 ( \35739 , \35738 , \35735 );
nor \U$35494 ( \35740 , \35737 , \35739 );
not \U$35495 ( \35741 , \35740 );
not \U$35496 ( \35742 , \35741 );
or \U$35497 ( \35743 , \35708 , \35742 );
nand \U$35498 ( \35744 , \35740 , \35706 );
nand \U$35499 ( \35745 , \35743 , \35744 );
not \U$35500 ( \35746 , \35745 );
nand \U$35501 ( \35747 , \35690 , \35746 );
not \U$35502 ( \35748 , \35729 );
not \U$35503 ( \35749 , \35748 );
not \U$35504 ( \35750 , \35734 );
or \U$35505 ( \35751 , \35749 , \35750 );
not \U$35506 ( \35752 , \35725 );
nand \U$35507 ( \35753 , \35752 , \35721 );
nand \U$35508 ( \35754 , \35751 , \35753 );
not \U$35509 ( \35755 , \35691 );
not \U$35510 ( \35756 , \35755 );
not \U$35511 ( \35757 , \35698 );
or \U$35512 ( \35758 , \35756 , \35757 );
or \U$35513 ( \35759 , \35698 , \35755 );
nand \U$35514 ( \35760 , \35759 , \35705 );
nand \U$35515 ( \35761 , \35758 , \35760 );
xor \U$35516 ( \35762 , \35754 , \35761 );
not \U$35517 ( \35763 , \35762 );
not \U$35518 ( \35764 , \33850 );
not \U$35519 ( \35765 , \33686 );
not \U$35520 ( \35766 , \35765 );
and \U$35521 ( \35767 , \35764 , \35766 );
and \U$35522 ( \35768 , \33850 , \35765 );
nor \U$35523 ( \35769 , \35767 , \35768 );
not \U$35524 ( \35770 , \35769 );
buf \U$35525 ( \35771 , \33534 );
not \U$35526 ( \35772 , \35771 );
not \U$35527 ( \35773 , \33508 );
not \U$35528 ( \35774 , \35773 );
and \U$35529 ( \35775 , \35772 , \35774 );
and \U$35530 ( \35776 , \35771 , \35773 );
nor \U$35531 ( \35777 , \35775 , \35776 );
and \U$35532 ( \35778 , \33617 , \33612 );
not \U$35533 ( \35779 , \33617 );
not \U$35534 ( \35780 , \33612 );
and \U$35535 ( \35781 , \35779 , \35780 );
nor \U$35536 ( \35782 , \35778 , \35781 );
xor \U$35537 ( \35783 , \35782 , \33614 );
and \U$35538 ( \35784 , \35777 , \35783 );
not \U$35539 ( \35785 , \35777 );
not \U$35540 ( \35786 , \35783 );
and \U$35541 ( \35787 , \35785 , \35786 );
nor \U$35542 ( \35788 , \35784 , \35787 );
not \U$35543 ( \35789 , \35788 );
and \U$35544 ( \35790 , \35770 , \35789 );
and \U$35545 ( \35791 , \35769 , \35788 );
nor \U$35546 ( \35792 , \35790 , \35791 );
not \U$35547 ( \35793 , \35792 );
or \U$35548 ( \35794 , \35763 , \35793 );
or \U$35549 ( \35795 , \35792 , \35762 );
nand \U$35550 ( \35796 , \35794 , \35795 );
not \U$35551 ( \35797 , \35707 );
not \U$35552 ( \35798 , \35740 );
or \U$35553 ( \35799 , \35797 , \35798 );
not \U$35554 ( \35800 , \35717 );
nand \U$35555 ( \35801 , \35800 , \35735 );
nand \U$35556 ( \35802 , \35799 , \35801 );
not \U$35557 ( \35803 , \35802 );
nand \U$35558 ( \35804 , \35796 , \35803 );
nand \U$35559 ( \35805 , \35747 , \35804 );
not \U$35560 ( \35806 , \35805 );
xor \U$35561 ( \35807 , \33437 , \33620 );
xnor \U$35562 ( \35808 , \35807 , \33539 );
not \U$35563 ( \35809 , \33869 );
not \U$35564 ( \35810 , \35809 );
not \U$35565 ( \35811 , \33855 );
and \U$35566 ( \35812 , \35810 , \35811 );
not \U$35567 ( \35813 , \33869 );
and \U$35568 ( \35814 , \35813 , \33855 );
nor \U$35569 ( \35815 , \35812 , \35814 );
xor \U$35570 ( \35816 , \35808 , \35815 );
not \U$35571 ( \35817 , \35777 );
not \U$35572 ( \35818 , \35769 );
or \U$35573 ( \35819 , \35817 , \35818 );
nand \U$35574 ( \35820 , \35819 , \35783 );
not \U$35575 ( \35821 , \35777 );
not \U$35576 ( \35822 , \35769 );
nand \U$35577 ( \35823 , \35821 , \35822 );
and \U$35578 ( \35824 , \35820 , \35823 );
xor \U$35579 ( \35825 , \35816 , \35824 );
or \U$35580 ( \35826 , \35761 , \35754 );
and \U$35581 ( \35827 , \35792 , \35826 );
and \U$35582 ( \35828 , \35754 , \35761 );
nor \U$35583 ( \35829 , \35827 , \35828 );
nand \U$35584 ( \35830 , \35825 , \35829 );
xor \U$35585 ( \35831 , \33875 , \33874 );
xnor \U$35586 ( \35832 , \35831 , \33877 );
xor \U$35587 ( \35833 , \35808 , \35815 );
and \U$35588 ( \35834 , \35833 , \35824 );
and \U$35589 ( \35835 , \35808 , \35815 );
or \U$35590 ( \35836 , \35834 , \35835 );
nand \U$35591 ( \35837 , \35832 , \35836 );
nand \U$35592 ( \35838 , \35806 , \35830 , \35837 );
nor \U$35593 ( \35839 , \35681 , \35838 );
buf \U$35594 ( \35840 , \35663 );
not \U$35595 ( \35841 , \35646 );
and \U$35596 ( \35842 , \35840 , \35841 );
not \U$35597 ( \35843 , \35840 );
and \U$35598 ( \35844 , \35843 , \35646 );
nor \U$35599 ( \35845 , \35842 , \35844 );
not \U$35600 ( \35846 , \35845 );
not \U$35601 ( \35847 , \35846 );
xor \U$35602 ( \35848 , \35638 , \35640 );
xor \U$35603 ( \35849 , \35848 , \35643 );
not \U$35604 ( \35850 , \35849 );
not \U$35605 ( \35851 , \35495 );
not \U$35606 ( \35852 , \35535 );
not \U$35607 ( \35853 , \35852 );
or \U$35608 ( \35854 , \35851 , \35853 );
not \U$35609 ( \35855 , \35495 );
nand \U$35610 ( \35856 , \35855 , \35535 );
nand \U$35611 ( \35857 , \35854 , \35856 );
not \U$35612 ( \35858 , \35857 );
xor \U$35613 ( \35859 , \35456 , \35446 );
xor \U$35614 ( \35860 , \35859 , \35438 );
not \U$35615 ( \35861 , \35860 );
xnor \U$35616 ( \35862 , \35465 , \35483 );
not \U$35617 ( \35863 , \35862 );
and \U$35618 ( \35864 , \35378 , \35391 );
not \U$35619 ( \35865 , \35378 );
and \U$35620 ( \35866 , \35865 , \35392 );
or \U$35621 ( \35867 , \35864 , \35866 );
not \U$35622 ( \35868 , \35867 );
or \U$35623 ( \35869 , \35863 , \35868 );
or \U$35624 ( \35870 , \35867 , \35862 );
nand \U$35625 ( \35871 , \35869 , \35870 );
not \U$35626 ( \35872 , \35871 );
or \U$35627 ( \35873 , \35861 , \35872 );
not \U$35628 ( \35874 , \35862 );
nand \U$35629 ( \35875 , \35874 , \35867 );
nand \U$35630 ( \35876 , \35873 , \35875 );
not \U$35631 ( \35877 , \35876 );
not \U$35632 ( \35878 , \35877 );
or \U$35633 ( \35879 , \35858 , \35878 );
not \U$35634 ( \35880 , \35876 );
or \U$35635 ( \35881 , \35880 , \35857 );
nand \U$35636 ( \35882 , \35879 , \35881 );
not \U$35637 ( \35883 , \35882 );
or \U$35638 ( \35884 , \35850 , \35883 );
nand \U$35639 ( \35885 , \35876 , \35857 );
nand \U$35640 ( \35886 , \35884 , \35885 );
not \U$35641 ( \35887 , \35550 );
not \U$35642 ( \35888 , \35491 );
and \U$35643 ( \35889 , \35887 , \35888 );
and \U$35644 ( \35890 , \35550 , \35491 );
nor \U$35645 ( \35891 , \35889 , \35890 );
and \U$35646 ( \35892 , \35886 , \35891 );
not \U$35647 ( \35893 , \35886 );
not \U$35648 ( \35894 , \35891 );
and \U$35649 ( \35895 , \35893 , \35894 );
or \U$35650 ( \35896 , \35892 , \35895 );
not \U$35651 ( \35897 , \35896 );
or \U$35652 ( \35898 , \35847 , \35897 );
nand \U$35653 ( \35899 , \35886 , \35894 );
nand \U$35654 ( \35900 , \35898 , \35899 );
not \U$35655 ( \35901 , \35555 );
not \U$35656 ( \35902 , \35669 );
or \U$35657 ( \35903 , \35901 , \35902 );
nand \U$35658 ( \35904 , \35668 , \35556 );
nand \U$35659 ( \35905 , \35903 , \35904 );
and \U$35660 ( \35906 , \35905 , \35429 );
not \U$35661 ( \35907 , \35905 );
and \U$35662 ( \35908 , \35907 , \35430 );
nor \U$35663 ( \35909 , \35906 , \35908 );
nor \U$35664 ( \35910 , \35900 , \35909 );
not \U$35665 ( \35911 , \35845 );
not \U$35666 ( \35912 , \35896 );
or \U$35667 ( \35913 , \35911 , \35912 );
or \U$35668 ( \35914 , \35896 , \35845 );
nand \U$35669 ( \35915 , \35913 , \35914 );
not \U$35670 ( \35916 , \35625 );
nand \U$35671 ( \35917 , \35916 , \35635 );
not \U$35672 ( \35918 , \35917 );
not \U$35673 ( \35919 , \35632 );
and \U$35674 ( \35920 , \35918 , \35919 );
and \U$35675 ( \35921 , \35917 , \35632 );
nor \U$35676 ( \35922 , \35920 , \35921 );
not \U$35677 ( \35923 , \35922 );
not \U$35678 ( \35924 , \35923 );
not \U$35679 ( \35925 , \35586 );
not \U$35680 ( \35926 , \35925 );
not \U$35681 ( \35927 , \35605 );
or \U$35682 ( \35928 , \35926 , \35927 );
or \U$35683 ( \35929 , \35605 , \35925 );
nand \U$35684 ( \35930 , \35928 , \35929 );
not \U$35685 ( \35931 , \35930 );
and \U$35686 ( \35932 , \8794 , RIbe2ae38_110);
xor \U$35687 ( \35933 , RIbe2a550_91, RIbe2b450_123);
not \U$35688 ( \35934 , \35933 );
not \U$35689 ( \35935 , \18635 );
or \U$35690 ( \35936 , \35934 , \35935 );
nand \U$35691 ( \35937 , \32080 , \35562 );
nand \U$35692 ( \35938 , \35936 , \35937 );
xor \U$35693 ( \35939 , \35932 , \35938 );
and \U$35694 ( \35940 , RIbe2adc0_109, RIbe2af28_112);
nor \U$35695 ( \35941 , RIbe2adc0_109, RIbe2af28_112);
nor \U$35696 ( \35942 , \35940 , \35941 );
not \U$35697 ( \35943 , \35942 );
not \U$35698 ( \35944 , \35366 );
or \U$35699 ( \35945 , \35943 , \35944 );
nand \U$35700 ( \35946 , \17811 , \35596 );
nand \U$35701 ( \35947 , \35945 , \35946 );
and \U$35702 ( \35948 , \35939 , \35947 );
and \U$35703 ( \35949 , \35932 , \35938 );
nor \U$35704 ( \35950 , \35948 , \35949 );
not \U$35705 ( \35951 , \35950 );
or \U$35706 ( \35952 , \35931 , \35951 );
or \U$35707 ( \35953 , \35950 , \35930 );
nand \U$35708 ( \35954 , \35952 , \35953 );
not \U$35709 ( \35955 , \35954 );
or \U$35710 ( \35956 , \35924 , \35955 );
not \U$35711 ( \35957 , \35950 );
nand \U$35712 ( \35958 , \35957 , \35930 );
nand \U$35713 ( \35959 , \35956 , \35958 );
not \U$35714 ( \35960 , \35959 );
xor \U$35715 ( \35961 , \35515 , \35521 );
xnor \U$35716 ( \35962 , \35961 , \35509 );
not \U$35717 ( \35963 , \35962 );
not \U$35718 ( \35964 , \16812 );
not \U$35719 ( \35965 , \35964 );
not \U$35720 ( \35966 , RIbe2b018_114);
not \U$35721 ( \35967 , RIbe2a4d8_90);
or \U$35722 ( \35968 , \35966 , \35967 );
or \U$35723 ( \35969 , RIbe2a4d8_90, RIbe2b018_114);
nand \U$35724 ( \35970 , \35968 , \35969 );
not \U$35725 ( \35971 , \35970 );
and \U$35726 ( \35972 , \35965 , \35971 );
and \U$35727 ( \35973 , \20583 , \35588 );
nor \U$35728 ( \35974 , \35972 , \35973 );
not \U$35729 ( \35975 , \35974 );
not \U$35730 ( \35976 , \35975 );
xor \U$35731 ( \35977 , RIbe2aaf0_103, RIbe2b360_121);
and \U$35732 ( \35978 , \34608 , \35977 );
not \U$35733 ( \35979 , RIbe2ab68_104);
nor \U$35734 ( \35980 , \35979 , \35568 );
nor \U$35735 ( \35981 , \35978 , \35980 );
not \U$35736 ( \35982 , \35981 );
xor \U$35737 ( \35983 , RIbe2b108_116, RIbe2a6b8_94);
not \U$35738 ( \35984 , \35983 );
not \U$35739 ( \35985 , \14297 );
or \U$35740 ( \35986 , \35984 , \35985 );
nand \U$35741 ( \35987 , \16875 , \35581 );
nand \U$35742 ( \35988 , \35986 , \35987 );
not \U$35743 ( \35989 , \35988 );
or \U$35744 ( \35990 , \35982 , \35989 );
or \U$35745 ( \35991 , \35988 , \35981 );
nand \U$35746 ( \35992 , \35990 , \35991 );
not \U$35747 ( \35993 , \35992 );
or \U$35748 ( \35994 , \35976 , \35993 );
not \U$35749 ( \35995 , \35981 );
nand \U$35750 ( \35996 , \35995 , \35988 );
nand \U$35751 ( \35997 , \35994 , \35996 );
not \U$35752 ( \35998 , \35997 );
xor \U$35753 ( \35999 , \35508 , \35501 );
not \U$35754 ( \36000 , \35999 );
not \U$35755 ( \36001 , \11396 );
xor \U$35756 ( \36002 , RIbe2a7a8_96, RIbe2a190_83);
not \U$35757 ( \36003 , \36002 );
or \U$35758 ( \36004 , \36001 , \36003 );
nand \U$35759 ( \36005 , \31948 , \35626 );
nand \U$35760 ( \36006 , \36004 , \36005 );
not \U$35761 ( \36007 , \36006 );
xor \U$35762 ( \36008 , RIbe2ac58_106, RIbe2a280_85);
not \U$35763 ( \36009 , \36008 );
buf \U$35764 ( \36010 , \27992 );
not \U$35765 ( \36011 , \36010 );
or \U$35766 ( \36012 , \36009 , \36011 );
nand \U$35767 ( \36013 , \14649 , \35573 );
nand \U$35768 ( \36014 , \36012 , \36013 );
not \U$35769 ( \36015 , \36014 );
or \U$35770 ( \36016 , \36007 , \36015 );
or \U$35771 ( \36017 , \36014 , \36006 );
xor \U$35772 ( \36018 , RIbe2a910_99, RIbe2aeb0_111);
not \U$35773 ( \36019 , \36018 );
not \U$35774 ( \36020 , \9738 );
or \U$35775 ( \36021 , \36019 , \36020 );
nand \U$35776 ( \36022 , \10401 , \35503 );
nand \U$35777 ( \36023 , \36021 , \36022 );
nand \U$35778 ( \36024 , \36017 , \36023 );
nand \U$35779 ( \36025 , \36016 , \36024 );
not \U$35780 ( \36026 , \36025 );
or \U$35781 ( \36027 , \36000 , \36026 );
or \U$35782 ( \36028 , \36025 , \35999 );
nand \U$35783 ( \36029 , \36027 , \36028 );
not \U$35784 ( \36030 , \36029 );
or \U$35785 ( \36031 , \35998 , \36030 );
not \U$35786 ( \36032 , \35999 );
nand \U$35787 ( \36033 , \36032 , \36025 );
nand \U$35788 ( \36034 , \36031 , \36033 );
not \U$35789 ( \36035 , \36034 );
not \U$35790 ( \36036 , \36035 );
or \U$35791 ( \36037 , \35963 , \36036 );
not \U$35792 ( \36038 , \35962 );
nand \U$35793 ( \36039 , \36038 , \36034 );
nand \U$35794 ( \36040 , \36037 , \36039 );
not \U$35795 ( \36041 , \36040 );
or \U$35796 ( \36042 , \35960 , \36041 );
nand \U$35797 ( \36043 , \36034 , \35962 );
nand \U$35798 ( \36044 , \36042 , \36043 );
xor \U$35799 ( \36045 , \35849 , \35882 );
xor \U$35800 ( \36046 , \36044 , \36045 );
not \U$35801 ( \36047 , \35636 );
not \U$35802 ( \36048 , \35609 );
not \U$35803 ( \36049 , \35579 );
not \U$35804 ( \36050 , \36049 );
and \U$35805 ( \36051 , \36048 , \36050 );
and \U$35806 ( \36052 , \35609 , \36049 );
nor \U$35807 ( \36053 , \36051 , \36052 );
not \U$35808 ( \36054 , \36053 );
or \U$35809 ( \36055 , \36047 , \36054 );
or \U$35810 ( \36056 , \36053 , \35636 );
nand \U$35811 ( \36057 , \36055 , \36056 );
not \U$35812 ( \36058 , \36057 );
buf \U$35813 ( \36059 , \35871 );
not \U$35814 ( \36060 , \35860 );
and \U$35815 ( \36061 , \36059 , \36060 );
not \U$35816 ( \36062 , \36059 );
and \U$35817 ( \36063 , \36062 , \35860 );
nor \U$35818 ( \36064 , \36061 , \36063 );
not \U$35819 ( \36065 , \36064 );
or \U$35820 ( \36066 , \36058 , \36065 );
or \U$35821 ( \36067 , \36064 , \36057 );
nand \U$35822 ( \36068 , \36066 , \36067 );
not \U$35823 ( \36069 , \36068 );
not \U$35824 ( \36070 , \35959 );
not \U$35825 ( \36071 , \36070 );
not \U$35826 ( \36072 , \36040 );
or \U$35827 ( \36073 , \36071 , \36072 );
or \U$35828 ( \36074 , \36040 , \36070 );
nand \U$35829 ( \36075 , \36073 , \36074 );
not \U$35830 ( \36076 , \36075 );
or \U$35831 ( \36077 , \36069 , \36076 );
not \U$35832 ( \36078 , \36064 );
nand \U$35833 ( \36079 , \36078 , \36057 );
nand \U$35834 ( \36080 , \36077 , \36079 );
and \U$35835 ( \36081 , \36046 , \36080 );
and \U$35836 ( \36082 , \36044 , \36045 );
or \U$35837 ( \36083 , \36081 , \36082 );
nor \U$35838 ( \36084 , \35915 , \36083 );
nor \U$35839 ( \36085 , \35910 , \36084 );
xor \U$35840 ( \36086 , \36044 , \36045 );
xor \U$35841 ( \36087 , \36086 , \36080 );
xor \U$35842 ( \36088 , \36068 , \36075 );
not \U$35843 ( \36089 , \36088 );
not \U$35844 ( \36090 , \15353 );
not \U$35845 ( \36091 , RIbe2b540_125);
not \U$35846 ( \36092 , RIbe2b180_117);
or \U$35847 ( \36093 , \36091 , \36092 );
or \U$35848 ( \36094 , RIbe2b180_117, RIbe2b540_125);
nand \U$35849 ( \36095 , \36093 , \36094 );
nor \U$35850 ( \36096 , \36090 , \36095 );
and \U$35851 ( \36097 , \21759 , \35613 );
nor \U$35852 ( \36098 , \36096 , \36097 );
not \U$35853 ( \36099 , \36098 );
not \U$35854 ( \36100 , RIbe2a550_91);
not \U$35855 ( \36101 , RIbe2b3d8_122);
and \U$35856 ( \36102 , \36100 , \36101 );
and \U$35857 ( \36103 , RIbe2a550_91, RIbe2b3d8_122);
nor \U$35858 ( \36104 , \36102 , \36103 );
not \U$35859 ( \36105 , \36104 );
not \U$35860 ( \36106 , \10434 );
or \U$35861 ( \36107 , \36105 , \36106 );
nand \U$35862 ( \36108 , \10440 , \35933 );
nand \U$35863 ( \36109 , \36107 , \36108 );
not \U$35864 ( \36110 , RIbe2ae38_110);
nand \U$35865 ( \36111 , \36110 , \9729 , RIbe2a910_99);
and \U$35866 ( \36112 , \36111 , \9734 );
not \U$35867 ( \36113 , \36112 );
and \U$35868 ( \36114 , \36109 , \36113 );
not \U$35869 ( \36115 , \36114 );
or \U$35870 ( \36116 , \36099 , \36115 );
or \U$35871 ( \36117 , \36114 , \36098 );
nand \U$35872 ( \36118 , \36116 , \36117 );
not \U$35873 ( \36119 , \36118 );
and \U$35874 ( \36120 , RIbe2ad48_108, RIbe2af28_112);
nor \U$35875 ( \36121 , RIbe2ad48_108, RIbe2af28_112);
nor \U$35876 ( \36122 , \36120 , \36121 );
and \U$35877 ( \36123 , \18649 , \36122 );
and \U$35878 ( \36124 , \15348 , \35942 );
nor \U$35879 ( \36125 , \36123 , \36124 );
not \U$35880 ( \36126 , \36125 );
not \U$35881 ( \36127 , \36126 );
xor \U$35882 ( \36128 , RIbe2a280_85, RIbe2abe0_105);
not \U$35883 ( \36129 , \36128 );
not \U$35884 ( \36130 , \27993 );
or \U$35885 ( \36131 , \36129 , \36130 );
nand \U$35886 ( \36132 , \11348 , \36008 );
nand \U$35887 ( \36133 , \36131 , \36132 );
not \U$35888 ( \36134 , \36133 );
and \U$35889 ( \36135 , RIbe2a910_99, RIbe2ae38_110);
not \U$35890 ( \36136 , RIbe2a910_99);
and \U$35891 ( \36137 , \36136 , \24871 );
nor \U$35892 ( \36138 , \36135 , \36137 );
not \U$35893 ( \36139 , \36138 );
not \U$35894 ( \36140 , \9738 );
or \U$35895 ( \36141 , \36139 , \36140 );
nand \U$35896 ( \36142 , \11456 , \36018 );
nand \U$35897 ( \36143 , \36141 , \36142 );
not \U$35898 ( \36144 , \36143 );
not \U$35899 ( \36145 , \36144 );
or \U$35900 ( \36146 , \36134 , \36145 );
not \U$35901 ( \36147 , \36133 );
nand \U$35902 ( \36148 , \36147 , \36143 );
nand \U$35903 ( \36149 , \36146 , \36148 );
not \U$35904 ( \36150 , \36149 );
or \U$35905 ( \36151 , \36127 , \36150 );
nand \U$35906 ( \36152 , \36143 , \36133 );
nand \U$35907 ( \36153 , \36151 , \36152 );
not \U$35908 ( \36154 , \36153 );
or \U$35909 ( \36155 , \36119 , \36154 );
not \U$35910 ( \36156 , \36098 );
nand \U$35911 ( \36157 , \36156 , \36114 );
nand \U$35912 ( \36158 , \36155 , \36157 );
not \U$35913 ( \36159 , \36158 );
not \U$35914 ( \36160 , \35572 );
nand \U$35915 ( \36161 , \36160 , \35578 );
and \U$35916 ( \36162 , \36161 , \35576 );
not \U$35917 ( \36163 , \36161 );
not \U$35918 ( \36164 , \35576 );
and \U$35919 ( \36165 , \36163 , \36164 );
or \U$35920 ( \36166 , \36162 , \36165 );
not \U$35921 ( \36167 , \36166 );
and \U$35922 ( \36168 , \36159 , \36167 );
and \U$35923 ( \36169 , \36158 , \36166 );
nor \U$35924 ( \36170 , \36168 , \36169 );
not \U$35925 ( \36171 , \36170 );
buf \U$35926 ( \36172 , \36029 );
and \U$35927 ( \36173 , \36172 , \35997 );
not \U$35928 ( \36174 , \36172 );
not \U$35929 ( \36175 , \35997 );
and \U$35930 ( \36176 , \36174 , \36175 );
nor \U$35931 ( \36177 , \36173 , \36176 );
and \U$35932 ( \36178 , \36171 , \36177 );
not \U$35933 ( \36179 , \36158 );
nor \U$35934 ( \36180 , \36179 , \36166 );
nor \U$35935 ( \36181 , \36178 , \36180 );
not \U$35936 ( \36182 , \36181 );
xor \U$35937 ( \36183 , \36153 , \36118 );
not \U$35938 ( \36184 , \36183 );
xor \U$35939 ( \36185 , \36014 , \36006 );
xnor \U$35940 ( \36186 , \36185 , \36023 );
not \U$35941 ( \36187 , \36186 );
and \U$35942 ( \36188 , \36109 , \36113 );
not \U$35943 ( \36189 , \36109 );
and \U$35944 ( \36190 , \36189 , \36112 );
nor \U$35945 ( \36191 , \36188 , \36190 );
not \U$35946 ( \36192 , \36191 );
not \U$35947 ( \36193 , \34558 );
or \U$35948 ( \36194 , RIbe2a460_89, RIbe2b018_114);
nand \U$35949 ( \36195 , RIbe2a460_89, RIbe2b018_114);
nand \U$35950 ( \36196 , \36194 , \36195 );
not \U$35951 ( \36197 , \36196 );
and \U$35952 ( \36198 , \36193 , \36197 );
not \U$35953 ( \36199 , \20583 );
nor \U$35954 ( \36200 , \36199 , \35970 );
nor \U$35955 ( \36201 , \36198 , \36200 );
not \U$35956 ( \36202 , \36201 );
and \U$35957 ( \36203 , RIbe2b180_117, RIbe2b4c8_124);
nor \U$35958 ( \36204 , RIbe2b180_117, RIbe2b4c8_124);
nor \U$35959 ( \36205 , \36203 , \36204 );
not \U$35960 ( \36206 , \36205 );
not \U$35961 ( \36207 , \34588 );
or \U$35962 ( \36208 , \36206 , \36207 );
not \U$35963 ( \36209 , \36095 );
nand \U$35964 ( \36210 , \36209 , \21759 );
nand \U$35965 ( \36211 , \36208 , \36210 );
not \U$35966 ( \36212 , \36211 );
or \U$35967 ( \36213 , \36202 , \36212 );
or \U$35968 ( \36214 , \36211 , \36201 );
nand \U$35969 ( \36215 , \36213 , \36214 );
not \U$35970 ( \36216 , \36215 );
or \U$35971 ( \36217 , \36192 , \36216 );
not \U$35972 ( \36218 , \36201 );
nand \U$35973 ( \36219 , \36218 , \36211 );
nand \U$35974 ( \36220 , \36217 , \36219 );
not \U$35975 ( \36221 , \36220 );
or \U$35976 ( \36222 , \36187 , \36221 );
or \U$35977 ( \36223 , \36220 , \36186 );
nand \U$35978 ( \36224 , \36222 , \36223 );
not \U$35979 ( \36225 , \36224 );
or \U$35980 ( \36226 , \36184 , \36225 );
not \U$35981 ( \36227 , \36186 );
nand \U$35982 ( \36228 , \36227 , \36220 );
nand \U$35983 ( \36229 , \36226 , \36228 );
not \U$35984 ( \36230 , \36229 );
not \U$35985 ( \36231 , \35923 );
not \U$35986 ( \36232 , \35954 );
not \U$35987 ( \36233 , \36232 );
or \U$35988 ( \36234 , \36231 , \36233 );
nand \U$35989 ( \36235 , \35954 , \35922 );
nand \U$35990 ( \36236 , \36234 , \36235 );
not \U$35991 ( \36237 , \36236 );
xor \U$35992 ( \36238 , \35939 , \35947 );
not \U$35993 ( \36239 , \36238 );
not \U$35994 ( \36240 , RIbe2a640_93);
not \U$35995 ( \36241 , RIbe2b108_116);
and \U$35996 ( \36242 , \36240 , \36241 );
and \U$35997 ( \36243 , RIbe2a640_93, RIbe2b108_116);
nor \U$35998 ( \36244 , \36242 , \36243 );
not \U$35999 ( \36245 , \36244 );
not \U$36000 ( \36246 , \23582 );
or \U$36001 ( \36247 , \36245 , \36246 );
nand \U$36002 ( \36248 , \16875 , \35983 );
nand \U$36003 ( \36249 , \36247 , \36248 );
not \U$36004 ( \36250 , \36249 );
not \U$36005 ( \36251 , RIbe2aaf0_103);
not \U$36006 ( \36252 , RIbe2b2e8_120);
and \U$36007 ( \36253 , \36251 , \36252 );
and \U$36008 ( \36254 , RIbe2aaf0_103, RIbe2b2e8_120);
nor \U$36009 ( \36255 , \36253 , \36254 );
and \U$36010 ( \36256 , \28282 , \36255 );
and \U$36011 ( \36257 , \35977 , RIbe2ab68_104);
nor \U$36012 ( \36258 , \36256 , \36257 );
not \U$36013 ( \36259 , \36258 );
xor \U$36014 ( \36260 , RIbe2a730_95, RIbe2a190_83);
not \U$36015 ( \36261 , \36260 );
not \U$36016 ( \36262 , \14730 );
or \U$36017 ( \36263 , \36261 , \36262 );
nand \U$36018 ( \36264 , \13278 , \36002 );
nand \U$36019 ( \36265 , \36263 , \36264 );
not \U$36020 ( \36266 , \36265 );
or \U$36021 ( \36267 , \36259 , \36266 );
or \U$36022 ( \36268 , \36265 , \36258 );
nand \U$36023 ( \36269 , \36267 , \36268 );
not \U$36024 ( \36270 , \36269 );
or \U$36025 ( \36271 , \36250 , \36270 );
not \U$36026 ( \36272 , \36258 );
nand \U$36027 ( \36273 , \36272 , \36265 );
nand \U$36028 ( \36274 , \36271 , \36273 );
not \U$36029 ( \36275 , \36274 );
not \U$36030 ( \36276 , \35992 );
not \U$36031 ( \36277 , \35974 );
and \U$36032 ( \36278 , \36276 , \36277 );
and \U$36033 ( \36279 , \35992 , \35974 );
nor \U$36034 ( \36280 , \36278 , \36279 );
not \U$36035 ( \36281 , \36280 );
or \U$36036 ( \36282 , \36275 , \36281 );
or \U$36037 ( \36283 , \36280 , \36274 );
nand \U$36038 ( \36284 , \36282 , \36283 );
not \U$36039 ( \36285 , \36284 );
or \U$36040 ( \36286 , \36239 , \36285 );
not \U$36041 ( \36287 , \36280 );
nand \U$36042 ( \36288 , \36287 , \36274 );
nand \U$36043 ( \36289 , \36286 , \36288 );
not \U$36044 ( \36290 , \36289 );
not \U$36045 ( \36291 , \36290 );
or \U$36046 ( \36292 , \36237 , \36291 );
or \U$36047 ( \36293 , \36290 , \36236 );
nand \U$36048 ( \36294 , \36292 , \36293 );
not \U$36049 ( \36295 , \36294 );
or \U$36050 ( \36296 , \36230 , \36295 );
nand \U$36051 ( \36297 , \36289 , \36236 );
nand \U$36052 ( \36298 , \36296 , \36297 );
not \U$36053 ( \36299 , \36298 );
or \U$36054 ( \36300 , \36182 , \36299 );
or \U$36055 ( \36301 , \36298 , \36181 );
nand \U$36056 ( \36302 , \36300 , \36301 );
not \U$36057 ( \36303 , \36302 );
or \U$36058 ( \36304 , \36089 , \36303 );
not \U$36059 ( \36305 , \36181 );
nand \U$36060 ( \36306 , \36305 , \36298 );
nand \U$36061 ( \36307 , \36304 , \36306 );
nor \U$36062 ( \36308 , \36087 , \36307 );
not \U$36063 ( \36309 , \36308 );
xor \U$36064 ( \36310 , \36294 , \36229 );
not \U$36065 ( \36311 , \36177 );
not \U$36066 ( \36312 , \36311 );
not \U$36067 ( \36313 , \36170 );
not \U$36068 ( \36314 , \36313 );
or \U$36069 ( \36315 , \36312 , \36314 );
nand \U$36070 ( \36316 , \36170 , \36177 );
nand \U$36071 ( \36317 , \36315 , \36316 );
or \U$36072 ( \36318 , \36310 , \36317 );
xor \U$36073 ( \36319 , \36215 , \36191 );
not \U$36074 ( \36320 , \36319 );
xor \U$36075 ( \36321 , \36269 , \36249 );
not \U$36076 ( \36322 , \36125 );
not \U$36077 ( \36323 , \36149 );
or \U$36078 ( \36324 , \36322 , \36323 );
or \U$36079 ( \36325 , \36149 , \36125 );
nand \U$36080 ( \36326 , \36324 , \36325 );
xor \U$36081 ( \36327 , \36321 , \36326 );
not \U$36082 ( \36328 , \36327 );
or \U$36083 ( \36329 , \36320 , \36328 );
nand \U$36084 ( \36330 , \36326 , \36321 );
nand \U$36085 ( \36331 , \36329 , \36330 );
not \U$36086 ( \36332 , \36331 );
xor \U$36087 ( \36333 , RIbe2adc0_109, RIbe2b018_114);
not \U$36088 ( \36334 , \36333 );
not \U$36089 ( \36335 , \25897 );
or \U$36090 ( \36336 , \36334 , \36335 );
not \U$36091 ( \36337 , \36196 );
nand \U$36092 ( \36338 , \36337 , \19371 );
nand \U$36093 ( \36339 , \36336 , \36338 );
not \U$36094 ( \36340 , \36339 );
nand \U$36095 ( \36341 , \11456 , RIbe2ae38_110);
not \U$36096 ( \36342 , \36341 );
not \U$36097 ( \36343 , \36342 );
xor \U$36098 ( \36344 , RIbe2b450_123, RIbe2a190_83);
and \U$36099 ( \36345 , \36344 , \15690 );
and \U$36100 ( \36346 , \11400 , \36260 );
nor \U$36101 ( \36347 , \36345 , \36346 );
not \U$36102 ( \36348 , \36347 );
or \U$36103 ( \36349 , \36343 , \36348 );
not \U$36104 ( \36350 , \36341 );
or \U$36105 ( \36351 , \36347 , \36350 );
nand \U$36106 ( \36352 , \36349 , \36351 );
not \U$36107 ( \36353 , \36352 );
or \U$36108 ( \36354 , \36340 , \36353 );
not \U$36109 ( \36355 , \36347 );
nand \U$36110 ( \36356 , \36355 , \36350 );
nand \U$36111 ( \36357 , \36354 , \36356 );
xor \U$36112 ( \36358 , RIbe2af28_112, RIbe2b540_125);
not \U$36113 ( \36359 , \36358 );
not \U$36114 ( \36360 , \15345 );
or \U$36115 ( \36361 , \36359 , \36360 );
nand \U$36116 ( \36362 , \16917 , \36122 );
nand \U$36117 ( \36363 , \36361 , \36362 );
xor \U$36118 ( \36364 , RIbe2a550_91, RIbe2aeb0_111);
not \U$36119 ( \36365 , \36364 );
not \U$36120 ( \36366 , \22975 );
or \U$36121 ( \36367 , \36365 , \36366 );
nand \U$36122 ( \36368 , \10440 , \36104 );
nand \U$36123 ( \36369 , \36367 , \36368 );
or \U$36124 ( \36370 , \36363 , \36369 );
xor \U$36125 ( \36371 , RIbe2b180_117, RIbe2a6b8_94);
not \U$36126 ( \36372 , \36371 );
not \U$36127 ( \36373 , \15353 );
or \U$36128 ( \36374 , \36372 , \36373 );
nand \U$36129 ( \36375 , \14966 , \36205 );
nand \U$36130 ( \36376 , \36374 , \36375 );
nand \U$36131 ( \36377 , \36370 , \36376 );
nand \U$36132 ( \36378 , \36363 , \36369 );
and \U$36133 ( \36379 , \36377 , \36378 );
not \U$36134 ( \36380 , \36379 );
or \U$36135 ( \36381 , \36357 , \36380 );
xnor \U$36136 ( \36382 , RIbe2a7a8_96, RIbe2a280_85);
not \U$36137 ( \36383 , \36382 );
not \U$36138 ( \36384 , \36383 );
not \U$36139 ( \36385 , \14383 );
or \U$36140 ( \36386 , \36384 , \36385 );
nand \U$36141 ( \36387 , \11348 , \36128 );
nand \U$36142 ( \36388 , \36386 , \36387 );
not \U$36143 ( \36389 , \36388 );
not \U$36144 ( \36390 , \19580 );
xnor \U$36145 ( \36391 , RIbe2aaf0_103, RIbe2a4d8_90);
not \U$36146 ( \36392 , \36391 );
and \U$36147 ( \36393 , \36390 , \36392 );
and \U$36148 ( \36394 , \36255 , RIbe2ab68_104);
nor \U$36149 ( \36395 , \36393 , \36394 );
not \U$36150 ( \36396 , \36395 );
xor \U$36151 ( \36397 , RIbe2ac58_106, RIbe2b108_116);
not \U$36152 ( \36398 , \36397 );
not \U$36153 ( \36399 , \25617 );
or \U$36154 ( \36400 , \36398 , \36399 );
nand \U$36155 ( \36401 , \23015 , \36244 );
nand \U$36156 ( \36402 , \36400 , \36401 );
not \U$36157 ( \36403 , \36402 );
or \U$36158 ( \36404 , \36396 , \36403 );
or \U$36159 ( \36405 , \36402 , \36395 );
nand \U$36160 ( \36406 , \36404 , \36405 );
not \U$36161 ( \36407 , \36406 );
or \U$36162 ( \36408 , \36389 , \36407 );
not \U$36163 ( \36409 , \36395 );
nand \U$36164 ( \36410 , \36409 , \36402 );
nand \U$36165 ( \36411 , \36408 , \36410 );
nand \U$36166 ( \36412 , \36381 , \36411 );
nand \U$36167 ( \36413 , \36357 , \36380 );
and \U$36168 ( \36414 , \36412 , \36413 );
not \U$36169 ( \36415 , \36414 );
not \U$36170 ( \36416 , \36238 );
not \U$36171 ( \36417 , \36284 );
not \U$36172 ( \36418 , \36417 );
or \U$36173 ( \36419 , \36416 , \36418 );
not \U$36174 ( \36420 , \36238 );
nand \U$36175 ( \36421 , \36420 , \36284 );
nand \U$36176 ( \36422 , \36419 , \36421 );
not \U$36177 ( \36423 , \36422 );
or \U$36178 ( \36424 , \36415 , \36423 );
or \U$36179 ( \36425 , \36422 , \36414 );
nand \U$36180 ( \36426 , \36424 , \36425 );
not \U$36181 ( \36427 , \36426 );
or \U$36182 ( \36428 , \36332 , \36427 );
not \U$36183 ( \36429 , \36414 );
nand \U$36184 ( \36430 , \36429 , \36422 );
nand \U$36185 ( \36431 , \36428 , \36430 );
nand \U$36186 ( \36432 , \36318 , \36431 );
nand \U$36187 ( \36433 , \36310 , \36317 );
nand \U$36188 ( \36434 , \36432 , \36433 );
not \U$36189 ( \36435 , \36088 );
not \U$36190 ( \36436 , \36435 );
not \U$36191 ( \36437 , \36302 );
or \U$36192 ( \36438 , \36436 , \36437 );
or \U$36193 ( \36439 , \36302 , \36435 );
nand \U$36194 ( \36440 , \36438 , \36439 );
or \U$36195 ( \36441 , \36434 , \36440 );
and \U$36196 ( \36442 , \36085 , \36309 , \36441 );
not \U$36197 ( \36443 , \36442 );
not \U$36198 ( \36444 , \36331 );
and \U$36199 ( \36445 , \36426 , \36444 );
not \U$36200 ( \36446 , \36426 );
and \U$36201 ( \36447 , \36446 , \36331 );
nor \U$36202 ( \36448 , \36445 , \36447 );
not \U$36203 ( \36449 , \36448 );
not \U$36204 ( \36450 , \36449 );
xor \U$36205 ( \36451 , \36224 , \36183 );
not \U$36206 ( \36452 , \36451 );
xor \U$36207 ( \36453 , \36379 , \36357 );
xnor \U$36208 ( \36454 , \36453 , \36411 );
not \U$36209 ( \36455 , \36454 );
not \U$36210 ( \36456 , \36406 );
and \U$36211 ( \36457 , \36388 , \36456 );
not \U$36212 ( \36458 , \36388 );
and \U$36213 ( \36459 , \36458 , \36406 );
nor \U$36214 ( \36460 , \36457 , \36459 );
not \U$36215 ( \36461 , \36460 );
not \U$36216 ( \36462 , \36461 );
not \U$36217 ( \36463 , \36352 );
not \U$36218 ( \36464 , \36339 );
not \U$36219 ( \36465 , \36464 );
and \U$36220 ( \36466 , \36463 , \36465 );
and \U$36221 ( \36467 , \36352 , \36464 );
nor \U$36222 ( \36468 , \36466 , \36467 );
not \U$36223 ( \36469 , \36468 );
not \U$36224 ( \36470 , \36469 );
or \U$36225 ( \36471 , \36462 , \36470 );
not \U$36226 ( \36472 , \36468 );
not \U$36227 ( \36473 , \36460 );
or \U$36228 ( \36474 , \36472 , \36473 );
xor \U$36229 ( \36475 , \36363 , \36369 );
xor \U$36230 ( \36476 , \36475 , \36376 );
nand \U$36231 ( \36477 , \36474 , \36476 );
nand \U$36232 ( \36478 , \36471 , \36477 );
not \U$36233 ( \36479 , \36478 );
not \U$36234 ( \36480 , \36479 );
not \U$36235 ( \36481 , \36358 );
not \U$36236 ( \36482 , \15348 );
or \U$36237 ( \36483 , \36481 , \36482 );
and \U$36238 ( \36484 , RIbe2af28_112, RIbe2b4c8_124);
nor \U$36239 ( \36485 , RIbe2af28_112, RIbe2b4c8_124);
nor \U$36240 ( \36486 , \36484 , \36485 );
nand \U$36241 ( \36487 , \18649 , \36486 );
nand \U$36242 ( \36488 , \36483 , \36487 );
not \U$36243 ( \36489 , \36488 );
xor \U$36244 ( \36490 , RIbe2a730_95, RIbe2a280_85);
and \U$36245 ( \36491 , \27993 , \36490 );
not \U$36246 ( \36492 , \11348 );
nor \U$36247 ( \36493 , \36492 , \36382 );
nor \U$36248 ( \36494 , \36491 , \36493 );
not \U$36249 ( \36495 , \36494 );
xor \U$36250 ( \36496 , RIbe2b180_117, RIbe2a640_93);
not \U$36251 ( \36497 , \36496 );
not \U$36252 ( \36498 , \14852 );
or \U$36253 ( \36499 , \36497 , \36498 );
nand \U$36254 ( \36500 , \21759 , \36371 );
nand \U$36255 ( \36501 , \36499 , \36500 );
not \U$36256 ( \36502 , \36501 );
and \U$36257 ( \36503 , \36495 , \36502 );
and \U$36258 ( \36504 , \36501 , \36494 );
nor \U$36259 ( \36505 , \36503 , \36504 );
not \U$36260 ( \36506 , \36505 );
not \U$36261 ( \36507 , \36506 );
or \U$36262 ( \36508 , \36489 , \36507 );
not \U$36263 ( \36509 , \36494 );
nand \U$36264 ( \36510 , \36509 , \36501 );
nand \U$36265 ( \36511 , \36508 , \36510 );
not \U$36266 ( \36512 , \36511 );
not \U$36267 ( \36513 , \34550 );
not \U$36268 ( \36514 , \36513 );
xor \U$36269 ( \36515 , RIbe2aaf0_103, RIbe2a460_89);
not \U$36270 ( \36516 , \36515 );
or \U$36271 ( \36517 , \36514 , \36516 );
or \U$36272 ( \36518 , \18830 , \36391 );
nand \U$36273 ( \36519 , \36517 , \36518 );
not \U$36274 ( \36520 , \36519 );
xor \U$36275 ( \36521 , RIbe2ad48_108, RIbe2b018_114);
not \U$36276 ( \36522 , \36521 );
not \U$36277 ( \36523 , \22763 );
or \U$36278 ( \36524 , \36522 , \36523 );
nand \U$36279 ( \36525 , \15953 , \36333 );
nand \U$36280 ( \36526 , \36524 , \36525 );
not \U$36281 ( \36527 , \36526 );
not \U$36282 ( \36528 , \36527 );
not \U$36283 ( \36529 , RIbe2abe0_105);
not \U$36284 ( \36530 , RIbe2b108_116);
and \U$36285 ( \36531 , \36529 , \36530 );
and \U$36286 ( \36532 , RIbe2abe0_105, RIbe2b108_116);
nor \U$36287 ( \36533 , \36531 , \36532 );
not \U$36288 ( \36534 , \36533 );
not \U$36289 ( \36535 , \14297 );
or \U$36290 ( \36536 , \36534 , \36535 );
nand \U$36291 ( \36537 , \16898 , \36397 );
nand \U$36292 ( \36538 , \36536 , \36537 );
not \U$36293 ( \36539 , \36538 );
or \U$36294 ( \36540 , \36528 , \36539 );
not \U$36295 ( \36541 , \36526 );
or \U$36296 ( \36542 , \36538 , \36541 );
nand \U$36297 ( \36543 , \36540 , \36542 );
not \U$36298 ( \36544 , \36543 );
or \U$36299 ( \36545 , \36520 , \36544 );
nand \U$36300 ( \36546 , \36538 , \36526 );
nand \U$36301 ( \36547 , \36545 , \36546 );
xor \U$36302 ( \36548 , RIbe2b3d8_122, RIbe2a190_83);
not \U$36303 ( \36549 , \36548 );
not \U$36304 ( \36550 , \15690 );
or \U$36305 ( \36551 , \36549 , \36550 );
nand \U$36306 ( \36552 , \11400 , \36344 );
nand \U$36307 ( \36553 , \36551 , \36552 );
or \U$36308 ( \36554 , RIbe2a190_83, RIbe2a5c8_92);
nand \U$36309 ( \36555 , \36554 , RIbe2ae38_110);
nand \U$36310 ( \36556 , RIbe2a190_83, RIbe2a5c8_92);
and \U$36311 ( \36557 , \36555 , \36556 , RIbe2a550_91);
nand \U$36312 ( \36558 , \36553 , \36557 );
not \U$36313 ( \36559 , \36558 );
and \U$36314 ( \36560 , \36547 , \36559 );
not \U$36315 ( \36561 , \36547 );
and \U$36316 ( \36562 , \36561 , \36558 );
nor \U$36317 ( \36563 , \36560 , \36562 );
not \U$36318 ( \36564 , \36563 );
or \U$36319 ( \36565 , \36512 , \36564 );
nand \U$36320 ( \36566 , \36547 , \36559 );
nand \U$36321 ( \36567 , \36565 , \36566 );
not \U$36322 ( \36568 , \36567 );
or \U$36323 ( \36569 , \36480 , \36568 );
or \U$36324 ( \36570 , \36567 , \36479 );
nand \U$36325 ( \36571 , \36569 , \36570 );
not \U$36326 ( \36572 , \36571 );
or \U$36327 ( \36573 , \36455 , \36572 );
not \U$36328 ( \36574 , \36479 );
nand \U$36329 ( \36575 , \36574 , \36567 );
nand \U$36330 ( \36576 , \36573 , \36575 );
not \U$36331 ( \36577 , \36576 );
not \U$36332 ( \36578 , \36577 );
or \U$36333 ( \36579 , \36452 , \36578 );
not \U$36334 ( \36580 , \36451 );
nand \U$36335 ( \36581 , \36580 , \36576 );
nand \U$36336 ( \36582 , \36579 , \36581 );
not \U$36337 ( \36583 , \36582 );
or \U$36338 ( \36584 , \36450 , \36583 );
nand \U$36339 ( \36585 , \36576 , \36451 );
nand \U$36340 ( \36586 , \36584 , \36585 );
not \U$36341 ( \36587 , \36586 );
xor \U$36342 ( \36588 , \36317 , \36431 );
xnor \U$36343 ( \36589 , \36588 , \36310 );
nand \U$36344 ( \36590 , \36587 , \36589 );
not \U$36345 ( \36591 , \36582 );
not \U$36346 ( \36592 , \36448 );
and \U$36347 ( \36593 , \36591 , \36592 );
and \U$36348 ( \36594 , \36582 , \36448 );
nor \U$36349 ( \36595 , \36593 , \36594 );
buf \U$36350 ( \36596 , \36571 );
not \U$36351 ( \36597 , \36454 );
and \U$36352 ( \36598 , \36596 , \36597 );
not \U$36353 ( \36599 , \36596 );
and \U$36354 ( \36600 , \36599 , \36454 );
nor \U$36355 ( \36601 , \36598 , \36600 );
not \U$36356 ( \36602 , \36601 );
not \U$36357 ( \36603 , \36602 );
xor \U$36358 ( \36604 , \36327 , \36319 );
not \U$36359 ( \36605 , \36604 );
buf \U$36360 ( \36606 , \36563 );
and \U$36361 ( \36607 , \36606 , \36511 );
not \U$36362 ( \36608 , \36606 );
not \U$36363 ( \36609 , \36511 );
and \U$36364 ( \36610 , \36608 , \36609 );
nor \U$36365 ( \36611 , \36607 , \36610 );
not \U$36366 ( \36612 , \36611 );
not \U$36367 ( \36613 , \36543 );
not \U$36368 ( \36614 , \36519 );
not \U$36369 ( \36615 , \36614 );
and \U$36370 ( \36616 , \36613 , \36615 );
and \U$36371 ( \36617 , \36543 , \36614 );
nor \U$36372 ( \36618 , \36616 , \36617 );
not \U$36373 ( \36619 , \36618 );
not \U$36374 ( \36620 , \20396 );
xnor \U$36375 ( \36621 , RIbe2b540_125, RIbe2b018_114);
or \U$36376 ( \36622 , \36620 , \36621 );
not \U$36377 ( \36623 , \36521 );
or \U$36378 ( \36624 , \25891 , \36623 );
nand \U$36379 ( \36625 , \36622 , \36624 );
not \U$36380 ( \36626 , \36625 );
not \U$36381 ( \36627 , \19580 );
xnor \U$36382 ( \36628 , RIbe2aaf0_103, RIbe2adc0_109);
not \U$36383 ( \36629 , \36628 );
and \U$36384 ( \36630 , \36627 , \36629 );
and \U$36385 ( \36631 , \36515 , RIbe2ab68_104);
nor \U$36386 ( \36632 , \36630 , \36631 );
not \U$36387 ( \36633 , \36632 );
xor \U$36388 ( \36634 , RIbe2b108_116, RIbe2a7a8_96);
not \U$36389 ( \36635 , \36634 );
not \U$36390 ( \36636 , \14297 );
or \U$36391 ( \36637 , \36635 , \36636 );
nand \U$36392 ( \36638 , \13534 , \36533 );
nand \U$36393 ( \36639 , \36637 , \36638 );
not \U$36394 ( \36640 , \36639 );
or \U$36395 ( \36641 , \36633 , \36640 );
or \U$36396 ( \36642 , \36639 , \36632 );
nand \U$36397 ( \36643 , \36641 , \36642 );
not \U$36398 ( \36644 , \36643 );
or \U$36399 ( \36645 , \36626 , \36644 );
not \U$36400 ( \36646 , \36632 );
nand \U$36401 ( \36647 , \36646 , \36639 );
nand \U$36402 ( \36648 , \36645 , \36647 );
not \U$36403 ( \36649 , \36648 );
not \U$36404 ( \36650 , \36649 );
or \U$36405 ( \36651 , \36619 , \36650 );
not \U$36406 ( \36652 , \36488 );
not \U$36407 ( \36653 , \36505 );
or \U$36408 ( \36654 , \36652 , \36653 );
or \U$36409 ( \36655 , \36505 , \36488 );
nand \U$36410 ( \36656 , \36654 , \36655 );
nand \U$36411 ( \36657 , \36651 , \36656 );
not \U$36412 ( \36658 , \36618 );
nand \U$36413 ( \36659 , \36648 , \36658 );
and \U$36414 ( \36660 , \36657 , \36659 );
not \U$36415 ( \36661 , RIbe2a6b8_94);
not \U$36416 ( \36662 , RIbe2af28_112);
and \U$36417 ( \36663 , \36661 , \36662 );
and \U$36418 ( \36664 , RIbe2a6b8_94, RIbe2af28_112);
nor \U$36419 ( \36665 , \36663 , \36664 );
not \U$36420 ( \36666 , \36665 );
not \U$36421 ( \36667 , \35366 );
or \U$36422 ( \36668 , \36666 , \36667 );
nand \U$36423 ( \36669 , \19721 , \36486 );
nand \U$36424 ( \36670 , \36668 , \36669 );
not \U$36425 ( \36671 , \36670 );
nand \U$36426 ( \36672 , \11228 , RIbe2ae38_110);
not \U$36427 ( \36673 , \36672 );
xor \U$36428 ( \36674 , RIbe2b450_123, RIbe2a280_85);
not \U$36429 ( \36675 , \36674 );
not \U$36430 ( \36676 , \24028 );
or \U$36431 ( \36677 , \36675 , \36676 );
nand \U$36432 ( \36678 , \11348 , \36490 );
nand \U$36433 ( \36679 , \36677 , \36678 );
not \U$36434 ( \36680 , \36679 );
or \U$36435 ( \36681 , \36673 , \36680 );
or \U$36436 ( \36682 , \36679 , \36672 );
nand \U$36437 ( \36683 , \36681 , \36682 );
not \U$36438 ( \36684 , \36683 );
or \U$36439 ( \36685 , \36671 , \36684 );
not \U$36440 ( \36686 , \36672 );
nand \U$36441 ( \36687 , \36686 , \36679 );
nand \U$36442 ( \36688 , \36685 , \36687 );
not \U$36443 ( \36689 , \36688 );
xor \U$36444 ( \36690 , \36557 , \36553 );
not \U$36445 ( \36691 , \36690 );
xor \U$36446 ( \36692 , RIbe2a550_91, RIbe2ae38_110);
not \U$36447 ( \36693 , \36692 );
not \U$36448 ( \36694 , \10434 );
or \U$36449 ( \36695 , \36693 , \36694 );
nand \U$36450 ( \36696 , \11228 , \36364 );
nand \U$36451 ( \36697 , \36695 , \36696 );
not \U$36452 ( \36698 , \36697 );
nand \U$36453 ( \36699 , \36691 , \36698 );
not \U$36454 ( \36700 , \36699 );
or \U$36455 ( \36701 , \36689 , \36700 );
not \U$36456 ( \36702 , \36698 );
nand \U$36457 ( \36703 , \36702 , \36690 );
nand \U$36458 ( \36704 , \36701 , \36703 );
not \U$36459 ( \36705 , \36704 );
and \U$36460 ( \36706 , \36660 , \36705 );
not \U$36461 ( \36707 , \36660 );
and \U$36462 ( \36708 , \36707 , \36704 );
nor \U$36463 ( \36709 , \36706 , \36708 );
not \U$36464 ( \36710 , \36709 );
or \U$36465 ( \36711 , \36612 , \36710 );
not \U$36466 ( \36712 , \36660 );
nand \U$36467 ( \36713 , \36712 , \36704 );
nand \U$36468 ( \36714 , \36711 , \36713 );
not \U$36469 ( \36715 , \36714 );
not \U$36470 ( \36716 , \36715 );
or \U$36471 ( \36717 , \36605 , \36716 );
not \U$36472 ( \36718 , \36714 );
or \U$36473 ( \36719 , \36718 , \36604 );
nand \U$36474 ( \36720 , \36717 , \36719 );
not \U$36475 ( \36721 , \36720 );
or \U$36476 ( \36722 , \36603 , \36721 );
not \U$36477 ( \36723 , \36718 );
nand \U$36478 ( \36724 , \36723 , \36604 );
nand \U$36479 ( \36725 , \36722 , \36724 );
not \U$36480 ( \36726 , \36725 );
nand \U$36481 ( \36727 , \36595 , \36726 );
nand \U$36482 ( \36728 , \36590 , \36727 );
not \U$36483 ( \36729 , \36728 );
xnor \U$36484 ( \36730 , RIbe2b540_125, RIbe2aaf0_103);
not \U$36485 ( \36731 , \36730 );
not \U$36486 ( \36732 , \36731 );
not \U$36487 ( \36733 , \36513 );
or \U$36488 ( \36734 , \36732 , \36733 );
xor \U$36489 ( \36735 , RIbe2ad48_108, RIbe2aaf0_103);
nand \U$36490 ( \36736 , \36735 , RIbe2ab68_104);
nand \U$36491 ( \36737 , \36734 , \36736 );
not \U$36492 ( \36738 , \36737 );
xor \U$36493 ( \36739 , RIbe2ac58_106, RIbe2af28_112);
not \U$36494 ( \36740 , \36739 );
not \U$36495 ( \36741 , \16914 );
or \U$36496 ( \36742 , \36740 , \36741 );
xor \U$36497 ( \36743 , RIbe2af28_112, RIbe2a640_93);
nand \U$36498 ( \36744 , \16917 , \36743 );
nand \U$36499 ( \36745 , \36742 , \36744 );
not \U$36500 ( \36746 , \36745 );
or \U$36501 ( \36747 , \36738 , \36746 );
or \U$36502 ( \36748 , \36745 , \36737 );
xor \U$36503 ( \36749 , RIbe2a280_85, RIbe2aeb0_111);
not \U$36504 ( \36750 , \36749 );
not \U$36505 ( \36751 , \36010 );
or \U$36506 ( \36752 , \36750 , \36751 );
xor \U$36507 ( \36753 , RIbe2a280_85, RIbe2b3d8_122);
nand \U$36508 ( \36754 , \11348 , \36753 );
nand \U$36509 ( \36755 , \36752 , \36754 );
nand \U$36510 ( \36756 , \36748 , \36755 );
nand \U$36511 ( \36757 , \36747 , \36756 );
not \U$36512 ( \36758 , \36753 );
not \U$36513 ( \36759 , \36010 );
or \U$36514 ( \36760 , \36758 , \36759 );
nand \U$36515 ( \36761 , \14649 , \36674 );
nand \U$36516 ( \36762 , \36760 , \36761 );
or \U$36517 ( \36763 , RIbe2a208_84, RIbe2a280_85);
nand \U$36518 ( \36764 , \36763 , RIbe2ae38_110);
nand \U$36519 ( \36765 , RIbe2a208_84, RIbe2a280_85);
and \U$36520 ( \36766 , \36764 , \36765 , RIbe2a190_83);
or \U$36521 ( \36767 , \36762 , \36766 );
nand \U$36522 ( \36768 , \36762 , \36766 );
and \U$36523 ( \36769 , \36767 , \36768 );
xor \U$36524 ( \36770 , \36757 , \36769 );
xor \U$36525 ( \36771 , RIbe2b180_117, RIbe2a7a8_96);
not \U$36526 ( \36772 , \36771 );
buf \U$36527 ( \36773 , \15353 );
not \U$36528 ( \36774 , \36773 );
or \U$36529 ( \36775 , \36772 , \36774 );
xnor \U$36530 ( \36776 , RIbe2abe0_105, RIbe2b180_117);
not \U$36531 ( \36777 , \36776 );
nand \U$36532 ( \36778 , \36777 , \14966 );
nand \U$36533 ( \36779 , \36775 , \36778 );
not \U$36534 ( \36780 , \36779 );
nand \U$36535 ( \36781 , \31948 , RIbe2ae38_110);
not \U$36536 ( \36782 , \36781 );
and \U$36537 ( \36783 , \36780 , \36782 );
and \U$36538 ( \36784 , \36779 , \36781 );
nor \U$36539 ( \36785 , \36783 , \36784 );
xor \U$36540 ( \36786 , RIbe2b108_116, RIbe2b450_123);
not \U$36541 ( \36787 , \36786 );
not \U$36542 ( \36788 , \23582 );
or \U$36543 ( \36789 , \36787 , \36788 );
xor \U$36544 ( \36790 , RIbe2a730_95, RIbe2b108_116);
nand \U$36545 ( \36791 , \13534 , \36790 );
nand \U$36546 ( \36792 , \36789 , \36791 );
not \U$36547 ( \36793 , \36792 );
or \U$36548 ( \36794 , \36785 , \36793 );
not \U$36549 ( \36795 , \36781 );
nand \U$36550 ( \36796 , \36795 , \36779 );
nand \U$36551 ( \36797 , \36794 , \36796 );
and \U$36552 ( \36798 , \36770 , \36797 );
and \U$36553 ( \36799 , \36757 , \36769 );
or \U$36554 ( \36800 , \36798 , \36799 );
xnor \U$36555 ( \36801 , \36643 , \36625 );
not \U$36556 ( \36802 , \36801 );
not \U$36557 ( \36803 , \14730 );
not \U$36558 ( \36804 , \36803 );
xnor \U$36559 ( \36805 , RIbe2aeb0_111, RIbe2a190_83);
not \U$36560 ( \36806 , \36805 );
and \U$36561 ( \36807 , \36804 , \36806 );
and \U$36562 ( \36808 , \15693 , \36548 );
nor \U$36563 ( \36809 , \36807 , \36808 );
not \U$36564 ( \36810 , \36809 );
xnor \U$36565 ( \36811 , RIbe2b180_117, RIbe2ac58_106);
not \U$36566 ( \36812 , \36811 );
not \U$36567 ( \36813 , \36812 );
not \U$36568 ( \36814 , \32900 );
or \U$36569 ( \36815 , \36813 , \36814 );
nand \U$36570 ( \36816 , \21759 , \36496 );
nand \U$36571 ( \36817 , \36815 , \36816 );
not \U$36572 ( \36818 , \36817 );
or \U$36573 ( \36819 , \36810 , \36818 );
or \U$36574 ( \36820 , \36817 , \36809 );
nand \U$36575 ( \36821 , \36819 , \36820 );
and \U$36576 ( \36822 , \36821 , \36768 );
not \U$36577 ( \36823 , \36821 );
not \U$36578 ( \36824 , \36768 );
and \U$36579 ( \36825 , \36823 , \36824 );
or \U$36580 ( \36826 , \36822 , \36825 );
not \U$36581 ( \36827 , \36826 );
or \U$36582 ( \36828 , \36802 , \36827 );
or \U$36583 ( \36829 , \36826 , \36801 );
nand \U$36584 ( \36830 , \36828 , \36829 );
not \U$36585 ( \36831 , \36830 );
and \U$36586 ( \36832 , \36800 , \36831 );
not \U$36587 ( \36833 , \36800 );
and \U$36588 ( \36834 , \36833 , \36830 );
nor \U$36589 ( \36835 , \36832 , \36834 );
not \U$36590 ( \36836 , \36835 );
not \U$36591 ( \36837 , \15690 );
and \U$36592 ( \36838 , \24871 , RIbe2a190_83);
not \U$36593 ( \36839 , RIbe2a190_83);
and \U$36594 ( \36840 , \36839 , RIbe2ae38_110);
nor \U$36595 ( \36841 , \36838 , \36840 );
or \U$36596 ( \36842 , \36837 , \36841 );
or \U$36597 ( \36843 , \11971 , \36805 );
nand \U$36598 ( \36844 , \36842 , \36843 );
not \U$36599 ( \36845 , \36844 );
or \U$36600 ( \36846 , \24450 , \36776 );
not \U$36601 ( \36847 , \14966 );
or \U$36602 ( \36848 , \36847 , \36811 );
nand \U$36603 ( \36849 , \36846 , \36848 );
not \U$36604 ( \36850 , \36849 );
xor \U$36605 ( \36851 , RIbe2b4c8_124, RIbe2b018_114);
not \U$36606 ( \36852 , \36851 );
not \U$36607 ( \36853 , \15967 );
or \U$36608 ( \36854 , \36852 , \36853 );
not \U$36609 ( \36855 , \36621 );
nand \U$36610 ( \36856 , \36855 , \20583 );
nand \U$36611 ( \36857 , \36854 , \36856 );
not \U$36612 ( \36858 , \36857 );
and \U$36613 ( \36859 , \36850 , \36858 );
not \U$36614 ( \36860 , \36850 );
and \U$36615 ( \36861 , \36860 , \36857 );
nor \U$36616 ( \36862 , \36859 , \36861 );
not \U$36617 ( \36863 , \36862 );
or \U$36618 ( \36864 , \36845 , \36863 );
nand \U$36619 ( \36865 , \36849 , \36857 );
nand \U$36620 ( \36866 , \36864 , \36865 );
not \U$36621 ( \36867 , \36866 );
not \U$36622 ( \36868 , \36670 );
not \U$36623 ( \36869 , \36868 );
not \U$36624 ( \36870 , \36683 );
or \U$36625 ( \36871 , \36869 , \36870 );
or \U$36626 ( \36872 , \36683 , \36868 );
nand \U$36627 ( \36873 , \36871 , \36872 );
not \U$36628 ( \36874 , \36873 );
not \U$36629 ( \36875 , \36874 );
or \U$36630 ( \36876 , \36867 , \36875 );
not \U$36631 ( \36877 , \36866 );
nand \U$36632 ( \36878 , \36877 , \36873 );
nand \U$36633 ( \36879 , \36876 , \36878 );
not \U$36634 ( \36880 , \36879 );
not \U$36635 ( \36881 , \36735 );
not \U$36636 ( \36882 , \19581 );
or \U$36637 ( \36883 , \36881 , \36882 );
not \U$36638 ( \36884 , \36628 );
nand \U$36639 ( \36885 , \36884 , RIbe2ab68_104);
nand \U$36640 ( \36886 , \36883 , \36885 );
not \U$36641 ( \36887 , \36743 );
not \U$36642 ( \36888 , \15345 );
or \U$36643 ( \36889 , \36887 , \36888 );
nand \U$36644 ( \36890 , \17811 , \36665 );
nand \U$36645 ( \36891 , \36889 , \36890 );
xor \U$36646 ( \36892 , \36886 , \36891 );
not \U$36647 ( \36893 , \36790 );
not \U$36648 ( \36894 , \21852 );
or \U$36649 ( \36895 , \36893 , \36894 );
nand \U$36650 ( \36896 , \13534 , \36634 );
nand \U$36651 ( \36897 , \36895 , \36896 );
and \U$36652 ( \36898 , \36892 , \36897 );
and \U$36653 ( \36899 , \36886 , \36891 );
or \U$36654 ( \36900 , \36898 , \36899 );
not \U$36655 ( \36901 , \36900 );
not \U$36656 ( \36902 , \36901 );
and \U$36657 ( \36903 , \36880 , \36902 );
and \U$36658 ( \36904 , \36879 , \36901 );
nor \U$36659 ( \36905 , \36903 , \36904 );
not \U$36660 ( \36906 , \36905 );
or \U$36661 ( \36907 , \36836 , \36906 );
xor \U$36662 ( \36908 , \36886 , \36891 );
xor \U$36663 ( \36909 , \36908 , \36897 );
xor \U$36664 ( \36910 , \36844 , \36862 );
xor \U$36665 ( \36911 , \36909 , \36910 );
not \U$36666 ( \36912 , \15345 );
xnor \U$36667 ( \36913 , RIbe2abe0_105, RIbe2af28_112);
or \U$36668 ( \36914 , \36912 , \36913 );
not \U$36669 ( \36915 , \17811 );
not \U$36670 ( \36916 , \36739 );
or \U$36671 ( \36917 , \36915 , \36916 );
nand \U$36672 ( \36918 , \36914 , \36917 );
not \U$36673 ( \36919 , \36918 );
and \U$36674 ( \36920 , RIbe2a280_85, RIbe2ae38_110);
not \U$36675 ( \36921 , RIbe2a280_85);
and \U$36676 ( \36922 , \36921 , \24871 );
nor \U$36677 ( \36923 , \36920 , \36922 );
not \U$36678 ( \36924 , \36923 );
not \U$36679 ( \36925 , \36010 );
or \U$36680 ( \36926 , \36924 , \36925 );
nand \U$36681 ( \36927 , \14649 , \36749 );
nand \U$36682 ( \36928 , \36926 , \36927 );
not \U$36683 ( \36929 , \36928 );
xor \U$36684 ( \36930 , RIbe2b180_117, RIbe2a730_95);
not \U$36685 ( \36931 , \36930 );
nor \U$36686 ( \36932 , \36931 , \14853 );
not \U$36687 ( \36933 , \36771 );
nor \U$36688 ( \36934 , \36933 , \36847 );
nor \U$36689 ( \36935 , \36932 , \36934 );
not \U$36690 ( \36936 , \36935 );
or \U$36691 ( \36937 , \36929 , \36936 );
or \U$36692 ( \36938 , \36935 , \36928 );
nand \U$36693 ( \36939 , \36937 , \36938 );
not \U$36694 ( \36940 , \36939 );
or \U$36695 ( \36941 , \36919 , \36940 );
not \U$36696 ( \36942 , \36935 );
nand \U$36697 ( \36943 , \36942 , \36928 );
nand \U$36698 ( \36944 , \36941 , \36943 );
not \U$36699 ( \36945 , \36944 );
not \U$36700 ( \36946 , \34558 );
not \U$36701 ( \36947 , RIbe2a6b8_94);
not \U$36702 ( \36948 , RIbe2b018_114);
and \U$36703 ( \36949 , \36947 , \36948 );
and \U$36704 ( \36950 , RIbe2a6b8_94, RIbe2b018_114);
nor \U$36705 ( \36951 , \36949 , \36950 );
not \U$36706 ( \36952 , \36951 );
not \U$36707 ( \36953 , \36952 );
and \U$36708 ( \36954 , \36946 , \36953 );
buf \U$36709 ( \36955 , \19371 );
and \U$36710 ( \36956 , \36955 , \36851 );
nor \U$36711 ( \36957 , \36954 , \36956 );
not \U$36712 ( \36958 , \36957 );
xor \U$36713 ( \36959 , RIbe2b108_116, RIbe2b3d8_122);
not \U$36714 ( \36960 , \36959 );
not \U$36715 ( \36961 , \13543 );
or \U$36716 ( \36962 , \36960 , \36961 );
nand \U$36717 ( \36963 , \23015 , \36786 );
nand \U$36718 ( \36964 , \36962 , \36963 );
or \U$36719 ( \36965 , RIbe2ae38_110, RIbe2b090_115);
nand \U$36720 ( \36966 , \36965 , RIbe2b108_116);
nand \U$36721 ( \36967 , RIbe2ae38_110, RIbe2b090_115);
and \U$36722 ( \36968 , \36966 , \36967 , RIbe2a280_85);
and \U$36723 ( \36969 , \36964 , \36968 );
not \U$36724 ( \36970 , \36969 );
or \U$36725 ( \36971 , \36958 , \36970 );
or \U$36726 ( \36972 , \36969 , \36957 );
nand \U$36727 ( \36973 , \36971 , \36972 );
not \U$36728 ( \36974 , \36973 );
or \U$36729 ( \36975 , \36945 , \36974 );
not \U$36730 ( \36976 , \36957 );
nand \U$36731 ( \36977 , \36976 , \36969 );
nand \U$36732 ( \36978 , \36975 , \36977 );
and \U$36733 ( \36979 , \36911 , \36978 );
and \U$36734 ( \36980 , \36909 , \36910 );
or \U$36735 ( \36981 , \36979 , \36980 );
nand \U$36736 ( \36982 , \36907 , \36981 );
or \U$36737 ( \36983 , \36905 , \36835 );
nand \U$36738 ( \36984 , \36982 , \36983 );
not \U$36739 ( \36985 , \36984 );
buf \U$36740 ( \36986 , \36658 );
not \U$36741 ( \36987 , \36986 );
not \U$36742 ( \36988 , \36649 );
not \U$36743 ( \36989 , \36656 );
or \U$36744 ( \36990 , \36988 , \36989 );
or \U$36745 ( \36991 , \36656 , \36649 );
nand \U$36746 ( \36992 , \36990 , \36991 );
not \U$36747 ( \36993 , \36992 );
or \U$36748 ( \36994 , \36987 , \36993 );
or \U$36749 ( \36995 , \36992 , \36986 );
nand \U$36750 ( \36996 , \36994 , \36995 );
not \U$36751 ( \36997 , \36996 );
not \U$36752 ( \36998 , \36830 );
not \U$36753 ( \36999 , \36800 );
or \U$36754 ( \37000 , \36998 , \36999 );
not \U$36755 ( \37001 , \36801 );
nand \U$36756 ( \37002 , \37001 , \36826 );
nand \U$36757 ( \37003 , \37000 , \37002 );
not \U$36758 ( \37004 , \37003 );
or \U$36759 ( \37005 , \36997 , \37004 );
or \U$36760 ( \37006 , \37003 , \36996 );
nand \U$36761 ( \37007 , \37005 , \37006 );
not \U$36762 ( \37008 , \37007 );
not \U$36763 ( \37009 , \36900 );
not \U$36764 ( \37010 , \36879 );
or \U$36765 ( \37011 , \37009 , \37010 );
nand \U$36766 ( \37012 , \36873 , \36866 );
nand \U$36767 ( \37013 , \37011 , \37012 );
not \U$36768 ( \37014 , \37013 );
and \U$36769 ( \37015 , \36690 , \36697 );
not \U$36770 ( \37016 , \36690 );
and \U$36771 ( \37017 , \37016 , \36698 );
nor \U$36772 ( \37018 , \37015 , \37017 );
not \U$36773 ( \37019 , \37018 );
not \U$36774 ( \37020 , \36688 );
and \U$36775 ( \37021 , \37019 , \37020 );
and \U$36776 ( \37022 , \37018 , \36688 );
nor \U$36777 ( \37023 , \37021 , \37022 );
not \U$36778 ( \37024 , \37023 );
not \U$36779 ( \37025 , \36824 );
not \U$36780 ( \37026 , \36821 );
or \U$36781 ( \37027 , \37025 , \37026 );
not \U$36782 ( \37028 , \36809 );
nand \U$36783 ( \37029 , \37028 , \36817 );
nand \U$36784 ( \37030 , \37027 , \37029 );
not \U$36785 ( \37031 , \37030 );
nand \U$36786 ( \37032 , \37024 , \37031 );
not \U$36787 ( \37033 , \37031 );
nand \U$36788 ( \37034 , \37033 , \37023 );
nand \U$36789 ( \37035 , \37032 , \37034 );
not \U$36790 ( \37036 , \37035 );
not \U$36791 ( \37037 , \37036 );
and \U$36792 ( \37038 , \37014 , \37037 );
not \U$36793 ( \37039 , \37035 );
and \U$36794 ( \37040 , \37013 , \37039 );
nor \U$36795 ( \37041 , \37038 , \37040 );
not \U$36796 ( \37042 , \37041 );
or \U$36797 ( \37043 , \37008 , \37042 );
or \U$36798 ( \37044 , \37041 , \37007 );
nand \U$36799 ( \37045 , \37043 , \37044 );
nand \U$36800 ( \37046 , \36985 , \37045 );
xor \U$36801 ( \37047 , \36981 , \36905 );
xnor \U$36802 ( \37048 , \37047 , \36835 );
and \U$36803 ( \37049 , \36785 , \36792 );
not \U$36804 ( \37050 , \36785 );
and \U$36805 ( \37051 , \37050 , \36793 );
nor \U$36806 ( \37052 , \37049 , \37051 );
not \U$36807 ( \37053 , \37052 );
not \U$36808 ( \37054 , \37053 );
not \U$36809 ( \37055 , RIbe2b4c8_124);
not \U$36810 ( \37056 , RIbe2aaf0_103);
or \U$36811 ( \37057 , \37055 , \37056 );
or \U$36812 ( \37058 , RIbe2aaf0_103, RIbe2b4c8_124);
nand \U$36813 ( \37059 , \37057 , \37058 );
or \U$36814 ( \37060 , \19580 , \37059 );
or \U$36815 ( \37061 , \18830 , \36730 );
nand \U$36816 ( \37062 , \37060 , \37061 );
not \U$36817 ( \37063 , \37062 );
not \U$36818 ( \37064 , \15968 );
xnor \U$36819 ( \37065 , RIbe2a640_93, RIbe2b018_114);
not \U$36820 ( \37066 , \37065 );
and \U$36821 ( \37067 , \37064 , \37066 );
and \U$36822 ( \37068 , \36955 , \36951 );
nor \U$36823 ( \37069 , \37067 , \37068 );
not \U$36824 ( \37070 , \37069 );
or \U$36825 ( \37071 , \37063 , \37070 );
or \U$36826 ( \37072 , \37069 , \37062 );
nand \U$36827 ( \37073 , \37071 , \37072 );
not \U$36828 ( \37074 , \37073 );
xor \U$36829 ( \37075 , \36968 , \36964 );
not \U$36830 ( \37076 , \37075 );
or \U$36831 ( \37077 , \37074 , \37076 );
not \U$36832 ( \37078 , \37069 );
nand \U$36833 ( \37079 , \37078 , \37062 );
nand \U$36834 ( \37080 , \37077 , \37079 );
not \U$36835 ( \37081 , \37080 );
or \U$36836 ( \37082 , \37054 , \37081 );
or \U$36837 ( \37083 , \37080 , \37053 );
not \U$36838 ( \37084 , \36755 );
not \U$36839 ( \37085 , \36737 );
not \U$36840 ( \37086 , \37085 );
and \U$36841 ( \37087 , \37084 , \37086 );
and \U$36842 ( \37088 , \36755 , \37085 );
nor \U$36843 ( \37089 , \37087 , \37088 );
buf \U$36844 ( \37090 , \36745 );
xnor \U$36845 ( \37091 , \37089 , \37090 );
nand \U$36846 ( \37092 , \37083 , \37091 );
nand \U$36847 ( \37093 , \37082 , \37092 );
xor \U$36848 ( \37094 , \36757 , \36769 );
xor \U$36849 ( \37095 , \37094 , \36797 );
xor \U$36850 ( \37096 , \37093 , \37095 );
xor \U$36851 ( \37097 , \36909 , \36910 );
xor \U$36852 ( \37098 , \37097 , \36978 );
and \U$36853 ( \37099 , \37096 , \37098 );
and \U$36854 ( \37100 , \37093 , \37095 );
or \U$36855 ( \37101 , \37099 , \37100 );
not \U$36856 ( \37102 , \37101 );
nand \U$36857 ( \37103 , \37048 , \37102 );
nand \U$36858 ( \37104 , \37046 , \37103 );
xor \U$36859 ( \37105 , RIbe2af28_112, RIbe2b3d8_122);
not \U$36860 ( \37106 , \37105 );
not \U$36861 ( \37107 , \18649 );
or \U$36862 ( \37108 , \37106 , \37107 );
xor \U$36863 ( \37109 , RIbe2af28_112, RIbe2b450_123);
nand \U$36864 ( \37110 , \19721 , \37109 );
nand \U$36865 ( \37111 , \37108 , \37110 );
or \U$36866 ( \37112 , RIbe2ae38_110, RIbe2af28_112);
nand \U$36867 ( \37113 , \37112 , RIbe2b1f8_118);
nand \U$36868 ( \37114 , RIbe2ae38_110, RIbe2af28_112);
nand \U$36869 ( \37115 , \37113 , \37114 , RIbe2b180_117);
xor \U$36870 ( \37116 , \37111 , \37115 );
not \U$36871 ( \37117 , \37116 );
not \U$36872 ( \37118 , \37117 );
and \U$36873 ( \37119 , RIbe2b018_114, RIbe2b450_123);
not \U$36874 ( \37120 , RIbe2b018_114);
not \U$36875 ( \37121 , RIbe2b450_123);
and \U$36876 ( \37122 , \37120 , \37121 );
nor \U$36877 ( \37123 , \37119 , \37122 );
not \U$36878 ( \37124 , \37123 );
not \U$36879 ( \37125 , \17571 );
or \U$36880 ( \37126 , \37124 , \37125 );
and \U$36881 ( \37127 , RIbe2b018_114, RIbe2a730_95);
not \U$36882 ( \37128 , RIbe2b018_114);
not \U$36883 ( \37129 , RIbe2a730_95);
and \U$36884 ( \37130 , \37128 , \37129 );
nor \U$36885 ( \37131 , \37127 , \37130 );
nand \U$36886 ( \37132 , \15953 , \37131 );
nand \U$36887 ( \37133 , \37126 , \37132 );
not \U$36888 ( \37134 , \37133 );
nand \U$36889 ( \37135 , \14966 , RIbe2ae38_110);
not \U$36890 ( \37136 , \37135 );
xor \U$36891 ( \37137 , RIbe2af28_112, RIbe2aeb0_111);
not \U$36892 ( \37138 , \37137 );
not \U$36893 ( \37139 , \16913 );
or \U$36894 ( \37140 , \37138 , \37139 );
nand \U$36895 ( \37141 , \17810 , \37105 );
nand \U$36896 ( \37142 , \37140 , \37141 );
not \U$36897 ( \37143 , \37142 );
or \U$36898 ( \37144 , \37136 , \37143 );
or \U$36899 ( \37145 , \37142 , \37135 );
nand \U$36900 ( \37146 , \37144 , \37145 );
not \U$36901 ( \37147 , \37146 );
or \U$36902 ( \37148 , \37134 , \37147 );
not \U$36903 ( \37149 , \37135 );
nand \U$36904 ( \37150 , \37149 , \37142 );
nand \U$36905 ( \37151 , \37148 , \37150 );
not \U$36906 ( \37152 , \37151 );
not \U$36907 ( \37153 , \37152 );
or \U$36908 ( \37154 , \37118 , \37153 );
nand \U$36909 ( \37155 , \37151 , \37116 );
nand \U$36910 ( \37156 , \37154 , \37155 );
not \U$36911 ( \37157 , \36773 );
and \U$36912 ( \37158 , RIbe2b180_117, \24871 );
not \U$36913 ( \37159 , RIbe2b180_117);
and \U$36914 ( \37160 , \37159 , RIbe2ae38_110);
nor \U$36915 ( \37161 , \37158 , \37160 );
or \U$36916 ( \37162 , \37157 , \37161 );
xor \U$36917 ( \37163 , RIbe2aeb0_111, RIbe2b180_117);
not \U$36918 ( \37164 , \37163 );
or \U$36919 ( \37165 , \36847 , \37164 );
nand \U$36920 ( \37166 , \37162 , \37165 );
not \U$36921 ( \37167 , \37166 );
not \U$36922 ( \37168 , \37167 );
not \U$36923 ( \37169 , RIbe2aaf0_103);
not \U$36924 ( \37170 , RIbe2abe0_105);
and \U$36925 ( \37171 , \37169 , \37170 );
and \U$36926 ( \37172 , RIbe2aaf0_103, RIbe2abe0_105);
nor \U$36927 ( \37173 , \37171 , \37172 );
not \U$36928 ( \37174 , \37173 );
not \U$36929 ( \37175 , \28282 );
or \U$36930 ( \37176 , \37174 , \37175 );
xor \U$36931 ( \37177 , RIbe2aaf0_103, RIbe2ac58_106);
nand \U$36932 ( \37178 , \37177 , RIbe2ab68_104);
nand \U$36933 ( \37179 , \37176 , \37178 );
not \U$36934 ( \37180 , \37179 );
not \U$36935 ( \37181 , \37131 );
not \U$36936 ( \37182 , \22763 );
or \U$36937 ( \37183 , \37181 , \37182 );
not \U$36938 ( \37184 , RIbe2b018_114);
not \U$36939 ( \37185 , RIbe2a7a8_96);
or \U$36940 ( \37186 , \37184 , \37185 );
or \U$36941 ( \37187 , RIbe2a7a8_96, RIbe2b018_114);
nand \U$36942 ( \37188 , \37186 , \37187 );
not \U$36943 ( \37189 , \37188 );
nand \U$36944 ( \37190 , \37189 , \20583 );
nand \U$36945 ( \37191 , \37183 , \37190 );
not \U$36946 ( \37192 , \37191 );
not \U$36947 ( \37193 , \37192 );
or \U$36948 ( \37194 , \37180 , \37193 );
or \U$36949 ( \37195 , \37192 , \37179 );
nand \U$36950 ( \37196 , \37194 , \37195 );
not \U$36951 ( \37197 , \37196 );
or \U$36952 ( \37198 , \37168 , \37197 );
not \U$36953 ( \37199 , \37196 );
nand \U$36954 ( \37200 , \37199 , \37166 );
nand \U$36955 ( \37201 , \37198 , \37200 );
and \U$36956 ( \37202 , \37156 , \37201 );
not \U$36957 ( \37203 , \37156 );
not \U$36958 ( \37204 , \37201 );
and \U$36959 ( \37205 , \37203 , \37204 );
nor \U$36960 ( \37206 , \37202 , \37205 );
not \U$36961 ( \37207 , \37206 );
xor \U$36962 ( \37208 , RIbe2a7a8_96, RIbe2aaf0_103);
not \U$36963 ( \37209 , \37208 );
not \U$36964 ( \37210 , \35178 );
or \U$36965 ( \37211 , \37209 , \37210 );
nand \U$36966 ( \37212 , \37173 , RIbe2ab68_104);
nand \U$36967 ( \37213 , \37211 , \37212 );
not \U$36968 ( \37214 , \37213 );
or \U$36969 ( \37215 , \14417 , \24871 );
nand \U$36970 ( \37216 , RIbe2afa0_113, RIbe2b018_114);
and \U$36971 ( \37217 , \37216 , RIbe2af28_112);
nand \U$36972 ( \37218 , \37215 , \37217 );
not \U$36973 ( \37219 , \37218 );
and \U$36974 ( \37220 , RIbe2aaf0_103, RIbe2a730_95);
not \U$36975 ( \37221 , RIbe2aaf0_103);
and \U$36976 ( \37222 , \37221 , \37129 );
nor \U$36977 ( \37223 , \37220 , \37222 );
not \U$36978 ( \37224 , \37223 );
not \U$36979 ( \37225 , \23169 );
or \U$36980 ( \37226 , \37224 , \37225 );
nand \U$36981 ( \37227 , \37208 , RIbe2ab68_104);
nand \U$36982 ( \37228 , \37226 , \37227 );
nand \U$36983 ( \37229 , \37219 , \37228 );
or \U$36984 ( \37230 , \37214 , \37229 );
not \U$36985 ( \37231 , \37229 );
not \U$36986 ( \37232 , \37214 );
or \U$36987 ( \37233 , \37231 , \37232 );
and \U$36988 ( \37234 , \37146 , \37133 );
not \U$36989 ( \37235 , \37146 );
not \U$36990 ( \37236 , \37133 );
and \U$36991 ( \37237 , \37235 , \37236 );
nor \U$36992 ( \37238 , \37234 , \37237 );
nand \U$36993 ( \37239 , \37233 , \37238 );
nand \U$36994 ( \37240 , \37230 , \37239 );
not \U$36995 ( \37241 , \37240 );
nand \U$36996 ( \37242 , \37207 , \37241 );
not \U$36997 ( \37243 , \37242 );
not \U$36998 ( \37244 , \37240 );
not \U$36999 ( \37245 , \37206 );
or \U$37000 ( \37246 , \37244 , \37245 );
not \U$37001 ( \37247 , \25897 );
not \U$37002 ( \37248 , RIbe2b018_114);
not \U$37003 ( \37249 , RIbe2aeb0_111);
or \U$37004 ( \37250 , \37248 , \37249 );
or \U$37005 ( \37251 , RIbe2aeb0_111, RIbe2b018_114);
nand \U$37006 ( \37252 , \37250 , \37251 );
or \U$37007 ( \37253 , \37247 , \37252 );
xnor \U$37008 ( \37254 , RIbe2b018_114, RIbe2b3d8_122);
or \U$37009 ( \37255 , \25891 , \37254 );
nand \U$37010 ( \37256 , \37253 , \37255 );
and \U$37011 ( \37257 , RIbe2aaf0_103, RIbe2b450_123);
not \U$37012 ( \37258 , RIbe2aaf0_103);
and \U$37013 ( \37259 , \37258 , \37121 );
nor \U$37014 ( \37260 , \37257 , \37259 );
not \U$37015 ( \37261 , \37260 );
or \U$37016 ( \37262 , \34550 , \37261 );
not \U$37017 ( \37263 , \37223 );
or \U$37018 ( \37264 , \37263 , \18830 );
nand \U$37019 ( \37265 , \37262 , \37264 );
not \U$37020 ( \37266 , \37265 );
nand \U$37021 ( \37267 , \15348 , RIbe2ae38_110);
nand \U$37022 ( \37268 , \37266 , \37267 );
nand \U$37023 ( \37269 , \37256 , \37268 );
not \U$37024 ( \37270 , \37267 );
nand \U$37025 ( \37271 , \37270 , \37265 );
nand \U$37026 ( \37272 , \37269 , \37271 );
not \U$37027 ( \37273 , \37272 );
not \U$37028 ( \37274 , \37218 );
not \U$37029 ( \37275 , \37228 );
not \U$37030 ( \37276 , \37275 );
or \U$37031 ( \37277 , \37274 , \37276 );
nand \U$37032 ( \37278 , \37277 , \37229 );
nor \U$37033 ( \37279 , \34558 , \37254 );
and \U$37034 ( \37280 , \19371 , \37123 );
nor \U$37035 ( \37281 , \37279 , \37280 );
xor \U$37036 ( \37282 , \37278 , \37281 );
or \U$37037 ( \37283 , \24871 , RIbe2af28_112);
not \U$37038 ( \37284 , RIbe2af28_112);
or \U$37039 ( \37285 , \37284 , RIbe2ae38_110);
nand \U$37040 ( \37286 , \37283 , \37285 );
and \U$37041 ( \37287 , \35366 , \37286 );
and \U$37042 ( \37288 , \19721 , \37137 );
nor \U$37043 ( \37289 , \37287 , \37288 );
xor \U$37044 ( \37290 , \37282 , \37289 );
not \U$37045 ( \37291 , \37290 );
not \U$37046 ( \37292 , \37291 );
or \U$37047 ( \37293 , \37273 , \37292 );
not \U$37048 ( \37294 , \22763 );
and \U$37049 ( \37295 , \15958 , RIbe2ae38_110);
and \U$37050 ( \37296 , \24871 , RIbe2b018_114);
nor \U$37051 ( \37297 , \37295 , \37296 );
or \U$37052 ( \37298 , \37294 , \37297 );
not \U$37053 ( \37299 , \20583 );
or \U$37054 ( \37300 , \37299 , \37252 );
nand \U$37055 ( \37301 , \37298 , \37300 );
not \U$37056 ( \37302 , \37301 );
not \U$37057 ( \37303 , RIbe2aaf0_103);
nand \U$37058 ( \37304 , \37303 , \24871 );
and \U$37059 ( \37305 , \37304 , RIbe2b630_127);
nand \U$37060 ( \37306 , RIbe2aaf0_103, RIbe2ae38_110);
nand \U$37061 ( \37307 , \37306 , RIbe2b018_114);
nor \U$37062 ( \37308 , \37305 , \37307 );
not \U$37063 ( \37309 , RIbe2ab68_104);
not \U$37064 ( \37310 , \37260 );
or \U$37065 ( \37311 , \37309 , \37310 );
xnor \U$37066 ( \37312 , RIbe2b3d8_122, RIbe2aaf0_103);
or \U$37067 ( \37313 , \19580 , \37312 );
nand \U$37068 ( \37314 , \37311 , \37313 );
xor \U$37069 ( \37315 , \37308 , \37314 );
not \U$37070 ( \37316 , \37315 );
or \U$37071 ( \37317 , \37302 , \37316 );
or \U$37072 ( \37318 , \37315 , \37301 );
nand \U$37073 ( \37319 , \25891 , RIbe2ae38_110);
or \U$37074 ( \37320 , \37312 , \18830 );
not \U$37075 ( \37321 , \35178 );
nand \U$37076 ( \37322 , \37320 , \37321 );
not \U$37077 ( \37323 , RIbe2ae38_110);
not \U$37078 ( \37324 , RIbe2ab68_104);
or \U$37079 ( \37325 , \37323 , \37324 );
nand \U$37080 ( \37326 , \37325 , RIbe2aeb0_111);
and \U$37081 ( \37327 , \37319 , \37322 , \37304 , \37326 );
nand \U$37082 ( \37328 , \37318 , \37327 );
nand \U$37083 ( \37329 , \37317 , \37328 );
and \U$37084 ( \37330 , \37308 , \37314 );
nand \U$37085 ( \37331 , \37329 , \37330 );
nand \U$37086 ( \37332 , \37268 , \37271 );
and \U$37087 ( \37333 , \37332 , \37256 );
not \U$37088 ( \37334 , \37332 );
not \U$37089 ( \37335 , \37256 );
and \U$37090 ( \37336 , \37334 , \37335 );
nor \U$37091 ( \37337 , \37333 , \37336 );
and \U$37092 ( \37338 , \37331 , \37337 );
nor \U$37093 ( \37339 , \37329 , \37330 );
nor \U$37094 ( \37340 , \37338 , \37339 );
not \U$37095 ( \37341 , \37272 );
nand \U$37096 ( \37342 , \37341 , \37290 );
nand \U$37097 ( \37343 , \37340 , \37342 );
nand \U$37098 ( \37344 , \37293 , \37343 );
not \U$37099 ( \37345 , \37238 );
not \U$37100 ( \37346 , \37229 );
not \U$37101 ( \37347 , \37213 );
or \U$37102 ( \37348 , \37346 , \37347 );
or \U$37103 ( \37349 , \37213 , \37229 );
nand \U$37104 ( \37350 , \37348 , \37349 );
nand \U$37105 ( \37351 , \37345 , \37350 );
not \U$37106 ( \37352 , \37350 );
nand \U$37107 ( \37353 , \37352 , \37238 );
xor \U$37108 ( \37354 , \37278 , \37281 );
and \U$37109 ( \37355 , \37354 , \37289 );
and \U$37110 ( \37356 , \37278 , \37281 );
or \U$37111 ( \37357 , \37355 , \37356 );
nand \U$37112 ( \37358 , \37351 , \37353 , \37357 );
and \U$37113 ( \37359 , \37344 , \37358 );
and \U$37114 ( \37360 , \37353 , \37351 );
nor \U$37115 ( \37361 , \37360 , \37357 );
nor \U$37116 ( \37362 , \37359 , \37361 );
nand \U$37117 ( \37363 , \37246 , \37362 );
not \U$37118 ( \37364 , \37363 );
or \U$37119 ( \37365 , \37243 , \37364 );
not \U$37120 ( \37366 , \34558 );
not \U$37121 ( \37367 , \37188 );
and \U$37122 ( \37368 , \37366 , \37367 );
not \U$37123 ( \37369 , \36199 );
xor \U$37124 ( \37370 , RIbe2abe0_105, RIbe2b018_114);
and \U$37125 ( \37371 , \37369 , \37370 );
nor \U$37126 ( \37372 , \37368 , \37371 );
not \U$37127 ( \37373 , \37163 );
not \U$37128 ( \37374 , \36773 );
or \U$37129 ( \37375 , \37373 , \37374 );
xnor \U$37130 ( \37376 , RIbe2b3d8_122, RIbe2b180_117);
not \U$37131 ( \37377 , \37376 );
nand \U$37132 ( \37378 , \37377 , \21759 );
nand \U$37133 ( \37379 , \37375 , \37378 );
xor \U$37134 ( \37380 , \37372 , \37379 );
not \U$37135 ( \37381 , \37115 );
and \U$37136 ( \37382 , \37111 , \37381 );
xor \U$37137 ( \37383 , \37380 , \37382 );
not \U$37138 ( \37384 , \37383 );
and \U$37139 ( \37385 , \30236 , \37177 );
xor \U$37140 ( \37386 , RIbe2aaf0_103, RIbe2a640_93);
and \U$37141 ( \37387 , \37386 , RIbe2ab68_104);
nor \U$37142 ( \37388 , \37385 , \37387 );
not \U$37143 ( \37389 , \37388 );
nand \U$37144 ( \37390 , \23015 , RIbe2ae38_110);
not \U$37145 ( \37391 , \37390 );
not \U$37146 ( \37392 , \37391 );
and \U$37147 ( \37393 , \37389 , \37392 );
and \U$37148 ( \37394 , \37388 , \37391 );
nor \U$37149 ( \37395 , \37393 , \37394 );
not \U$37150 ( \37396 , \37395 );
xor \U$37151 ( \37397 , RIbe2a730_95, RIbe2af28_112);
not \U$37152 ( \37398 , \37397 );
not \U$37153 ( \37399 , \15348 );
or \U$37154 ( \37400 , \37398 , \37399 );
nand \U$37155 ( \37401 , \18649 , \37109 );
nand \U$37156 ( \37402 , \37400 , \37401 );
not \U$37157 ( \37403 , \37402 );
and \U$37158 ( \37404 , \37396 , \37403 );
and \U$37159 ( \37405 , \37395 , \37402 );
nor \U$37160 ( \37406 , \37404 , \37405 );
not \U$37161 ( \37407 , \37406 );
not \U$37162 ( \37408 , \37407 );
not \U$37163 ( \37409 , \37166 );
not \U$37164 ( \37410 , \37196 );
or \U$37165 ( \37411 , \37409 , \37410 );
nand \U$37166 ( \37412 , \37191 , \37179 );
nand \U$37167 ( \37413 , \37411 , \37412 );
not \U$37168 ( \37414 , \37413 );
not \U$37169 ( \37415 , \37414 );
or \U$37170 ( \37416 , \37408 , \37415 );
nand \U$37171 ( \37417 , \37406 , \37413 );
nand \U$37172 ( \37418 , \37416 , \37417 );
not \U$37173 ( \37419 , \37418 );
or \U$37174 ( \37420 , \37384 , \37419 );
or \U$37175 ( \37421 , \37418 , \37383 );
nand \U$37176 ( \37422 , \37420 , \37421 );
not \U$37177 ( \37423 , \37422 );
nand \U$37178 ( \37424 , \37365 , \37423 );
nand \U$37179 ( \37425 , \37363 , \37242 , \37422 );
and \U$37180 ( \37426 , \37156 , \37201 );
and \U$37181 ( \37427 , \37151 , \37117 );
nor \U$37182 ( \37428 , \37426 , \37427 );
nand \U$37183 ( \37429 , \37425 , \37428 );
not \U$37184 ( \37430 , \37386 );
not \U$37185 ( \37431 , \35178 );
or \U$37186 ( \37432 , \37430 , \37431 );
xor \U$37187 ( \37433 , RIbe2aaf0_103, RIbe2a6b8_94);
nand \U$37188 ( \37434 , \37433 , RIbe2ab68_104);
nand \U$37189 ( \37435 , \37432 , \37434 );
not \U$37190 ( \37436 , \37370 );
not \U$37191 ( \37437 , \25897 );
or \U$37192 ( \37438 , \37436 , \37437 );
xnor \U$37193 ( \37439 , RIbe2b018_114, RIbe2ac58_106);
not \U$37194 ( \37440 , \37439 );
nand \U$37195 ( \37441 , \37440 , \19371 );
nand \U$37196 ( \37442 , \37438 , \37441 );
xor \U$37197 ( \37443 , \37435 , \37442 );
not \U$37198 ( \37444 , \37397 );
not \U$37199 ( \37445 , \15345 );
or \U$37200 ( \37446 , \37444 , \37445 );
and \U$37201 ( \37447 , \37284 , RIbe2a7a8_96);
and \U$37202 ( \37448 , \15634 , RIbe2af28_112);
nor \U$37203 ( \37449 , \37447 , \37448 );
not \U$37204 ( \37450 , \37449 );
nand \U$37205 ( \37451 , \37450 , \17811 );
nand \U$37206 ( \37452 , \37446 , \37451 );
xnor \U$37207 ( \37453 , \37443 , \37452 );
not \U$37208 ( \37454 , \37372 );
and \U$37209 ( \37455 , \37454 , \37379 );
not \U$37210 ( \37456 , \37379 );
nand \U$37211 ( \37457 , \37456 , \37372 );
and \U$37212 ( \37458 , \37382 , \37457 );
nor \U$37213 ( \37459 , \37455 , \37458 );
xor \U$37214 ( \37460 , \37453 , \37459 );
not \U$37215 ( \37461 , \37460 );
and \U$37216 ( \37462 , RIbe2b108_116, \24871 );
not \U$37217 ( \37463 , RIbe2b108_116);
and \U$37218 ( \37464 , \37463 , RIbe2ae38_110);
nor \U$37219 ( \37465 , \37462 , \37464 );
or \U$37220 ( \37466 , \13544 , \37465 );
not \U$37221 ( \37467 , RIbe2aeb0_111);
not \U$37222 ( \37468 , RIbe2b108_116);
and \U$37223 ( \37469 , \37467 , \37468 );
and \U$37224 ( \37470 , RIbe2aeb0_111, RIbe2b108_116);
nor \U$37225 ( \37471 , \37469 , \37470 );
not \U$37226 ( \37472 , \37471 );
or \U$37227 ( \37473 , \16876 , \37472 );
nand \U$37228 ( \37474 , \37466 , \37473 );
nand \U$37229 ( \37475 , RIbe2ae38_110, RIbe2b180_117);
or \U$37230 ( \37476 , RIbe2ae38_110, RIbe2b180_117);
nand \U$37231 ( \37477 , \37476 , RIbe2b270_119);
nand \U$37232 ( \37478 , \37475 , RIbe2b108_116, \37477 );
not \U$37233 ( \37479 , \37478 );
or \U$37234 ( \37480 , \14853 , \37376 );
xor \U$37235 ( \37481 , RIbe2b450_123, RIbe2b180_117);
not \U$37236 ( \37482 , \37481 );
or \U$37237 ( \37483 , \25254 , \37482 );
nand \U$37238 ( \37484 , \37480 , \37483 );
not \U$37239 ( \37485 , \37484 );
or \U$37240 ( \37486 , \37479 , \37485 );
or \U$37241 ( \37487 , \37484 , \37478 );
nand \U$37242 ( \37488 , \37486 , \37487 );
xor \U$37243 ( \37489 , \37474 , \37488 );
not \U$37244 ( \37490 , \37402 );
or \U$37245 ( \37491 , \37395 , \37490 );
not \U$37246 ( \37492 , \37388 );
nand \U$37247 ( \37493 , \37492 , \37391 );
nand \U$37248 ( \37494 , \37491 , \37493 );
xor \U$37249 ( \37495 , \37489 , \37494 );
not \U$37250 ( \37496 , \37495 );
or \U$37251 ( \37497 , \37461 , \37496 );
or \U$37252 ( \37498 , \37495 , \37460 );
nand \U$37253 ( \37499 , \37497 , \37498 );
not \U$37254 ( \37500 , \37383 );
and \U$37255 ( \37501 , \37418 , \37500 );
and \U$37256 ( \37502 , \37407 , \37413 );
nor \U$37257 ( \37503 , \37501 , \37502 );
nand \U$37258 ( \37504 , \37499 , \37503 );
nand \U$37259 ( \37505 , \37424 , \37429 , \37504 );
not \U$37260 ( \37506 , \37478 );
nand \U$37261 ( \37507 , \37506 , \37484 );
not \U$37262 ( \37508 , \37435 );
not \U$37263 ( \37509 , \37442 );
or \U$37264 ( \37510 , \37508 , \37509 );
or \U$37265 ( \37511 , \37442 , \37435 );
nand \U$37266 ( \37512 , \37511 , \37452 );
nand \U$37267 ( \37513 , \37510 , \37512 );
xor \U$37268 ( \37514 , \37507 , \37513 );
and \U$37269 ( \37515 , \13543 , \37471 );
and \U$37270 ( \37516 , \23015 , \36959 );
nor \U$37271 ( \37517 , \37515 , \37516 );
not \U$37272 ( \37518 , \37517 );
not \U$37273 ( \37519 , \37481 );
not \U$37274 ( \37520 , \15353 );
or \U$37275 ( \37521 , \37519 , \37520 );
nand \U$37276 ( \37522 , \14966 , \36930 );
nand \U$37277 ( \37523 , \37521 , \37522 );
nand \U$37278 ( \37524 , \14649 , RIbe2ae38_110);
not \U$37279 ( \37525 , \37524 );
and \U$37280 ( \37526 , \37523 , \37525 );
not \U$37281 ( \37527 , \37523 );
and \U$37282 ( \37528 , \37527 , \37524 );
nor \U$37283 ( \37529 , \37526 , \37528 );
not \U$37284 ( \37530 , \37529 );
or \U$37285 ( \37531 , \37518 , \37530 );
or \U$37286 ( \37532 , \37529 , \37517 );
nand \U$37287 ( \37533 , \37531 , \37532 );
xnor \U$37288 ( \37534 , \37514 , \37533 );
xor \U$37289 ( \37535 , \37474 , \37488 );
and \U$37290 ( \37536 , \37535 , \37494 );
and \U$37291 ( \37537 , \37474 , \37488 );
or \U$37292 ( \37538 , \37536 , \37537 );
not \U$37293 ( \37539 , \37433 );
or \U$37294 ( \37540 , \19580 , \37539 );
or \U$37295 ( \37541 , \18830 , \37059 );
nand \U$37296 ( \37542 , \37540 , \37541 );
or \U$37297 ( \37543 , \37294 , \37439 );
or \U$37298 ( \37544 , \15954 , \37065 );
nand \U$37299 ( \37545 , \37543 , \37544 );
xor \U$37300 ( \37546 , \37542 , \37545 );
or \U$37301 ( \37547 , \14424 , \37449 );
not \U$37302 ( \37548 , \15348 );
or \U$37303 ( \37549 , \37548 , \36913 );
nand \U$37304 ( \37550 , \37547 , \37549 );
xor \U$37305 ( \37551 , \37546 , \37550 );
nor \U$37306 ( \37552 , \37538 , \37551 );
not \U$37307 ( \37553 , \37552 );
nand \U$37308 ( \37554 , \37538 , \37551 );
nand \U$37309 ( \37555 , \37553 , \37554 );
not \U$37310 ( \37556 , \37555 );
and \U$37311 ( \37557 , \37534 , \37556 );
not \U$37312 ( \37558 , \37534 );
and \U$37313 ( \37559 , \37558 , \37555 );
nor \U$37314 ( \37560 , \37557 , \37559 );
not \U$37315 ( \37561 , \37495 );
and \U$37316 ( \37562 , \37453 , \37459 );
or \U$37317 ( \37563 , \37561 , \37562 );
or \U$37318 ( \37564 , \37459 , \37453 );
nand \U$37319 ( \37565 , \37563 , \37564 );
nand \U$37320 ( \37566 , \37560 , \37565 );
or \U$37321 ( \37567 , \37499 , \37503 );
nand \U$37322 ( \37568 , \37505 , \37566 , \37567 );
not \U$37323 ( \37569 , \37552 );
not \U$37324 ( \37570 , \37569 );
not \U$37325 ( \37571 , \37534 );
or \U$37326 ( \37572 , \37570 , \37571 );
nand \U$37327 ( \37573 , \37572 , \37554 );
not \U$37328 ( \37574 , \37573 );
not \U$37329 ( \37575 , \37073 );
and \U$37330 ( \37576 , \37075 , \37575 );
not \U$37331 ( \37577 , \37075 );
and \U$37332 ( \37578 , \37577 , \37073 );
nor \U$37333 ( \37579 , \37576 , \37578 );
not \U$37334 ( \37580 , \37513 );
not \U$37335 ( \37581 , \37507 );
not \U$37336 ( \37582 , \37533 );
or \U$37337 ( \37583 , \37581 , \37582 );
or \U$37338 ( \37584 , \37533 , \37507 );
nand \U$37339 ( \37585 , \37583 , \37584 );
not \U$37340 ( \37586 , \37585 );
or \U$37341 ( \37587 , \37580 , \37586 );
not \U$37342 ( \37588 , \37507 );
nand \U$37343 ( \37589 , \37588 , \37533 );
nand \U$37344 ( \37590 , \37587 , \37589 );
xor \U$37345 ( \37591 , \37579 , \37590 );
xor \U$37346 ( \37592 , \37542 , \37545 );
and \U$37347 ( \37593 , \37592 , \37550 );
and \U$37348 ( \37594 , \37542 , \37545 );
or \U$37349 ( \37595 , \37593 , \37594 );
not \U$37350 ( \37596 , \37595 );
not \U$37351 ( \37597 , \37517 );
not \U$37352 ( \37598 , \37597 );
not \U$37353 ( \37599 , \37529 );
or \U$37354 ( \37600 , \37598 , \37599 );
nand \U$37355 ( \37601 , \37523 , \37525 );
nand \U$37356 ( \37602 , \37600 , \37601 );
not \U$37357 ( \37603 , \37602 );
not \U$37358 ( \37604 , \37603 );
or \U$37359 ( \37605 , \37596 , \37604 );
or \U$37360 ( \37606 , \37603 , \37595 );
nand \U$37361 ( \37607 , \37605 , \37606 );
xor \U$37362 ( \37608 , \36939 , \36918 );
xor \U$37363 ( \37609 , \37607 , \37608 );
xor \U$37364 ( \37610 , \37591 , \37609 );
nand \U$37365 ( \37611 , \37574 , \37610 );
not \U$37366 ( \37612 , \37560 );
not \U$37367 ( \37613 , \37565 );
nand \U$37368 ( \37614 , \37612 , \37613 );
nand \U$37369 ( \37615 , \37568 , \37611 , \37614 );
not \U$37370 ( \37616 , \37610 );
nand \U$37371 ( \37617 , \37616 , \37573 );
nand \U$37372 ( \37618 , \37615 , \37617 );
xor \U$37373 ( \37619 , \36973 , \36944 );
not \U$37374 ( \37620 , \37091 );
not \U$37375 ( \37621 , \37620 );
not \U$37376 ( \37622 , \37053 );
or \U$37377 ( \37623 , \37621 , \37622 );
nand \U$37378 ( \37624 , \37052 , \37091 );
nand \U$37379 ( \37625 , \37623 , \37624 );
and \U$37380 ( \37626 , \37625 , \37080 );
not \U$37381 ( \37627 , \37625 );
not \U$37382 ( \37628 , \37080 );
and \U$37383 ( \37629 , \37627 , \37628 );
nor \U$37384 ( \37630 , \37626 , \37629 );
xor \U$37385 ( \37631 , \37619 , \37630 );
not \U$37386 ( \37632 , \37608 );
not \U$37387 ( \37633 , \37607 );
or \U$37388 ( \37634 , \37632 , \37633 );
nand \U$37389 ( \37635 , \37602 , \37595 );
nand \U$37390 ( \37636 , \37634 , \37635 );
and \U$37391 ( \37637 , \37631 , \37636 );
and \U$37392 ( \37638 , \37619 , \37630 );
or \U$37393 ( \37639 , \37637 , \37638 );
xor \U$37394 ( \37640 , \37093 , \37095 );
xor \U$37395 ( \37641 , \37640 , \37098 );
nor \U$37396 ( \37642 , \37639 , \37641 );
xor \U$37397 ( \37643 , \37619 , \37630 );
xor \U$37398 ( \37644 , \37643 , \37636 );
not \U$37399 ( \37645 , \37579 );
not \U$37400 ( \37646 , \37645 );
not \U$37401 ( \37647 , \37609 );
or \U$37402 ( \37648 , \37646 , \37647 );
not \U$37403 ( \37649 , \37609 );
nand \U$37404 ( \37650 , \37649 , \37579 );
nand \U$37405 ( \37651 , \37650 , \37590 );
nand \U$37406 ( \37652 , \37648 , \37651 );
nor \U$37407 ( \37653 , \37644 , \37652 );
nor \U$37408 ( \37654 , \37642 , \37653 );
nand \U$37409 ( \37655 , \37618 , \37654 );
or \U$37410 ( \37656 , \37104 , \37655 );
and \U$37411 ( \37657 , \37652 , \37644 );
not \U$37412 ( \37658 , \37642 );
and \U$37413 ( \37659 , \37657 , \37658 );
and \U$37414 ( \37660 , \37641 , \37639 );
nor \U$37415 ( \37661 , \37659 , \37660 );
or \U$37416 ( \37662 , \37104 , \37661 );
not \U$37417 ( \37663 , \37046 );
not \U$37418 ( \37664 , \37048 );
nand \U$37419 ( \37665 , \37664 , \37101 );
or \U$37420 ( \37666 , \37663 , \37665 );
not \U$37421 ( \37667 , \37045 );
nand \U$37422 ( \37668 , \37667 , \36984 );
nand \U$37423 ( \37669 , \37666 , \37668 );
not \U$37424 ( \37670 , \37669 );
nand \U$37425 ( \37671 , \37656 , \37662 , \37670 );
not \U$37426 ( \37672 , \36601 );
not \U$37427 ( \37673 , \36720 );
or \U$37428 ( \37674 , \37672 , \37673 );
or \U$37429 ( \37675 , \36720 , \36601 );
nand \U$37430 ( \37676 , \37674 , \37675 );
not \U$37431 ( \37677 , \37032 );
not \U$37432 ( \37678 , \37013 );
or \U$37433 ( \37679 , \37677 , \37678 );
nand \U$37434 ( \37680 , \37679 , \37034 );
not \U$37435 ( \37681 , \37680 );
not \U$37436 ( \37682 , \36469 );
not \U$37437 ( \37683 , \36460 );
or \U$37438 ( \37684 , \37682 , \37683 );
nand \U$37439 ( \37685 , \36461 , \36468 );
nand \U$37440 ( \37686 , \37684 , \37685 );
not \U$37441 ( \37687 , \37686 );
not \U$37442 ( \37688 , \36476 );
not \U$37443 ( \37689 , \37688 );
and \U$37444 ( \37690 , \37687 , \37689 );
and \U$37445 ( \37691 , \37686 , \37688 );
nor \U$37446 ( \37692 , \37690 , \37691 );
and \U$37447 ( \37693 , \37681 , \37692 );
not \U$37448 ( \37694 , \37681 );
not \U$37449 ( \37695 , \37692 );
and \U$37450 ( \37696 , \37694 , \37695 );
nor \U$37451 ( \37697 , \37693 , \37696 );
not \U$37452 ( \37698 , \37697 );
xnor \U$37453 ( \37699 , \36611 , \36709 );
or \U$37454 ( \37700 , \37698 , \37699 );
nand \U$37455 ( \37701 , \37680 , \37695 );
nand \U$37456 ( \37702 , \37700 , \37701 );
nor \U$37457 ( \37703 , \37676 , \37702 );
not \U$37458 ( \37704 , \37699 );
not \U$37459 ( \37705 , \37697 );
or \U$37460 ( \37706 , \37704 , \37705 );
or \U$37461 ( \37707 , \37697 , \37699 );
nand \U$37462 ( \37708 , \37706 , \37707 );
not \U$37463 ( \37709 , \36996 );
not \U$37464 ( \37710 , \37709 );
not \U$37465 ( \37711 , \37003 );
or \U$37466 ( \37712 , \37710 , \37711 );
not \U$37467 ( \37713 , \37003 );
nand \U$37468 ( \37714 , \37713 , \36996 );
nand \U$37469 ( \37715 , \37041 , \37714 );
nand \U$37470 ( \37716 , \37712 , \37715 );
nor \U$37471 ( \37717 , \37708 , \37716 );
nor \U$37472 ( \37718 , \37703 , \37717 );
nand \U$37473 ( \37719 , \36729 , \37671 , \37718 );
nand \U$37474 ( \37720 , \37708 , \37716 );
or \U$37475 ( \37721 , \37703 , \37720 );
nand \U$37476 ( \37722 , \37676 , \37702 );
nand \U$37477 ( \37723 , \37721 , \37722 );
nand \U$37478 ( \37724 , \36729 , \37723 );
nor \U$37479 ( \37725 , \36595 , \36726 );
and \U$37480 ( \37726 , \36590 , \37725 );
nor \U$37481 ( \37727 , \36587 , \36589 );
nor \U$37482 ( \37728 , \37726 , \37727 );
nand \U$37483 ( \37729 , \37719 , \37724 , \37728 );
not \U$37484 ( \37730 , \37729 );
or \U$37485 ( \37731 , \36443 , \37730 );
nand \U$37486 ( \37732 , \36440 , \36434 );
or \U$37487 ( \37733 , \36308 , \37732 );
nand \U$37488 ( \37734 , \36087 , \36307 );
nand \U$37489 ( \37735 , \37733 , \37734 );
not \U$37490 ( \37736 , \37735 );
not \U$37491 ( \37737 , \36085 );
or \U$37492 ( \37738 , \37736 , \37737 );
not \U$37493 ( \37739 , \35910 );
and \U$37494 ( \37740 , \35915 , \36083 );
and \U$37495 ( \37741 , \37739 , \37740 );
and \U$37496 ( \37742 , \35900 , \35909 );
nor \U$37497 ( \37743 , \37741 , \37742 );
nand \U$37498 ( \37744 , \37738 , \37743 );
not \U$37499 ( \37745 , \37744 );
nand \U$37500 ( \37746 , \37731 , \37745 );
nand \U$37501 ( \37747 , \35839 , \37746 );
not \U$37502 ( \37748 , \35671 );
nand \U$37503 ( \37749 , \35423 , \37748 );
or \U$37504 ( \37750 , \37749 , \35679 );
nand \U$37505 ( \37751 , \35674 , \35678 );
nand \U$37506 ( \37752 , \37750 , \37751 );
nor \U$37507 ( \37753 , \35138 , \35334 );
or \U$37508 ( \37754 , \37752 , \37753 );
nand \U$37509 ( \37755 , \37754 , \35337 );
nand \U$37510 ( \37756 , \35052 , \35127 );
nand \U$37511 ( \37757 , \37755 , \37756 );
not \U$37512 ( \37758 , \35838 );
nand \U$37513 ( \37759 , \37757 , \37758 );
not \U$37514 ( \37760 , \35830 );
nand \U$37515 ( \37761 , \35745 , \35689 );
not \U$37516 ( \37762 , \37761 );
nand \U$37517 ( \37763 , \37762 , \35804 );
not \U$37518 ( \37764 , \35796 );
nand \U$37519 ( \37765 , \37764 , \35802 );
nand \U$37520 ( \37766 , \37763 , \37765 );
not \U$37521 ( \37767 , \37766 );
or \U$37522 ( \37768 , \37760 , \37767 );
not \U$37523 ( \37769 , \35825 );
not \U$37524 ( \37770 , \35829 );
nand \U$37525 ( \37771 , \37769 , \37770 );
nand \U$37526 ( \37772 , \37768 , \37771 );
buf \U$37527 ( \37773 , \35837 );
nand \U$37528 ( \37774 , \37772 , \37773 );
or \U$37529 ( \37775 , \35832 , \35836 );
nand \U$37530 ( \37776 , \37747 , \37759 , \37774 , \37775 );
nand \U$37531 ( \37777 , \34307 , \34308 , \34294 , \37776 );
not \U$37532 ( \37778 , \34294 );
not \U$37533 ( \37779 , \34263 );
nor \U$37534 ( \37780 , \34295 , \34300 );
not \U$37535 ( \37781 , \37780 );
or \U$37536 ( \37782 , \37779 , \37781 );
or \U$37537 ( \37783 , \34262 , \34204 );
nand \U$37538 ( \37784 , \37782 , \37783 );
not \U$37539 ( \37785 , \37784 );
or \U$37540 ( \37786 , \37778 , \37785 );
not \U$37541 ( \37787 , \34293 );
and \U$37542 ( \37788 , \34285 , \34278 );
and \U$37543 ( \37789 , \37787 , \37788 );
and \U$37544 ( \37790 , \34290 , \34292 );
nor \U$37545 ( \37791 , \37789 , \37790 );
nand \U$37546 ( \37792 , \37786 , \37791 );
not \U$37547 ( \37793 , \37792 );
nand \U$37548 ( \37794 , \34303 , \37777 , \37793 );
not \U$37549 ( \37795 , \29271 );
not \U$37550 ( \37796 , \25797 );
not \U$37551 ( \37797 , \25389 );
or \U$37552 ( \37798 , \25354 , \25385 );
and \U$37553 ( \37799 , \37796 , \37797 , \37798 , \28103 );
not \U$37554 ( \37800 , \28155 );
and \U$37555 ( \37801 , \37799 , \37800 , \28165 );
nand \U$37556 ( \37802 , \37794 , \37795 , \37801 );
nand \U$37557 ( \37803 , \29306 , \37802 );
not \U$37558 ( \37804 , \37803 );
or \U$37559 ( \37805 , \22680 , \37804 );
nor \U$37560 ( \37806 , \22677 , \22643 );
not \U$37561 ( \37807 , \37806 );
not \U$37562 ( \37808 , \21681 );
and \U$37563 ( \37809 , \21687 , \22158 );
not \U$37564 ( \37810 , \37809 );
or \U$37565 ( \37811 , \37808 , \37810 );
not \U$37566 ( \37812 , \21680 );
nand \U$37567 ( \37813 , \37812 , \21177 );
nand \U$37568 ( \37814 , \37811 , \37813 );
not \U$37569 ( \37815 , \37814 );
not \U$37570 ( \37816 , \22514 );
or \U$37571 ( \37817 , \37815 , \37816 );
not \U$37572 ( \37818 , \22513 );
nor \U$37573 ( \37819 , \22381 , \22368 );
not \U$37574 ( \37820 , \37819 );
or \U$37575 ( \37821 , \37818 , \37820 );
not \U$37576 ( \37822 , \22512 );
nand \U$37577 ( \37823 , \37822 , \22392 , \22383 );
nand \U$37578 ( \37824 , \37821 , \37823 );
not \U$37579 ( \37825 , \37824 );
nand \U$37580 ( \37826 , \37817 , \37825 );
not \U$37581 ( \37827 , \37826 );
or \U$37582 ( \37828 , \37807 , \37827 );
nor \U$37583 ( \37829 , \22664 , \22668 );
not \U$37584 ( \37830 , \37829 );
not \U$37585 ( \37831 , \22676 );
or \U$37586 ( \37832 , \37830 , \37831 );
not \U$37587 ( \37833 , \22671 );
not \U$37588 ( \37834 , \22675 );
nand \U$37589 ( \37835 , \37833 , \37834 );
nand \U$37590 ( \37836 , \37832 , \37835 );
nor \U$37591 ( \37837 , \22585 , \22631 );
or \U$37592 ( \37838 , \37836 , \37837 );
nand \U$37593 ( \37839 , \37838 , \22644 );
or \U$37594 ( \37840 , \22637 , \22641 );
nand \U$37595 ( \37841 , \37839 , \37840 );
not \U$37596 ( \37842 , \37841 );
nand \U$37597 ( \37843 , \37828 , \37842 );
not \U$37598 ( \37844 , \37843 );
nand \U$37599 ( \37845 , \37805 , \37844 );
nand \U$37600 ( \37846 , \18576 , \37845 , \7202 );
nand \U$37601 ( \37847 , \7192 , \18568 , \37846 );
not \U$37602 ( \37848 , \37847 );
or \U$37603 ( \37849 , \855 , \37848 );
not \U$37604 ( \37850 , \837 );
not \U$37605 ( \37851 , \638 );
nand \U$37606 ( \37852 , \37851 , \585 );
not \U$37607 ( \37853 , \37852 );
and \U$37608 ( \37854 , \37853 , \686 );
nor \U$37609 ( \37855 , \643 , \685 );
nor \U$37610 ( \37856 , \37854 , \37855 );
or \U$37611 ( \37857 , \37856 , \737 );
not \U$37612 ( \37858 , \692 );
nand \U$37613 ( \37859 , \37858 , \736 );
nand \U$37614 ( \37860 , \37857 , \37859 );
and \U$37615 ( \37861 , \37860 , \774 );
nor \U$37616 ( \37862 , \744 , \773 );
nor \U$37617 ( \37863 , \37861 , \37862 );
nor \U$37618 ( \37864 , \37850 , \37863 );
not \U$37619 ( \37865 , \836 );
not \U$37620 ( \37866 , \804 );
nor \U$37621 ( \37867 , \37866 , \809 );
not \U$37622 ( \37868 , \37867 );
or \U$37623 ( \37869 , \37865 , \37868 );
or \U$37624 ( \37870 , \829 , \835 );
nand \U$37625 ( \37871 , \37869 , \37870 );
or \U$37626 ( \37872 , \37864 , \37871 );
and \U$37627 ( \37873 , \37872 , \853 );
nor \U$37628 ( \37874 , \840 , \852 );
nor \U$37629 ( \37875 , \37873 , \37874 );
nand \U$37630 ( \37876 , \37849 , \37875 );
not \U$37631 ( \37877 , \783 );
or \U$37632 ( \37878 , \413 , \446 );
nand \U$37633 ( \37879 , \37878 , RIbe27b98_2);
not \U$37634 ( \37880 , \37879 );
not \U$37635 ( \37881 , \824 );
and \U$37636 ( \37882 , \37880 , \37881 );
and \U$37637 ( \37883 , \37879 , \824 );
nor \U$37638 ( \37884 , \37882 , \37883 );
not \U$37639 ( \37885 , \37884 );
or \U$37640 ( \37886 , \37877 , \37885 );
or \U$37641 ( \37887 , \37884 , \783 );
nand \U$37642 ( \37888 , \37886 , \37887 );
not \U$37643 ( \37889 , \37888 );
or \U$37644 ( \37890 , \843 , \851 );
or \U$37645 ( \37891 , \848 , \783 );
nand \U$37646 ( \37892 , \37890 , \37891 );
not \U$37647 ( \37893 , \37892 );
or \U$37648 ( \37894 , \37889 , \37893 );
or \U$37649 ( \37895 , \37892 , \37888 );
nand \U$37650 ( \37896 , \37894 , \37895 );
not \U$37651 ( \37897 , \37896 );
and \U$37652 ( \37898 , \37876 , \37897 );
not \U$37653 ( \37899 , \37876 );
and \U$37654 ( \37900 , \37899 , \37896 );
nor \U$37655 ( \37901 , \37898 , \37900 );
buf \U$37656 ( \37902 , \37901 );
not \U$37657 ( \37903 , \837 );
and \U$37658 ( \37904 , \18571 , \18572 , \18574 );
nand \U$37659 ( \37905 , \37843 , \37904 , \18565 , \18570 );
not \U$37660 ( \37906 , \37905 );
not \U$37661 ( \37907 , \14234 );
or \U$37662 ( \37908 , \37906 , \37907 );
nand \U$37663 ( \37909 , \37908 , \7201 );
not \U$37664 ( \37910 , \18566 );
nand \U$37665 ( \37911 , \37803 , \18575 , \18565 , \22679 );
not \U$37666 ( \37912 , \37911 );
or \U$37667 ( \37913 , \37910 , \37912 );
nand \U$37668 ( \37914 , \37913 , \7201 );
buf \U$37669 ( \37915 , \7157 );
not \U$37670 ( \37916 , \37915 );
nand \U$37671 ( \37917 , \37909 , \37914 , \37916 );
and \U$37672 ( \37918 , \2202 , \775 );
and \U$37673 ( \37919 , \37917 , \37918 );
not \U$37674 ( \37920 , \37919 );
or \U$37675 ( \37921 , \37903 , \37920 );
nand \U$37676 ( \37922 , \7189 , \775 );
nand \U$37677 ( \37923 , \37922 , \37863 );
and \U$37678 ( \37924 , \37923 , \837 );
nor \U$37679 ( \37925 , \37924 , \37871 );
nand \U$37680 ( \37926 , \37921 , \37925 );
not \U$37681 ( \37927 , \37874 );
nand \U$37682 ( \37928 , \37927 , \853 );
not \U$37683 ( \37929 , \37928 );
and \U$37684 ( \37930 , \37926 , \37929 );
not \U$37685 ( \37931 , \37926 );
and \U$37686 ( \37932 , \37931 , \37928 );
nor \U$37687 ( \37933 , \37930 , \37932 );
buf \U$37688 ( \37934 , \37933 );
not \U$37689 ( \37935 , \810 );
not \U$37690 ( \37936 , \37919 );
or \U$37691 ( \37937 , \37935 , \37936 );
and \U$37692 ( \37938 , \37923 , \810 );
nor \U$37693 ( \37939 , \37938 , \37867 );
nand \U$37694 ( \37940 , \37937 , \37939 );
nand \U$37695 ( \37941 , \37870 , \836 );
not \U$37696 ( \37942 , \37941 );
and \U$37697 ( \37943 , \37940 , \37942 );
not \U$37698 ( \37944 , \37940 );
and \U$37699 ( \37945 , \37944 , \37941 );
nor \U$37700 ( \37946 , \37943 , \37945 );
buf \U$37701 ( \37947 , \37946 );
not \U$37702 ( \37948 , \775 );
not \U$37703 ( \37949 , \37847 );
or \U$37704 ( \37950 , \37948 , \37949 );
buf \U$37705 ( \37951 , \37863 );
nand \U$37706 ( \37952 , \37950 , \37951 );
not \U$37707 ( \37953 , \37867 );
nand \U$37708 ( \37954 , \37953 , \810 );
not \U$37709 ( \37955 , \37954 );
and \U$37710 ( \37956 , \37952 , \37955 );
not \U$37711 ( \37957 , \37952 );
and \U$37712 ( \37958 , \37957 , \37954 );
nor \U$37713 ( \37959 , \37956 , \37958 );
buf \U$37714 ( \37960 , \37959 );
not \U$37715 ( \37961 , \738 );
not \U$37716 ( \37962 , \7191 );
nand \U$37717 ( \37963 , \37962 , \18568 , \37846 );
not \U$37718 ( \37964 , \37963 );
or \U$37719 ( \37965 , \37961 , \37964 );
not \U$37720 ( \37966 , \37860 );
nand \U$37721 ( \37967 , \37965 , \37966 );
not \U$37722 ( \37968 , \37862 );
nand \U$37723 ( \37969 , \37968 , \774 );
not \U$37724 ( \37970 , \37969 );
and \U$37725 ( \37971 , \37967 , \37970 );
not \U$37726 ( \37972 , \37967 );
and \U$37727 ( \37973 , \37972 , \37969 );
nor \U$37728 ( \37974 , \37971 , \37973 );
buf \U$37729 ( \37975 , \37974 );
not \U$37730 ( \37976 , \687 );
not \U$37731 ( \37977 , \37847 );
or \U$37732 ( \37978 , \37976 , \37977 );
nand \U$37733 ( \37979 , \37978 , \37856 );
not \U$37734 ( \37980 , \737 );
nand \U$37735 ( \37981 , \37980 , \37859 );
not \U$37736 ( \37982 , \37981 );
and \U$37737 ( \37983 , \37979 , \37982 );
not \U$37738 ( \37984 , \37979 );
and \U$37739 ( \37985 , \37984 , \37981 );
nor \U$37740 ( \37986 , \37983 , \37985 );
buf \U$37741 ( \37987 , \37986 );
not \U$37742 ( \37988 , \639 );
not \U$37743 ( \37989 , \37847 );
or \U$37744 ( \37990 , \37988 , \37989 );
nand \U$37745 ( \37991 , \37990 , \37852 );
not \U$37746 ( \37992 , \37855 );
nand \U$37747 ( \37993 , \37992 , \686 );
not \U$37748 ( \37994 , \37993 );
and \U$37749 ( \37995 , \37991 , \37994 );
not \U$37750 ( \37996 , \37991 );
and \U$37751 ( \37997 , \37996 , \37993 );
nor \U$37752 ( \37998 , \37995 , \37997 );
buf \U$37753 ( \37999 , \37998 );
nand \U$37754 ( \38000 , \639 , \37852 );
xnor \U$37755 ( \38001 , \38000 , \37963 );
buf \U$37756 ( \38002 , \38001 );
not \U$37757 ( \38003 , \2194 );
and \U$37758 ( \38004 , \7201 , \2101 );
nand \U$37759 ( \38005 , \37845 , \18576 , \38004 );
not \U$37760 ( \38006 , \18566 );
not \U$37761 ( \38007 , \14234 );
or \U$37762 ( \38008 , \38006 , \38007 );
nand \U$37763 ( \38009 , \38008 , \38004 );
nand \U$37764 ( \38010 , \7157 , \2101 );
nand \U$37765 ( \38011 , \38005 , \38009 , \38010 );
not \U$37766 ( \38012 , \38011 );
or \U$37767 ( \38013 , \38003 , \38012 );
not \U$37768 ( \38014 , \7184 );
nand \U$37769 ( \38015 , \38013 , \38014 );
nand \U$37770 ( \38016 , \2201 , \7188 );
not \U$37771 ( \38017 , \38016 );
and \U$37772 ( \38018 , \38015 , \38017 );
not \U$37773 ( \38019 , \38015 );
and \U$37774 ( \38020 , \38019 , \38016 );
nor \U$37775 ( \38021 , \38018 , \38020 );
buf \U$37776 ( \38022 , \38021 );
not \U$37777 ( \38023 , \2173 );
not \U$37778 ( \38024 , \7172 );
nand \U$37779 ( \38025 , \38024 , \38010 , \38005 , \38009 );
not \U$37780 ( \38026 , \38025 );
or \U$37781 ( \38027 , \38023 , \38026 );
nand \U$37782 ( \38028 , \38027 , \7179 );
not \U$37783 ( \38029 , \7182 );
nand \U$37784 ( \38030 , \38029 , \2193 );
not \U$37785 ( \38031 , \38030 );
and \U$37786 ( \38032 , \38028 , \38031 );
not \U$37787 ( \38033 , \38028 );
and \U$37788 ( \38034 , \38033 , \38030 );
nor \U$37789 ( \38035 , \38032 , \38034 );
buf \U$37790 ( \38036 , \38035 );
buf \U$37791 ( \38037 , \2148 );
not \U$37792 ( \38038 , \38037 );
not \U$37793 ( \38039 , \38025 );
or \U$37794 ( \38040 , \38038 , \38039 );
not \U$37795 ( \38041 , \7176 );
nand \U$37796 ( \38042 , \38040 , \38041 );
not \U$37797 ( \38043 , \7178 );
nand \U$37798 ( \38044 , \38043 , \2172 );
not \U$37799 ( \38045 , \38044 );
and \U$37800 ( \38046 , \38042 , \38045 );
not \U$37801 ( \38047 , \38042 );
and \U$37802 ( \38048 , \38047 , \38044 );
nor \U$37803 ( \38049 , \38046 , \38048 );
buf \U$37804 ( \38050 , \38049 );
nand \U$37805 ( \38051 , \38041 , \38037 );
not \U$37806 ( \38052 , \38051 );
not \U$37807 ( \38053 , \38025 );
or \U$37808 ( \38054 , \38052 , \38053 );
or \U$37809 ( \38055 , \38051 , \38025 );
nand \U$37810 ( \38056 , \38054 , \38055 );
buf \U$37811 ( \38057 , \38056 );
and \U$37812 ( \38058 , \37911 , \37905 , \18566 , \14234 );
not \U$37813 ( \38059 , \38058 );
and \U$37814 ( \38060 , \7201 , \1872 );
nand \U$37815 ( \38061 , \38059 , \38060 );
nand \U$37816 ( \38062 , \2094 , \7171 );
nand \U$37817 ( \38063 , \38062 , \2100 );
or \U$37818 ( \38064 , \38061 , \38063 );
not \U$37819 ( \38065 , \38060 );
not \U$37820 ( \38066 , \38059 );
or \U$37821 ( \38067 , \38065 , \38066 );
not \U$37822 ( \38068 , \1872 );
not \U$37823 ( \38069 , \37915 );
or \U$37824 ( \38070 , \38068 , \38069 );
not \U$37825 ( \38071 , \7164 );
nand \U$37826 ( \38072 , \38070 , \38071 );
not \U$37827 ( \38073 , \38062 );
nand \U$37828 ( \38074 , \38073 , \7166 );
nor \U$37829 ( \38075 , \38072 , \38074 );
nand \U$37830 ( \38076 , \38067 , \38075 );
not \U$37831 ( \38077 , \38062 );
not \U$37832 ( \38078 , \2100 );
and \U$37833 ( \38079 , \38077 , \38078 );
not \U$37834 ( \38080 , \2100 );
not \U$37835 ( \38081 , \38072 );
or \U$37836 ( \38082 , \38080 , \38081 );
nand \U$37837 ( \38083 , \38082 , \7166 );
and \U$37838 ( \38084 , \38083 , \38062 );
nor \U$37839 ( \38085 , \38079 , \38084 );
nand \U$37840 ( \38086 , \38064 , \38076 , \38085 );
buf \U$37841 ( \38087 , \38086 );
not \U$37842 ( \38088 , \38060 );
not \U$37843 ( \38089 , \38058 );
not \U$37844 ( \38090 , \38089 );
or \U$37845 ( \38091 , \38088 , \38090 );
not \U$37846 ( \38092 , \38072 );
nand \U$37847 ( \38093 , \38091 , \38092 );
nand \U$37848 ( \38094 , \2100 , \7166 );
not \U$37849 ( \38095 , \38094 );
and \U$37850 ( \38096 , \38093 , \38095 );
not \U$37851 ( \38097 , \38093 );
and \U$37852 ( \38098 , \38097 , \38094 );
nor \U$37853 ( \38099 , \38096 , \38098 );
buf \U$37854 ( \38100 , \38099 );
not \U$37855 ( \38101 , \1871 );
buf \U$37856 ( \38102 , \37917 );
not \U$37857 ( \38103 , \38102 );
or \U$37858 ( \38104 , \38101 , \38103 );
nand \U$37859 ( \38105 , \38104 , \7161 );
nand \U$37860 ( \38106 , \1669 , \7163 );
not \U$37861 ( \38107 , \38106 );
and \U$37862 ( \38108 , \38105 , \38107 );
not \U$37863 ( \38109 , \38105 );
and \U$37864 ( \38110 , \38109 , \38106 );
nor \U$37865 ( \38111 , \38108 , \38110 );
buf \U$37866 ( \38112 , \38111 );
nand \U$37867 ( \38113 , \7161 , \1871 );
not \U$37868 ( \38114 , \38113 );
and \U$37869 ( \38115 , \38102 , \38114 );
not \U$37870 ( \38116 , \38102 );
and \U$37871 ( \38117 , \38116 , \38113 );
nor \U$37872 ( \38118 , \38115 , \38117 );
buf \U$37873 ( \38119 , \38118 );
not \U$37874 ( \38120 , \7153 );
not \U$37875 ( \38121 , \7199 );
nand \U$37876 ( \38122 , \38059 , \38121 , \7122 );
nand \U$37877 ( \38123 , \38120 , \38122 );
nand \U$37878 ( \38124 , \2360 , \7156 );
not \U$37879 ( \38125 , \38124 );
and \U$37880 ( \38126 , \38123 , \38125 );
not \U$37881 ( \38127 , \38123 );
and \U$37882 ( \38128 , \38127 , \38124 );
nor \U$37883 ( \38129 , \38126 , \38128 );
buf \U$37884 ( \38130 , \38129 );
not \U$37885 ( \38131 , \7124 );
and \U$37886 ( \38132 , \38121 , \7053 );
and \U$37887 ( \38133 , \38089 , \38132 );
not \U$37888 ( \38134 , \38133 );
or \U$37889 ( \38135 , \38131 , \38134 );
not \U$37890 ( \38136 , \7142 );
not \U$37891 ( \38137 , \6431 );
not \U$37892 ( \38138 , \38137 );
nand \U$37893 ( \38139 , \38138 , \7053 );
nand \U$37894 ( \38140 , \38136 , \38139 );
and \U$37895 ( \38141 , \38140 , \7124 );
not \U$37896 ( \38142 , \7148 );
nor \U$37897 ( \38143 , \38141 , \38142 );
nand \U$37898 ( \38144 , \38135 , \38143 );
nand \U$37899 ( \38145 , \7150 , \7152 );
not \U$37900 ( \38146 , \38145 );
and \U$37901 ( \38147 , \38144 , \38146 );
not \U$37902 ( \38148 , \38144 );
and \U$37903 ( \38149 , \38148 , \38145 );
nor \U$37904 ( \38150 , \38147 , \38149 );
buf \U$37905 ( \38151 , \38150 );
buf \U$37906 ( \38152 , \7112 );
not \U$37907 ( \38153 , \38152 );
not \U$37908 ( \38154 , \38133 );
or \U$37909 ( \38155 , \38153 , \38154 );
and \U$37910 ( \38156 , \38140 , \38152 );
nor \U$37911 ( \38157 , \38156 , \7145 );
nand \U$37912 ( \38158 , \38155 , \38157 );
not \U$37913 ( \38159 , \7147 );
nand \U$37914 ( \38160 , \38159 , \7099 );
not \U$37915 ( \38161 , \38160 );
and \U$37916 ( \38162 , \38158 , \38161 );
not \U$37917 ( \38163 , \38158 );
and \U$37918 ( \38164 , \38163 , \38160 );
nor \U$37919 ( \38165 , \38162 , \38164 );
buf \U$37920 ( \38166 , \38165 );
not \U$37921 ( \38167 , \38132 );
not \U$37922 ( \38168 , \38059 );
or \U$37923 ( \38169 , \38167 , \38168 );
not \U$37924 ( \38170 , \38140 );
nand \U$37925 ( \38171 , \38169 , \38170 );
not \U$37926 ( \38172 , \7145 );
nand \U$37927 ( \38173 , \38172 , \38152 );
not \U$37928 ( \38174 , \38173 );
and \U$37929 ( \38175 , \38171 , \38174 );
not \U$37930 ( \38176 , \38171 );
and \U$37931 ( \38177 , \38176 , \38173 );
nor \U$37932 ( \38178 , \38175 , \38177 );
buf \U$37933 ( \38179 , \38178 );
not \U$37934 ( \38180 , \6966 );
not \U$37935 ( \38181 , \38180 );
not \U$37936 ( \38182 , \6973 );
nor \U$37937 ( \38183 , \7199 , \38182 );
and \U$37938 ( \38184 , \38089 , \38183 );
not \U$37939 ( \38185 , \38184 );
or \U$37940 ( \38186 , \38181 , \38185 );
not \U$37941 ( \38187 , \6941 );
not \U$37942 ( \38188 , \6965 );
nor \U$37943 ( \38189 , \38137 , \38182 );
not \U$37944 ( \38190 , \38189 );
or \U$37945 ( \38191 , \38188 , \38190 );
not \U$37946 ( \38192 , \7134 );
nand \U$37947 ( \38193 , \38191 , \38192 );
not \U$37948 ( \38194 , \38193 );
or \U$37949 ( \38195 , \38187 , \38194 );
nand \U$37950 ( \38196 , \38195 , \7138 );
not \U$37951 ( \38197 , \38196 );
nand \U$37952 ( \38198 , \38186 , \38197 );
nand \U$37953 ( \38199 , \7051 , \7141 );
not \U$37954 ( \38200 , \38199 );
and \U$37955 ( \38201 , \38198 , \38200 );
not \U$37956 ( \38202 , \38198 );
and \U$37957 ( \38203 , \38202 , \38199 );
nor \U$37958 ( \38204 , \38201 , \38203 );
buf \U$37959 ( \38205 , \38204 );
not \U$37960 ( \38206 , \6965 );
not \U$37961 ( \38207 , \38184 );
or \U$37962 ( \38208 , \38206 , \38207 );
not \U$37963 ( \38209 , \38193 );
nand \U$37964 ( \38210 , \38208 , \38209 );
nand \U$37965 ( \38211 , \6941 , \7138 );
not \U$37966 ( \38212 , \38211 );
and \U$37967 ( \38213 , \38210 , \38212 );
not \U$37968 ( \38214 , \38210 );
and \U$37969 ( \38215 , \38214 , \38211 );
nor \U$37970 ( \38216 , \38213 , \38215 );
buf \U$37971 ( \38217 , \38216 );
not \U$37972 ( \38218 , \38183 );
not \U$37973 ( \38219 , \38089 );
or \U$37974 ( \38220 , \38218 , \38219 );
buf \U$37975 ( \38221 , \7128 );
nor \U$37976 ( \38222 , \38189 , \38221 );
nand \U$37977 ( \38223 , \38220 , \38222 );
nand \U$37978 ( \38224 , \7133 , \6965 );
not \U$37979 ( \38225 , \38224 );
and \U$37980 ( \38226 , \38223 , \38225 );
not \U$37981 ( \38227 , \38223 );
and \U$37982 ( \38228 , \38227 , \38224 );
nor \U$37983 ( \38229 , \38226 , \38228 );
buf \U$37984 ( \38230 , \38229 );
not \U$37985 ( \38231 , \38121 );
not \U$37986 ( \38232 , \38089 );
or \U$37987 ( \38233 , \38231 , \38232 );
not \U$37988 ( \38234 , \38138 );
nand \U$37989 ( \38235 , \38233 , \38234 );
nor \U$37990 ( \38236 , \38221 , \38182 );
and \U$37991 ( \38237 , \38235 , \38236 );
not \U$37992 ( \38238 , \38235 );
not \U$37993 ( \38239 , \38236 );
and \U$37994 ( \38240 , \38238 , \38239 );
nor \U$37995 ( \38241 , \38237 , \38240 );
buf \U$37996 ( \38242 , \38241 );
buf \U$37997 ( \38243 , \5900 );
and \U$37998 ( \38244 , \7198 , \38243 );
not \U$37999 ( \38245 , \38244 );
not \U$38000 ( \38246 , \38059 );
or \U$38001 ( \38247 , \38245 , \38246 );
not \U$38002 ( \38248 , \38243 );
not \U$38003 ( \38249 , \7195 );
not \U$38004 ( \38250 , \4308 );
not \U$38005 ( \38251 , \5110 );
buf \U$38006 ( \38252 , \4753 );
nand \U$38007 ( \38253 , \38251 , \38252 );
nand \U$38008 ( \38254 , \38253 , \5113 );
not \U$38009 ( \38255 , \38254 );
or \U$38010 ( \38256 , \38250 , \38255 );
buf \U$38011 ( \38257 , \5116 );
nand \U$38012 ( \38258 , \38256 , \38257 );
not \U$38013 ( \38259 , \38258 );
or \U$38014 ( \38260 , \38249 , \38259 );
buf \U$38015 ( \38261 , \5376 );
nand \U$38016 ( \38262 , \38260 , \38261 );
not \U$38017 ( \38263 , \38262 );
or \U$38018 ( \38264 , \38248 , \38263 );
not \U$38019 ( \38265 , \6425 );
nand \U$38020 ( \38266 , \38264 , \38265 );
not \U$38021 ( \38267 , \38266 );
nand \U$38022 ( \38268 , \38247 , \38267 );
and \U$38023 ( \38269 , \6412 , \6430 );
nand \U$38024 ( \38270 , \38269 , \6417 );
or \U$38025 ( \38271 , \38268 , \38270 );
not \U$38026 ( \38272 , \6164 );
nor \U$38027 ( \38273 , \38269 , \38272 );
and \U$38028 ( \38274 , \38059 , \38244 , \38273 );
and \U$38029 ( \38275 , \38269 , \38272 );
not \U$38030 ( \38276 , \38269 );
not \U$38031 ( \38277 , \6164 );
not \U$38032 ( \38278 , \38266 );
or \U$38033 ( \38279 , \38277 , \38278 );
nand \U$38034 ( \38280 , \38279 , \6417 );
and \U$38035 ( \38281 , \38276 , \38280 );
or \U$38036 ( \38282 , \38275 , \38281 );
nor \U$38037 ( \38283 , \38274 , \38282 );
nand \U$38038 ( \38284 , \38271 , \38283 );
buf \U$38039 ( \38285 , \38284 );
nand \U$38040 ( \38286 , \6164 , \6417 );
not \U$38041 ( \38287 , \38286 );
and \U$38042 ( \38288 , \38268 , \38287 );
not \U$38043 ( \38289 , \38268 );
and \U$38044 ( \38290 , \38289 , \38286 );
nor \U$38045 ( \38291 , \38288 , \38290 );
buf \U$38046 ( \38292 , \38291 );
not \U$38047 ( \38293 , \7198 );
not \U$38048 ( \38294 , \38059 );
or \U$38049 ( \38295 , \38293 , \38294 );
not \U$38050 ( \38296 , \38262 );
nand \U$38051 ( \38297 , \38295 , \38296 );
not \U$38052 ( \38298 , \6419 );
nand \U$38053 ( \38299 , \38298 , \6424 );
not \U$38054 ( \38300 , \38299 );
nand \U$38055 ( \38301 , \38300 , \6422 );
or \U$38056 ( \38302 , \38297 , \38301 );
and \U$38057 ( \38303 , \38299 , \5634 );
and \U$38058 ( \38304 , \38059 , \38303 , \7198 );
or \U$38059 ( \38305 , \38299 , \5634 );
not \U$38060 ( \38306 , \5634 );
not \U$38061 ( \38307 , \38262 );
or \U$38062 ( \38308 , \38306 , \38307 );
nand \U$38063 ( \38309 , \38308 , \6422 );
nand \U$38064 ( \38310 , \38309 , \38299 );
nand \U$38065 ( \38311 , \38305 , \38310 );
nor \U$38066 ( \38312 , \38304 , \38311 );
nand \U$38067 ( \38313 , \38302 , \38312 );
buf \U$38068 ( \38314 , \38313 );
nand \U$38069 ( \38315 , \5634 , \6422 );
not \U$38070 ( \38316 , \38315 );
and \U$38071 ( \38317 , \38297 , \38316 );
not \U$38072 ( \38318 , \38297 );
and \U$38073 ( \38319 , \38318 , \38315 );
nor \U$38074 ( \38320 , \38317 , \38319 );
buf \U$38075 ( \38321 , \38320 );
not \U$38076 ( \38322 , \7197 );
not \U$38077 ( \38323 , \38322 );
and \U$38078 ( \38324 , \38089 , \7194 );
not \U$38079 ( \38325 , \38324 );
or \U$38080 ( \38326 , \38323 , \38325 );
not \U$38081 ( \38327 , \38258 );
nand \U$38082 ( \38328 , \38326 , \38327 );
nand \U$38083 ( \38329 , \7195 , \38261 );
not \U$38084 ( \38330 , \38329 );
and \U$38085 ( \38331 , \38328 , \38330 );
not \U$38086 ( \38332 , \38328 );
and \U$38087 ( \38333 , \38332 , \38329 );
nor \U$38088 ( \38334 , \38331 , \38333 );
buf \U$38089 ( \38335 , \38334 );
not \U$38090 ( \38336 , \38252 );
not \U$38091 ( \38337 , \38324 );
or \U$38092 ( \38338 , \38336 , \38337 );
not \U$38093 ( \38339 , \38254 );
nand \U$38094 ( \38340 , \38338 , \38339 );
nand \U$38095 ( \38341 , \4308 , \38257 );
not \U$38096 ( \38342 , \38341 );
and \U$38097 ( \38343 , \38340 , \38342 );
not \U$38098 ( \38344 , \38340 );
and \U$38099 ( \38345 , \38344 , \38341 );
nor \U$38100 ( \38346 , \38343 , \38345 );
buf \U$38101 ( \38347 , \38346 );
not \U$38102 ( \38348 , \7194 );
not \U$38103 ( \38349 , \38089 );
or \U$38104 ( \38350 , \38348 , \38349 );
buf \U$38105 ( \38351 , \5110 );
nand \U$38106 ( \38352 , \38350 , \38351 );
nand \U$38107 ( \38353 , \5113 , \38252 );
not \U$38108 ( \38354 , \38353 );
and \U$38109 ( \38355 , \38352 , \38354 );
not \U$38110 ( \38356 , \38352 );
and \U$38111 ( \38357 , \38356 , \38353 );
nor \U$38112 ( \38358 , \38355 , \38357 );
buf \U$38113 ( \38359 , \38358 );
nand \U$38114 ( \38360 , \7194 , \38351 );
not \U$38115 ( \38361 , \38059 );
and \U$38116 ( \38362 , \38360 , \38361 );
not \U$38117 ( \38363 , \38360 );
not \U$38118 ( \38364 , \38361 );
and \U$38119 ( \38365 , \38363 , \38364 );
nor \U$38120 ( \38366 , \38362 , \38365 );
buf \U$38121 ( \38367 , \38366 );
buf \U$38122 ( \38368 , \14154 );
and \U$38123 ( \38369 , \18563 , \38368 );
not \U$38124 ( \38370 , \38369 );
not \U$38125 ( \38371 , \18558 );
nand \U$38126 ( \38372 , \37803 , \18575 , \22679 );
nand \U$38127 ( \38373 , \37843 , \18575 );
nand \U$38128 ( \38374 , \38371 , \38372 , \38373 );
not \U$38129 ( \38375 , \38374 );
or \U$38130 ( \38376 , \38370 , \38375 );
not \U$38131 ( \38377 , \14189 );
not \U$38132 ( \38378 , \13975 );
buf \U$38133 ( \38379 , \13707 );
not \U$38134 ( \38380 , \38379 );
or \U$38135 ( \38381 , \38378 , \38380 );
not \U$38136 ( \38382 , \14190 );
nand \U$38137 ( \38383 , \38381 , \38382 );
not \U$38138 ( \38384 , \38383 );
or \U$38139 ( \38385 , \38377 , \38384 );
buf \U$38140 ( \38386 , \14187 );
nand \U$38141 ( \38387 , \38385 , \38386 );
and \U$38142 ( \38388 , \38387 , \38368 );
nor \U$38143 ( \38389 , \38388 , \14214 );
nand \U$38144 ( \38390 , \38376 , \38389 );
nand \U$38145 ( \38391 , \14229 , \14160 );
not \U$38146 ( \38392 , \14173 );
nor \U$38147 ( \38393 , \38391 , \38392 );
not \U$38148 ( \38394 , \38393 );
or \U$38149 ( \38395 , \38390 , \38394 );
not \U$38150 ( \38396 , \14216 );
and \U$38151 ( \38397 , \38393 , \38396 );
nor \U$38152 ( \38398 , \38392 , \8520 );
nor \U$38153 ( \38399 , \38397 , \38398 );
nand \U$38154 ( \38400 , \38395 , \38399 );
nand \U$38155 ( \38401 , \14184 , \14233 );
and \U$38156 ( \38402 , \38400 , \38401 );
not \U$38157 ( \38403 , \38400 );
not \U$38158 ( \38404 , \38401 );
and \U$38159 ( \38405 , \38403 , \38404 );
nor \U$38160 ( \38406 , \38402 , \38405 );
buf \U$38161 ( \38407 , \38406 );
not \U$38162 ( \38408 , \8519 );
nor \U$38163 ( \38409 , \38408 , \14164 );
not \U$38164 ( \38410 , \38409 );
not \U$38165 ( \38411 , \18564 );
buf \U$38166 ( \38412 , \38374 );
not \U$38167 ( \38413 , \38412 );
or \U$38168 ( \38414 , \38411 , \38413 );
buf \U$38169 ( \38415 , \14230 );
buf \U$38170 ( \38416 , \14161 );
nor \U$38171 ( \38417 , \38415 , \38416 );
nand \U$38172 ( \38418 , \38414 , \38417 );
not \U$38173 ( \38419 , \38418 );
or \U$38174 ( \38420 , \38410 , \38419 );
not \U$38175 ( \38421 , \14170 );
nand \U$38176 ( \38422 , \38420 , \38421 );
not \U$38177 ( \38423 , \14172 );
nand \U$38178 ( \38424 , \38423 , \8128 );
not \U$38179 ( \38425 , \38424 );
and \U$38180 ( \38426 , \38422 , \38425 );
not \U$38181 ( \38427 , \38422 );
and \U$38182 ( \38428 , \38427 , \38424 );
nor \U$38183 ( \38429 , \38426 , \38428 );
buf \U$38184 ( \38430 , \38429 );
not \U$38185 ( \38431 , \38418 );
not \U$38186 ( \38432 , \8519 );
or \U$38187 ( \38433 , \38431 , \38432 );
nand \U$38188 ( \38434 , \38433 , \14167 );
nand \U$38189 ( \38435 , \8103 , \14169 );
not \U$38190 ( \38436 , \38435 );
and \U$38191 ( \38437 , \38434 , \38436 );
not \U$38192 ( \38438 , \38434 );
and \U$38193 ( \38439 , \38438 , \38435 );
nor \U$38194 ( \38440 , \38437 , \38439 );
buf \U$38195 ( \38441 , \38440 );
nand \U$38196 ( \38442 , \14167 , \8519 );
not \U$38197 ( \38443 , \38442 );
not \U$38198 ( \38444 , \38418 );
or \U$38199 ( \38445 , \38443 , \38444 );
or \U$38200 ( \38446 , \38442 , \38418 );
nand \U$38201 ( \38447 , \38445 , \38446 );
buf \U$38202 ( \38448 , \38447 );
not \U$38203 ( \38449 , \14159 );
nand \U$38204 ( \38450 , \38449 , \14157 );
and \U$38205 ( \38451 , \38450 , \10382 );
not \U$38206 ( \38452 , \38451 );
not \U$38207 ( \38453 , \10346 );
not \U$38208 ( \38454 , \38453 );
not \U$38209 ( \38455 , \38390 );
or \U$38210 ( \38456 , \38454 , \38455 );
not \U$38211 ( \38457 , \14228 );
nand \U$38212 ( \38458 , \38456 , \38457 );
not \U$38213 ( \38459 , \38458 );
or \U$38214 ( \38460 , \38452 , \38459 );
nor \U$38215 ( \38461 , \14228 , \38450 , \14156 );
not \U$38216 ( \38462 , \38461 );
nand \U$38217 ( \38463 , \38390 , \38453 );
not \U$38218 ( \38464 , \38463 );
or \U$38219 ( \38465 , \38462 , \38464 );
not \U$38220 ( \38466 , \38450 );
not \U$38221 ( \38467 , \10382 );
and \U$38222 ( \38468 , \38466 , \38467 );
and \U$38223 ( \38469 , \38450 , \14156 );
nor \U$38224 ( \38470 , \38468 , \38469 );
nand \U$38225 ( \38471 , \38465 , \38470 );
not \U$38226 ( \38472 , \38471 );
nand \U$38227 ( \38473 , \38460 , \38472 );
buf \U$38228 ( \38474 , \38473 );
not \U$38229 ( \38475 , \14156 );
nand \U$38230 ( \38476 , \38475 , \10382 );
not \U$38231 ( \38477 , \38476 );
not \U$38232 ( \38478 , \38458 );
or \U$38233 ( \38479 , \38477 , \38478 );
or \U$38234 ( \38480 , \38458 , \38476 );
nand \U$38235 ( \38481 , \38479 , \38480 );
buf \U$38236 ( \38482 , \38481 );
not \U$38237 ( \38483 , \10289 );
not \U$38238 ( \38484 , \38390 );
or \U$38239 ( \38485 , \38483 , \38484 );
nand \U$38240 ( \38486 , \38485 , \14223 );
not \U$38241 ( \38487 , \14219 );
nand \U$38242 ( \38488 , \38487 , \14227 );
not \U$38243 ( \38489 , \38488 );
and \U$38244 ( \38490 , \38486 , \38489 );
not \U$38245 ( \38491 , \38486 );
and \U$38246 ( \38492 , \38491 , \38488 );
nor \U$38247 ( \38493 , \38490 , \38492 );
buf \U$38248 ( \38494 , \38493 );
nand \U$38249 ( \38495 , \10289 , \14223 );
not \U$38250 ( \38496 , \38495 );
and \U$38251 ( \38497 , \38390 , \38496 );
not \U$38252 ( \38498 , \38390 );
and \U$38253 ( \38499 , \38498 , \38495 );
nor \U$38254 ( \38500 , \38497 , \38499 );
buf \U$38255 ( \38501 , \38500 );
not \U$38256 ( \38502 , \18563 );
not \U$38257 ( \38503 , \38412 );
or \U$38258 ( \38504 , \38502 , \38503 );
not \U$38259 ( \38505 , \38387 );
nand \U$38260 ( \38506 , \38504 , \38505 );
not \U$38261 ( \38507 , \14110 );
nand \U$38262 ( \38508 , \38506 , \38507 );
not \U$38263 ( \38509 , \14152 );
not \U$38264 ( \38510 , \38509 );
nand \U$38265 ( \38511 , \14131 , \14212 );
nand \U$38266 ( \38512 , \38510 , \38511 );
or \U$38267 ( \38513 , \38508 , \38512 );
nor \U$38268 ( \38514 , \38511 , \14209 , \14204 );
nand \U$38269 ( \38515 , \38508 , \38514 );
not \U$38270 ( \38516 , \14204 );
or \U$38271 ( \38517 , \38516 , \38509 );
nand \U$38272 ( \38518 , \38517 , \14208 );
and \U$38273 ( \38519 , \38511 , \38518 );
not \U$38274 ( \38520 , \38511 );
and \U$38275 ( \38521 , \38520 , \38509 );
nor \U$38276 ( \38522 , \38519 , \38521 );
nand \U$38277 ( \38523 , \38513 , \38515 , \38522 );
buf \U$38278 ( \38524 , \38523 );
nand \U$38279 ( \38525 , \38508 , \38516 );
nand \U$38280 ( \38526 , \14152 , \14208 );
not \U$38281 ( \38527 , \38526 );
and \U$38282 ( \38528 , \38525 , \38527 );
not \U$38283 ( \38529 , \38525 );
and \U$38284 ( \38530 , \38529 , \38526 );
nor \U$38285 ( \38531 , \38528 , \38530 );
buf \U$38286 ( \38532 , \38531 );
not \U$38287 ( \38533 , \14109 );
not \U$38288 ( \38534 , \38506 );
or \U$38289 ( \38535 , \38533 , \38534 );
nand \U$38290 ( \38536 , \38535 , \14200 );
not \U$38291 ( \38537 , \14201 );
nand \U$38292 ( \38538 , \38537 , \14203 );
not \U$38293 ( \38539 , \38538 );
and \U$38294 ( \38540 , \38536 , \38539 );
not \U$38295 ( \38541 , \38536 );
and \U$38296 ( \38542 , \38541 , \38538 );
nor \U$38297 ( \38543 , \38540 , \38542 );
buf \U$38298 ( \38544 , \38543 );
nand \U$38299 ( \38545 , \14109 , \14200 );
not \U$38300 ( \38546 , \38545 );
and \U$38301 ( \38547 , \38506 , \38546 );
not \U$38302 ( \38548 , \38506 );
and \U$38303 ( \38549 , \38548 , \38545 );
nor \U$38304 ( \38550 , \38547 , \38549 );
buf \U$38305 ( \38551 , \38550 );
not \U$38306 ( \38552 , \13975 );
not \U$38307 ( \38553 , \18562 );
and \U$38308 ( \38554 , \38412 , \38553 );
not \U$38309 ( \38555 , \38554 );
or \U$38310 ( \38556 , \38552 , \38555 );
not \U$38311 ( \38557 , \38383 );
nand \U$38312 ( \38558 , \38556 , \38557 );
nand \U$38313 ( \38559 , \14189 , \38386 );
not \U$38314 ( \38560 , \38559 );
and \U$38315 ( \38561 , \38558 , \38560 );
not \U$38316 ( \38562 , \38558 );
and \U$38317 ( \38563 , \38562 , \38559 );
nor \U$38318 ( \38564 , \38561 , \38563 );
buf \U$38319 ( \38565 , \38564 );
not \U$38320 ( \38566 , \38553 );
not \U$38321 ( \38567 , \38412 );
or \U$38322 ( \38568 , \38566 , \38567 );
not \U$38323 ( \38569 , \38379 );
nand \U$38324 ( \38570 , \38568 , \38569 );
nand \U$38325 ( \38571 , \38382 , \13975 );
not \U$38326 ( \38572 , \38571 );
and \U$38327 ( \38573 , \38570 , \38572 );
not \U$38328 ( \38574 , \38570 );
and \U$38329 ( \38575 , \38574 , \38571 );
nor \U$38330 ( \38576 , \38573 , \38575 );
buf \U$38331 ( \38577 , \38576 );
not \U$38332 ( \38578 , \18561 );
not \U$38333 ( \38579 , \38412 );
or \U$38334 ( \38580 , \38578 , \38579 );
nand \U$38335 ( \38581 , \38580 , \13701 );
nand \U$38336 ( \38582 , \13706 , \18560 );
not \U$38337 ( \38583 , \38582 );
and \U$38338 ( \38584 , \38581 , \38583 );
not \U$38339 ( \38585 , \38581 );
and \U$38340 ( \38586 , \38585 , \38582 );
nor \U$38341 ( \38587 , \38584 , \38586 );
buf \U$38342 ( \38588 , \38587 );
nand \U$38343 ( \38589 , \18561 , \13701 );
not \U$38344 ( \38590 , \38589 );
not \U$38345 ( \38591 , \38412 );
or \U$38346 ( \38592 , \38590 , \38591 );
or \U$38347 ( \38593 , \38589 , \38412 );
nand \U$38348 ( \38594 , \38592 , \38593 );
buf \U$38349 ( \38595 , \38594 );
not \U$38350 ( \38596 , \18556 );
nand \U$38351 ( \38597 , \38596 , \18538 );
buf \U$38352 ( \38598 , \18522 );
nand \U$38353 ( \38599 , \38597 , \38598 );
not \U$38354 ( \38600 , \37904 );
not \U$38355 ( \38601 , \37845 );
or \U$38356 ( \38602 , \38600 , \38601 );
and \U$38357 ( \38603 , \18355 , \18357 , \18492 );
not \U$38358 ( \38604 , \16622 );
nor \U$38359 ( \38605 , \38603 , \38604 );
nand \U$38360 ( \38606 , \38602 , \38605 );
nand \U$38361 ( \38607 , \38606 , \18490 );
or \U$38362 ( \38608 , \38599 , \38607 );
nor \U$38363 ( \38609 , \18554 , \38597 );
nand \U$38364 ( \38610 , \38607 , \38609 );
not \U$38365 ( \38611 , \18551 );
nand \U$38366 ( \38612 , \38611 , \38598 );
nand \U$38367 ( \38613 , \38612 , \18553 );
and \U$38368 ( \38614 , \38597 , \38613 );
not \U$38369 ( \38615 , \38597 );
not \U$38370 ( \38616 , \38598 );
and \U$38371 ( \38617 , \38615 , \38616 );
nor \U$38372 ( \38618 , \38614 , \38617 );
nand \U$38373 ( \38619 , \38608 , \38610 , \38618 );
buf \U$38374 ( \38620 , \38619 );
not \U$38375 ( \38621 , \38611 );
nand \U$38376 ( \38622 , \38607 , \38621 );
nand \U$38377 ( \38623 , \38598 , \18553 );
not \U$38378 ( \38624 , \38623 );
and \U$38379 ( \38625 , \38622 , \38624 );
not \U$38380 ( \38626 , \38622 );
and \U$38381 ( \38627 , \38626 , \38623 );
nor \U$38382 ( \38628 , \38625 , \38627 );
buf \U$38383 ( \38629 , \38628 );
buf \U$38384 ( \38630 , \18440 );
not \U$38385 ( \38631 , \38630 );
not \U$38386 ( \38632 , \38606 );
or \U$38387 ( \38633 , \38631 , \38632 );
buf \U$38388 ( \38634 , \18543 );
nand \U$38389 ( \38635 , \38633 , \38634 );
nor \U$38390 ( \38636 , \18550 , \18545 );
and \U$38391 ( \38637 , \38635 , \38636 );
not \U$38392 ( \38638 , \38635 );
not \U$38393 ( \38639 , \38636 );
and \U$38394 ( \38640 , \38638 , \38639 );
nor \U$38395 ( \38641 , \38637 , \38640 );
buf \U$38396 ( \38642 , \38641 );
nand \U$38397 ( \38643 , \38630 , \38634 );
not \U$38398 ( \38644 , \38643 );
and \U$38399 ( \38645 , \38606 , \38644 );
not \U$38400 ( \38646 , \38606 );
and \U$38401 ( \38647 , \38646 , \38643 );
nor \U$38402 ( \38648 , \38645 , \38647 );
buf \U$38403 ( \38649 , \38648 );
nand \U$38404 ( \38650 , \18571 , \18574 );
nor \U$38405 ( \38651 , \38650 , \18356 );
not \U$38406 ( \38652 , \38651 );
buf \U$38407 ( \38653 , \37845 );
not \U$38408 ( \38654 , \38653 );
or \U$38409 ( \38655 , \38652 , \38654 );
nand \U$38410 ( \38656 , \38655 , \18358 );
nand \U$38411 ( \38657 , \18492 , \16622 );
not \U$38412 ( \38658 , \38657 );
and \U$38413 ( \38659 , \38656 , \38658 );
not \U$38414 ( \38660 , \38656 );
and \U$38415 ( \38661 , \38660 , \38657 );
nor \U$38416 ( \38662 , \38659 , \38661 );
buf \U$38417 ( \38663 , \38662 );
not \U$38418 ( \38664 , \38650 );
not \U$38419 ( \38665 , \38664 );
not \U$38420 ( \38666 , \38653 );
or \U$38421 ( \38667 , \38665 , \38666 );
buf \U$38422 ( \38668 , \18305 );
not \U$38423 ( \38669 , \38668 );
buf \U$38424 ( \38670 , \18352 );
nand \U$38425 ( \38671 , \38669 , \38670 );
nand \U$38426 ( \38672 , \38671 , \18571 );
nand \U$38427 ( \38673 , \38667 , \38672 );
not \U$38428 ( \38674 , \18356 );
nand \U$38429 ( \38675 , \38674 , \18348 );
not \U$38430 ( \38676 , \38675 );
and \U$38431 ( \38677 , \38673 , \38676 );
not \U$38432 ( \38678 , \38673 );
and \U$38433 ( \38679 , \38678 , \38675 );
nor \U$38434 ( \38680 , \38677 , \38679 );
buf \U$38435 ( \38681 , \38680 );
not \U$38436 ( \38682 , \18574 );
not \U$38437 ( \38683 , \38653 );
or \U$38438 ( \38684 , \38682 , \38683 );
buf \U$38439 ( \38685 , \38669 );
nand \U$38440 ( \38686 , \38684 , \38685 );
nand \U$38441 ( \38687 , \38670 , \18571 );
not \U$38442 ( \38688 , \38687 );
and \U$38443 ( \38689 , \38686 , \38688 );
not \U$38444 ( \38690 , \38686 );
and \U$38445 ( \38691 , \38690 , \38687 );
nor \U$38446 ( \38692 , \38689 , \38691 );
buf \U$38447 ( \38693 , \38692 );
not \U$38448 ( \38694 , \38668 );
nand \U$38449 ( \38695 , \38694 , \18574 );
not \U$38450 ( \38696 , \38695 );
not \U$38451 ( \38697 , \38653 );
or \U$38452 ( \38698 , \38696 , \38697 );
or \U$38453 ( \38699 , \38653 , \38695 );
nand \U$38454 ( \38700 , \38698 , \38699 );
buf \U$38455 ( \38701 , \38700 );
not \U$38456 ( \38702 , \22632 );
not \U$38457 ( \38703 , \22678 );
not \U$38458 ( \38704 , \22514 );
not \U$38459 ( \38705 , \22160 );
nor \U$38460 ( \38706 , \38704 , \38705 );
not \U$38461 ( \38707 , \38706 );
buf \U$38462 ( \38708 , \37803 );
not \U$38463 ( \38709 , \38708 );
or \U$38464 ( \38710 , \38707 , \38709 );
not \U$38465 ( \38711 , \37826 );
nand \U$38466 ( \38712 , \38710 , \38711 );
not \U$38467 ( \38713 , \38712 );
or \U$38468 ( \38714 , \38703 , \38713 );
not \U$38469 ( \38715 , \37836 );
nand \U$38470 ( \38716 , \38714 , \38715 );
not \U$38471 ( \38717 , \38716 );
or \U$38472 ( \38718 , \38702 , \38717 );
not \U$38473 ( \38719 , \37837 );
nand \U$38474 ( \38720 , \38718 , \38719 );
nand \U$38475 ( \38721 , \37840 , \22642 );
not \U$38476 ( \38722 , \38721 );
and \U$38477 ( \38723 , \38720 , \38722 );
not \U$38478 ( \38724 , \38720 );
and \U$38479 ( \38725 , \38724 , \38721 );
nor \U$38480 ( \38726 , \38723 , \38725 );
buf \U$38481 ( \38727 , \38726 );
nand \U$38482 ( \38728 , \38719 , \22632 );
not \U$38483 ( \38729 , \38728 );
and \U$38484 ( \38730 , \38716 , \38729 );
not \U$38485 ( \38731 , \38716 );
and \U$38486 ( \38732 , \38731 , \38728 );
nor \U$38487 ( \38733 , \38730 , \38732 );
buf \U$38488 ( \38734 , \38733 );
not \U$38489 ( \38735 , \22669 );
not \U$38490 ( \38736 , \38712 );
or \U$38491 ( \38737 , \38735 , \38736 );
not \U$38492 ( \38738 , \37829 );
nand \U$38493 ( \38739 , \38737 , \38738 );
nand \U$38494 ( \38740 , \37835 , \22676 );
not \U$38495 ( \38741 , \38740 );
and \U$38496 ( \38742 , \38739 , \38741 );
not \U$38497 ( \38743 , \38739 );
and \U$38498 ( \38744 , \38743 , \38740 );
nor \U$38499 ( \38745 , \38742 , \38744 );
buf \U$38500 ( \38746 , \38745 );
nand \U$38501 ( \38747 , \22669 , \38738 );
not \U$38502 ( \38748 , \38747 );
and \U$38503 ( \38749 , \38712 , \38748 );
not \U$38504 ( \38750 , \38712 );
and \U$38505 ( \38751 , \38750 , \38747 );
nor \U$38506 ( \38752 , \38749 , \38751 );
buf \U$38507 ( \38753 , \38752 );
buf \U$38508 ( \38754 , \22382 );
not \U$38509 ( \38755 , \38754 );
not \U$38510 ( \38756 , \38705 );
not \U$38511 ( \38757 , \38756 );
not \U$38512 ( \38758 , \38708 );
or \U$38513 ( \38759 , \38757 , \38758 );
not \U$38514 ( \38760 , \37814 );
nand \U$38515 ( \38761 , \38759 , \38760 );
not \U$38516 ( \38762 , \38761 );
or \U$38517 ( \38763 , \38755 , \38762 );
buf \U$38518 ( \38764 , \37819 );
not \U$38519 ( \38765 , \38764 );
nand \U$38520 ( \38766 , \38763 , \38765 );
nand \U$38521 ( \38767 , \37823 , \22513 );
not \U$38522 ( \38768 , \38767 );
and \U$38523 ( \38769 , \38766 , \38768 );
not \U$38524 ( \38770 , \38766 );
and \U$38525 ( \38771 , \38770 , \38767 );
nor \U$38526 ( \38772 , \38769 , \38771 );
buf \U$38527 ( \38773 , \38772 );
not \U$38528 ( \38774 , \38764 );
nand \U$38529 ( \38775 , \38774 , \38754 );
not \U$38530 ( \38776 , \38775 );
and \U$38531 ( \38777 , \38761 , \38776 );
not \U$38532 ( \38778 , \38761 );
and \U$38533 ( \38779 , \38778 , \38775 );
nor \U$38534 ( \38780 , \38777 , \38779 );
buf \U$38535 ( \38781 , \38780 );
not \U$38536 ( \38782 , \22159 );
not \U$38537 ( \38783 , \38708 );
or \U$38538 ( \38784 , \38782 , \38783 );
not \U$38539 ( \38785 , \37809 );
nand \U$38540 ( \38786 , \38784 , \38785 );
nand \U$38541 ( \38787 , \21682 , \37813 );
not \U$38542 ( \38788 , \38787 );
and \U$38543 ( \38789 , \38786 , \38788 );
not \U$38544 ( \38790 , \38786 );
and \U$38545 ( \38791 , \38790 , \38787 );
nor \U$38546 ( \38792 , \38789 , \38791 );
buf \U$38547 ( \38793 , \38792 );
nand \U$38548 ( \38794 , \38785 , \22159 );
not \U$38549 ( \38795 , \38794 );
not \U$38550 ( \38796 , \38708 );
or \U$38551 ( \38797 , \38795 , \38796 );
or \U$38552 ( \38798 , \38794 , \38708 );
nand \U$38553 ( \38799 , \38797 , \38798 );
buf \U$38554 ( \38800 , \38799 );
not \U$38555 ( \38801 , \29295 );
not \U$38556 ( \38802 , \29270 );
not \U$38557 ( \38803 , \37801 );
not \U$38558 ( \38804 , \37794 );
or \U$38559 ( \38805 , \38803 , \38804 );
not \U$38560 ( \38806 , \28180 );
nand \U$38561 ( \38807 , \38805 , \38806 );
not \U$38562 ( \38808 , \38807 );
or \U$38563 ( \38809 , \38802 , \38808 );
not \U$38564 ( \38810 , \29289 );
nand \U$38565 ( \38811 , \38809 , \38810 );
buf \U$38566 ( \38812 , \29101 );
nand \U$38567 ( \38813 , \38811 , \38812 );
not \U$38568 ( \38814 , \38813 );
or \U$38569 ( \38815 , \38801 , \38814 );
buf \U$38570 ( \38816 , \28949 );
nand \U$38571 ( \38817 , \38815 , \38816 );
not \U$38572 ( \38818 , \38817 );
buf \U$38573 ( \38819 , \28769 );
and \U$38574 ( \38820 , \38818 , \38819 );
not \U$38575 ( \38821 , \29299 );
nor \U$38576 ( \38822 , \38820 , \38821 );
nand \U$38577 ( \38823 , \29300 , \29303 );
and \U$38578 ( \38824 , \38822 , \38823 );
not \U$38579 ( \38825 , \38822 );
not \U$38580 ( \38826 , \38823 );
and \U$38581 ( \38827 , \38825 , \38826 );
nor \U$38582 ( \38828 , \38824 , \38827 );
buf \U$38583 ( \38829 , \38828 );
nand \U$38584 ( \38830 , \38819 , \29299 );
and \U$38585 ( \38831 , \38817 , \38830 );
not \U$38586 ( \38832 , \38817 );
not \U$38587 ( \38833 , \38830 );
and \U$38588 ( \38834 , \38832 , \38833 );
nor \U$38589 ( \38835 , \38831 , \38834 );
buf \U$38590 ( \38836 , \38835 );
nand \U$38591 ( \38837 , \38813 , \29293 );
nand \U$38592 ( \38838 , \38816 , \29294 );
not \U$38593 ( \38839 , \38838 );
and \U$38594 ( \38840 , \38837 , \38839 );
not \U$38595 ( \38841 , \38837 );
and \U$38596 ( \38842 , \38841 , \38838 );
nor \U$38597 ( \38843 , \38840 , \38842 );
buf \U$38598 ( \38844 , \38843 );
nand \U$38599 ( \38845 , \29293 , \38812 );
not \U$38600 ( \38846 , \38845 );
and \U$38601 ( \38847 , \38811 , \38846 );
not \U$38602 ( \38848 , \38811 );
and \U$38603 ( \38849 , \38848 , \38845 );
nor \U$38604 ( \38850 , \38847 , \38849 );
buf \U$38605 ( \38851 , \38850 );
not \U$38606 ( \38852 , \29218 );
buf \U$38607 ( \38853 , \29262 );
and \U$38608 ( \38854 , \38853 , \29269 );
not \U$38609 ( \38855 , \38854 );
not \U$38610 ( \38856 , \38807 );
or \U$38611 ( \38857 , \38855 , \38856 );
nand \U$38612 ( \38858 , \29281 , \38853 );
nand \U$38613 ( \38859 , \38857 , \38858 );
not \U$38614 ( \38860 , \38859 );
or \U$38615 ( \38861 , \38852 , \38860 );
not \U$38616 ( \38862 , \29283 );
nand \U$38617 ( \38863 , \38861 , \38862 );
nand \U$38618 ( \38864 , \29239 , \29286 );
not \U$38619 ( \38865 , \38864 );
and \U$38620 ( \38866 , \38863 , \38865 );
not \U$38621 ( \38867 , \38863 );
and \U$38622 ( \38868 , \38867 , \38864 );
nor \U$38623 ( \38869 , \38866 , \38868 );
buf \U$38624 ( \38870 , \38869 );
nand \U$38625 ( \38871 , \29218 , \38862 );
not \U$38626 ( \38872 , \38871 );
and \U$38627 ( \38873 , \38859 , \38872 );
not \U$38628 ( \38874 , \38859 );
and \U$38629 ( \38875 , \38874 , \38871 );
nor \U$38630 ( \38876 , \38873 , \38875 );
buf \U$38631 ( \38877 , \38876 );
not \U$38632 ( \38878 , \29269 );
not \U$38633 ( \38879 , \38807 );
or \U$38634 ( \38880 , \38878 , \38879 );
nand \U$38635 ( \38881 , \38880 , \29280 );
not \U$38636 ( \38882 , \29260 );
not \U$38637 ( \38883 , \29249 );
or \U$38638 ( \38884 , \38882 , \38883 );
nand \U$38639 ( \38885 , \38884 , \38853 );
not \U$38640 ( \38886 , \38885 );
and \U$38641 ( \38887 , \38881 , \38886 );
not \U$38642 ( \38888 , \38881 );
and \U$38643 ( \38889 , \38888 , \38885 );
nor \U$38644 ( \38890 , \38887 , \38889 );
buf \U$38645 ( \38891 , \38890 );
nand \U$38646 ( \38892 , \29269 , \29280 );
not \U$38647 ( \38893 , \38892 );
and \U$38648 ( \38894 , \38807 , \38893 );
not \U$38649 ( \38895 , \38807 );
and \U$38650 ( \38896 , \38895 , \38892 );
nor \U$38651 ( \38897 , \38894 , \38896 );
buf \U$38652 ( \38898 , \38897 );
not \U$38653 ( \38899 , \28163 );
not \U$38654 ( \38900 , \38899 );
not \U$38655 ( \38901 , \37800 );
not \U$38656 ( \38902 , \37799 );
buf \U$38657 ( \38903 , \37794 );
not \U$38658 ( \38904 , \38903 );
or \U$38659 ( \38905 , \38902 , \38904 );
nand \U$38660 ( \38906 , \26275 , \28103 );
nand \U$38661 ( \38907 , \38905 , \38906 );
not \U$38662 ( \38908 , \38907 );
or \U$38663 ( \38909 , \38901 , \38908 );
not \U$38664 ( \38910 , \28162 );
nand \U$38665 ( \38911 , \38909 , \38910 );
not \U$38666 ( \38912 , \38911 );
or \U$38667 ( \38913 , \38900 , \38912 );
nand \U$38668 ( \38914 , \38913 , \28174 );
nand \U$38669 ( \38915 , \28101 , \28168 );
not \U$38670 ( \38916 , \38915 );
and \U$38671 ( \38917 , \38914 , \38916 );
not \U$38672 ( \38918 , \38914 );
and \U$38673 ( \38919 , \38918 , \38915 );
nor \U$38674 ( \38920 , \38917 , \38919 );
buf \U$38675 ( \38921 , \38920 );
nand \U$38676 ( \38922 , \38899 , \28174 );
not \U$38677 ( \38923 , \38922 );
and \U$38678 ( \38924 , \38911 , \38923 );
not \U$38679 ( \38925 , \38911 );
and \U$38680 ( \38926 , \38925 , \38922 );
nor \U$38681 ( \38927 , \38924 , \38926 );
buf \U$38682 ( \38928 , \38927 );
not \U$38683 ( \38929 , \28140 );
not \U$38684 ( \38930 , \38907 );
or \U$38685 ( \38931 , \38929 , \38930 );
buf \U$38686 ( \38932 , \28160 );
nand \U$38687 ( \38933 , \38931 , \38932 );
nand \U$38688 ( \38934 , \28154 , \28159 );
not \U$38689 ( \38935 , \38934 );
and \U$38690 ( \38936 , \38933 , \38935 );
not \U$38691 ( \38937 , \38933 );
and \U$38692 ( \38938 , \38937 , \38934 );
nor \U$38693 ( \38939 , \38936 , \38938 );
buf \U$38694 ( \38940 , \38939 );
nand \U$38695 ( \38941 , \38932 , \28140 );
not \U$38696 ( \38942 , \38941 );
and \U$38697 ( \38943 , \38907 , \38942 );
not \U$38698 ( \38944 , \38907 );
and \U$38699 ( \38945 , \38944 , \38941 );
nor \U$38700 ( \38946 , \38943 , \38945 );
buf \U$38701 ( \38947 , \38946 );
not \U$38702 ( \38948 , \25387 );
not \U$38703 ( \38949 , \38948 );
nand \U$38704 ( \38950 , \37794 , \37798 );
not \U$38705 ( \38951 , \38950 );
or \U$38706 ( \38952 , \38949 , \38951 );
buf \U$38707 ( \38953 , \37797 );
nand \U$38708 ( \38954 , \38952 , \38953 );
not \U$38709 ( \38955 , \37796 );
or \U$38710 ( \38956 , \38954 , \38955 );
buf \U$38711 ( \38957 , \25801 );
nand \U$38712 ( \38958 , \38956 , \38957 );
nand \U$38713 ( \38959 , \26273 , \28103 );
not \U$38714 ( \38960 , \38959 );
and \U$38715 ( \38961 , \38958 , \38960 );
not \U$38716 ( \38962 , \38958 );
and \U$38717 ( \38963 , \38962 , \38959 );
nor \U$38718 ( \38964 , \38961 , \38963 );
buf \U$38719 ( \38965 , \38964 );
nand \U$38720 ( \38966 , \37796 , \38957 );
and \U$38721 ( \38967 , \38954 , \38966 );
not \U$38722 ( \38968 , \38954 );
not \U$38723 ( \38969 , \38966 );
and \U$38724 ( \38970 , \38968 , \38969 );
nor \U$38725 ( \38971 , \38967 , \38970 );
buf \U$38726 ( \38972 , \38971 );
nand \U$38727 ( \38973 , \25386 , \38950 );
nand \U$38728 ( \38974 , \38953 , \25349 );
not \U$38729 ( \38975 , \38974 );
and \U$38730 ( \38976 , \38973 , \38975 );
not \U$38731 ( \38977 , \38973 );
and \U$38732 ( \38978 , \38977 , \38974 );
nor \U$38733 ( \38979 , \38976 , \38978 );
buf \U$38734 ( \38980 , \38979 );
nand \U$38735 ( \38981 , \25386 , \37798 );
not \U$38736 ( \38982 , \38981 );
and \U$38737 ( \38983 , \38903 , \38982 );
not \U$38738 ( \38984 , \38903 );
and \U$38739 ( \38985 , \38984 , \38981 );
nor \U$38740 ( \38986 , \38983 , \38985 );
buf \U$38741 ( \38987 , \38986 );
not \U$38742 ( \38988 , \34286 );
not \U$38743 ( \38989 , \38988 );
not \U$38744 ( \38990 , \34308 );
not \U$38745 ( \38991 , \31902 );
buf \U$38746 ( \38992 , \34092 );
and \U$38747 ( \38993 , \37776 , \34306 );
nor \U$38748 ( \38994 , \38992 , \38993 );
not \U$38749 ( \38995 , \38994 );
not \U$38750 ( \38996 , \38995 );
or \U$38751 ( \38997 , \38991 , \38996 );
buf \U$38752 ( \38998 , \34110 );
nand \U$38753 ( \38999 , \38997 , \38998 );
not \U$38754 ( \39000 , \38999 );
or \U$38755 ( \39001 , \38990 , \39000 );
not \U$38756 ( \39002 , \37784 );
nand \U$38757 ( \39003 , \39001 , \39002 );
not \U$38758 ( \39004 , \39003 );
or \U$38759 ( \39005 , \38989 , \39004 );
not \U$38760 ( \39006 , \37788 );
nand \U$38761 ( \39007 , \39005 , \39006 );
nor \U$38762 ( \39008 , \37790 , \34293 );
and \U$38763 ( \39009 , \39007 , \39008 );
not \U$38764 ( \39010 , \39007 );
not \U$38765 ( \39011 , \39008 );
and \U$38766 ( \39012 , \39010 , \39011 );
nor \U$38767 ( \39013 , \39009 , \39012 );
buf \U$38768 ( \39014 , \39013 );
nand \U$38769 ( \39015 , \38988 , \39006 );
not \U$38770 ( \39016 , \39015 );
and \U$38771 ( \39017 , \39003 , \39016 );
not \U$38772 ( \39018 , \39003 );
and \U$38773 ( \39019 , \39018 , \39015 );
nor \U$38774 ( \39020 , \39017 , \39019 );
buf \U$38775 ( \39021 , \39020 );
not \U$38776 ( \39022 , \34301 );
not \U$38777 ( \39023 , \38999 );
or \U$38778 ( \39024 , \39022 , \39023 );
not \U$38779 ( \39025 , \37780 );
nand \U$38780 ( \39026 , \39024 , \39025 );
nand \U$38781 ( \39027 , \34263 , \37783 );
not \U$38782 ( \39028 , \39027 );
and \U$38783 ( \39029 , \39026 , \39028 );
not \U$38784 ( \39030 , \39026 );
and \U$38785 ( \39031 , \39030 , \39027 );
nor \U$38786 ( \39032 , \39029 , \39031 );
buf \U$38787 ( \39033 , \39032 );
nand \U$38788 ( \39034 , \39025 , \34301 );
not \U$38789 ( \39035 , \39034 );
and \U$38790 ( \39036 , \38999 , \39035 );
not \U$38791 ( \39037 , \38999 );
and \U$38792 ( \39038 , \39037 , \39034 );
nor \U$38793 ( \39039 , \39036 , \39038 );
buf \U$38794 ( \39040 , \39039 );
not \U$38795 ( \39041 , \34095 );
not \U$38796 ( \39042 , \31901 );
not \U$38797 ( \39043 , \31891 );
not \U$38798 ( \39044 , \38995 );
or \U$38799 ( \39045 , \39043 , \39044 );
buf \U$38800 ( \39046 , \34097 );
not \U$38801 ( \39047 , \39046 );
nand \U$38802 ( \39048 , \39045 , \39047 );
not \U$38803 ( \39049 , \39048 );
or \U$38804 ( \39050 , \39042 , \39049 );
nand \U$38805 ( \39051 , \39050 , \34103 );
not \U$38806 ( \39052 , \39051 );
or \U$38807 ( \39053 , \39041 , \39052 );
nand \U$38808 ( \39054 , \39053 , \34101 );
nand \U$38809 ( \39055 , \34109 , \34107 );
not \U$38810 ( \39056 , \39055 );
and \U$38811 ( \39057 , \39054 , \39056 );
not \U$38812 ( \39058 , \39054 );
and \U$38813 ( \39059 , \39058 , \39055 );
nor \U$38814 ( \39060 , \39057 , \39059 );
buf \U$38815 ( \39061 , \39060 );
nand \U$38816 ( \39062 , \34101 , \34095 );
not \U$38817 ( \39063 , \39062 );
and \U$38818 ( \39064 , \39051 , \39063 );
not \U$38819 ( \39065 , \39051 );
and \U$38820 ( \39066 , \39065 , \39062 );
nor \U$38821 ( \39067 , \39064 , \39066 );
buf \U$38822 ( \39068 , \39067 );
nand \U$38823 ( \39069 , \31901 , \34103 );
not \U$38824 ( \39070 , \39069 );
and \U$38825 ( \39071 , \39048 , \39070 );
not \U$38826 ( \39072 , \39048 );
and \U$38827 ( \39073 , \39072 , \39069 );
nor \U$38828 ( \39074 , \39071 , \39073 );
buf \U$38829 ( \39075 , \39074 );
not \U$38830 ( \39076 , \38994 );
not \U$38831 ( \39077 , \31891 );
nor \U$38832 ( \39078 , \39077 , \39046 );
not \U$38833 ( \39079 , \39078 );
or \U$38834 ( \39080 , \39076 , \39079 );
or \U$38835 ( \39081 , \39078 , \38994 );
nand \U$38836 ( \39082 , \39080 , \39081 );
buf \U$38837 ( \39083 , \39082 );
buf \U$38838 ( \39084 , \34030 );
not \U$38839 ( \39085 , \39084 );
and \U$38840 ( \39086 , \33640 , \34305 );
not \U$38841 ( \39087 , \39086 );
not \U$38842 ( \39088 , \37776 );
or \U$38843 ( \39089 , \39087 , \39088 );
buf \U$38844 ( \39090 , \33888 );
nand \U$38845 ( \39091 , \39089 , \39090 );
buf \U$38846 ( \39092 , \34073 );
nand \U$38847 ( \39093 , \39091 , \39092 );
buf \U$38848 ( \39094 , \34053 );
not \U$38849 ( \39095 , \39094 );
or \U$38850 ( \39096 , \39093 , \39095 );
not \U$38851 ( \39097 , \34086 );
nand \U$38852 ( \39098 , \39096 , \39097 );
not \U$38853 ( \39099 , \39098 );
or \U$38854 ( \39100 , \39085 , \39099 );
nand \U$38855 ( \39101 , \39100 , \34089 );
nand \U$38856 ( \39102 , \34088 , \33961 );
not \U$38857 ( \39103 , \39102 );
and \U$38858 ( \39104 , \39101 , \39103 );
not \U$38859 ( \39105 , \39101 );
and \U$38860 ( \39106 , \39105 , \39102 );
nor \U$38861 ( \39107 , \39104 , \39106 );
buf \U$38862 ( \39108 , \39107 );
nand \U$38863 ( \39109 , \39084 , \34089 );
not \U$38864 ( \39110 , \39109 );
and \U$38865 ( \39111 , \39098 , \39110 );
not \U$38866 ( \39112 , \39098 );
and \U$38867 ( \39113 , \39112 , \39109 );
nor \U$38868 ( \39114 , \39111 , \39113 );
buf \U$38869 ( \39115 , \39114 );
buf \U$38870 ( \39116 , \34080 );
nand \U$38871 ( \39117 , \39093 , \39116 );
nand \U$38872 ( \39118 , \34085 , \39094 );
not \U$38873 ( \39119 , \39118 );
and \U$38874 ( \39120 , \39117 , \39119 );
not \U$38875 ( \39121 , \39117 );
and \U$38876 ( \39122 , \39121 , \39118 );
nor \U$38877 ( \39123 , \39120 , \39122 );
buf \U$38878 ( \39124 , \39123 );
nand \U$38879 ( \39125 , \39092 , \39116 );
not \U$38880 ( \39126 , \39125 );
and \U$38881 ( \39127 , \39091 , \39126 );
not \U$38882 ( \39128 , \39091 );
and \U$38883 ( \39129 , \39128 , \39125 );
nor \U$38884 ( \39130 , \39127 , \39129 );
buf \U$38885 ( \39131 , \39130 );
not \U$38886 ( \39132 , \33225 );
not \U$38887 ( \39133 , \39132 );
not \U$38888 ( \39134 , \33639 );
not \U$38889 ( \39135 , \39134 );
not \U$38890 ( \39136 , \34304 );
and \U$38891 ( \39137 , \37776 , \39136 );
not \U$38892 ( \39138 , \39137 );
or \U$38893 ( \39139 , \39135 , \39138 );
nand \U$38894 ( \39140 , \33882 , \39134 );
nand \U$38895 ( \39141 , \39139 , \39140 );
not \U$38896 ( \39142 , \39141 );
or \U$38897 ( \39143 , \39133 , \39142 );
nand \U$38898 ( \39144 , \39143 , \33221 );
nand \U$38899 ( \39145 , \33887 , \33182 );
not \U$38900 ( \39146 , \39145 );
and \U$38901 ( \39147 , \39144 , \39146 );
not \U$38902 ( \39148 , \39144 );
and \U$38903 ( \39149 , \39148 , \39145 );
nor \U$38904 ( \39150 , \39147 , \39149 );
buf \U$38905 ( \39151 , \39150 );
nand \U$38906 ( \39152 , \39132 , \33221 );
not \U$38907 ( \39153 , \39152 );
and \U$38908 ( \39154 , \39141 , \39153 );
not \U$38909 ( \39155 , \39141 );
and \U$38910 ( \39156 , \39155 , \39152 );
nor \U$38911 ( \39157 , \39154 , \39156 );
buf \U$38912 ( \39158 , \39157 );
not \U$38913 ( \39159 , \39137 );
nand \U$38914 ( \39160 , \39159 , \33881 );
nand \U$38915 ( \39161 , \39134 , \33641 );
not \U$38916 ( \39162 , \39161 );
and \U$38917 ( \39163 , \39160 , \39162 );
not \U$38918 ( \39164 , \39160 );
and \U$38919 ( \39165 , \39164 , \39161 );
nor \U$38920 ( \39166 , \39163 , \39165 );
buf \U$38921 ( \39167 , \39166 );
nand \U$38922 ( \39168 , \33881 , \39136 );
not \U$38923 ( \39169 , \39168 );
and \U$38924 ( \39170 , \37776 , \39169 );
not \U$38925 ( \39171 , \37776 );
and \U$38926 ( \39172 , \39171 , \39168 );
nor \U$38927 ( \39173 , \39170 , \39172 );
buf \U$38928 ( \39174 , \39173 );
not \U$38929 ( \39175 , \35830 );
not \U$38930 ( \39176 , \35805 );
not \U$38931 ( \39177 , \39176 );
not \U$38932 ( \39178 , \35681 );
not \U$38933 ( \39179 , \39178 );
not \U$38934 ( \39180 , \37746 );
or \U$38935 ( \39181 , \39179 , \39180 );
not \U$38936 ( \39182 , \37757 );
nand \U$38937 ( \39183 , \39181 , \39182 );
not \U$38938 ( \39184 , \39183 );
or \U$38939 ( \39185 , \39177 , \39184 );
not \U$38940 ( \39186 , \37766 );
nand \U$38941 ( \39187 , \39185 , \39186 );
not \U$38942 ( \39188 , \39187 );
or \U$38943 ( \39189 , \39175 , \39188 );
nand \U$38944 ( \39190 , \39189 , \37771 );
nand \U$38945 ( \39191 , \37775 , \37773 );
not \U$38946 ( \39192 , \39191 );
and \U$38947 ( \39193 , \39190 , \39192 );
not \U$38948 ( \39194 , \39190 );
and \U$38949 ( \39195 , \39194 , \39191 );
nor \U$38950 ( \39196 , \39193 , \39195 );
buf \U$38951 ( \39197 , \39196 );
nand \U$38952 ( \39198 , \35830 , \37771 );
not \U$38953 ( \39199 , \39198 );
and \U$38954 ( \39200 , \39187 , \39199 );
not \U$38955 ( \39201 , \39187 );
and \U$38956 ( \39202 , \39201 , \39198 );
nor \U$38957 ( \39203 , \39200 , \39202 );
buf \U$38958 ( \39204 , \39203 );
not \U$38959 ( \39205 , \35747 );
not \U$38960 ( \39206 , \39183 );
or \U$38961 ( \39207 , \39205 , \39206 );
nand \U$38962 ( \39208 , \39207 , \37761 );
nand \U$38963 ( \39209 , \35804 , \37765 );
not \U$38964 ( \39210 , \39209 );
and \U$38965 ( \39211 , \39208 , \39210 );
not \U$38966 ( \39212 , \39208 );
and \U$38967 ( \39213 , \39212 , \39209 );
nor \U$38968 ( \39214 , \39211 , \39213 );
buf \U$38969 ( \39215 , \39214 );
nand \U$38970 ( \39216 , \35747 , \37761 );
not \U$38971 ( \39217 , \39216 );
and \U$38972 ( \39218 , \39183 , \39217 );
not \U$38973 ( \39219 , \39183 );
and \U$38974 ( \39220 , \39219 , \39216 );
nor \U$38975 ( \39221 , \39218 , \39220 );
buf \U$38976 ( \39222 , \39221 );
not \U$38977 ( \39223 , \35336 );
not \U$38978 ( \39224 , \39223 );
nand \U$38979 ( \39225 , \37746 , \35672 );
not \U$38980 ( \39226 , \35680 );
or \U$38981 ( \39227 , \39225 , \39226 );
not \U$38982 ( \39228 , \37752 );
nand \U$38983 ( \39229 , \39227 , \39228 );
not \U$38984 ( \39230 , \39229 );
or \U$38985 ( \39231 , \39224 , \39230 );
not \U$38986 ( \39232 , \37753 );
nand \U$38987 ( \39233 , \39231 , \39232 );
not \U$38988 ( \39234 , \35128 );
nand \U$38989 ( \39235 , \39234 , \37756 );
not \U$38990 ( \39236 , \39235 );
and \U$38991 ( \39237 , \39233 , \39236 );
not \U$38992 ( \39238 , \39233 );
and \U$38993 ( \39239 , \39238 , \39235 );
nor \U$38994 ( \39240 , \39237 , \39239 );
buf \U$38995 ( \39241 , \39240 );
nand \U$38996 ( \39242 , \39232 , \39223 );
not \U$38997 ( \39243 , \39242 );
and \U$38998 ( \39244 , \39229 , \39243 );
not \U$38999 ( \39245 , \39229 );
and \U$39000 ( \39246 , \39245 , \39242 );
nor \U$39001 ( \39247 , \39244 , \39246 );
buf \U$39002 ( \39248 , \39247 );
nand \U$39003 ( \39249 , \39225 , \37749 );
nand \U$39004 ( \39250 , \35680 , \37751 );
not \U$39005 ( \39251 , \39250 );
and \U$39006 ( \39252 , \39249 , \39251 );
not \U$39007 ( \39253 , \39249 );
and \U$39008 ( \39254 , \39253 , \39250 );
nor \U$39009 ( \39255 , \39252 , \39254 );
buf \U$39010 ( \39256 , \39255 );
nand \U$39011 ( \39257 , \35672 , \37749 );
not \U$39012 ( \39258 , \39257 );
and \U$39013 ( \39259 , \37746 , \39258 );
not \U$39014 ( \39260 , \37746 );
and \U$39015 ( \39261 , \39260 , \39257 );
nor \U$39016 ( \39262 , \39259 , \39261 );
buf \U$39017 ( \39263 , \39262 );
not \U$39018 ( \39264 , \36084 );
not \U$39019 ( \39265 , \39264 );
not \U$39020 ( \39266 , \36309 );
and \U$39021 ( \39267 , \37729 , \36441 );
not \U$39022 ( \39268 , \39267 );
or \U$39023 ( \39269 , \39266 , \39268 );
not \U$39024 ( \39270 , \37735 );
nand \U$39025 ( \39271 , \39269 , \39270 );
not \U$39026 ( \39272 , \39271 );
or \U$39027 ( \39273 , \39265 , \39272 );
not \U$39028 ( \39274 , \37740 );
nand \U$39029 ( \39275 , \39273 , \39274 );
nor \U$39030 ( \39276 , \35910 , \37742 );
and \U$39031 ( \39277 , \39275 , \39276 );
not \U$39032 ( \39278 , \39275 );
not \U$39033 ( \39279 , \39276 );
and \U$39034 ( \39280 , \39278 , \39279 );
nor \U$39035 ( \39281 , \39277 , \39280 );
buf \U$39036 ( \39282 , \39281 );
nand \U$39037 ( \39283 , \39274 , \39264 );
not \U$39038 ( \39284 , \39283 );
and \U$39039 ( \39285 , \39271 , \39284 );
not \U$39040 ( \39286 , \39271 );
and \U$39041 ( \39287 , \39286 , \39283 );
nor \U$39042 ( \39288 , \39285 , \39287 );
buf \U$39043 ( \39289 , \39288 );
not \U$39044 ( \39290 , \39267 );
buf \U$39045 ( \39291 , \37732 );
nand \U$39046 ( \39292 , \39290 , \39291 );
nand \U$39047 ( \39293 , \36309 , \37734 );
not \U$39048 ( \39294 , \39293 );
and \U$39049 ( \39295 , \39292 , \39294 );
not \U$39050 ( \39296 , \39292 );
and \U$39051 ( \39297 , \39296 , \39293 );
nor \U$39052 ( \39298 , \39295 , \39297 );
buf \U$39053 ( \39299 , \39298 );
nand \U$39054 ( \39300 , \39291 , \36441 );
xnor \U$39055 ( \39301 , \37729 , \39300 );
buf \U$39056 ( \39302 , \39301 );
not \U$39057 ( \39303 , \36727 );
not \U$39058 ( \39304 , \37718 );
buf \U$39059 ( \39305 , \37671 );
not \U$39060 ( \39306 , \39305 );
or \U$39061 ( \39307 , \39304 , \39306 );
not \U$39062 ( \39308 , \37723 );
nand \U$39063 ( \39309 , \39307 , \39308 );
not \U$39064 ( \39310 , \39309 );
or \U$39065 ( \39311 , \39303 , \39310 );
not \U$39066 ( \39312 , \37725 );
nand \U$39067 ( \39313 , \39311 , \39312 );
not \U$39068 ( \39314 , \37727 );
nand \U$39069 ( \39315 , \39314 , \36590 );
not \U$39070 ( \39316 , \39315 );
and \U$39071 ( \39317 , \39313 , \39316 );
not \U$39072 ( \39318 , \39313 );
and \U$39073 ( \39319 , \39318 , \39315 );
nor \U$39074 ( \39320 , \39317 , \39319 );
buf \U$39075 ( \39321 , \39320 );
nand \U$39076 ( \39322 , \39312 , \36727 );
not \U$39077 ( \39323 , \39322 );
not \U$39078 ( \39324 , \39309 );
or \U$39079 ( \39325 , \39323 , \39324 );
or \U$39080 ( \39326 , \39322 , \39309 );
nand \U$39081 ( \39327 , \39325 , \39326 );
buf \U$39082 ( \39328 , \39327 );
not \U$39083 ( \39329 , \37717 );
not \U$39084 ( \39330 , \39329 );
not \U$39085 ( \39331 , \39305 );
or \U$39086 ( \39332 , \39330 , \39331 );
nand \U$39087 ( \39333 , \39332 , \37720 );
not \U$39088 ( \39334 , \37703 );
nand \U$39089 ( \39335 , \39334 , \37722 );
not \U$39090 ( \39336 , \39335 );
and \U$39091 ( \39337 , \39333 , \39336 );
not \U$39092 ( \39338 , \39333 );
and \U$39093 ( \39339 , \39338 , \39335 );
nor \U$39094 ( \39340 , \39337 , \39339 );
buf \U$39095 ( \39341 , \39340 );
nand \U$39096 ( \39342 , \37720 , \39329 );
not \U$39097 ( \39343 , \39342 );
and \U$39098 ( \39344 , \39305 , \39343 );
not \U$39099 ( \39345 , \39305 );
and \U$39100 ( \39346 , \39345 , \39342 );
nor \U$39101 ( \39347 , \39344 , \39346 );
buf \U$39102 ( \39348 , \39347 );
not \U$39103 ( \39349 , \37103 );
nand \U$39104 ( \39350 , \37655 , \37661 );
not \U$39105 ( \39351 , \39350 );
or \U$39106 ( \39352 , \39349 , \39351 );
nand \U$39107 ( \39353 , \39352 , \37665 );
not \U$39108 ( \39354 , \37663 );
nand \U$39109 ( \39355 , \39354 , \37668 );
not \U$39110 ( \39356 , \39355 );
and \U$39111 ( \39357 , \39353 , \39356 );
not \U$39112 ( \39358 , \39353 );
and \U$39113 ( \39359 , \39358 , \39355 );
nor \U$39114 ( \39360 , \39357 , \39359 );
buf \U$39115 ( \39361 , \39360 );
nand \U$39116 ( \39362 , \37665 , \37103 );
not \U$39117 ( \39363 , \39362 );
and \U$39118 ( \39364 , \39350 , \39363 );
not \U$39119 ( \39365 , \39350 );
and \U$39120 ( \39366 , \39365 , \39362 );
nor \U$39121 ( \39367 , \39364 , \39366 );
buf \U$39122 ( \39368 , \39367 );
not \U$39123 ( \39369 , \37653 );
not \U$39124 ( \39370 , \39369 );
not \U$39125 ( \39371 , \37618 );
or \U$39126 ( \39372 , \39370 , \39371 );
not \U$39127 ( \39373 , \37657 );
nand \U$39128 ( \39374 , \39372 , \39373 );
nor \U$39129 ( \39375 , \37660 , \37642 );
and \U$39130 ( \39376 , \39374 , \39375 );
not \U$39131 ( \39377 , \39374 );
not \U$39132 ( \39378 , \39375 );
and \U$39133 ( \39379 , \39377 , \39378 );
nor \U$39134 ( \39380 , \39376 , \39379 );
buf \U$39135 ( \39381 , \39380 );
endmodule

