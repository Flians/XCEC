//
// Conformal-LEC Version 20.10-d215 (04-Sep-2020)
//
module top(RIae9a408_1,RIae9a480_2,RIae9a4f8_3,RIae9a570_4,RIae9a5e8_5,RIae9a660_6,RIae9a6d8_7,RIae9a750_8,RIae9a7c8_9,
        RIae9a840_10,RIae9a8b8_11,RIae9a930_12,RIae9a9a8_13,RIae9aa20_14,RIae9aa98_15,RIae9ab10_16,RIae9ab88_17,RIae9ac00_18,RIae9ac78_19,
        RIae9acf0_20,RIae9ad68_21,RIae9ade0_22,RIae9ae58_23,RIae9aed0_24,RIae9af48_25,RIae9afc0_26,RIae9b038_27,RIae9b0b0_28,RIae9b128_29,
        RIae9b1a0_30,RIae9b218_31,RIae9b290_32,RIae9b308_33,RIae9b380_34,RIae9b3f8_35,RIae9b470_36,RIae9b4e8_37,RIae9b560_38,RIae9b5d8_39,
        RIae9b650_40,RIae9b6c8_41,RIae9b740_42,RIae9b7b8_43,RIae9b830_44,RIae9b8a8_45,RIae9b920_46,RIae9b998_47,RIae9ba10_48,RIae9ba88_49,
        RIae9bb00_50,RIae9bb78_51,RIae9bbf0_52,RIae9bc68_53,RIae9bce0_54,RIae9bd58_55,RIae9bdd0_56,RIae9be48_57,RIae9bec0_58,RIae9bf38_59,
        RIae9bfb0_60,RIae9c028_61,RIae9c0a0_62,RIae9c118_63,RIae9c190_64,RIae9c208_65,RIae9c280_66,RIae9c2f8_67,RIae9c370_68,RIae9c3e8_69,
        RIae9c460_70,RIae9c4d8_71,RIae9c550_72,RIae9c5c8_73,RIae9c640_74,RIae9c6b8_75,RIae9c730_76,RIae9c7a8_77,RIae9c820_78,RIae9c898_79,
        RIae9c910_80,RIae9c988_81,RIae9ca00_82,RIae9ca78_83,RIae9caf0_84,RIae9cb68_85,RIae9cbe0_86,RIae9cc58_87,RIae9ccd0_88,RIae9cd48_89,
        RIae9cdc0_90,RIae9ce38_91,RIae9ceb0_92,RIae9cf28_93,RIae9cfa0_94,RIae9d018_95,RIae9d090_96,RIae9d108_97,RIae9d180_98,RIae9d1f8_99,
        RIae9d270_100,RIae9d2e8_101,RIae9d360_102,RIae9d3d8_103,RIae9d450_104,RIae9d4c8_105,RIae9d540_106,RIae9d5b8_107,RIae9d630_108,RIae9d6a8_109,
        RIae9d720_110,RIae9d798_111,RIae9d810_112,RIae9d888_113,RIae9d900_114,RIae9d978_115,RIae9d9f0_116,RIae9da68_117,RIae9dae0_118,RIae9db58_119,
        RIae9dbd0_120,RIae9dc48_121,RIae9dcc0_122,RIae9dd38_123,RIae9ddb0_124,RIae9de28_125,RIae9dea0_126,RIae9df18_127,RIae9df90_128,RIae9e008_129,
        RIae9e080_130,RIae9e0f8_131,RIae9e170_132,RIae9e1e8_133,RIae9e260_134,RIae9e2d8_135,RIae9e350_136,RIae9e3c8_137,RIae9e440_138,RIae9e4b8_139,
        RIae9e530_140,RIae9e5a8_141,RIae9e620_142,RIae9e698_143,RIae9e710_144,RIae9e788_145,RIae9e800_146,RIae9e878_147,RIae9e8f0_148,RIae9e968_149,
        RIae9e9e0_150,RIae9ea58_151,RIae9ead0_152,RIae9eb48_153,RIae9ebc0_154,RIae9ec38_155,RIae9ecb0_156,RIae9ed28_157,RIae9eda0_158,RIae9ee18_159,
        RIae9ee90_160,RIae9ef08_161,RIae9ef80_162,RIae9eff8_163,RIae9f070_164,RIae9f0e8_165,RIae9f160_166,RIae9f1d8_167,RIae9f250_168,RIae9f2c8_169,
        RIae9f340_170,RIae9f3b8_171,RIae9f430_172,RIae9f4a8_173,RIae9f520_174,RIae9f598_175,RIae9f610_176,RIae9f688_177,RIae9f700_178,RIae9f778_179,
        RIae9f7f0_180,RIae9f868_181,RIae9f8e0_182,RIae9f958_183,RIae9f9d0_184,RIae9fa48_185,RIae9fac0_186,RIae9fb38_187,RIae9fbb0_188,RIae9fc28_189,
        RIae9fca0_190,RIae9fd18_191,RIae9fd90_192,RIae9fe08_193,RIae9fe80_194,RIae9fef8_195,RIae9ff70_196,RIae9ffe8_197,RIaea0060_198,RIaea00d8_199,
        RIaea0150_200,RIaea01c8_201,RIaea0240_202,RIaea02b8_203,RIaea0330_204,RIaea03a8_205,RIaea0420_206,RIaea0498_207,RIaea0510_208,RIaea0588_209,
        RIaea0600_210,RIaea0678_211,RIaea06f0_212,RIaea0768_213,RIaea07e0_214,RIaea0858_215,RIaea08d0_216,RIaea0948_217,RIaea09c0_218,RIaea0a38_219,
        RIaea0ab0_220,RIaea0b28_221,RIaea0ba0_222,RIaea0c18_223,RIaea0c90_224,RIaea0d08_225,RIaea0d80_226,RIaea0df8_227,RIaea0e70_228,RIaea0ee8_229,
        RIaea0f60_230,RIaea0fd8_231,RIaea1050_232,RIaea10c8_233,RIaea1140_234,RIaea11b8_235,RIaea1230_236,RIaea12a8_237,RIaea1320_238,RIaea1398_239,
        RIaea1410_240,RIaea1488_241,RIaea1500_242,RIaea1578_243,RIaea15f0_244,RIaea1668_245,RIaea16e0_246,RIaea1758_247,RIaea17d0_248,RIaea1848_249,
        RIaea18c0_250,RIaea1938_251,RIaea19b0_252,RIaea1a28_253,RIaea1aa0_254,RIaea1b18_255,RIaea1b90_256,RIaea1c08_257,RIaea1c80_258,RIaea1cf8_259,
        RIaea1d70_260,RIaea1de8_261,RIaea1e60_262,RIaea1ed8_263,RIaea1f50_264,RIaea1fc8_265,RIaea2040_266,RIaea20b8_267,RIaea2130_268,RIaea21a8_269,
        RIaea2220_270,RIaea2298_271,RIaea2310_272,RIaea2388_273,RIaea2400_274,RIaea2478_275,RIaea24f0_276,RIaea2568_277,RIaea25e0_278,RIaea2658_279,
        RIaea26d0_280,RIaea2748_281,RIaea27c0_282,RIaea2838_283,RIaea28b0_284,RIaea2928_285,RIaea29a0_286,RIaea2a18_287,RIaea2a90_288,RIaea2b08_289,
        RIaea2b80_290,RIaea2bf8_291,RIaea2c70_292,RIaea2ce8_293,RIaea2d60_294,RIaea2dd8_295,RIaea2e50_296,RIaea2ec8_297,RIaea2f40_298,RIaea2fb8_299,
        RIaea3030_300,RIaea30a8_301,RIaea3120_302,RIaea3198_303,RIaea3210_304,RIaea3288_305,RIaea3300_306,RIaea3378_307,RIaea33f0_308,RIaea3468_309,
        RIaea34e0_310,RIaea3558_311,RIaea35d0_312,RIaea3648_313,RIaea36c0_314,RIaea3738_315,RIaea37b0_316,RIaea3828_317,RIaea38a0_318,RIaea3918_319,
        RIaea3990_320,RIaea3a08_321,RIaea3a80_322,RIaea3af8_323,RIaea3b70_324,RIaea3be8_325,RIaea3c60_326,RIaea3cd8_327,RIaea3d50_328,RIaea3dc8_329,
        RIaea3e40_330,RIaea3eb8_331,RIaea3f30_332,RIaea3fa8_333,RIaea4020_334,RIaea4098_335,RIaea4110_336,RIaea4188_337,RIaea4200_338,RIaea4278_339,
        RIaea42f0_340,RIaea4368_341,RIaea43e0_342,RIaea4458_343,RIaea44d0_344,RIaea4548_345,RIaea45c0_346,RIaea4638_347,RIaea46b0_348,RIaea4728_349,
        RIaea47a0_350,RIaea4818_351,RIaea4890_352,RIaea4908_353,RIaea4980_354,RIaea49f8_355,RIaea4a70_356,RIaea4ae8_357,RIaea4b60_358,RIaea4bd8_359,
        RIaea4c50_360,RIaea4cc8_361,RIaea4d40_362,RIaea4db8_363,RIaea4e30_364,RIaea4ea8_365,RIaea4f20_366,RIaea4f98_367,RIaea5010_368,RIaea5088_369,
        RIaea5100_370,RIaea5178_371,RIaea51f0_372,RIaea5268_373,RIaea52e0_374,RIaea5358_375,RIaea53d0_376,RIaea5448_377,RIaea54c0_378,RIaea5538_379,
        RIaea55b0_380,RIaea5628_381,RIaea56a0_382,RIaea5718_383,RIaea5790_384,RIaea5808_385,RIaea5880_386,RIaea58f8_387,RIaea5970_388,RIaea59e8_389,
        RIaea5a60_390,RIaea5ad8_391,RIaea5b50_392,RIaea5bc8_393,RIaea5c40_394,RIaea5cb8_395,RIaea5d30_396,RIaea5da8_397,RIaea5e20_398,RIaea5e98_399,
        RIaea5f10_400,RIaea5f88_401,RIaea6000_402,RIaea6078_403,RIaea60f0_404,RIaea6168_405,RIaea61e0_406,RIaea6258_407,RIaea62d0_408,RIaea6348_409,
        RIaea63c0_410,RIaea6438_411,RIaea64b0_412,RIaea6528_413,RIaea65a0_414,RIaea6618_415,RIaea6690_416,RIaea6708_417,RIaea6780_418,RIaea67f8_419,
        RIaea6870_420,RIaea68e8_421,RIaea6960_422,RIaea69d8_423,RIaea6a50_424,RIaea6ac8_425,RIaea6b40_426,RIaea6bb8_427,RIaea6c30_428,RIaea6ca8_429,
        RIaea6d20_430,RIaea6d98_431,RIaea6e10_432,RIaea6e88_433,RIaea6f00_434,RIaea6f78_435,RIaea6ff0_436,RIaea7068_437,RIaea70e0_438,RIaea7158_439,
        RIaea71d0_440,RIaea7248_441,RIaea72c0_442,RIaea7338_443,RIaea73b0_444,RIaea7428_445,RIaea74a0_446,RIaea7518_447,RIaea7590_448,RIaea7608_449,
        RIaea7680_450,RIaea76f8_451,RIaea7770_452,RIaea77e8_453,RIaea7860_454,RIaea78d8_455,RIaea7950_456,RIaea79c8_457,RIaea7a40_458,RIaea7ab8_459,
        RIaea7b30_460,RIaea7ba8_461,RIaea7c20_462,RIaea7c98_463,RIaea7d10_464,RIaea7d88_465,RIaea7e00_466,RIaea7e78_467,RIaea7ef0_468,RIaea7f68_469,
        RIaea7fe0_470,RIaea8058_471,RIaea80d0_472,RIaea8148_473,RIaea81c0_474,RIaea8238_475,RIaea82b0_476,RIaea8328_477,RIaea83a0_478,RIaea8418_479,
        RIaea8490_480,RIaea8508_481,RIaea8580_482,RIaea85f8_483,RIaea8670_484,RIaea86e8_485,RIaea8760_486,RIaea87d8_487,RIaea8850_488,RIaea88c8_489,
        RIaea8940_490,RIaea89b8_491,RIaea8a30_492,RIaea8aa8_493,RIaea8b20_494,RIaea8b98_495,RIaea8c10_496,RIaea8c88_497,RIaea8d00_498,RIaea8d78_499,
        RIaea8df0_500,RIaea8e68_501,RIaea8ee0_502,RIaea8f58_503,RIaea8fd0_504,RIaea9048_505,RIaea90c0_506,RIaea9138_507,RIaea91b0_508,RIaea9228_509,
        RIaea92a0_510,RIaea9318_511,RIaea9390_512,RIaea9408_513,RIaea9480_514,RIaea94f8_515,RIaea9570_516,RIaea95e8_517,RIaea9660_518,RIaea96d8_519,
        RIaea9750_520,RIaea97c8_521,RIaea9840_522,RIaea98b8_523,RIaea9930_524,RIaea99a8_525,RIaea9a20_526,RIaea9a98_527,RIaea9b10_528,RIaea9b88_529,
        RIaea9c00_530,RIaea9c78_531,RIaea9cf0_532,RIaea9d68_533,RIaea9de0_534,RIaea9e58_535,RIaea9ed0_536,RIaea9f48_537,RIaea9fc0_538,RIaeaa038_539,
        RIaeaa0b0_540,RIaeaa128_541,RIaeaa1a0_542,RIaeaa218_543,RIaeaa290_544,RIaeaa308_545,RIaeaa380_546,RIaeaa3f8_547,RIaeaa470_548,RIaeaa4e8_549,
        RIaeaa560_550,RIaeaa5d8_551,RIaeaa650_552,RIaeaa6c8_553,RIaeaa740_554,RIaeaa7b8_555,RIaeaa830_556,RIaeaa8a8_557,RIaeaa920_558,RIaeaa998_559,
        RIaeaaa10_560,RIaeaaa88_561,RIaeaab00_562,RIaeaab78_563,RIaeaabf0_564,RIaeaac68_565,RIaeaace0_566,RIaeaad58_567,RIaeaadd0_568,RIaeaae48_569,
        RIaeaaec0_570,RIaeaaf38_571,RIaeaafb0_572,RIaeab028_573,RIaeab0a0_574,RIaeab118_575,RIaeab190_576,RIaeab208_577,RIaeab280_578,RIaeab2f8_579,
        RIaeab370_580,RIaeab3e8_581,RIaeab460_582,RIaeab4d8_583,RIaeab550_584,RIaeab5c8_585,RIaeab640_586,RIaeab6b8_587,RIaeab730_588,RIaeab7a8_589,
        RIaeab820_590,RIaeab898_591,RIaeab910_592,RIaeab988_593,RIaeaba00_594,RIaeaba78_595,RIaeabaf0_596,RIaeabb68_597,RIaeabbe0_598,RIaeabc58_599,
        RIaeabcd0_600,RIaeabd48_601,RIaeabdc0_602,RIaeabe38_603,RIaeabeb0_604,RIaeabf28_605,RIaeabfa0_606,RIaeac018_607,RIaeac090_608,RIaeac108_609,
        RIaeac180_610,RIaeac1f8_611,RIaeac270_612,RIaeac2e8_613,RIaeac360_614,RIaeac3d8_615,RIaeac450_616,RIaeac4c8_617,RIaeac540_618,RIaeac5b8_619,
        RIaeac630_620,RIaeac6a8_621,RIaeac720_622,RIaeac798_623,RIaeac810_624,RIaeac888_625,RIaeac900_626,RIaeac978_627,RIaeac9f0_628,RIaeaca68_629,
        RIaeacae0_630,RIaeacb58_631,RIaeacbd0_632,RIaeacc48_633,RIaeaccc0_634,RIaeacd38_635,RIaeacdb0_636,RIaeace28_637,RIaeacea0_638,RIaeacf18_639,
        RIaeacf90_640,RIaead008_641,RIaead080_642,RIaead0f8_643,RIaead170_644,RIaead1e8_645,RIaead260_646,RIaead2d8_647,RIaead350_648,RIaead3c8_649,
        RIaead440_650,RIaead4b8_651,RIaead530_652,RIaead5a8_653,RIaead620_654,RIaead698_655,RIaead710_656,RIaead788_657,RIaead800_658,RIaead878_659,
        RIaead8f0_660,RIaead968_661,RIaead9e0_662,RIaeada58_663,RIaeadad0_664,RIaeadb48_665,RIaeadbc0_666,RIaeadc38_667,RIaeadcb0_668,RIaeadd28_669,
        RIaeadda0_670,RIaeade18_671,RIaeade90_672,RIaeadf08_673,RIaeadf80_674,RIaeadff8_675,RIaeae070_676,RIaeae0e8_677,RIaeae160_678,RIaeae1d8_679,
        RIaeae250_680,RIaeae2c8_681,RIaeae340_682,RIaeae3b8_683,RIaeae430_684,RIaeae4a8_685,RIaeae520_686,RIaeae598_687,RIaeae610_688,RIaeae688_689,
        RIaeae700_690,RIaeae778_691,RIaeae7f0_692,RIaeae868_693,RIaeae8e0_694,RIaeae958_695,RIaeae9d0_696,RIaeaea48_697,RIaeaeac0_698,RIaeaeb38_699,
        RIaeaebb0_700,RIaeaec28_701,RIaeaeca0_702,RIaeaed18_703,RIaeaed90_704,RIaeaee08_705,RIaeaee80_706,RIaeaeef8_707,RIaeaef70_708,RIaeaefe8_709,
        RIaeaf060_710,RIaeaf0d8_711,RIaeaf150_712,RIaeaf1c8_713,RIaeaf240_714,RIaeaf2b8_715,RIaeaf330_716,RIaeaf3a8_717,RIaeaf420_718,RIaeaf498_719,
        RIaeaf510_720,RIaeaf588_721,RIaeaf600_722,RIaeaf678_723,RIaeaf6f0_724,RIaeaf768_725,RIaeaf7e0_726,RIaeaf858_727,RIaeaf8d0_728,RIaeaf948_729,
        RIaeaf9c0_730,RIaeafa38_731,RIaeafab0_732,RIaeafb28_733,RIaeafba0_734,RIaeafc18_735,RIaeafc90_736,RIaeafd08_737,RIaeafd80_738,RIaeafdf8_739,
        RIaeafe70_740,RIaeafee8_741,RIaeaff60_742,RIaeaffd8_743,RIaeb0050_744,RIaeb00c8_745,RIaeb0140_746,RIaeb01b8_747,RIaeb0230_748,RIaeb02a8_749,
        RIaeb0320_750,RIaeb0398_751,RIaeb0410_752,RIaeb0488_753,RIaeb0500_754,RIaeb0578_755,RIaeb05f0_756,RIaeb0668_757,RIaeb06e0_758,RIaeb0758_759,
        RIaeb07d0_760,RIaeb0848_761,RIaeb08c0_762,RIaeb0938_763,RIaeb09b0_764,RIaeb0a28_765,RIaeb0aa0_766,RIaeb0b18_767,RIaeb0b90_768,RIaeb0c08_769,
        RIaeb0c80_770,RIaeb0cf8_771,RIaeb0d70_772,RIaeb0de8_773,RIaeb0e60_774,RIaeb0ed8_775,RIaeb0f50_776,RIaeb0fc8_777,RIaeb1040_778,RIaeb10b8_779,
        RIaeb1130_780,RIaeb11a8_781,RIaeb1220_782,RIaeb1298_783,RIaeb1310_784,RIaeb1388_785,RIaeb1400_786,RIaeb1478_787,RIaeb14f0_788,RIaeb1568_789,
        RIaeb15e0_790,RIaeb1658_791,RIaeb16d0_792,RIaeb1748_793,RIaeb17c0_794,RIaeb1838_795,RIaeb18b0_796,RIaeb1928_797,RIaeb19a0_798,RIaeb1a18_799,
        RIaeb1a90_800,RIaeb1b08_801,RIaeb1b80_802,RIaeb1bf8_803,RIaeb1c70_804,RIaeb1ce8_805,RIaeb1d60_806,RIaeb1dd8_807,RIaeb1e50_808,RIaeb1ec8_809,
        RIaeb1f40_810,RIaeb1fb8_811,RIaeb2030_812,RIaeb20a8_813,RIaeb2120_814,RIaeb2198_815,RIaeb2210_816,RIaeb2288_817,RIaeb2300_818,RIaeb2378_819,
        RIaeb23f0_820,RIaeb2468_821,RIaeb24e0_822,RIaeb2558_823,RIaeb25d0_824,RIaeb2648_825,RIaeb26c0_826,RIaeb2738_827,RIaeb27b0_828,RIaeb2828_829,
        RIaeb28a0_830,RIaeb2918_831,RIaeb2990_832,RIaeb2a08_833,RIaeb2a80_834,RIaeb2af8_835,RIaeb2b70_836,RIaeb2be8_837,RIaeb2c60_838,RIaeb2cd8_839,
        RIaeb2d50_840,RIaeb2dc8_841,RIaeb2e40_842,RIaeb2eb8_843,RIaeb2f30_844,RIaeb2fa8_845,RIaeb3020_846,RIaeb3098_847,RIaeb3110_848,RIaeb3188_849,
        RIaeb3200_850,RIaeb3278_851,RIaeb32f0_852,RIaeb3368_853,RIaeb33e0_854,RIaeb3458_855,RIaeb34d0_856,RIaeb3548_857,RIaeb35c0_858,RIaeb3638_859,
        RIaeb36b0_860,RIaeb3728_861,RIaeb37a0_862,RIaeb3818_863,RIaeb3890_864,RIaeb3908_865,RIaeb3980_866,RIaeb39f8_867,RIaeb3a70_868,RIaeb3ae8_869,
        RIaeb3b60_870,RIaeb3bd8_871,RIaeb3c50_872,RIaeb3cc8_873,RIaeb3d40_874,RIaeb3db8_875,RIaeb3e30_876,RIaeb3ea8_877,RIaeb3f20_878,RIaeb3f98_879,
        RIaeb4010_880,RIaeb4088_881,RIaeb4100_882,RIaeb4178_883,RIaeb41f0_884,RIaeb4268_885,RIaeb42e0_886,RIaeb4358_887,RIaeb43d0_888,RIaeb4448_889,
        RIaeb44c0_890,RIaeb4538_891,RIaeb45b0_892,RIaeb4628_893,RIaeb46a0_894,RIaeb4718_895,RIaeb4790_896,RIaeb4808_897,RIaeb4880_898,RIaeb48f8_899,
        RIaeb4970_900,RIaeb49e8_901,RIaeb4a60_902,RIaeb4ad8_903,RIaeb4b50_904,RIaeb4bc8_905,RIaeb4c40_906,RIaeb4cb8_907,RIaeb4d30_908,RIaeb4da8_909,
        RIaeb4e20_910,RIaeb4e98_911,RIaeb4f10_912,RIaeb4f88_913,RIaeb5000_914,RIaeb5078_915,RIaeb50f0_916,RIaeb5168_917,RIaeb51e0_918,RIaeb5258_919,
        RIaeb52d0_920,RIaeb5348_921,RIaeb53c0_922,RIaeb5438_923,RIaeb54b0_924,RIaeb5528_925,RIaeb55a0_926,RIaeb5618_927,RIaeb5690_928,RIaeb5708_929,
        RIaeb5780_930,RIaeb57f8_931,RIaeb5870_932,RIaeb58e8_933,RIaeb5960_934,RIaeb59d8_935,RIaeb5a50_936,RIaeb5ac8_937,RIaeb5b40_938,RIaeb5bb8_939,
        RIaeb5c30_940,RIaeb5ca8_941,RIaeb5d20_942,RIaeb5d98_943,RIaeb5e10_944,RIaeb5e88_945,RIaeb5f00_946,RIaeb5f78_947,RIaeb5ff0_948,RIaeb6068_949,
        RIaeb60e0_950,RIaeb6158_951,RIaeb61d0_952,RIaeb6248_953,RIaeb62c0_954,RIaeb6338_955,RIaeb63b0_956,RIaeb6428_957,RIaeb64a0_958,RIaeb6518_959,
        RIaeb6590_960,RIaeb6608_961,RIaeb6680_962,RIaeb66f8_963,RIaeb6770_964,RIaeb67e8_965,RIaeb6860_966,RIaeb68d8_967,RIaeb6950_968,RIaeb69c8_969,
        RIaeb6a40_970,RIaeb6ab8_971,RIaeb6b30_972,RIaeb6ba8_973,RIaeb6c20_974,RIaeb6c98_975,RIaeb6d10_976,RIaeb6d88_977,RIaeb6e00_978,RIaeb6e78_979,
        RIaeb6ef0_980,RIaeb6f68_981,RIaeb6fe0_982,RIaeb7058_983,RIaeb70d0_984,RIaeb7148_985,RIaeb71c0_986,RIaeb7238_987,RIaeb72b0_988,RIaeb7328_989,
        RIaeb73a0_990,RIaeb7418_991,RIaeb7490_992,RIaeb7508_993,RIaeb7580_994,RIaeb75f8_995,RIaeb7670_996,RIaeb76e8_997,RIaeb7760_998,RIaeb77d8_999,
        RIaeb7850_1000,RIaeb78c8_1001,RIaeb7940_1002,RIaeb79b8_1003,RIaeb7a30_1004,RIaeb7aa8_1005,RIaeb7b20_1006,RIaeb7b98_1007,RIaeb7c10_1008,RIaeb7c88_1009,
        RIaeb7d00_1010,RIaeb7d78_1011,RIaeb7df0_1012,RIaeb7e68_1013,RIaeb7ee0_1014,RIaeb7f58_1015,RIaeb7fd0_1016,RIaeb8048_1017,RIaeb80c0_1018,RIaeb8138_1019,
        RIaeb81b0_1020,RIaeb8228_1021,RIaeb82a0_1022,RIaeb8318_1023,RIaeb8390_1024,RIaeb8408_1025,RIaeb8480_1026,RIaeb84f8_1027,RIaeb8570_1028,RIaeb85e8_1029,
        RIaeb8660_1030,RIaeb86d8_1031,RIaeb8750_1032,RIaeb87c8_1033,RIaeb8840_1034,RIaeb88b8_1035,RIaeb8930_1036,RIaeb89a8_1037,RIaeb8a20_1038,RIaeb8a98_1039,
        RIaeb8b10_1040,RIaeb8b88_1041,RIaeb8c00_1042,RIaeb8c78_1043,RIaeb8cf0_1044,RIaeb8d68_1045,RIaeb8de0_1046,RIaeb8e58_1047,RIaeb8ed0_1048,RIaeb8f48_1049,
        RIaeb8fc0_1050,RIaeb9038_1051,RIaeb90b0_1052,RIaeb9128_1053,RIaeb91a0_1054,RIaeb9218_1055,RIaeb9290_1056,RIaeb9308_1057,RIaeb9380_1058,RIaeb93f8_1059,
        RIaeb9470_1060,RIaeb94e8_1061,RIaeb9560_1062,RIaeb95d8_1063,RIaeb9650_1064,RIaeb96c8_1065,RIaeb9740_1066,RIaeb97b8_1067,RIaeb9830_1068,RIaeb98a8_1069,
        RIaeb9920_1070,RIaeb9998_1071,RIaeb9a10_1072,RIaeb9a88_1073,RIaeb9b00_1074,RIaeb9b78_1075,RIaeb9bf0_1076,RIaeb9c68_1077,RIaeb9ce0_1078,RIaeb9d58_1079,
        RIaeb9dd0_1080,RIaeb9e48_1081,RIaeb9ec0_1082,RIaeb9f38_1083,RIaeb9fb0_1084,RIaeba028_1085,RIaeba0a0_1086,RIaeba118_1087,RIaeba190_1088,RIaeba208_1089,
        RIaeba280_1090,RIaeba2f8_1091,RIaeba370_1092,RIaeba3e8_1093,RIaeba460_1094,RIaeba4d8_1095,RIaeba550_1096,RIaeba5c8_1097,RIaeba640_1098,RIaeba6b8_1099,
        RIaeba730_1100,RIaeba7a8_1101,RIaeba820_1102,RIaeba898_1103,RIaeba910_1104,RIaeba988_1105,RIaebaa00_1106,RIaebaa78_1107,RIaebaaf0_1108,RIaebab68_1109,
        RIaebabe0_1110,RIaebac58_1111,RIaebacd0_1112,RIaebad48_1113,RIaebadc0_1114,RIaebae38_1115,RIaebaeb0_1116,RIaebaf28_1117,RIaebafa0_1118,RIaebb018_1119,
        RIaebb090_1120,RIaebb108_1121,RIaebb180_1122,RIaebb1f8_1123,RIaebb270_1124,RIaebb2e8_1125,RIaebb360_1126,RIaebb3d8_1127,RIaebb450_1128,RIaebb4c8_1129,
        RIaebb540_1130,RIaebb5b8_1131,RIaebb630_1132,RIaebb6a8_1133,RIaebb720_1134,RIaebb798_1135,RIaebb810_1136,RIaebb888_1137,RIaebb900_1138,RIaebb978_1139,
        RIaebb9f0_1140,RIaebba68_1141,RIaebbae0_1142,RIaebbb58_1143,RIaebbbd0_1144,RIaebbc48_1145,RIaebbcc0_1146,RIaebbd38_1147,RIaebbdb0_1148,RIaebbe28_1149,
        RIaebbea0_1150,RIaebbf18_1151,RIaebbf90_1152,RIaebc008_1153,RIaebc080_1154,RIaebc0f8_1155,RIaebc170_1156,RIaebc1e8_1157,RIaebc260_1158,RIaebc2d8_1159,
        RIaebc350_1160,RIaebc3c8_1161,RIaebc440_1162,RIaebc4b8_1163,RIaebc530_1164,RIaebc5a8_1165,RIaebc620_1166,RIaebc698_1167,RIaebc710_1168,RIaebc788_1169,
        RIaebc800_1170,RIaebc878_1171,RIaebc8f0_1172,RIaebc968_1173,RIaebc9e0_1174,RIaebca58_1175,RIaebcad0_1176,RIaebcb48_1177,RIaebcbc0_1178,RIaebcc38_1179,
        RIaebccb0_1180,RIaebcd28_1181,RIaebcda0_1182,RIaebce18_1183,RIaebce90_1184,RIaebcf08_1185,RIaebcf80_1186,RIaebcff8_1187,RIaebd070_1188,RIaebd0e8_1189,
        RIaebd160_1190,RIaebd1d8_1191,RIaebd250_1192,RIaebd2c8_1193,RIaebd340_1194,RIaebd3b8_1195,RIaebd430_1196,RIaebd4a8_1197,RIaebd520_1198,RIaebd598_1199,
        RIaebd610_1200,RIaebd688_1201,RIaebd700_1202,RIaebd778_1203,RIaebd7f0_1204,RIaebd868_1205,RIaebd8e0_1206,RIaebd958_1207,RIaebd9d0_1208,RIaebda48_1209,
        RIaebdac0_1210,RIaebdb38_1211,RIaebdbb0_1212,RIaebdc28_1213,RIaebdca0_1214,RIaebdd18_1215,RIaebdd90_1216,RIaebde08_1217,RIaebde80_1218,RIaebdef8_1219,
        RIaebdf70_1220,RIaebdfe8_1221,RIaebe060_1222,RIaebe0d8_1223,RIaebe150_1224,RIaebe1c8_1225,RIaebe240_1226,RIaebe2b8_1227,RIaebe330_1228,RIaebe3a8_1229,
        RIaebe420_1230,RIaebe498_1231,RIaebe510_1232,RIaebe588_1233,RIaebe600_1234,RIaebe678_1235,RIaebe6f0_1236,RIaebe768_1237,RIaebe7e0_1238,RIaebe858_1239,
        RIaebe8d0_1240,RIaebe948_1241,RIaebe9c0_1242,RIaebea38_1243,RIaebeab0_1244,RIaebeb28_1245,RIaebeba0_1246,RIaebec18_1247,RIaebec90_1248,RIaebed08_1249,
        RIaebed80_1250,RIaebedf8_1251,RIaebee70_1252,RIaebeee8_1253,RIaebef60_1254,RIaebefd8_1255,RIaebf050_1256,RIaebf0c8_1257,RIaebf140_1258,RIaebf1b8_1259,
        RIaebf230_1260,RIaebf2a8_1261,RIaebf320_1262,RIaebf398_1263,RIaebf410_1264,RIaebf488_1265,RIaebf500_1266,RIaebf578_1267,RIaebf5f0_1268,RIaebf668_1269,
        RIaebf6e0_1270,RIaebf758_1271,RIaebf7d0_1272,RIaebf848_1273,RIaebf8c0_1274,RIaebf938_1275,RIaebf9b0_1276,RIaebfa28_1277,RIaebfaa0_1278,RIaebfb18_1279,
        RIaebfb90_1280,RIaebfc08_1281,RIaebfc80_1282,RIaebfcf8_1283,RIaebfd70_1284,RIaebfde8_1285,RIaebfe60_1286,RIaebfed8_1287,RIaebff50_1288,RIaebffc8_1289,
        RIaec0040_1290,RIaec00b8_1291,RIaec0130_1292,RIaec01a8_1293,RIaec0220_1294,RIaec0298_1295,RIaec0310_1296,RIaec0388_1297,RIaec0400_1298,RIaec0478_1299,
        RIaec04f0_1300,RIaec0568_1301,RIaec05e0_1302,RIaec0658_1303,RIaec06d0_1304,RIaec0748_1305,RIaec07c0_1306,RIaec0838_1307,RIaec08b0_1308,RIaec0928_1309,
        RIaec09a0_1310,RIaec0a18_1311,RIaec0a90_1312,RIaec0b08_1313,RIaec0b80_1314,RIaec0bf8_1315,RIaec0c70_1316,RIaec0ce8_1317,RIaec0d60_1318,RIaec0dd8_1319,
        RIaec0e50_1320,RIaec0ec8_1321,RIaec0f40_1322,RIaec0fb8_1323,RIaec1030_1324,RIaec10a8_1325,RIaec1120_1326,RIaec1198_1327,RIaec1210_1328,RIaec1288_1329,
        RIaec1300_1330,RIaec1378_1331,RIaec13f0_1332,RIaec1468_1333,RIaec14e0_1334,RIaec1558_1335,RIaec15d0_1336,RIaec1648_1337,RIaec16c0_1338,RIaec1738_1339,
        RIaec17b0_1340,RIaec1828_1341,RIaec18a0_1342,RIaec1918_1343,RIaec1990_1344,RIaec1a08_1345,RIaec1a80_1346,RIaec1af8_1347,RIaec1b70_1348,RIaec1be8_1349,
        RIaec1c60_1350,RIaec1cd8_1351,RIaec1d50_1352,RIaec1dc8_1353,RIaec1e40_1354,RIaec1eb8_1355,RIaec1f30_1356,RIaec1fa8_1357,RIaec2020_1358,RIaec2098_1359,
        RIaec2110_1360,RIaec2188_1361,RIaec2200_1362,RIaec2278_1363,RIaec22f0_1364,RIaec2368_1365,RIaec23e0_1366,RIaec2458_1367,RIaec24d0_1368,RIaec2548_1369,
        RIaec25c0_1370,RIaec2638_1371,RIaec26b0_1372,RIaec2728_1373,RIaec27a0_1374,RIaec2818_1375,RIaec2890_1376,RIaec2908_1377,RIaec2980_1378,RIaec29f8_1379,
        RIaec2a70_1380,RIaec2ae8_1381,RIaec2b60_1382,RIaec2bd8_1383,RIaec2c50_1384,RIaec2cc8_1385,RIaec2d40_1386,RIaec2db8_1387,RIaec2e30_1388,RIaec2ea8_1389,
        RIaec2f20_1390,RIaec2f98_1391,RIaec3010_1392,RIaec3088_1393,RIaec3100_1394,RIaec3178_1395,RIaec31f0_1396,RIaec3268_1397,RIaec32e0_1398,RIaec3358_1399,
        RIaec33d0_1400,RIaec3448_1401,RIaec34c0_1402,RIaec3538_1403,RIaec35b0_1404,RIaec3628_1405,RIaec36a0_1406,RIaec3718_1407,RIaec3790_1408,RIaec3808_1409,
        RIaec3880_1410,RIaec38f8_1411,RIaec3970_1412,RIaec39e8_1413,RIaec3a60_1414,RIaec3ad8_1415,RIaec3b50_1416,RIaec3bc8_1417,RIaec3c40_1418,RIaec3cb8_1419,
        RIaec3d30_1420,RIaec3da8_1421,RIaec3e20_1422,RIaec3e98_1423,RIaec3f10_1424,RIaec3f88_1425,RIaec4000_1426,RIaec4078_1427,RIaec40f0_1428,RIaec4168_1429,
        RIaec41e0_1430,RIaec4258_1431,RIaec42d0_1432,RIaec4348_1433,RIaec43c0_1434,RIaec4438_1435,RIaec44b0_1436,RIaec4528_1437,RIaec45a0_1438,RIaec4618_1439,
        RIaec4690_1440,RIaec4708_1441,RIaec4780_1442,RIaec47f8_1443,RIaec4870_1444,RIaec48e8_1445,RIaec4960_1446,RIaec49d8_1447,RIaec4a50_1448,RIaec4ac8_1449,
        RIaec4b40_1450,RIaec4bb8_1451,RIaec4c30_1452,RIaec4ca8_1453,RIaec4d20_1454,RIaec4d98_1455,RIaec4e10_1456,RIaec4e88_1457,RIaec4f00_1458,RIaec4f78_1459,
        RIaec4ff0_1460,RIaec5068_1461,RIaec50e0_1462,RIaec5158_1463,RIaec51d0_1464,RIaec5248_1465,RIaec52c0_1466,RIaec5338_1467,RIaec53b0_1468,RIaec5428_1469,
        RIaec54a0_1470,RIaec5518_1471,RIaec5590_1472,RIaec5608_1473,RIaec5680_1474,RIaec56f8_1475,RIaec5770_1476,RIaec57e8_1477,RIaec5860_1478,RIaec58d8_1479,
        RIaec5950_1480,RIaec59c8_1481,RIaec5a40_1482,RIaec5ab8_1483,RIaec5b30_1484,RIaec5ba8_1485,RIaec5c20_1486,RIaec5c98_1487,RIaec5d10_1488,RIaec5d88_1489,
        RIaec5e00_1490,RIaec5e78_1491,RIaec5ef0_1492,RIaec5f68_1493,RIaec5fe0_1494,RIaec6058_1495,RIaec60d0_1496,RIaec6148_1497,RIaec61c0_1498,RIaec6238_1499,
        RIaec62b0_1500,RIaec6328_1501,RIaec63a0_1502,RIaec6418_1503,RIaec6490_1504,RIaec6508_1505,RIaec6580_1506,RIaec65f8_1507,RIaec6670_1508,RIaec66e8_1509,
        RIaec6760_1510,RIaec67d8_1511,RIaec6850_1512,RIaec68c8_1513,RIaec6940_1514,RIaec69b8_1515,RIaec6a30_1516,RIaec6aa8_1517,RIaec6b20_1518,RIaec6b98_1519,
        RIaec6c10_1520,RIaec6c88_1521,RIaec6d00_1522,RIaec6d78_1523,RIaec6df0_1524,RIaec6e68_1525,RIaec6ee0_1526,RIaec6f58_1527,RIaec6fd0_1528,RIaec7048_1529,
        RIaec70c0_1530,RIaec7138_1531,RIaec71b0_1532,RIaec7228_1533,RIaec72a0_1534,RIaec7318_1535,RIaec7390_1536,RIaec7408_1537,RIaec7480_1538,RIaec74f8_1539,
        RIaec7570_1540,RIaec75e8_1541,RIaec7660_1542,RIaec76d8_1543,RIaec7750_1544,RIaec77c8_1545,RIaec7840_1546,RIaec78b8_1547,RIaec7930_1548,RIaec79a8_1549,
        RIaec7a20_1550,RIaec7a98_1551,RIaec7b10_1552,RIaec7b88_1553,RIaec7c00_1554,RIaec7c78_1555,RIaec7cf0_1556,RIaec7d68_1557,RIaec7de0_1558,RIaec7e58_1559,
        RIaec7ed0_1560,RIaec7f48_1561,RIaec7fc0_1562,RIaec8038_1563,RIaec80b0_1564,RIaec8128_1565,RIaec81a0_1566,RIaec8218_1567,RIaec8290_1568,RIaec8308_1569,
        RIaec8380_1570,RIaec83f8_1571,RIaec8470_1572,RIaec84e8_1573,RIaec8560_1574,RIaec85d8_1575,RIaec8650_1576,RIaec86c8_1577,RIaec8740_1578,RIaec87b8_1579,
        RIaec8830_1580,RIaec88a8_1581,RIaec8920_1582,RIaec8998_1583,RIaec8a10_1584,RIaec8a88_1585,RIaec8b00_1586,RIaec8b78_1587,RIaec8bf0_1588,RIaec8c68_1589,
        RIaec8ce0_1590,RIaec8d58_1591,RIaec8dd0_1592,RIaec8e48_1593,RIaec8ec0_1594,RIaec8f38_1595,RIaec8fb0_1596,RIaec9028_1597,RIaec90a0_1598,RIaec9118_1599,
        RIaec9190_1600,RIaec9208_1601,RIaec9280_1602,RIaec92f8_1603,RIaec9370_1604,RIaec93e8_1605,RIaec9460_1606,RIaec94d8_1607,RIaec9550_1608,RIaec95c8_1609,
        RIaec9640_1610,RIaec96b8_1611,RIaec9730_1612,RIaec97a8_1613,RIaec9820_1614,RIaec9898_1615,RIaec9910_1616,RIaec9988_1617,RIaec9a00_1618,RIaec9a78_1619,
        RIaec9af0_1620,RIaec9b68_1621,RIaec9be0_1622,RIaec9c58_1623,RIaec9cd0_1624,RIaec9d48_1625,RIaec9dc0_1626,RIaec9e38_1627,RIaec9eb0_1628,RIaec9f28_1629,
        RIaec9fa0_1630,RIaeca018_1631,RIaeca090_1632,RIaeca108_1633,RIaeca180_1634,RIaeca1f8_1635,RIaeca270_1636,RIaeca2e8_1637,RIaeca360_1638,RIaeca3d8_1639,
        RIaeca450_1640,RIaeca4c8_1641,RIaeca540_1642,RIaeca5b8_1643,RIaeca630_1644,RIaeca6a8_1645,RIaeca720_1646,RIaeca798_1647,RIaeca810_1648,RIaeca888_1649,
        RIaeca900_1650,RIaeca978_1651,RIaeca9f0_1652,RIaecaa68_1653,RIaecaae0_1654,RIaecab58_1655,RIaecabd0_1656,RIaecac48_1657,RIaecacc0_1658,RIaecad38_1659,
        RIaecadb0_1660,RIaecae28_1661,RIaecaea0_1662,RIaecaf18_1663,RIaecaf90_1664,RIaecb008_1665,RIaecb080_1666,RIaecb0f8_1667,RIaecb170_1668,RIaecb1e8_1669,
        RIaecb260_1670,RIaecb2d8_1671,RIaecb350_1672,RIaecb3c8_1673,RIaecb440_1674,RIaecb4b8_1675,RIaecb530_1676,RIaecb5a8_1677,RIaecb620_1678,RIaecb698_1679,
        RIaecb710_1680,RIaecb788_1681,RIaecb800_1682,RIaecb878_1683,RIaecb8f0_1684,RIaecb968_1685,RIaecb9e0_1686,RIaecba58_1687,RIaecbad0_1688,RIaecbb48_1689,
        RIaecbbc0_1690,RIaecbc38_1691,RIaecbcb0_1692,RIaecbd28_1693,RIaecbda0_1694,RIaecbe18_1695,RIaecbe90_1696,RIaecbf08_1697,RIaecbf80_1698,RIaecbff8_1699,
        RIaecc070_1700,RIaecc0e8_1701,RIaecc160_1702,RIaecc1d8_1703,RIaecc250_1704,RIaecc2c8_1705,RIaecc340_1706,RIaecc3b8_1707,RIaecc430_1708,RIaecc4a8_1709,
        RIaecc520_1710,RIaecc598_1711,RIaecc610_1712,RIaecc688_1713,RIaecc700_1714,RIaecc778_1715,RIaecc7f0_1716,RIaecc868_1717,RIaecc8e0_1718,RIaecc958_1719,
        RIaecc9d0_1720,RIaecca48_1721,RIaeccac0_1722,RIaeccb38_1723,RIaeccbb0_1724,RIaeccc28_1725,RIaeccca0_1726,RIaeccd18_1727,RIaeccd90_1728,RIaecce08_1729,
        RIaecce80_1730,RIaeccef8_1731,RIaeccf70_1732,RIaeccfe8_1733,RIaecd060_1734,RIaecd0d8_1735,RIaecd150_1736,RIaecd1c8_1737,RIaecd240_1738,RIaecd2b8_1739,
        RIaecd330_1740,RIaecd3a8_1741,RIaecd420_1742,RIaecd498_1743,RIaecd510_1744,RIaecd588_1745,RIaecd600_1746,RIaecd678_1747,RIaecd6f0_1748,RIaecd768_1749,
        RIaecd7e0_1750,RIaecd858_1751,RIaecd8d0_1752,RIaecd948_1753,RIaecd9c0_1754,RIaecda38_1755,RIaecdab0_1756,RIaecdb28_1757,RIaecdba0_1758,RIaecdc18_1759,
        RIaecdc90_1760,RIaecdd08_1761,RIaecdd80_1762,RIaecddf8_1763,RIaecde70_1764,RIaecdee8_1765,RIaecdf60_1766,RIaecdfd8_1767,RIaece050_1768,RIaece0c8_1769,
        RIaece140_1770,RIaece1b8_1771,RIaece230_1772,RIaece2a8_1773,RIaece320_1774,RIaece398_1775,RIaece410_1776,RIaece488_1777,RIaece500_1778,RIaece578_1779,
        RIaece5f0_1780,RIaece668_1781,RIaece6e0_1782,RIaece758_1783,RIaece7d0_1784,RIaece848_1785,RIaece8c0_1786,RIaece938_1787,RIaece9b0_1788,RIaecea28_1789,
        RIaeceaa0_1790,RIaeceb18_1791,RIaeceb90_1792,RIaecec08_1793,RIaecec80_1794,RIaececf8_1795,RIaeced70_1796,RIaecede8_1797,RIaecee60_1798,RIaeceed8_1799,
        RIaecef50_1800,RIaecefc8_1801,RIaecf040_1802,RIaecf0b8_1803,RIaecf130_1804,RIaecf1a8_1805,RIaecf220_1806,RIaecf298_1807,RIaecf310_1808,RIaecf388_1809,
        RIaecf400_1810,RIaecf478_1811,RIaecf4f0_1812,RIaecf568_1813,RIaecf5e0_1814,RIaecf658_1815,RIaecf6d0_1816,RIaecf748_1817,RIaecf7c0_1818,RIaecf838_1819,
        RIaecf8b0_1820,RIaecf928_1821,RIaecf9a0_1822,RIaecfa18_1823,RIaecfa90_1824,RIaecfb08_1825,RIaecfb80_1826,RIaecfbf8_1827,RIaecfc70_1828,RIaecfce8_1829,
        RIaecfd60_1830,RIaecfdd8_1831,RIaecfe50_1832,RIaecfec8_1833,RIaecff40_1834,RIaecffb8_1835,RIaed0030_1836,RIaed00a8_1837,RIaed0120_1838,RIaed0198_1839,
        RIaed0210_1840,RIaed0288_1841,RIaed0300_1842,RIaed0378_1843,RIaed03f0_1844,RIaed0468_1845,RIaed04e0_1846,RIaed0558_1847,RIaed05d0_1848,RIaed0648_1849,
        RIaed06c0_1850,RIaed0738_1851,RIaed07b0_1852,RIaed0828_1853,RIaed08a0_1854,RIaed0918_1855,RIaed0990_1856,RIaed0a08_1857,RIaed0a80_1858,RIaed0af8_1859,
        RIaed0b70_1860,RIaed0be8_1861,RIaed0c60_1862,RIaed0cd8_1863,RIaed0d50_1864,RIaed0dc8_1865,RIaed0e40_1866,RIaed0eb8_1867,RIaed0f30_1868,RIaed0fa8_1869,
        RIaed1020_1870,RIaed1098_1871,RIaed1110_1872,RIaed1188_1873,RIaed1200_1874,RIaed1278_1875,RIaed12f0_1876,RIaed1368_1877,RIaed13e0_1878,RIaed1458_1879,
        RIaed14d0_1880,RIaed1548_1881,RIaed15c0_1882,RIaed1638_1883,RIaed16b0_1884,RIaed1728_1885,RIaed17a0_1886,RIaed1818_1887,RIaed1890_1888,RIaed1908_1889,
        RIaed1980_1890,RIaed19f8_1891,RIaed1a70_1892,RIaed1ae8_1893,RIaed1b60_1894,RIaed1bd8_1895,RIaed1c50_1896,RIaed1cc8_1897,RIaed1d40_1898,RIaed1db8_1899,
        RIaed1e30_1900,RIaed1ea8_1901,RIaed1f20_1902,RIaed1f98_1903,RIaed2010_1904,RIaed2088_1905,RIaed2100_1906,RIaed2178_1907,RIaed21f0_1908,RIaed2268_1909,
        RIaed22e0_1910,RIaed2358_1911,RIaed23d0_1912,RIaed2448_1913,RIaed24c0_1914,RIaed2538_1915,RIaed25b0_1916,RIaed2628_1917,RIaed26a0_1918,RIaed2718_1919,
        RIaed2790_1920,RIaed2808_1921,RIaed2880_1922,RIaed28f8_1923,RIaed2970_1924,RIaed29e8_1925,RIaed2a60_1926,RIaed2ad8_1927,RIaed2b50_1928,RIaed2bc8_1929,
        RIaed2c40_1930,RIaed2cb8_1931,RIaed2d30_1932,RIaed2da8_1933,RIaed2e20_1934,RIaed2e98_1935,RIaed2f10_1936,RIaed2f88_1937,RIaed3000_1938,RIaed3078_1939,
        RIaed30f0_1940,RIaed3168_1941,RIaed31e0_1942,RIaed3258_1943,RIaed32d0_1944,RIaed3348_1945,RIaed33c0_1946,RIaed3438_1947,RIaed34b0_1948,RIaed3528_1949,
        RIaed35a0_1950,RIaed3618_1951,RIaed3690_1952,RIaed3708_1953,RIaed3780_1954,RIaed37f8_1955,RIaed3870_1956,RIaed38e8_1957,RIaed3960_1958,RIaed39d8_1959,
        RIaed3a50_1960,RIaed3ac8_1961,RIaed3b40_1962,RIaed3bb8_1963,RIaed3c30_1964,RIaed3ca8_1965,RIaed3d20_1966,RIaed3d98_1967,RIaed3e10_1968,RIaed3e88_1969,
        RIaed3f00_1970,RIaed3f78_1971,RIaed3ff0_1972,RIaed4068_1973,RIaed40e0_1974,RIaed4158_1975,RIaed41d0_1976,RIaed4248_1977,RIaed42c0_1978,RIaed4338_1979,
        RIaed43b0_1980,RIaed4428_1981,RIaed44a0_1982,RIaed4518_1983,RIaed4590_1984,RIaed4608_1985,RIaed4680_1986,RIaed46f8_1987,RIaed4770_1988,RIaed47e8_1989,
        RIaed4860_1990,RIaed48d8_1991,RIaed4950_1992,RIaed49c8_1993,RIaed4a40_1994,RIaed4ab8_1995,RIaed4b30_1996,RIaed4ba8_1997,RIaed4c20_1998,RIaed4c98_1999,
        RIaed4d10_2000,RIaed4d88_2001,RIaed4e00_2002,RIaed4e78_2003,RIaed4ef0_2004,RIaed4f68_2005,RIaed4fe0_2006,RIaed5058_2007,RIaed50d0_2008,RIaed5148_2009,
        RIaed51c0_2010,RIaed5238_2011,RIaed52b0_2012,RIaed5328_2013,RIaed53a0_2014,RIaed5418_2015,RIaed5490_2016,RIaed5508_2017,RIaed5580_2018,RIaed55f8_2019,
        RIaed5670_2020,RIaed56e8_2021,RIaed5760_2022,RIaed57d8_2023,RIaed5850_2024,RIaed58c8_2025,RIaed5940_2026,RIaed59b8_2027,RIaed5a30_2028,RIaed5aa8_2029,
        RIaed5b20_2030,RIaed5b98_2031,RIaed5c10_2032,RIaed5c88_2033,RIaed5d00_2034,RIaed5d78_2035,RIaed5df0_2036,RIaed5e68_2037,RIaed5ee0_2038,RIaed5f58_2039,
        RIaed5fd0_2040,RIaed6048_2041,RIaed60c0_2042,RIaed6138_2043,RIaed61b0_2044,RIaed6228_2045,RIaed62a0_2046,RIaed6318_2047,RIaed6390_2048,RIaed6408_2049,
        RIaed6480_2050,RIaed64f8_2051,RIaed6570_2052,RIaed65e8_2053,RIaed6660_2054,RIaed66d8_2055,RIaed6750_2056,RIaed67c8_2057,RIaed6840_2058,RIaed68b8_2059,
        RIaed6930_2060,RIaed69a8_2061,RIaed6a20_2062,RIaed6a98_2063,RIaed6b10_2064,RIaed6b88_2065,RIaed6c00_2066,RIaed6c78_2067,RIaed6cf0_2068,RIaed6d68_2069,
        RIaed6de0_2070,RIaed6e58_2071,RIaed6ed0_2072,RIaed6f48_2073,RIaed6fc0_2074,RIaed7038_2075,RIaed70b0_2076,RIaed7128_2077,RIaed71a0_2078,RIaed7218_2079,
        RIaed7290_2080,RIaed7308_2081,RIaed7380_2082,RIaed73f8_2083,RIaed7470_2084,RIaed74e8_2085,RIaed7560_2086,RIaed75d8_2087,RIaed7650_2088,RIaed76c8_2089,
        RIaed7740_2090,RIaed77b8_2091,RIaed7830_2092,RIaed78a8_2093,RIaed7920_2094,RIaed7998_2095,RIaed7a10_2096,RIaed7a88_2097,RIaed7b00_2098,RIaed7b78_2099,
        RIaed7bf0_2100,RIaed7c68_2101,RIaed7ce0_2102,RIaed7d58_2103,RIaed7dd0_2104,RIaed7e48_2105,RIaed7ec0_2106,RIaed7f38_2107,RIaed7fb0_2108,RIaed8028_2109,
        RIaed80a0_2110,RIaed8118_2111,RIaed8190_2112,RIaed8208_2113,RIaed8280_2114,RIaed82f8_2115,RIaed8370_2116,RIaed83e8_2117,RIaed8460_2118,RIaed84d8_2119,
        RIaed8550_2120,RIaed85c8_2121,RIaed8640_2122,RIaed86b8_2123,RIaed8730_2124,RIaed87a8_2125,RIaed8820_2126,RIaed8898_2127,RIaed8910_2128,RIaed8988_2129,
        RIaed8a00_2130,RIaed8a78_2131,RIaed8af0_2132,RIaed8b68_2133,RIaed8be0_2134,RIaed8c58_2135,RIaed8cd0_2136,RIaed8d48_2137,RIaed8dc0_2138,RIaed8e38_2139,
        RIaed8eb0_2140,RIaed8f28_2141,RIaed8fa0_2142,RIaed9018_2143,RIaed9090_2144,RIaed9108_2145,RIaed9180_2146,RIaed91f8_2147,RIaed9270_2148,RIaed92e8_2149,
        RIaed9360_2150,RIaed93d8_2151,RIaed9450_2152,RIaed94c8_2153,RIaed9540_2154,RIaed95b8_2155,RIaed9630_2156,RIaed96a8_2157,RIaed9720_2158,RIaed9798_2159,
        RIaed9810_2160,RIaed9888_2161,RIaed9900_2162,RIaed9978_2163,RIaed99f0_2164,RIaed9a68_2165,RIaed9ae0_2166,RIaed9b58_2167,RIaed9bd0_2168,RIaed9c48_2169,
        RIaed9cc0_2170,RIaed9d38_2171,RIaed9db0_2172,RIaed9e28_2173,RIaed9ea0_2174,RIaed9f18_2175,RIaed9f90_2176,RIaeda008_2177,RIaeda080_2178,RIaeda0f8_2179,
        RIaeda170_2180,RIaeda1e8_2181,RIaeda260_2182,RIaeda2d8_2183,RIaeda350_2184,RIaeda3c8_2185,RIaeda440_2186,RIaeda4b8_2187,RIaeda530_2188,RIaeda5a8_2189,
        RIaeda620_2190,RIaeda698_2191,RIaeda710_2192,RIaeda788_2193,RIaeda800_2194,RIaeda878_2195,RIaeda8f0_2196,RIaeda968_2197,RIaeda9e0_2198,RIaedaa58_2199,
        RIaedaad0_2200,RIaedab48_2201,RIaedabc0_2202,RIaedac38_2203,RIaedacb0_2204,RIaedad28_2205,RIaedada0_2206,RIaedae18_2207,RIaedae90_2208,RIaedaf08_2209,
        RIaedaf80_2210,RIaedaff8_2211,RIaedb070_2212,RIaedb0e8_2213,RIaedb160_2214,RIaedb1d8_2215,RIaedb250_2216,RIaedb2c8_2217,RIaedb340_2218,RIaedb3b8_2219,
        RIaedb430_2220,RIaedb4a8_2221,RIaedb520_2222,RIaedb598_2223,RIaedb610_2224,RIaedb688_2225,RIaedb700_2226,RIaedb778_2227,RIaedb7f0_2228,RIaedb868_2229,
        RIaedb8e0_2230,RIaedb958_2231,RIaedb9d0_2232,RIaedba48_2233,RIaedbac0_2234,RIaedbb38_2235,RIaedbbb0_2236,RIaedbc28_2237,RIaedbca0_2238,RIaedbd18_2239,
        RIaedbd90_2240,RIaedbe08_2241,RIaedbe80_2242,RIaedbef8_2243,RIaedbf70_2244,RIaedbfe8_2245,RIaedc060_2246,RIaedc0d8_2247,RIaedc150_2248,RIaedc1c8_2249,
        RIaedc240_2250,RIaedc2b8_2251,RIaedc330_2252,RIaedc3a8_2253,RIaedc420_2254,RIaedc498_2255,RIaedc510_2256,RIaedc588_2257,RIaedc600_2258,RIaedc678_2259,
        RIaedc6f0_2260,RIaedc768_2261,RIaedc7e0_2262,RIaedc858_2263,RIaedc8d0_2264,RIaedc948_2265,RIaedc9c0_2266,RIaedca38_2267,RIaedcab0_2268,RIaedcb28_2269,
        RIaedcba0_2270,RIaedcc18_2271,RIaedcc90_2272,RIaedcd08_2273,RIaedcd80_2274,RIaedcdf8_2275,RIaedce70_2276,RIaedcee8_2277,RIaedcf60_2278,RIaedcfd8_2279,
        RIaedd050_2280,RIaedd0c8_2281,RIaedd140_2282,RIaedd1b8_2283,RIaedd230_2284,RIaedd2a8_2285,RIaedd320_2286,RIaedd398_2287,RIaedd410_2288,RIaedd488_2289,
        RIaedd500_2290,RIaedd578_2291,RIaedd5f0_2292,RIaedd668_2293,RIaedd6e0_2294,RIaedd758_2295,RIaedd7d0_2296,RIaedd848_2297,RIaedd8c0_2298,RIaedd938_2299,
        RIaedd9b0_2300,RIaedda28_2301,RIaeddaa0_2302,RIaeddb18_2303,RIaeddb90_2304,RIaeddc08_2305,RIaeddc80_2306,RIaeddcf8_2307,RIaeddd70_2308,RIaeddde8_2309,
        RIaedde60_2310,RIaedded8_2311,RIaeddf50_2312,RIaeddfc8_2313,RIaede040_2314,RIaede0b8_2315,RIaede130_2316,RIaede1a8_2317,RIaede220_2318,RIaede298_2319,
        RIaede310_2320,RIaede388_2321,RIaede400_2322,RIaede478_2323,RIaede4f0_2324,RIaede568_2325,RIaede5e0_2326,RIaede658_2327,RIaede6d0_2328,RIaede748_2329,
        RIaede7c0_2330,RIaede838_2331,RIaede8b0_2332,RIaede928_2333,RIaede9a0_2334,RIaedea18_2335,RIaedea90_2336,RIaedeb08_2337,RIaedeb80_2338,RIaedebf8_2339,
        RIaedec70_2340,RIaedece8_2341,RIaeded60_2342,RIaededd8_2343,RIaedee50_2344,RIaedeec8_2345,RIaedef40_2346,RIaedefb8_2347,RIaedf030_2348,RIaedf0a8_2349,
        RIaedf120_2350,RIaedf198_2351,RIaedf210_2352,RIaedf288_2353,RIaedf300_2354,RIaedf378_2355,RIaedf3f0_2356,RIaedf468_2357,RIaedf4e0_2358,RIaedf558_2359,
        RIaedf5d0_2360,RIaedf648_2361,RIaedf6c0_2362,RIaedf738_2363,RIaedf7b0_2364,RIaedf828_2365,RIaedf8a0_2366,RIaedf918_2367,RIaedf990_2368,RIaedfa08_2369,
        RIaedfa80_2370,RIaedfaf8_2371,RIaedfb70_2372,RIaedfbe8_2373,RIaedfc60_2374,RIaedfcd8_2375,RIaedfd50_2376,RIaedfdc8_2377,RIaedfe40_2378,RIaedfeb8_2379,
        RIaedff30_2380,RIaedffa8_2381,RIaee0020_2382,RIaee0098_2383,RIaee0110_2384,RIaee0188_2385,RIaee0200_2386,RIaee0278_2387,RIaee02f0_2388,RIaee0368_2389,
        RIaee03e0_2390,RIaee0458_2391,RIaee04d0_2392,RIaee0548_2393,RIaee05c0_2394,RIaee0638_2395,RIaee06b0_2396,RIaee0728_2397,RIaee07a0_2398,RIaee0818_2399,
        RIaee0890_2400,RIaee0908_2401,RIaee0980_2402,RIaee09f8_2403,RIaee0a70_2404,RIaee0ae8_2405,RIaee0b60_2406,RIaee0bd8_2407,RIaee0c50_2408,RIaee0cc8_2409,
        RIaee0d40_2410,RIaee0db8_2411,RIaee0e30_2412,RIaee0ea8_2413,RIaee0f20_2414,RIaee0f98_2415,RIaee1010_2416,RIaee1088_2417,RIaee1100_2418,RIaee1178_2419,
        RIaee11f0_2420,RIaee1268_2421,RIaee12e0_2422,RIaee1358_2423,RIaee13d0_2424,RIaee1448_2425,RIaee14c0_2426,RIaee1538_2427,RIaee15b0_2428,RIaee1628_2429,
        RIaee16a0_2430,RIaee1718_2431,RIaee1790_2432,RIaee1808_2433,RIaee1880_2434,RIaee18f8_2435,RIaee1970_2436,RIaee19e8_2437,RIaee1a60_2438,RIaee1ad8_2439,
        RIaee1b50_2440,RIaee1bc8_2441,RIaee1c40_2442,RIaee1cb8_2443,RIaee1d30_2444,RIaee1da8_2445,RIaee1e20_2446,RIaee1e98_2447,RIaee1f10_2448,RIaee1f88_2449,
        RIaee2000_2450,RIaee2078_2451,RIaee20f0_2452,RIaee2168_2453,RIaee21e0_2454,RIaee2258_2455,RIaee22d0_2456,RIaee2348_2457,RIaee23c0_2458,RIaee2438_2459,
        RIaee24b0_2460,RIaee2528_2461,RIaee25a0_2462,RIaee2618_2463,RIaee2690_2464,RIaee2708_2465,RIaee2780_2466,RIaee27f8_2467,RIaee2870_2468,RIaee28e8_2469,
        RIaee2960_2470,RIaee29d8_2471,RIaee2a50_2472,RIaee2ac8_2473,RIaee2b40_2474,RIaee2bb8_2475,RIaee2c30_2476,RIaee2ca8_2477,RIaee2d20_2478,RIaee2d98_2479,
        RIaee2e10_2480,RIaee2e88_2481,RIaee2f00_2482,RIaee2f78_2483,RIaee2ff0_2484,RIaee3068_2485,RIaee30e0_2486,RIaee3158_2487,RIaee31d0_2488,RIaee3248_2489,
        RIaee32c0_2490,RIaee3338_2491,RIaee33b0_2492,RIaee3428_2493,RIaee34a0_2494,RIaee3518_2495,RIaee3590_2496,RIaee3608_2497,RIaee3680_2498,RIaee36f8_2499,
        RIaee3770_2500,RIaee37e8_2501,RIaee3860_2502,RIaee38d8_2503,RIaee3950_2504,RIaee39c8_2505,RIaee3a40_2506,RIaee3ab8_2507,RIaee3b30_2508,RIaee3ba8_2509,
        RIaee3c20_2510,RIaee3c98_2511,RIaee3d10_2512,RIaee3d88_2513,RIaee3e00_2514,RIaee3e78_2515,RIaee3ef0_2516,RIaee3f68_2517,RIaee3fe0_2518,RIaee4058_2519,
        RIaee40d0_2520,RIaee4148_2521,RIaee41c0_2522,RIaee4238_2523,RIaee42b0_2524,RIaee4328_2525,RIaee43a0_2526,RIaee4418_2527,RIaee4490_2528,RIaee4508_2529,
        RIaee4580_2530,RIaee45f8_2531,RIaee4670_2532,RIaee46e8_2533,RIaee4760_2534,RIaee47d8_2535,RIaee4850_2536,RIaee48c8_2537,RIaee4940_2538,RIaee49b8_2539,
        RIaee4a30_2540,RIaee4aa8_2541,RIaee4b20_2542,RIaee4b98_2543,RIaee4c10_2544,RIaee4c88_2545,RIaee4d00_2546,RIaee4d78_2547,RIaee4df0_2548,RIaee4e68_2549,
        RIaee4ee0_2550,RIaee4f58_2551,RIaee4fd0_2552,RIaee5048_2553,RIaee50c0_2554,RIaee5138_2555,RIaee51b0_2556,RIaee5228_2557,RIaee52a0_2558,RIaee5318_2559,
        RIaee5390_2560,RIaee5408_2561,RIaee5480_2562,RIaee54f8_2563,RIaee5570_2564,RIaee55e8_2565,RIaee5660_2566,RIaee56d8_2567,RIaee5750_2568,RIaee57c8_2569,
        RIaee5840_2570,RIaee58b8_2571,RIaee5930_2572,RIaee59a8_2573,RIaee5a20_2574,RIaee5a98_2575,RIaee5b10_2576,RIaee5b88_2577,RIaee5c00_2578,RIaee5c78_2579,
        RIaee5cf0_2580,RIaee5d68_2581,RIaee5de0_2582,RIaee5e58_2583,RIaee5ed0_2584,RIaee5f48_2585,RIaee5fc0_2586,RIaee6038_2587,RIaee60b0_2588,RIaee6128_2589,
        RIaee61a0_2590,RIaee6218_2591,RIaee6290_2592,RIaee6308_2593,RIaee6380_2594,RIaee63f8_2595,RIaee6470_2596,RIaee64e8_2597,RIaee6560_2598,RIaee65d8_2599,
        RIaee6650_2600,RIaee66c8_2601,RIaee6740_2602,RIaee67b8_2603,RIaee6830_2604,RIaee68a8_2605,RIaee6920_2606,RIaee6998_2607,RIaee6a10_2608,RIaee6a88_2609,
        RIaee6b00_2610,RIaee6b78_2611,RIaee6bf0_2612,RIaee6c68_2613,RIaee6ce0_2614,RIaee6d58_2615,RIaee6dd0_2616,RIaee6e48_2617,RIaee6ec0_2618,RIaee6f38_2619,
        RIaee6fb0_2620,RIaee7028_2621,RIaee70a0_2622,RIaee7118_2623,RIaee7190_2624,RIaee7208_2625,RIaee7280_2626,RIaee72f8_2627,RIaee7370_2628,RIaee73e8_2629,
        RIaee7460_2630,RIaee74d8_2631,RIaee7550_2632,RIaee75c8_2633,RIaee7640_2634,RIaee76b8_2635,RIaee7730_2636,RIaee77a8_2637,RIaee7820_2638,RIaee7898_2639,
        RIaee7910_2640,RIaee7988_2641,RIaee7a00_2642,RIaee7a78_2643,RIaee7af0_2644,RIaee7b68_2645,RIaee7be0_2646,RIaee7c58_2647,RIaee7cd0_2648,RIaee7d48_2649,
        RIaee7dc0_2650,RIaee7e38_2651,RIaee7eb0_2652,RIaee7f28_2653,RIaee7fa0_2654,RIaee8018_2655,RIaee8090_2656,RIaee8108_2657,RIaee8180_2658,RIaee81f8_2659,
        RIaee8270_2660,RIaee82e8_2661,RIaee8360_2662,RIaee83d8_2663,RIaee8450_2664,RIaee84c8_2665,RIaee8540_2666,RIaee85b8_2667,RIaee8630_2668,RIaee86a8_2669,
        RIaee8720_2670,RIaee8798_2671,RIaee8810_2672,RIaee8888_2673,RIaee8900_2674,RIaee8978_2675,RIaee89f0_2676,RIaee8a68_2677,RIaee8ae0_2678,RIaee8b58_2679,
        RIaee8bd0_2680,RIaee8c48_2681,RIaee8cc0_2682,RIaee8d38_2683,RIaee8db0_2684,RIaee8e28_2685,RIaee8ea0_2686,RIaee8f18_2687,RIaee8f90_2688,RIaee9008_2689,
        RIaee9080_2690,RIaee90f8_2691,RIaee9170_2692,RIaee91e8_2693,RIaee9260_2694,RIaee92d8_2695,RIaee9350_2696,RIaee93c8_2697,RIaee9440_2698,RIaee94b8_2699,
        RIaee9530_2700,RIaee95a8_2701,RIaee9620_2702,RIaee9698_2703,RIaee9710_2704,RIaee9788_2705,RIaee9800_2706,RIaee9878_2707,RIaee98f0_2708,RIaee9968_2709,
        RIaee99e0_2710,RIaee9a58_2711,RIaee9ad0_2712,RIaee9b48_2713,RIaee9bc0_2714,RIaee9c38_2715,RIaee9cb0_2716,RIaee9d28_2717,RIaee9da0_2718,RIaee9e18_2719,
        RIaee9e90_2720,RIaee9f08_2721,RIaee9f80_2722,RIaee9ff8_2723,RIaeea070_2724,RIaeea0e8_2725,RIaeea160_2726,RIaeea1d8_2727,RIaeea250_2728,RIaeea2c8_2729,
        RIaeea340_2730,RIaeea3b8_2731,RIaeea430_2732,RIaeea4a8_2733,RIaeea520_2734,RIaeea598_2735,RIaeea610_2736,RIaeea688_2737,RIaeea700_2738,RIaeea778_2739,
        RIaeea7f0_2740,RIaeea868_2741,RIaeea8e0_2742,RIaeea958_2743,RIaeea9d0_2744,RIaeeaa48_2745,RIaeeaac0_2746,RIaeeab38_2747,RIaeeabb0_2748,RIaeeac28_2749,
        RIaeeaca0_2750,RIaeead18_2751,RIaeead90_2752,RIaeeae08_2753,RIaeeae80_2754,RIaeeaef8_2755,RIaeeaf70_2756,RIaeeafe8_2757,RIaeeb060_2758,RIaeeb0d8_2759,
        RIaeeb150_2760,RIaeeb1c8_2761,RIaeeb240_2762,RIaeeb2b8_2763,RIaeeb330_2764,RIaeeb3a8_2765,RIaeeb420_2766,RIaeeb498_2767,RIaeeb510_2768,RIaeeb588_2769,
        RIaeeb600_2770,RIaeeb678_2771,RIaeeb6f0_2772,RIaeeb768_2773,RIaeeb7e0_2774,RIaeeb858_2775,RIaeeb8d0_2776,RIaeeb948_2777,RIaeeb9c0_2778,RIaeeba38_2779,
        RIaeebab0_2780,RIaeebb28_2781,RIaeebba0_2782,RIaeebc18_2783,RIaeebc90_2784,RIaeebd08_2785,RIaeebd80_2786,RIaeebdf8_2787,RIaeebe70_2788,RIaeebee8_2789,
        RIaeebf60_2790,RIaeebfd8_2791,RIaeec050_2792,RIaeec0c8_2793,RIaeec140_2794,RIaeec1b8_2795,RIaeec230_2796,RIaeec2a8_2797,RIaeec320_2798,RIaeec398_2799,
        RIaeec410_2800,RIaeec488_2801,RIaeec500_2802,RIaeec578_2803,RIaeec5f0_2804,RIaeec668_2805,RIaeec6e0_2806,RIaeec758_2807,RIaeec7d0_2808,RIaeec848_2809,
        RIaeec8c0_2810,RIaeec938_2811,RIaeec9b0_2812,RIaeeca28_2813,RIaeecaa0_2814,RIaeecb18_2815,RIaeecb90_2816,RIaeecc08_2817,RIaeecc80_2818,RIaeeccf8_2819,
        RIaeecd70_2820,RIaeecde8_2821,RIaeece60_2822,RIaeeced8_2823,RIaeecf50_2824,RIaeecfc8_2825,RIaeed040_2826,RIaeed0b8_2827,RIaeed130_2828,RIaeed1a8_2829,
        RIaeed220_2830,RIaeed298_2831,RIaeed310_2832,RIaeed388_2833,RIaeed400_2834,RIaeed478_2835,RIaeed4f0_2836,RIaeed568_2837,RIaeed5e0_2838,RIaeed658_2839,
        RIaeed6d0_2840,RIaeed748_2841,RIaeed7c0_2842,RIaeed838_2843,RIaeed8b0_2844,RIaeed928_2845,RIaeed9a0_2846,RIaeeda18_2847,RIaeeda90_2848,RIaeedb08_2849,
        RIaeedb80_2850,RIaeedbf8_2851,RIaeedc70_2852,RIaeedce8_2853,RIaeedd60_2854,RIaeeddd8_2855,RIaeede50_2856,RIaeedec8_2857,RIaeedf40_2858,RIaeedfb8_2859,
        RIaeee030_2860,RIaeee0a8_2861,RIaeee120_2862,RIaeee198_2863,RIaeee210_2864,RIaeee288_2865,RIaeee300_2866,RIaeee378_2867,RIaeee3f0_2868,RIaeee468_2869,
        RIaeee4e0_2870,RIaeee558_2871,RIaeee5d0_2872,RIaeee648_2873,RIaeee6c0_2874,RIaeee738_2875,RIaeee7b0_2876,RIaeee828_2877,RIaeee8a0_2878,RIaeee918_2879,
        RIaeee990_2880,RIaeeea08_2881,RIaeeea80_2882,RIaeeeaf8_2883,RIaeeeb70_2884,RIaeeebe8_2885,RIaeeec60_2886,RIaeeecd8_2887,RIaeeed50_2888,RIaeeedc8_2889,
        RIaeeee40_2890,RIaeeeeb8_2891,RIaeeef30_2892,RIaeeefa8_2893,RIaeef020_2894,RIaeef098_2895,RIaeef110_2896,RIaeef188_2897,RIaeef200_2898,RIaeef278_2899,
        RIaeef2f0_2900,RIaeef368_2901,RIaeef3e0_2902,RIaeef458_2903,RIaeef4d0_2904,RIaeef548_2905,RIaeef5c0_2906,RIaeef638_2907,RIaeef6b0_2908,RIaeef728_2909,
        RIaeef7a0_2910,RIaeef818_2911,RIaeef890_2912,RIaeef908_2913,RIaeef980_2914,RIaeef9f8_2915,RIaeefa70_2916,RIaeefae8_2917,RIaeefb60_2918,RIaeefbd8_2919,
        RIaeefc50_2920,RIaeefcc8_2921,RIaeefd40_2922,RIaeefdb8_2923,RIaeefe30_2924,RIaeefea8_2925,RIaeeff20_2926,RIaeeff98_2927,RIaef0010_2928,RIaef0088_2929,
        RIaef0100_2930,RIaef0178_2931,RIaef01f0_2932,RIaef0268_2933,RIaef02e0_2934,RIaef0358_2935,RIaef03d0_2936,RIaef0448_2937,RIaef04c0_2938,RIaef0538_2939,
        RIaef05b0_2940,RIaef0628_2941,RIaef06a0_2942,RIaef0718_2943,RIaef0790_2944,RIaef0808_2945,RIaef0880_2946,RIaef08f8_2947,RIaef0970_2948,RIaef09e8_2949,
        RIaef0a60_2950,RIaef0ad8_2951,RIaef0b50_2952,RIaef0bc8_2953,RIaef0c40_2954,RIaef0cb8_2955,RIaef0d30_2956,RIaef0da8_2957,RIaef0e20_2958,RIaef0e98_2959,
        RIaef0f10_2960,RIaef0f88_2961,RIaef1000_2962,RIaef1078_2963,RIaef10f0_2964,RIaef1168_2965,RIaef11e0_2966,RIaef1258_2967,RIaef12d0_2968,RIaef1348_2969,
        RIaef13c0_2970,RIaef1438_2971,RIaef14b0_2972,RIaef1528_2973,RIaef15a0_2974,RIaef1618_2975,RIaef1690_2976,RIaef1708_2977,RIaef1780_2978,RIaef17f8_2979,
        RIaef1870_2980,RIaef18e8_2981,RIaef1960_2982,RIaef19d8_2983,RIaef1a50_2984,RIaef1ac8_2985,RIaef1b40_2986,RIaef1bb8_2987,RIaef1c30_2988,RIaef1ca8_2989,
        RIaef1d20_2990,RIaef1d98_2991,RIaef1e10_2992,RIaef1e88_2993,RIaef1f00_2994,RIaef1f78_2995,RIaef1ff0_2996,RIaef2068_2997,RIaef20e0_2998,RIaef2158_2999,
        RIaef21d0_3000,RIaef2248_3001,RIaef22c0_3002,RIaef2338_3003,RIaef23b0_3004,RIaef2428_3005,RIaef24a0_3006,RIaef2518_3007,RIaef2590_3008,RIaef2608_3009,
        RIaef2680_3010,RIaef26f8_3011,RIaef2770_3012,RIaef27e8_3013,RIaef2860_3014,RIaef28d8_3015,RIaef2950_3016,RIaef29c8_3017,RIaef2a40_3018,RIaef2ab8_3019,
        RIaef2b30_3020,RIaef2ba8_3021,RIaef2c20_3022,RIaef2c98_3023,RIaef2d10_3024,RIaef2d88_3025,RIaef2e00_3026,RIaef2e78_3027,RIaef2ef0_3028,RIaef2f68_3029,
        RIaef2fe0_3030,RIaef3058_3031,RIaef30d0_3032,RIaef3148_3033,RIaef31c0_3034,RIaef3238_3035,RIaef32b0_3036,RIaef3328_3037,RIaef33a0_3038,RIaef3418_3039,
        RIaef3490_3040,RIaef3508_3041,RIaef3580_3042,RIaef35f8_3043,RIaef3670_3044,RIaef36e8_3045,RIaef3760_3046,RIaef37d8_3047,RIaef3850_3048,RIaef38c8_3049,
        RIaef3940_3050,RIaef39b8_3051,RIaef3a30_3052,RIaef3aa8_3053,RIaef3b20_3054,RIaef3b98_3055,RIaef3c10_3056,RIaef3c88_3057,RIaef3d00_3058,RIaef3d78_3059,
        RIaef3df0_3060,RIaef3e68_3061,RIaef3ee0_3062,RIaef3f58_3063,RIaef3fd0_3064,RIaef4048_3065,RIaef40c0_3066,RIaef4138_3067,RIaef41b0_3068,RIaef4228_3069,
        RIaef42a0_3070,RIaef4318_3071,RIaef4390_3072,RIaef4408_3073,RIaef4480_3074,RIaef44f8_3075,RIaef4570_3076,RIaef45e8_3077,RIaef4660_3078,RIaef46d8_3079,
        RIaef4750_3080,RIaef47c8_3081,RIaef4840_3082,RIaef48b8_3083,RIaef4930_3084,RIaef49a8_3085,RIaef4a20_3086,RIaef4a98_3087,RIaef4b10_3088,RIaef4b88_3089,
        RIaef4c00_3090,RIaef4c78_3091,RIaef4cf0_3092,RIaef4d68_3093,RIaef4de0_3094,RIaef4e58_3095,RIaef4ed0_3096,RIaef4f48_3097,RIaef4fc0_3098,RIaef5038_3099,
        RIaef50b0_3100,RIaef5128_3101,RIaef51a0_3102,RIaef5218_3103,RIaef5290_3104,RIaef5308_3105,RIaef5380_3106,RIaef53f8_3107,RIaef5470_3108,RIaef54e8_3109,
        RIaef5560_3110,RIaef55d8_3111,RIaef5650_3112,RIaef56c8_3113,RIaef5740_3114,RIaef57b8_3115,RIaef5830_3116,RIaef58a8_3117,RIaef5920_3118,RIaef5998_3119,
        RIaef5a10_3120,RIaef5a88_3121,RIaef5b00_3122,RIaef5b78_3123,RIaef5bf0_3124,RIaef5c68_3125,RIaef5ce0_3126,RIaef5d58_3127,RIaef5dd0_3128,RIaef5e48_3129,
        RIaef5ec0_3130,RIaef5f38_3131,RIaef5fb0_3132,RIaef6028_3133,RIaef60a0_3134,RIaef6118_3135,RIaef6190_3136,RIaef6208_3137,RIaef6280_3138,RIaef62f8_3139,
        RIaef6370_3140,RIaef63e8_3141,RIaef6460_3142,RIaef64d8_3143,RIaef6550_3144,RIaef65c8_3145,RIaef6640_3146,RIaef66b8_3147,RIaef6730_3148,RIaef67a8_3149,
        RIaef6820_3150,RIaef6898_3151,RIaef6910_3152,RIaef6988_3153,RIaef6a00_3154,RIaef6a78_3155,RIaef6af0_3156,RIaef6b68_3157,RIaef6be0_3158,RIaef6c58_3159,
        RIaef6cd0_3160,RIaef6d48_3161,RIaef6dc0_3162,RIaef6e38_3163,RIaef6eb0_3164,RIaef6f28_3165,RIaef6fa0_3166,RIaef7018_3167,RIaef7090_3168,RIaef7108_3169,
        RIaef7180_3170,RIaef71f8_3171,RIaef7270_3172,RIaef72e8_3173,RIaef7360_3174,RIaef73d8_3175,RIaef7450_3176,RIaef74c8_3177,RIaef7540_3178,RIaef75b8_3179,
        RIaef7630_3180,RIaef76a8_3181,RIaef7720_3182,RIaef7798_3183,RIaef7810_3184,RIaef7888_3185,RIaef7900_3186,RIaef7978_3187,RIaef79f0_3188,RIaef7a68_3189,
        RIaef7ae0_3190,RIaef7b58_3191,RIaef7bd0_3192,RIaef7c48_3193,RIaef7cc0_3194,RIaef7d38_3195,RIaef7db0_3196,RIaef7e28_3197,RIaef7ea0_3198,RIaef7f18_3199,
        RIaef7f90_3200,RIaef8008_3201,RIaef8080_3202,RIaef80f8_3203,RIaef8170_3204,RIaef81e8_3205,RIaef8260_3206,RIaef82d8_3207,RIaef8350_3208,RIaef83c8_3209,
        RIaef8440_3210,RIaef84b8_3211,RIaef8530_3212,RIaef85a8_3213,RIaef8620_3214,RIaef8698_3215,RIaef8710_3216,RIaef8788_3217,RIaef8800_3218,RIaef8878_3219,
        RIaef88f0_3220,RIaef8968_3221,RIaef89e0_3222,RIaef8a58_3223,RIaef8ad0_3224,RIaef8b48_3225,RIaef8bc0_3226,RIaef8c38_3227,RIaef8cb0_3228,RIaef8d28_3229,
        RIaef8da0_3230,RIaef8e18_3231,RIaef8e90_3232,RIaef8f08_3233,RIaef8f80_3234,RIaef8ff8_3235,RIaef9070_3236,RIaef90e8_3237,RIaef9160_3238,RIaef91d8_3239,
        RIaef9250_3240,RIaef92c8_3241,RIaef9340_3242,RIaef93b8_3243,RIaef9430_3244,RIaef94a8_3245,RIaef9520_3246,RIaef9598_3247,RIaef9610_3248,RIaef9688_3249,
        RIaef9700_3250,RIaef9778_3251,RIaef97f0_3252,RIaef9868_3253,RIaef98e0_3254,RIaef9958_3255,RIaef99d0_3256,RIaef9a48_3257,RIaef9ac0_3258,RIaef9b38_3259,
        RIaef9bb0_3260,RIaef9c28_3261,RIaef9ca0_3262,RIaef9d18_3263,RIaef9d90_3264,RIaef9e08_3265,RIaef9e80_3266,RIaef9ef8_3267,RIaef9f70_3268,RIaef9fe8_3269,
        RIaefa060_3270,RIaefa0d8_3271,RIaefa150_3272,RIaefa1c8_3273,RIaefa240_3274,RIaefa2b8_3275,RIaefa330_3276,RIaefa3a8_3277,RIaefa420_3278,RIaefa498_3279,
        RIaefa510_3280,RIaefa588_3281,RIaefa600_3282,RIaefa678_3283,RIaefa6f0_3284,RIaefa768_3285,RIaefa7e0_3286,RIaefa858_3287,RIaefa8d0_3288,RIaefa948_3289,
        RIaefa9c0_3290,RIaefaa38_3291,RIaefaab0_3292,RIaefab28_3293,RIaefaba0_3294,RIaefac18_3295,RIaefac90_3296,RIaefad08_3297,RIaefad80_3298,RIaefadf8_3299,
        RIaefae70_3300,RIaefaee8_3301,RIaefaf60_3302,RIaefafd8_3303,RIaefb050_3304,RIaefb0c8_3305,RIaefb140_3306,RIaefb1b8_3307,RIaefb230_3308,RIaefb2a8_3309,
        RIaefb320_3310,RIaefb398_3311,RIaefb410_3312,RIaefb488_3313,RIaefb500_3314,RIaefb578_3315,RIaefb5f0_3316,RIaefb668_3317,RIaefb6e0_3318,RIaefb758_3319,
        RIaefb7d0_3320,RIaefb848_3321,RIaefb8c0_3322,RIaefb938_3323,RIaefb9b0_3324,RIaefba28_3325,RIaefbaa0_3326,RIaefbb18_3327,RIaefbb90_3328,RIaefbc08_3329,
        RIaefbc80_3330,RIaefbcf8_3331,RIaefbd70_3332,RIaefbde8_3333,RIaefbe60_3334,RIaefbed8_3335,RIaefbf50_3336,RIaefbfc8_3337,RIaefc040_3338,RIaefc0b8_3339,
        RIaefc130_3340,RIaefc1a8_3341,RIaefc220_3342,RIaefc298_3343,RIaefc310_3344,RIaefc388_3345,RIaefc400_3346,RIaefc478_3347,RIaefc4f0_3348,RIaefc568_3349,
        RIaefc5e0_3350,RIaefc658_3351,RIaefc6d0_3352,RIaefc748_3353,RIaefc7c0_3354,RIaefc838_3355,RIaefc8b0_3356,RIaefc928_3357,RIaefc9a0_3358,RIaefca18_3359,
        RIaefca90_3360,RIaefcb08_3361,RIaefcb80_3362,RIaefcbf8_3363,RIaefcc70_3364,RIaefcce8_3365,RIaefcd60_3366,RIaefcdd8_3367,RIaefce50_3368,RIaefcec8_3369,
        RIaefcf40_3370,RIaefcfb8_3371,RIaefd030_3372,RIaefd0a8_3373,RIaefd120_3374,RIaefd198_3375,RIaefd210_3376,RIaefd288_3377,RIaefd300_3378,RIaefd378_3379,
        RIaefd3f0_3380,RIaefd468_3381,RIaefd4e0_3382,RIaefd558_3383,RIaefd5d0_3384,RIaefd648_3385,RIaefd6c0_3386,RIaefd738_3387,RIaefd7b0_3388,RIaefd828_3389,
        RIaefd8a0_3390,RIaefd918_3391,RIaefd990_3392,RIaefda08_3393,RIaefda80_3394,RIaefdaf8_3395,RIaefdb70_3396,RIaefdbe8_3397,RIaefdc60_3398,RIaefdcd8_3399,
        RIaefdd50_3400,RIaefddc8_3401,RIaefde40_3402,RIaefdeb8_3403,RIaefdf30_3404,RIaefdfa8_3405,RIaefe020_3406,RIaefe098_3407,RIaefe110_3408,RIaefe188_3409,
        RIaefe200_3410,RIaefe278_3411,RIaefe2f0_3412,RIaefe368_3413,RIaefe3e0_3414,RIaefe458_3415,RIaefe4d0_3416,RIaefe548_3417,RIaefe5c0_3418,RIaefe638_3419,
        RIaefe6b0_3420,RIaefe728_3421,RIaefe7a0_3422,RIaefe818_3423,RIaefe890_3424,RIaefe908_3425,RIaefe980_3426,RIaefe9f8_3427,RIaefea70_3428,RIaefeae8_3429,
        RIaefeb60_3430,RIaefebd8_3431,RIaefec50_3432,RIaefecc8_3433,RIaefed40_3434,RIaefedb8_3435,RIaefee30_3436,RIaefeea8_3437,RIaefef20_3438,RIaefef98_3439,
        RIaeff010_3440,RIaeff088_3441,RIaeff100_3442,RIaeff178_3443,RIaeff1f0_3444,RIaeff268_3445,RIaeff2e0_3446,RIaeff358_3447,RIaeff3d0_3448,RIaeff448_3449,
        RIaeff4c0_3450,RIaeff538_3451,RIaeff5b0_3452,RIaeff628_3453,RIaeff6a0_3454,RIaeff718_3455,RIaeff790_3456,RIaeff808_3457,RIaeff880_3458,RIaeff8f8_3459,
        RIaeff970_3460,RIaeff9e8_3461,RIaeffa60_3462,RIaeffad8_3463,RIaeffb50_3464,RIaeffbc8_3465,RIaeffc40_3466,RIaeffcb8_3467,RIaeffd30_3468,RIaeffda8_3469,
        RIaeffe20_3470,RIaeffe98_3471,RIaefff10_3472,RIaefff88_3473,RIaf00000_3474,RIaf00078_3475,RIaf000f0_3476,RIaf00168_3477,RIaf001e0_3478,RIaf00258_3479,
        RIaf002d0_3480,RIaf00348_3481,RIaf003c0_3482,RIaf00438_3483,RIaf004b0_3484,RIaf00528_3485,RIaf005a0_3486,RIaf00618_3487,RIaf00690_3488,RIaf00708_3489,
        RIaf00780_3490,RIaf007f8_3491,RIaf00870_3492,RIaf008e8_3493,RIaf00960_3494,RIaf009d8_3495,RIaf00a50_3496,RIaf00ac8_3497,RIaf00b40_3498,RIaf00bb8_3499,
        RIaf00c30_3500,RIaf00ca8_3501,RIaf00d20_3502,RIaf00d98_3503,RIaf00e10_3504,RIaf00e88_3505,RIaf00f00_3506,RIaf00f78_3507,RIaf00ff0_3508,RIaf01068_3509,
        RIaf010e0_3510,RIaf01158_3511,RIaf011d0_3512,RIaf01248_3513,RIaf012c0_3514,RIaf01338_3515,RIaf013b0_3516,RIaf01428_3517,RIaf014a0_3518,RIaf01518_3519,
        RIaf01590_3520,RIaf01608_3521,RIaf01680_3522,RIaf016f8_3523,RIaf01770_3524,RIaf017e8_3525,RIaf01860_3526,RIaf018d8_3527,RIaf01950_3528,RIaf019c8_3529,
        RIaf01a40_3530,RIaf01ab8_3531,RIaf01b30_3532,RIaf01ba8_3533,RIaf01c20_3534,RIaf01c98_3535,RIaf01d10_3536,RIaf01d88_3537,RIaf01e00_3538,RIaf01e78_3539,
        RIaf01ef0_3540,RIaf01f68_3541,RIaf01fe0_3542,RIaf02058_3543,RIaf020d0_3544,RIaf02148_3545,RIaf021c0_3546,RIaf02238_3547,RIaf022b0_3548,RIaf02328_3549,
        RIaf023a0_3550,RIaf02418_3551,RIaf02490_3552,RIaf02508_3553,RIaf02580_3554,RIaf025f8_3555,RIaf02670_3556,RIaf026e8_3557,RIaf02760_3558,RIaf027d8_3559,
        RIaf02850_3560,RIaf028c8_3561,RIaf02940_3562,RIaf029b8_3563,RIaf02a30_3564,RIaf02aa8_3565,RIaf02b20_3566,RIaf02b98_3567,RIaf02c10_3568,RIaf02c88_3569,
        RIaf02d00_3570,RIaf02d78_3571,RIaf02df0_3572,RIaf02e68_3573,RIaf02ee0_3574,RIaf02f58_3575,RIaf02fd0_3576,RIaf03048_3577,RIaf030c0_3578,RIaf03138_3579,
        RIaf031b0_3580,RIaf03228_3581,RIaf032a0_3582,RIaf03318_3583,RIaf03390_3584,RIaf03408_3585,RIaf03480_3586,RIaf034f8_3587,RIaf03570_3588,RIaf035e8_3589,
        RIaf03660_3590,RIaf036d8_3591,RIaf03750_3592,RIaf037c8_3593,RIaf03840_3594,RIaf038b8_3595,RIaf03930_3596,RIaf039a8_3597,RIaf03a20_3598,RIaf03a98_3599,
        RIaf03b10_3600,RIaf03b88_3601,RIaf03c00_3602,RIaf03c78_3603,RIaf03cf0_3604,RIaf03d68_3605,RIaf03de0_3606,RIaf03e58_3607,RIaf03ed0_3608,RIaf03f48_3609,
        RIaf03fc0_3610,RIaf04038_3611,RIaf040b0_3612,RIaf04128_3613,RIaf041a0_3614,RIaf04218_3615,RIaf04290_3616,RIaf04308_3617,RIaf04380_3618,RIaf043f8_3619,
        RIaf04470_3620,RIaf044e8_3621,RIaf04560_3622,RIaf045d8_3623,RIaf04650_3624,RIaf046c8_3625,RIaf04740_3626,RIaf047b8_3627,RIaf04830_3628,RIaf048a8_3629,
        RIaf04920_3630,RIaf04998_3631,RIaf04a10_3632,RIaf04a88_3633,RIaf04b00_3634,RIaf04b78_3635,RIaf04bf0_3636,RIaf04c68_3637,RIaf04ce0_3638,RIaf04d58_3639,
        RIaf04dd0_3640,RIaf04e48_3641,RIaf04ec0_3642,RIaf04f38_3643,RIaf04fb0_3644,RIaf05028_3645,RIaf050a0_3646,RIaf05118_3647,RIaf05190_3648,RIaf05208_3649,
        RIaf05280_3650,RIaf052f8_3651,RIaf05370_3652,RIaf053e8_3653,RIaf05460_3654,RIaf054d8_3655,RIaf05550_3656,RIaf055c8_3657,RIaf05640_3658,RIaf056b8_3659,
        RIaf05730_3660,RIaf057a8_3661,RIaf05820_3662,RIaf05898_3663,RIaf05910_3664,RIaf05988_3665,RIaf05a00_3666,RIaf05a78_3667,RIaf05af0_3668,RIaf05b68_3669,
        RIaf05be0_3670,RIaf05c58_3671,RIaf05cd0_3672,RIaf05d48_3673,RIaf05dc0_3674,RIaf05e38_3675,RIaf05eb0_3676,RIaf05f28_3677,RIaf05fa0_3678,RIaf06018_3679,
        RIaf06090_3680,RIaf06108_3681,RIaf06180_3682,RIaf061f8_3683,RIaf06270_3684,RIaf062e8_3685,RIaf06360_3686,RIaf063d8_3687,RIaf06450_3688,RIaf064c8_3689,
        RIaf06540_3690,RIaf065b8_3691,RIaf06630_3692,RIaf066a8_3693,RIaf06720_3694,RIaf06798_3695,RIaf06810_3696,RIaf06888_3697,RIaf06900_3698,RIaf06978_3699,
        RIaf069f0_3700,RIaf06a68_3701,RIaf06ae0_3702,RIaf06b58_3703,RIaf06bd0_3704,RIaf06c48_3705,RIaf06cc0_3706,RIaf06d38_3707,RIaf06db0_3708,RIaf06e28_3709,
        RIaf06ea0_3710,RIaf06f18_3711,RIaf06f90_3712,RIaf07008_3713,RIaf07080_3714,RIaf070f8_3715,RIaf07170_3716,RIaf071e8_3717,RIaf07260_3718,RIaf072d8_3719,
        RIaf07350_3720,RIaf073c8_3721,RIaf07440_3722,RIaf074b8_3723,RIaf07530_3724,RIaf075a8_3725,RIaf07620_3726,RIaf07698_3727,RIaf07710_3728,RIaf07788_3729,
        RIaf07800_3730,RIaf07878_3731,RIaf078f0_3732,RIaf07968_3733,RIaf079e0_3734,RIaf07a58_3735,RIaf07ad0_3736,RIaf07b48_3737,RIaf07bc0_3738,RIaf07c38_3739,
        RIaf07cb0_3740,RIaf07d28_3741,RIaf07da0_3742,RIaf07e18_3743,RIaf07e90_3744,RIaf07f08_3745,RIaf07f80_3746,RIaf07ff8_3747,RIaf08070_3748,RIaf080e8_3749,
        RIaf08160_3750,RIaf081d8_3751,RIaf08250_3752,RIaf082c8_3753,RIaf08340_3754,RIaf083b8_3755,RIaf08430_3756,RIaf084a8_3757,RIaf08520_3758,RIaf08598_3759,
        RIaf08610_3760,RIaf08688_3761,RIaf08700_3762,RIaf08778_3763,RIaf087f0_3764,RIaf08868_3765,RIaf088e0_3766,RIaf08958_3767,RIaf089d0_3768,RIaf08a48_3769,
        RIaf08ac0_3770,RIaf08b38_3771,RIaf08bb0_3772,RIaf08c28_3773,RIaf08ca0_3774,RIaf08d18_3775,RIaf08d90_3776,RIaf08e08_3777,RIaf08e80_3778,RIaf08ef8_3779,
        RIaf08f70_3780,RIaf08fe8_3781,RIaf09060_3782,RIaf090d8_3783,RIaf09150_3784,RIaf091c8_3785,RIaf09240_3786,RIaf092b8_3787,RIaf09330_3788,RIaf093a8_3789,
        RIaf09420_3790,RIaf09498_3791,RIaf09510_3792,RIaf09588_3793,RIaf09600_3794,RIaf09678_3795,RIaf096f0_3796,RIaf09768_3797,RIaf097e0_3798,RIaf09858_3799,
        RIaf098d0_3800,RIaf09948_3801,RIaf099c0_3802,RIaf09a38_3803,RIaf09ab0_3804,RIaf09b28_3805,RIaf09ba0_3806,RIaf09c18_3807,RIaf09c90_3808,RIaf09d08_3809,
        RIaf09d80_3810,RIaf09df8_3811,RIaf09e70_3812,RIaf09ee8_3813,RIaf09f60_3814,RIaf09fd8_3815,RIaf0a050_3816,RIaf0a0c8_3817,RIaf0a140_3818,RIaf0a1b8_3819,
        RIaf0a230_3820,RIaf0a2a8_3821,RIaf0a320_3822,RIaf0a398_3823,RIaf0a410_3824,RIaf0a488_3825,RIaf0a500_3826,RIaf0a578_3827,RIaf0a5f0_3828,RIaf0a668_3829,
        RIaf0a6e0_3830,RIaf0a758_3831,RIaf0a7d0_3832,RIaf0a848_3833,RIaf0a8c0_3834,RIaf0a938_3835,RIaf0a9b0_3836,RIaf0aa28_3837,RIaf0aaa0_3838,RIaf0ab18_3839,
        RIaf0ab90_3840,RIaf0ac08_3841,RIaf0ac80_3842,RIaf0acf8_3843,RIaf0ad70_3844,RIaf0ade8_3845,RIaf0ae60_3846,RIaf0aed8_3847,RIaf0af50_3848,RIaf0afc8_3849,
        RIaf0b040_3850,RIaf0b0b8_3851,RIaf0b130_3852,RIaf0b1a8_3853,RIaf0b220_3854,RIaf0b298_3855,RIaf0b310_3856,RIaf0b388_3857,RIaf0b400_3858,RIaf0b478_3859,
        RIaf0b4f0_3860,RIaf0b568_3861,RIaf0b5e0_3862,RIaf0b658_3863,RIaf0b6d0_3864,RIaf0b748_3865,RIaf0b7c0_3866,RIaf0b838_3867,RIaf0b8b0_3868,RIaf0b928_3869,
        RIaf0b9a0_3870,RIaf0ba18_3871,RIaf0ba90_3872,RIaf0bb08_3873,RIaf0bb80_3874,RIaf0bbf8_3875,RIaf0bc70_3876,RIaf0bce8_3877,RIaf0bd60_3878,RIaf0bdd8_3879,
        RIaf0be50_3880,RIaf0bec8_3881,RIaf0bf40_3882,RIaf0bfb8_3883,RIaf0c030_3884,RIaf0c0a8_3885,RIaf0c120_3886,RIaf0c198_3887,RIaf0c210_3888,RIaf0c288_3889,
        RIaf0c300_3890,RIaf0c378_3891,RIaf0c3f0_3892,RIaf0c468_3893,RIaf0c4e0_3894,RIaf0c558_3895,RIaf0c5d0_3896,RIaf0c648_3897,RIaf0c6c0_3898,RIaf0c738_3899,
        RIaf0c7b0_3900,RIaf0c828_3901,RIaf0c8a0_3902,RIaf0c918_3903,RIaf0c990_3904,RIaf0ca08_3905,RIaf0ca80_3906,RIaf0caf8_3907,RIaf0cb70_3908,RIaf0cbe8_3909,
        RIaf0cc60_3910,RIaf0ccd8_3911,RIaf0cd50_3912,RIaf0cdc8_3913,RIaf0ce40_3914,RIaf0ceb8_3915,RIaf0cf30_3916,RIaf0cfa8_3917,RIaf0d020_3918,RIaf0d098_3919,
        RIaf0d110_3920,RIaf0d188_3921,RIaf0d200_3922,RIaf0d278_3923,RIaf0d2f0_3924,RIaf0d368_3925,RIaf0d3e0_3926,RIaf0d458_3927,RIaf0d4d0_3928,RIaf0d548_3929,
        RIaf0d5c0_3930,RIaf0d638_3931,RIaf0d6b0_3932,RIaf0d728_3933,RIaf0d7a0_3934,RIaf0d818_3935,RIaf0d890_3936,RIaf0d908_3937,RIaf0d980_3938,RIaf0d9f8_3939,
        RIaf0da70_3940,RIaf0dae8_3941,RIaf0db60_3942,RIaf0dbd8_3943,RIaf0dc50_3944,RIaf0dcc8_3945,RIaf0dd40_3946,RIaf0ddb8_3947,RIaf0de30_3948,RIaf0dea8_3949,
        RIaf0df20_3950,RIaf0df98_3951,RIaf0e010_3952,RIaf0e088_3953,RIaf0e100_3954,RIaf0e178_3955,RIaf0e1f0_3956,RIaf0e268_3957,RIaf0e2e0_3958,RIaf0e358_3959,
        RIaf0e3d0_3960,RIaf0e448_3961,RIaf0e4c0_3962,RIaf0e538_3963,RIaf0e5b0_3964,RIaf0e628_3965,RIaf0e6a0_3966,RIaf0e718_3967,RIaf0e790_3968,RIaf0e808_3969,
        RIaf0e880_3970,RIaf0e8f8_3971,RIaf0e970_3972,RIaf0e9e8_3973,RIaf0ea60_3974,RIaf0ead8_3975,RIaf0eb50_3976,RIaf0ebc8_3977,RIaf0ec40_3978,RIaf0ecb8_3979,
        RIaf0ed30_3980,RIaf0eda8_3981,RIaf0ee20_3982,RIaf0ee98_3983,RIaf0ef10_3984,RIaf0ef88_3985,RIaf0f000_3986,RIaf0f078_3987,RIaf0f0f0_3988,RIaf0f168_3989,
        RIaf0f1e0_3990,RIaf0f258_3991,RIaf0f2d0_3992,RIaf0f348_3993,RIaf0f3c0_3994,RIaf0f438_3995,RIaf0f4b0_3996,RIaf0f528_3997,RIaf0f5a0_3998,RIaf0f618_3999,
        RIaf0f690_4000,RIaf0f708_4001,RIaf0f780_4002,RIaf0f7f8_4003,RIaf0f870_4004,RIaf0f8e8_4005,RIaf0f960_4006,RIaf0f9d8_4007,RIaf0fa50_4008,RIaf0fac8_4009,
        RIaf0fb40_4010,RIaf0fbb8_4011,RIaf0fc30_4012,RIaf0fca8_4013,RIaf0fd20_4014,RIaf0fd98_4015,RIaf0fe10_4016,RIaf0fe88_4017,RIaf0ff00_4018,RIaf0ff78_4019,
        RIaf0fff0_4020,RIaf10068_4021,RIaf100e0_4022,RIaf10158_4023,RIaf101d0_4024,RIaf10248_4025,RIaf102c0_4026,RIaf10338_4027,RIaf103b0_4028,RIaf10428_4029,
        RIaf104a0_4030,RIaf10518_4031,RIaf10590_4032,RIaf10608_4033,RIaf10680_4034,RIaf106f8_4035,RIaf10770_4036,RIaf107e8_4037,RIaf10860_4038,RIaf108d8_4039,
        RIaf10950_4040,RIaf109c8_4041,RIaf10a40_4042,RIaf10ab8_4043,RIaf10b30_4044,RIaf10ba8_4045,RIaf10c20_4046,RIaf10c98_4047,RIaf10d10_4048,RIaf10d88_4049,
        RIaf10e00_4050,RIaf10e78_4051,RIaf10ef0_4052,RIaf10f68_4053,RIaf10fe0_4054,RIaf11058_4055,RIaf110d0_4056,RIaf11148_4057,RIaf111c0_4058,RIaf11238_4059,
        RIaf112b0_4060,RIaf11328_4061,RIaf113a0_4062,RIaf11418_4063,RIaf11490_4064,RIaf11508_4065,RIaf11580_4066,RIaf115f8_4067,RIaf11670_4068,RIaf116e8_4069,
        RIaf11760_4070,RIaf117d8_4071,RIaf11850_4072,RIaf118c8_4073,RIaf11940_4074,RIaf119b8_4075,RIaf11a30_4076,RIaf11aa8_4077,RIaf11b20_4078,RIaf11b98_4079,
        RIaf11c10_4080,RIaf11c88_4081,RIaf11d00_4082,RIaf11d78_4083,RIaf11df0_4084,RIaf11e68_4085,RIaf11ee0_4086,RIaf11f58_4087,RIaf11fd0_4088,RIaf12048_4089,
        RIaf120c0_4090,RIaf12138_4091,RIaf121b0_4092,RIaf12228_4093,RIaf122a0_4094,RIaf12318_4095,RIaf12390_4096,RIaf12408_4097,RIaf12480_4098,RIaf124f8_4099,
        RIaf12570_4100,RIaf125e8_4101,RIaf12660_4102,RIaf126d8_4103,RIaf12750_4104,RIaf127c8_4105,RIaf12840_4106,RIaf128b8_4107,RIaf12930_4108,RIaf129a8_4109,
        RIaf12a20_4110,RIaf12a98_4111,RIaf12b10_4112,RIaf12b88_4113,RIaf12c00_4114,RIaf12c78_4115,RIaf12cf0_4116,RIaf12d68_4117,RIaf12de0_4118,RIaf12e58_4119,
        RIaf12ed0_4120,RIaf12f48_4121,RIaf12fc0_4122,RIaf13038_4123,RIaf130b0_4124,RIaf13128_4125,RIaf131a0_4126,RIaf13218_4127,RIaf13290_4128,RIaf13308_4129,
        RIaf13380_4130,RIaf133f8_4131,RIaf13470_4132,RIaf134e8_4133,RIaf13560_4134,RIaf135d8_4135,RIaf13650_4136,RIaf136c8_4137,RIaf13740_4138,RIaf137b8_4139,
        RIaf13830_4140,RIaf138a8_4141,RIaf13920_4142,RIaf13998_4143,RIaf13a10_4144,RIaf13a88_4145,RIaf13b00_4146,RIaf13b78_4147,RIaf13bf0_4148,RIaf13c68_4149,
        RIaf13ce0_4150,RIaf13d58_4151,RIaf13dd0_4152,RIaf13e48_4153,RIaf13ec0_4154,RIaf13f38_4155,RIaf13fb0_4156,RIaf14028_4157,RIaf140a0_4158,RIaf14118_4159,
        RIaf14190_4160,RIaf14208_4161,RIaf14280_4162,RIaf142f8_4163,RIaf14370_4164,RIaf143e8_4165,RIaf14460_4166,RIaf144d8_4167,RIaf14550_4168,RIaf145c8_4169,
        RIaf14640_4170,RIaf146b8_4171,RIaf14730_4172,RIaf147a8_4173,RIaf14820_4174,RIaf14898_4175,RIaf14910_4176,RIaf14988_4177,RIaf14a00_4178,RIaf14a78_4179,
        RIaf14af0_4180,RIaf14b68_4181,RIaf14be0_4182,RIaf14c58_4183,RIaf14cd0_4184,RIaf14d48_4185,RIaf14dc0_4186,RIaf14e38_4187,RIaf14eb0_4188,RIaf14f28_4189,
        RIaf14fa0_4190,RIaf15018_4191,RIaf15090_4192,RIaf15108_4193,RIaf15180_4194,RIaf151f8_4195,RIaf15270_4196,RIaf152e8_4197,RIaf15360_4198,RIaf153d8_4199,
        RIaf15450_4200,RIaf154c8_4201,RIaf15540_4202,RIaf155b8_4203,RIaf15630_4204,RIaf156a8_4205,RIaf15720_4206,RIaf15798_4207,RIaf15810_4208,RIaf15888_4209,
        RIaf15900_4210,RIaf15978_4211,RIaf159f0_4212,RIaf15a68_4213,RIaf15ae0_4214,RIaf15b58_4215,RIaf15bd0_4216,RIaf15c48_4217,RIaf15cc0_4218,RIaf15d38_4219,
        RIaf15db0_4220,RIaf15e28_4221,RIaf15ea0_4222,RIaf15f18_4223,RIaf15f90_4224,RIaf16008_4225,RIaf16080_4226,RIaf160f8_4227,RIaf16170_4228,RIaf161e8_4229,
        RIaf16260_4230,RIaf162d8_4231,RIaf16350_4232,RIaf163c8_4233,RIaf16440_4234,RIaf164b8_4235,RIaf16530_4236,RIaf165a8_4237,RIaf16620_4238,RIaf16698_4239,
        RIaf16710_4240,RIaf16788_4241,RIaf16800_4242,RIaf16878_4243,RIaf168f0_4244,RIaf16968_4245,RIaf169e0_4246,RIaf16a58_4247,RIaf16ad0_4248,RIaf16b48_4249,
        RIaf16bc0_4250,RIaf16c38_4251,RIaf16cb0_4252,RIaf16d28_4253,RIaf16da0_4254,RIaf16e18_4255,RIaf16e90_4256,RIaf16f08_4257,RIaf16f80_4258,RIaf16ff8_4259,
        RIaf17070_4260,RIaf170e8_4261,RIaf17160_4262,RIaf171d8_4263,RIaf17250_4264,RIaf172c8_4265,RIaf17340_4266,RIaf173b8_4267,RIaf17430_4268,RIaf174a8_4269,
        RIaf17520_4270,RIaf17598_4271,RIaf17610_4272,RIaf17688_4273,RIaf17700_4274,RIaf17778_4275,RIaf177f0_4276,RIaf17868_4277,RIaf178e0_4278,RIaf17958_4279,
        RIaf179d0_4280,RIaf17a48_4281,RIaf17ac0_4282,RIaf17b38_4283,RIaf17bb0_4284,RIaf17c28_4285,RIaf17ca0_4286,RIaf17d18_4287,RIaf17d90_4288,RIaf17e08_4289,
        RIaf17e80_4290,RIaf17ef8_4291,RIaf17f70_4292,RIaf17fe8_4293,RIaf18060_4294,RIaf180d8_4295,RIaf18150_4296,RIaf181c8_4297,RIaf18240_4298,RIaf182b8_4299,
        RIaf18330_4300,RIaf183a8_4301,RIaf18420_4302,RIaf18498_4303,RIaf18510_4304,RIaf18588_4305,RIaf18600_4306,RIaf18678_4307,RIaf186f0_4308,RIaf18768_4309,
        RIaf187e0_4310,RIaf18858_4311,RIaf188d0_4312,RIaf18948_4313,RIaf189c0_4314,RIaf18a38_4315,RIaf18ab0_4316,RIaf18b28_4317,RIaf18ba0_4318,RIaf18c18_4319,
        RIaf18c90_4320,RIaf18d08_4321,RIaf18d80_4322,RIaf18df8_4323,RIaf18e70_4324,RIaf18ee8_4325,RIaf18f60_4326,RIaf18fd8_4327,RIaf19050_4328,RIaf190c8_4329,
        RIaf19140_4330,RIaf191b8_4331,RIaf19230_4332,RIaf192a8_4333,RIaf19320_4334,RIaf19398_4335,RIaf19410_4336,RIaf19488_4337,RIaf19500_4338,RIaf19578_4339,
        RIaf195f0_4340,RIaf19668_4341,RIaf196e0_4342,RIaf19758_4343,RIaf197d0_4344,RIaf19848_4345,RIaf198c0_4346,RIaf19938_4347,RIaf199b0_4348,RIaf19a28_4349,
        RIaf19aa0_4350,RIaf19b18_4351,RIaf19b90_4352,RIaf19c08_4353,RIaf19c80_4354,RIaf19cf8_4355,RIaf19d70_4356,RIaf19de8_4357,RIaf19e60_4358,RIaf19ed8_4359,
        RIaf19f50_4360,RIaf19fc8_4361,RIaf1a040_4362,RIaf1a0b8_4363,RIaf1a130_4364,RIaf1a1a8_4365,RIaf1a220_4366,RIaf1a298_4367,RIaf1a310_4368,RIaf1a388_4369,
        RIaf1a400_4370,RIaf1a478_4371,RIaf1a4f0_4372,RIaf1a568_4373,RIaf1a5e0_4374,RIaf1a658_4375,RIaf1a6d0_4376,RIaf1a748_4377,RIaf1a7c0_4378,RIaf1a838_4379,
        RIaf1a8b0_4380,RIaf1a928_4381,RIaf1a9a0_4382,RIaf1aa18_4383,RIaf1aa90_4384,RIaf1ab08_4385,RIaf1ab80_4386,RIaf1abf8_4387,RIaf1ac70_4388,RIaf1ace8_4389,
        RIaf1ad60_4390,RIaf1add8_4391,RIaf1ae50_4392,RIaf1aec8_4393,RIaf1af40_4394,RIaf1afb8_4395,RIaf1b030_4396,RIaf1b0a8_4397,RIaf1b120_4398,RIaf1b198_4399,
        RIaf1b210_4400,RIaf1b288_4401,RIaf1b300_4402,RIaf1b378_4403,RIaf1b3f0_4404,RIaf1b468_4405,RIaf1b4e0_4406,RIaf1b558_4407,RIaf1b5d0_4408,RIaf1b648_4409,
        RIaf1b6c0_4410,RIaf1b738_4411,RIaf1b7b0_4412,RIaf1b828_4413,RIaf1b8a0_4414,RIaf1b918_4415,RIaf1b990_4416,RIaf1ba08_4417,RIaf1ba80_4418,RIaf1baf8_4419,
        RIaf1bb70_4420,RIaf1bbe8_4421,RIaf1bc60_4422,RIaf1bcd8_4423,RIaf1bd50_4424,RIaf1bdc8_4425,RIaf1be40_4426,RIaf1beb8_4427,RIaf1bf30_4428,RIaf1bfa8_4429,
        RIaf1c020_4430,RIaf1c098_4431,RIaf1c110_4432,RIaf1c188_4433,RIaf1c200_4434,RIaf1c278_4435,RIaf1c2f0_4436,RIaf1c368_4437,RIaf1c3e0_4438,RIaf1c458_4439,
        RIaf1c4d0_4440,RIaf1c548_4441,RIaf1c5c0_4442,RIaf1c638_4443,RIaf1c6b0_4444,RIaf1c728_4445,RIaf1c7a0_4446,RIaf1c818_4447,RIaf1c890_4448,RIaf1c908_4449,
        RIaf1c980_4450,RIaf1c9f8_4451,RIaf1ca70_4452,RIaf1cae8_4453,RIaf1cb60_4454,RIaf1cbd8_4455,RIaf1cc50_4456,RIaf1ccc8_4457,RIaf1cd40_4458,RIaf1cdb8_4459,
        RIaf1ce30_4460,RIaf1cea8_4461,RIaf1cf20_4462,RIaf1cf98_4463,RIaf1d010_4464,RIaf1d088_4465,RIaf1d100_4466,RIaf1d178_4467,RIaf1d1f0_4468,RIaf1d268_4469,
        RIaf1d2e0_4470,RIaf1d358_4471,RIaf1d3d0_4472,RIaf1d448_4473,RIaf1d4c0_4474,RIaf1d538_4475,RIaf1d5b0_4476,RIaf1d628_4477,RIaf1d6a0_4478,RIaf1d718_4479,
        RIaf1d790_4480,RIaf1d808_4481,RIaf1d880_4482,RIaf1d8f8_4483,RIaf1d970_4484,RIaf1d9e8_4485,RIaf1da60_4486,RIaf1dad8_4487,RIaf1db50_4488,RIaf1dbc8_4489,
        RIaf1dc40_4490,RIaf1dcb8_4491,RIaf1dd30_4492,RIaf1dda8_4493,RIaf1de20_4494,RIaf1de98_4495,RIaf1df10_4496,RIaf1df88_4497,RIaf1e000_4498,RIaf1e078_4499,
        RIaf1e0f0_4500,RIaf1e168_4501,RIaf1e1e0_4502,RIaf1e258_4503,RIaf1e2d0_4504,RIaf1e348_4505,RIaf1e3c0_4506,RIaf1e438_4507,RIaf1e4b0_4508,RIaf1e528_4509,
        RIaf1e5a0_4510,RIaf1e618_4511,RIaf1e690_4512,RIaf1e708_4513,RIaf1e780_4514,RIaf1e7f8_4515,RIaf1e870_4516,RIaf1e8e8_4517,RIaf1e960_4518,RIaf1e9d8_4519,
        RIaf1ea50_4520,RIaf1eac8_4521,RIaf1eb40_4522,RIaf1ebb8_4523,RIaf1ec30_4524,RIaf1eca8_4525,RIaf1ed20_4526,RIaf1ed98_4527,RIaf1ee10_4528,RIaf1ee88_4529,
        RIaf1ef00_4530,RIaf1ef78_4531,RIaf1eff0_4532,RIaf1f068_4533,RIaf1f0e0_4534,RIaf1f158_4535,RIaf1f1d0_4536,RIaf1f248_4537,RIaf1f2c0_4538,RIaf1f338_4539,
        RIaf1f3b0_4540,RIaf1f428_4541,RIaf1f4a0_4542,RIaf1f518_4543,RIaf1f590_4544,RIaf1f608_4545,RIaf1f680_4546,RIaf1f6f8_4547,RIaf1f770_4548,RIaf1f7e8_4549,
        RIaf1f860_4550,RIaf1f8d8_4551,RIaf1f950_4552,RIaf1f9c8_4553,RIaf1fa40_4554,RIaf1fab8_4555,RIaf1fb30_4556,RIaf1fba8_4557,RIaf1fc20_4558,RIaf1fc98_4559,
        RIaf1fd10_4560,RIaf1fd88_4561,RIaf1fe00_4562,RIaf1fe78_4563,RIaf1fef0_4564,RIaf1ff68_4565,RIaf1ffe0_4566,RIaf20058_4567,RIaf200d0_4568,RIaf20148_4569,
        RIaf201c0_4570,RIaf20238_4571,RIaf202b0_4572,RIaf20328_4573,RIaf203a0_4574,RIaf20418_4575,RIaf20490_4576,RIaf20508_4577,RIaf20580_4578,RIaf205f8_4579,
        RIaf20670_4580,RIaf206e8_4581,RIaf20760_4582,RIaf207d8_4583,RIaf20850_4584,RIaf208c8_4585,RIaf20940_4586,RIaf209b8_4587,RIaf20a30_4588,RIaf20aa8_4589,
        RIaf20b20_4590,RIaf20b98_4591,RIaf20c10_4592,RIaf20c88_4593,RIaf20d00_4594,RIaf20d78_4595,RIaf20df0_4596,RIaf20e68_4597,RIaf20ee0_4598,RIaf20f58_4599,
        RIaf20fd0_4600,RIaf21048_4601,RIaf210c0_4602,RIaf21138_4603,RIaf211b0_4604,RIaf21228_4605,RIaf212a0_4606,RIaf21318_4607,RIaf21390_4608,RIaf21408_4609,
        RIaf21480_4610,RIaf214f8_4611,RIaf21570_4612,RIaf215e8_4613,RIaf21660_4614,RIaf216d8_4615,RIaf21750_4616,RIaf217c8_4617,RIaf21840_4618,RIaf218b8_4619,
        RIaf21930_4620,RIaf219a8_4621,RIaf21a20_4622,RIaf21a98_4623,RIaf21b10_4624,RIaf21b88_4625,RIaf21c00_4626,RIaf21c78_4627,RIaf21cf0_4628,RIaf21d68_4629,
        RIaf21de0_4630,RIaf21e58_4631,RIaf21ed0_4632,RIaf21f48_4633,RIaf21fc0_4634,RIaf22038_4635,RIaf220b0_4636,RIaf22128_4637,RIaf221a0_4638,RIaf22218_4639,
        RIaf22290_4640,RIaf22308_4641,RIaf22380_4642,RIaf223f8_4643,RIaf22470_4644,RIaf224e8_4645,RIaf22560_4646,RIaf225d8_4647,RIaf22650_4648,RIaf226c8_4649,
        RIaf22740_4650,RIaf227b8_4651,RIaf22830_4652,RIaf228a8_4653,RIaf22920_4654,RIaf22998_4655,RIaf22a10_4656,RIaf22a88_4657,RIaf22b00_4658,RIaf22b78_4659,
        RIaf22bf0_4660,RIaf22c68_4661,RIaf22ce0_4662,RIaf22d58_4663,RIaf22dd0_4664,RIaf22e48_4665,RIaf22ec0_4666,RIaf22f38_4667,RIaf22fb0_4668,RIaf23028_4669,
        RIaf230a0_4670,RIaf23118_4671,RIaf23190_4672,RIaf23208_4673,RIaf23280_4674,RIaf232f8_4675,RIaf23370_4676,RIaf233e8_4677,RIaf23460_4678,RIaf234d8_4679,
        RIaf23550_4680,R_1249_9a72be0,R_124a_9a72c88,R_124b_9a72d30,R_124c_9a72dd8,R_124d_9a72e80,R_124e_9a72f28,R_124f_9a72fd0,R_1250_9a73078,R_1251_9a73120);
input RIae9a408_1,RIae9a480_2,RIae9a4f8_3,RIae9a570_4,RIae9a5e8_5,RIae9a660_6,RIae9a6d8_7,RIae9a750_8,RIae9a7c8_9,
        RIae9a840_10,RIae9a8b8_11,RIae9a930_12,RIae9a9a8_13,RIae9aa20_14,RIae9aa98_15,RIae9ab10_16,RIae9ab88_17,RIae9ac00_18,RIae9ac78_19,
        RIae9acf0_20,RIae9ad68_21,RIae9ade0_22,RIae9ae58_23,RIae9aed0_24,RIae9af48_25,RIae9afc0_26,RIae9b038_27,RIae9b0b0_28,RIae9b128_29,
        RIae9b1a0_30,RIae9b218_31,RIae9b290_32,RIae9b308_33,RIae9b380_34,RIae9b3f8_35,RIae9b470_36,RIae9b4e8_37,RIae9b560_38,RIae9b5d8_39,
        RIae9b650_40,RIae9b6c8_41,RIae9b740_42,RIae9b7b8_43,RIae9b830_44,RIae9b8a8_45,RIae9b920_46,RIae9b998_47,RIae9ba10_48,RIae9ba88_49,
        RIae9bb00_50,RIae9bb78_51,RIae9bbf0_52,RIae9bc68_53,RIae9bce0_54,RIae9bd58_55,RIae9bdd0_56,RIae9be48_57,RIae9bec0_58,RIae9bf38_59,
        RIae9bfb0_60,RIae9c028_61,RIae9c0a0_62,RIae9c118_63,RIae9c190_64,RIae9c208_65,RIae9c280_66,RIae9c2f8_67,RIae9c370_68,RIae9c3e8_69,
        RIae9c460_70,RIae9c4d8_71,RIae9c550_72,RIae9c5c8_73,RIae9c640_74,RIae9c6b8_75,RIae9c730_76,RIae9c7a8_77,RIae9c820_78,RIae9c898_79,
        RIae9c910_80,RIae9c988_81,RIae9ca00_82,RIae9ca78_83,RIae9caf0_84,RIae9cb68_85,RIae9cbe0_86,RIae9cc58_87,RIae9ccd0_88,RIae9cd48_89,
        RIae9cdc0_90,RIae9ce38_91,RIae9ceb0_92,RIae9cf28_93,RIae9cfa0_94,RIae9d018_95,RIae9d090_96,RIae9d108_97,RIae9d180_98,RIae9d1f8_99,
        RIae9d270_100,RIae9d2e8_101,RIae9d360_102,RIae9d3d8_103,RIae9d450_104,RIae9d4c8_105,RIae9d540_106,RIae9d5b8_107,RIae9d630_108,RIae9d6a8_109,
        RIae9d720_110,RIae9d798_111,RIae9d810_112,RIae9d888_113,RIae9d900_114,RIae9d978_115,RIae9d9f0_116,RIae9da68_117,RIae9dae0_118,RIae9db58_119,
        RIae9dbd0_120,RIae9dc48_121,RIae9dcc0_122,RIae9dd38_123,RIae9ddb0_124,RIae9de28_125,RIae9dea0_126,RIae9df18_127,RIae9df90_128,RIae9e008_129,
        RIae9e080_130,RIae9e0f8_131,RIae9e170_132,RIae9e1e8_133,RIae9e260_134,RIae9e2d8_135,RIae9e350_136,RIae9e3c8_137,RIae9e440_138,RIae9e4b8_139,
        RIae9e530_140,RIae9e5a8_141,RIae9e620_142,RIae9e698_143,RIae9e710_144,RIae9e788_145,RIae9e800_146,RIae9e878_147,RIae9e8f0_148,RIae9e968_149,
        RIae9e9e0_150,RIae9ea58_151,RIae9ead0_152,RIae9eb48_153,RIae9ebc0_154,RIae9ec38_155,RIae9ecb0_156,RIae9ed28_157,RIae9eda0_158,RIae9ee18_159,
        RIae9ee90_160,RIae9ef08_161,RIae9ef80_162,RIae9eff8_163,RIae9f070_164,RIae9f0e8_165,RIae9f160_166,RIae9f1d8_167,RIae9f250_168,RIae9f2c8_169,
        RIae9f340_170,RIae9f3b8_171,RIae9f430_172,RIae9f4a8_173,RIae9f520_174,RIae9f598_175,RIae9f610_176,RIae9f688_177,RIae9f700_178,RIae9f778_179,
        RIae9f7f0_180,RIae9f868_181,RIae9f8e0_182,RIae9f958_183,RIae9f9d0_184,RIae9fa48_185,RIae9fac0_186,RIae9fb38_187,RIae9fbb0_188,RIae9fc28_189,
        RIae9fca0_190,RIae9fd18_191,RIae9fd90_192,RIae9fe08_193,RIae9fe80_194,RIae9fef8_195,RIae9ff70_196,RIae9ffe8_197,RIaea0060_198,RIaea00d8_199,
        RIaea0150_200,RIaea01c8_201,RIaea0240_202,RIaea02b8_203,RIaea0330_204,RIaea03a8_205,RIaea0420_206,RIaea0498_207,RIaea0510_208,RIaea0588_209,
        RIaea0600_210,RIaea0678_211,RIaea06f0_212,RIaea0768_213,RIaea07e0_214,RIaea0858_215,RIaea08d0_216,RIaea0948_217,RIaea09c0_218,RIaea0a38_219,
        RIaea0ab0_220,RIaea0b28_221,RIaea0ba0_222,RIaea0c18_223,RIaea0c90_224,RIaea0d08_225,RIaea0d80_226,RIaea0df8_227,RIaea0e70_228,RIaea0ee8_229,
        RIaea0f60_230,RIaea0fd8_231,RIaea1050_232,RIaea10c8_233,RIaea1140_234,RIaea11b8_235,RIaea1230_236,RIaea12a8_237,RIaea1320_238,RIaea1398_239,
        RIaea1410_240,RIaea1488_241,RIaea1500_242,RIaea1578_243,RIaea15f0_244,RIaea1668_245,RIaea16e0_246,RIaea1758_247,RIaea17d0_248,RIaea1848_249,
        RIaea18c0_250,RIaea1938_251,RIaea19b0_252,RIaea1a28_253,RIaea1aa0_254,RIaea1b18_255,RIaea1b90_256,RIaea1c08_257,RIaea1c80_258,RIaea1cf8_259,
        RIaea1d70_260,RIaea1de8_261,RIaea1e60_262,RIaea1ed8_263,RIaea1f50_264,RIaea1fc8_265,RIaea2040_266,RIaea20b8_267,RIaea2130_268,RIaea21a8_269,
        RIaea2220_270,RIaea2298_271,RIaea2310_272,RIaea2388_273,RIaea2400_274,RIaea2478_275,RIaea24f0_276,RIaea2568_277,RIaea25e0_278,RIaea2658_279,
        RIaea26d0_280,RIaea2748_281,RIaea27c0_282,RIaea2838_283,RIaea28b0_284,RIaea2928_285,RIaea29a0_286,RIaea2a18_287,RIaea2a90_288,RIaea2b08_289,
        RIaea2b80_290,RIaea2bf8_291,RIaea2c70_292,RIaea2ce8_293,RIaea2d60_294,RIaea2dd8_295,RIaea2e50_296,RIaea2ec8_297,RIaea2f40_298,RIaea2fb8_299,
        RIaea3030_300,RIaea30a8_301,RIaea3120_302,RIaea3198_303,RIaea3210_304,RIaea3288_305,RIaea3300_306,RIaea3378_307,RIaea33f0_308,RIaea3468_309,
        RIaea34e0_310,RIaea3558_311,RIaea35d0_312,RIaea3648_313,RIaea36c0_314,RIaea3738_315,RIaea37b0_316,RIaea3828_317,RIaea38a0_318,RIaea3918_319,
        RIaea3990_320,RIaea3a08_321,RIaea3a80_322,RIaea3af8_323,RIaea3b70_324,RIaea3be8_325,RIaea3c60_326,RIaea3cd8_327,RIaea3d50_328,RIaea3dc8_329,
        RIaea3e40_330,RIaea3eb8_331,RIaea3f30_332,RIaea3fa8_333,RIaea4020_334,RIaea4098_335,RIaea4110_336,RIaea4188_337,RIaea4200_338,RIaea4278_339,
        RIaea42f0_340,RIaea4368_341,RIaea43e0_342,RIaea4458_343,RIaea44d0_344,RIaea4548_345,RIaea45c0_346,RIaea4638_347,RIaea46b0_348,RIaea4728_349,
        RIaea47a0_350,RIaea4818_351,RIaea4890_352,RIaea4908_353,RIaea4980_354,RIaea49f8_355,RIaea4a70_356,RIaea4ae8_357,RIaea4b60_358,RIaea4bd8_359,
        RIaea4c50_360,RIaea4cc8_361,RIaea4d40_362,RIaea4db8_363,RIaea4e30_364,RIaea4ea8_365,RIaea4f20_366,RIaea4f98_367,RIaea5010_368,RIaea5088_369,
        RIaea5100_370,RIaea5178_371,RIaea51f0_372,RIaea5268_373,RIaea52e0_374,RIaea5358_375,RIaea53d0_376,RIaea5448_377,RIaea54c0_378,RIaea5538_379,
        RIaea55b0_380,RIaea5628_381,RIaea56a0_382,RIaea5718_383,RIaea5790_384,RIaea5808_385,RIaea5880_386,RIaea58f8_387,RIaea5970_388,RIaea59e8_389,
        RIaea5a60_390,RIaea5ad8_391,RIaea5b50_392,RIaea5bc8_393,RIaea5c40_394,RIaea5cb8_395,RIaea5d30_396,RIaea5da8_397,RIaea5e20_398,RIaea5e98_399,
        RIaea5f10_400,RIaea5f88_401,RIaea6000_402,RIaea6078_403,RIaea60f0_404,RIaea6168_405,RIaea61e0_406,RIaea6258_407,RIaea62d0_408,RIaea6348_409,
        RIaea63c0_410,RIaea6438_411,RIaea64b0_412,RIaea6528_413,RIaea65a0_414,RIaea6618_415,RIaea6690_416,RIaea6708_417,RIaea6780_418,RIaea67f8_419,
        RIaea6870_420,RIaea68e8_421,RIaea6960_422,RIaea69d8_423,RIaea6a50_424,RIaea6ac8_425,RIaea6b40_426,RIaea6bb8_427,RIaea6c30_428,RIaea6ca8_429,
        RIaea6d20_430,RIaea6d98_431,RIaea6e10_432,RIaea6e88_433,RIaea6f00_434,RIaea6f78_435,RIaea6ff0_436,RIaea7068_437,RIaea70e0_438,RIaea7158_439,
        RIaea71d0_440,RIaea7248_441,RIaea72c0_442,RIaea7338_443,RIaea73b0_444,RIaea7428_445,RIaea74a0_446,RIaea7518_447,RIaea7590_448,RIaea7608_449,
        RIaea7680_450,RIaea76f8_451,RIaea7770_452,RIaea77e8_453,RIaea7860_454,RIaea78d8_455,RIaea7950_456,RIaea79c8_457,RIaea7a40_458,RIaea7ab8_459,
        RIaea7b30_460,RIaea7ba8_461,RIaea7c20_462,RIaea7c98_463,RIaea7d10_464,RIaea7d88_465,RIaea7e00_466,RIaea7e78_467,RIaea7ef0_468,RIaea7f68_469,
        RIaea7fe0_470,RIaea8058_471,RIaea80d0_472,RIaea8148_473,RIaea81c0_474,RIaea8238_475,RIaea82b0_476,RIaea8328_477,RIaea83a0_478,RIaea8418_479,
        RIaea8490_480,RIaea8508_481,RIaea8580_482,RIaea85f8_483,RIaea8670_484,RIaea86e8_485,RIaea8760_486,RIaea87d8_487,RIaea8850_488,RIaea88c8_489,
        RIaea8940_490,RIaea89b8_491,RIaea8a30_492,RIaea8aa8_493,RIaea8b20_494,RIaea8b98_495,RIaea8c10_496,RIaea8c88_497,RIaea8d00_498,RIaea8d78_499,
        RIaea8df0_500,RIaea8e68_501,RIaea8ee0_502,RIaea8f58_503,RIaea8fd0_504,RIaea9048_505,RIaea90c0_506,RIaea9138_507,RIaea91b0_508,RIaea9228_509,
        RIaea92a0_510,RIaea9318_511,RIaea9390_512,RIaea9408_513,RIaea9480_514,RIaea94f8_515,RIaea9570_516,RIaea95e8_517,RIaea9660_518,RIaea96d8_519,
        RIaea9750_520,RIaea97c8_521,RIaea9840_522,RIaea98b8_523,RIaea9930_524,RIaea99a8_525,RIaea9a20_526,RIaea9a98_527,RIaea9b10_528,RIaea9b88_529,
        RIaea9c00_530,RIaea9c78_531,RIaea9cf0_532,RIaea9d68_533,RIaea9de0_534,RIaea9e58_535,RIaea9ed0_536,RIaea9f48_537,RIaea9fc0_538,RIaeaa038_539,
        RIaeaa0b0_540,RIaeaa128_541,RIaeaa1a0_542,RIaeaa218_543,RIaeaa290_544,RIaeaa308_545,RIaeaa380_546,RIaeaa3f8_547,RIaeaa470_548,RIaeaa4e8_549,
        RIaeaa560_550,RIaeaa5d8_551,RIaeaa650_552,RIaeaa6c8_553,RIaeaa740_554,RIaeaa7b8_555,RIaeaa830_556,RIaeaa8a8_557,RIaeaa920_558,RIaeaa998_559,
        RIaeaaa10_560,RIaeaaa88_561,RIaeaab00_562,RIaeaab78_563,RIaeaabf0_564,RIaeaac68_565,RIaeaace0_566,RIaeaad58_567,RIaeaadd0_568,RIaeaae48_569,
        RIaeaaec0_570,RIaeaaf38_571,RIaeaafb0_572,RIaeab028_573,RIaeab0a0_574,RIaeab118_575,RIaeab190_576,RIaeab208_577,RIaeab280_578,RIaeab2f8_579,
        RIaeab370_580,RIaeab3e8_581,RIaeab460_582,RIaeab4d8_583,RIaeab550_584,RIaeab5c8_585,RIaeab640_586,RIaeab6b8_587,RIaeab730_588,RIaeab7a8_589,
        RIaeab820_590,RIaeab898_591,RIaeab910_592,RIaeab988_593,RIaeaba00_594,RIaeaba78_595,RIaeabaf0_596,RIaeabb68_597,RIaeabbe0_598,RIaeabc58_599,
        RIaeabcd0_600,RIaeabd48_601,RIaeabdc0_602,RIaeabe38_603,RIaeabeb0_604,RIaeabf28_605,RIaeabfa0_606,RIaeac018_607,RIaeac090_608,RIaeac108_609,
        RIaeac180_610,RIaeac1f8_611,RIaeac270_612,RIaeac2e8_613,RIaeac360_614,RIaeac3d8_615,RIaeac450_616,RIaeac4c8_617,RIaeac540_618,RIaeac5b8_619,
        RIaeac630_620,RIaeac6a8_621,RIaeac720_622,RIaeac798_623,RIaeac810_624,RIaeac888_625,RIaeac900_626,RIaeac978_627,RIaeac9f0_628,RIaeaca68_629,
        RIaeacae0_630,RIaeacb58_631,RIaeacbd0_632,RIaeacc48_633,RIaeaccc0_634,RIaeacd38_635,RIaeacdb0_636,RIaeace28_637,RIaeacea0_638,RIaeacf18_639,
        RIaeacf90_640,RIaead008_641,RIaead080_642,RIaead0f8_643,RIaead170_644,RIaead1e8_645,RIaead260_646,RIaead2d8_647,RIaead350_648,RIaead3c8_649,
        RIaead440_650,RIaead4b8_651,RIaead530_652,RIaead5a8_653,RIaead620_654,RIaead698_655,RIaead710_656,RIaead788_657,RIaead800_658,RIaead878_659,
        RIaead8f0_660,RIaead968_661,RIaead9e0_662,RIaeada58_663,RIaeadad0_664,RIaeadb48_665,RIaeadbc0_666,RIaeadc38_667,RIaeadcb0_668,RIaeadd28_669,
        RIaeadda0_670,RIaeade18_671,RIaeade90_672,RIaeadf08_673,RIaeadf80_674,RIaeadff8_675,RIaeae070_676,RIaeae0e8_677,RIaeae160_678,RIaeae1d8_679,
        RIaeae250_680,RIaeae2c8_681,RIaeae340_682,RIaeae3b8_683,RIaeae430_684,RIaeae4a8_685,RIaeae520_686,RIaeae598_687,RIaeae610_688,RIaeae688_689,
        RIaeae700_690,RIaeae778_691,RIaeae7f0_692,RIaeae868_693,RIaeae8e0_694,RIaeae958_695,RIaeae9d0_696,RIaeaea48_697,RIaeaeac0_698,RIaeaeb38_699,
        RIaeaebb0_700,RIaeaec28_701,RIaeaeca0_702,RIaeaed18_703,RIaeaed90_704,RIaeaee08_705,RIaeaee80_706,RIaeaeef8_707,RIaeaef70_708,RIaeaefe8_709,
        RIaeaf060_710,RIaeaf0d8_711,RIaeaf150_712,RIaeaf1c8_713,RIaeaf240_714,RIaeaf2b8_715,RIaeaf330_716,RIaeaf3a8_717,RIaeaf420_718,RIaeaf498_719,
        RIaeaf510_720,RIaeaf588_721,RIaeaf600_722,RIaeaf678_723,RIaeaf6f0_724,RIaeaf768_725,RIaeaf7e0_726,RIaeaf858_727,RIaeaf8d0_728,RIaeaf948_729,
        RIaeaf9c0_730,RIaeafa38_731,RIaeafab0_732,RIaeafb28_733,RIaeafba0_734,RIaeafc18_735,RIaeafc90_736,RIaeafd08_737,RIaeafd80_738,RIaeafdf8_739,
        RIaeafe70_740,RIaeafee8_741,RIaeaff60_742,RIaeaffd8_743,RIaeb0050_744,RIaeb00c8_745,RIaeb0140_746,RIaeb01b8_747,RIaeb0230_748,RIaeb02a8_749,
        RIaeb0320_750,RIaeb0398_751,RIaeb0410_752,RIaeb0488_753,RIaeb0500_754,RIaeb0578_755,RIaeb05f0_756,RIaeb0668_757,RIaeb06e0_758,RIaeb0758_759,
        RIaeb07d0_760,RIaeb0848_761,RIaeb08c0_762,RIaeb0938_763,RIaeb09b0_764,RIaeb0a28_765,RIaeb0aa0_766,RIaeb0b18_767,RIaeb0b90_768,RIaeb0c08_769,
        RIaeb0c80_770,RIaeb0cf8_771,RIaeb0d70_772,RIaeb0de8_773,RIaeb0e60_774,RIaeb0ed8_775,RIaeb0f50_776,RIaeb0fc8_777,RIaeb1040_778,RIaeb10b8_779,
        RIaeb1130_780,RIaeb11a8_781,RIaeb1220_782,RIaeb1298_783,RIaeb1310_784,RIaeb1388_785,RIaeb1400_786,RIaeb1478_787,RIaeb14f0_788,RIaeb1568_789,
        RIaeb15e0_790,RIaeb1658_791,RIaeb16d0_792,RIaeb1748_793,RIaeb17c0_794,RIaeb1838_795,RIaeb18b0_796,RIaeb1928_797,RIaeb19a0_798,RIaeb1a18_799,
        RIaeb1a90_800,RIaeb1b08_801,RIaeb1b80_802,RIaeb1bf8_803,RIaeb1c70_804,RIaeb1ce8_805,RIaeb1d60_806,RIaeb1dd8_807,RIaeb1e50_808,RIaeb1ec8_809,
        RIaeb1f40_810,RIaeb1fb8_811,RIaeb2030_812,RIaeb20a8_813,RIaeb2120_814,RIaeb2198_815,RIaeb2210_816,RIaeb2288_817,RIaeb2300_818,RIaeb2378_819,
        RIaeb23f0_820,RIaeb2468_821,RIaeb24e0_822,RIaeb2558_823,RIaeb25d0_824,RIaeb2648_825,RIaeb26c0_826,RIaeb2738_827,RIaeb27b0_828,RIaeb2828_829,
        RIaeb28a0_830,RIaeb2918_831,RIaeb2990_832,RIaeb2a08_833,RIaeb2a80_834,RIaeb2af8_835,RIaeb2b70_836,RIaeb2be8_837,RIaeb2c60_838,RIaeb2cd8_839,
        RIaeb2d50_840,RIaeb2dc8_841,RIaeb2e40_842,RIaeb2eb8_843,RIaeb2f30_844,RIaeb2fa8_845,RIaeb3020_846,RIaeb3098_847,RIaeb3110_848,RIaeb3188_849,
        RIaeb3200_850,RIaeb3278_851,RIaeb32f0_852,RIaeb3368_853,RIaeb33e0_854,RIaeb3458_855,RIaeb34d0_856,RIaeb3548_857,RIaeb35c0_858,RIaeb3638_859,
        RIaeb36b0_860,RIaeb3728_861,RIaeb37a0_862,RIaeb3818_863,RIaeb3890_864,RIaeb3908_865,RIaeb3980_866,RIaeb39f8_867,RIaeb3a70_868,RIaeb3ae8_869,
        RIaeb3b60_870,RIaeb3bd8_871,RIaeb3c50_872,RIaeb3cc8_873,RIaeb3d40_874,RIaeb3db8_875,RIaeb3e30_876,RIaeb3ea8_877,RIaeb3f20_878,RIaeb3f98_879,
        RIaeb4010_880,RIaeb4088_881,RIaeb4100_882,RIaeb4178_883,RIaeb41f0_884,RIaeb4268_885,RIaeb42e0_886,RIaeb4358_887,RIaeb43d0_888,RIaeb4448_889,
        RIaeb44c0_890,RIaeb4538_891,RIaeb45b0_892,RIaeb4628_893,RIaeb46a0_894,RIaeb4718_895,RIaeb4790_896,RIaeb4808_897,RIaeb4880_898,RIaeb48f8_899,
        RIaeb4970_900,RIaeb49e8_901,RIaeb4a60_902,RIaeb4ad8_903,RIaeb4b50_904,RIaeb4bc8_905,RIaeb4c40_906,RIaeb4cb8_907,RIaeb4d30_908,RIaeb4da8_909,
        RIaeb4e20_910,RIaeb4e98_911,RIaeb4f10_912,RIaeb4f88_913,RIaeb5000_914,RIaeb5078_915,RIaeb50f0_916,RIaeb5168_917,RIaeb51e0_918,RIaeb5258_919,
        RIaeb52d0_920,RIaeb5348_921,RIaeb53c0_922,RIaeb5438_923,RIaeb54b0_924,RIaeb5528_925,RIaeb55a0_926,RIaeb5618_927,RIaeb5690_928,RIaeb5708_929,
        RIaeb5780_930,RIaeb57f8_931,RIaeb5870_932,RIaeb58e8_933,RIaeb5960_934,RIaeb59d8_935,RIaeb5a50_936,RIaeb5ac8_937,RIaeb5b40_938,RIaeb5bb8_939,
        RIaeb5c30_940,RIaeb5ca8_941,RIaeb5d20_942,RIaeb5d98_943,RIaeb5e10_944,RIaeb5e88_945,RIaeb5f00_946,RIaeb5f78_947,RIaeb5ff0_948,RIaeb6068_949,
        RIaeb60e0_950,RIaeb6158_951,RIaeb61d0_952,RIaeb6248_953,RIaeb62c0_954,RIaeb6338_955,RIaeb63b0_956,RIaeb6428_957,RIaeb64a0_958,RIaeb6518_959,
        RIaeb6590_960,RIaeb6608_961,RIaeb6680_962,RIaeb66f8_963,RIaeb6770_964,RIaeb67e8_965,RIaeb6860_966,RIaeb68d8_967,RIaeb6950_968,RIaeb69c8_969,
        RIaeb6a40_970,RIaeb6ab8_971,RIaeb6b30_972,RIaeb6ba8_973,RIaeb6c20_974,RIaeb6c98_975,RIaeb6d10_976,RIaeb6d88_977,RIaeb6e00_978,RIaeb6e78_979,
        RIaeb6ef0_980,RIaeb6f68_981,RIaeb6fe0_982,RIaeb7058_983,RIaeb70d0_984,RIaeb7148_985,RIaeb71c0_986,RIaeb7238_987,RIaeb72b0_988,RIaeb7328_989,
        RIaeb73a0_990,RIaeb7418_991,RIaeb7490_992,RIaeb7508_993,RIaeb7580_994,RIaeb75f8_995,RIaeb7670_996,RIaeb76e8_997,RIaeb7760_998,RIaeb77d8_999,
        RIaeb7850_1000,RIaeb78c8_1001,RIaeb7940_1002,RIaeb79b8_1003,RIaeb7a30_1004,RIaeb7aa8_1005,RIaeb7b20_1006,RIaeb7b98_1007,RIaeb7c10_1008,RIaeb7c88_1009,
        RIaeb7d00_1010,RIaeb7d78_1011,RIaeb7df0_1012,RIaeb7e68_1013,RIaeb7ee0_1014,RIaeb7f58_1015,RIaeb7fd0_1016,RIaeb8048_1017,RIaeb80c0_1018,RIaeb8138_1019,
        RIaeb81b0_1020,RIaeb8228_1021,RIaeb82a0_1022,RIaeb8318_1023,RIaeb8390_1024,RIaeb8408_1025,RIaeb8480_1026,RIaeb84f8_1027,RIaeb8570_1028,RIaeb85e8_1029,
        RIaeb8660_1030,RIaeb86d8_1031,RIaeb8750_1032,RIaeb87c8_1033,RIaeb8840_1034,RIaeb88b8_1035,RIaeb8930_1036,RIaeb89a8_1037,RIaeb8a20_1038,RIaeb8a98_1039,
        RIaeb8b10_1040,RIaeb8b88_1041,RIaeb8c00_1042,RIaeb8c78_1043,RIaeb8cf0_1044,RIaeb8d68_1045,RIaeb8de0_1046,RIaeb8e58_1047,RIaeb8ed0_1048,RIaeb8f48_1049,
        RIaeb8fc0_1050,RIaeb9038_1051,RIaeb90b0_1052,RIaeb9128_1053,RIaeb91a0_1054,RIaeb9218_1055,RIaeb9290_1056,RIaeb9308_1057,RIaeb9380_1058,RIaeb93f8_1059,
        RIaeb9470_1060,RIaeb94e8_1061,RIaeb9560_1062,RIaeb95d8_1063,RIaeb9650_1064,RIaeb96c8_1065,RIaeb9740_1066,RIaeb97b8_1067,RIaeb9830_1068,RIaeb98a8_1069,
        RIaeb9920_1070,RIaeb9998_1071,RIaeb9a10_1072,RIaeb9a88_1073,RIaeb9b00_1074,RIaeb9b78_1075,RIaeb9bf0_1076,RIaeb9c68_1077,RIaeb9ce0_1078,RIaeb9d58_1079,
        RIaeb9dd0_1080,RIaeb9e48_1081,RIaeb9ec0_1082,RIaeb9f38_1083,RIaeb9fb0_1084,RIaeba028_1085,RIaeba0a0_1086,RIaeba118_1087,RIaeba190_1088,RIaeba208_1089,
        RIaeba280_1090,RIaeba2f8_1091,RIaeba370_1092,RIaeba3e8_1093,RIaeba460_1094,RIaeba4d8_1095,RIaeba550_1096,RIaeba5c8_1097,RIaeba640_1098,RIaeba6b8_1099,
        RIaeba730_1100,RIaeba7a8_1101,RIaeba820_1102,RIaeba898_1103,RIaeba910_1104,RIaeba988_1105,RIaebaa00_1106,RIaebaa78_1107,RIaebaaf0_1108,RIaebab68_1109,
        RIaebabe0_1110,RIaebac58_1111,RIaebacd0_1112,RIaebad48_1113,RIaebadc0_1114,RIaebae38_1115,RIaebaeb0_1116,RIaebaf28_1117,RIaebafa0_1118,RIaebb018_1119,
        RIaebb090_1120,RIaebb108_1121,RIaebb180_1122,RIaebb1f8_1123,RIaebb270_1124,RIaebb2e8_1125,RIaebb360_1126,RIaebb3d8_1127,RIaebb450_1128,RIaebb4c8_1129,
        RIaebb540_1130,RIaebb5b8_1131,RIaebb630_1132,RIaebb6a8_1133,RIaebb720_1134,RIaebb798_1135,RIaebb810_1136,RIaebb888_1137,RIaebb900_1138,RIaebb978_1139,
        RIaebb9f0_1140,RIaebba68_1141,RIaebbae0_1142,RIaebbb58_1143,RIaebbbd0_1144,RIaebbc48_1145,RIaebbcc0_1146,RIaebbd38_1147,RIaebbdb0_1148,RIaebbe28_1149,
        RIaebbea0_1150,RIaebbf18_1151,RIaebbf90_1152,RIaebc008_1153,RIaebc080_1154,RIaebc0f8_1155,RIaebc170_1156,RIaebc1e8_1157,RIaebc260_1158,RIaebc2d8_1159,
        RIaebc350_1160,RIaebc3c8_1161,RIaebc440_1162,RIaebc4b8_1163,RIaebc530_1164,RIaebc5a8_1165,RIaebc620_1166,RIaebc698_1167,RIaebc710_1168,RIaebc788_1169,
        RIaebc800_1170,RIaebc878_1171,RIaebc8f0_1172,RIaebc968_1173,RIaebc9e0_1174,RIaebca58_1175,RIaebcad0_1176,RIaebcb48_1177,RIaebcbc0_1178,RIaebcc38_1179,
        RIaebccb0_1180,RIaebcd28_1181,RIaebcda0_1182,RIaebce18_1183,RIaebce90_1184,RIaebcf08_1185,RIaebcf80_1186,RIaebcff8_1187,RIaebd070_1188,RIaebd0e8_1189,
        RIaebd160_1190,RIaebd1d8_1191,RIaebd250_1192,RIaebd2c8_1193,RIaebd340_1194,RIaebd3b8_1195,RIaebd430_1196,RIaebd4a8_1197,RIaebd520_1198,RIaebd598_1199,
        RIaebd610_1200,RIaebd688_1201,RIaebd700_1202,RIaebd778_1203,RIaebd7f0_1204,RIaebd868_1205,RIaebd8e0_1206,RIaebd958_1207,RIaebd9d0_1208,RIaebda48_1209,
        RIaebdac0_1210,RIaebdb38_1211,RIaebdbb0_1212,RIaebdc28_1213,RIaebdca0_1214,RIaebdd18_1215,RIaebdd90_1216,RIaebde08_1217,RIaebde80_1218,RIaebdef8_1219,
        RIaebdf70_1220,RIaebdfe8_1221,RIaebe060_1222,RIaebe0d8_1223,RIaebe150_1224,RIaebe1c8_1225,RIaebe240_1226,RIaebe2b8_1227,RIaebe330_1228,RIaebe3a8_1229,
        RIaebe420_1230,RIaebe498_1231,RIaebe510_1232,RIaebe588_1233,RIaebe600_1234,RIaebe678_1235,RIaebe6f0_1236,RIaebe768_1237,RIaebe7e0_1238,RIaebe858_1239,
        RIaebe8d0_1240,RIaebe948_1241,RIaebe9c0_1242,RIaebea38_1243,RIaebeab0_1244,RIaebeb28_1245,RIaebeba0_1246,RIaebec18_1247,RIaebec90_1248,RIaebed08_1249,
        RIaebed80_1250,RIaebedf8_1251,RIaebee70_1252,RIaebeee8_1253,RIaebef60_1254,RIaebefd8_1255,RIaebf050_1256,RIaebf0c8_1257,RIaebf140_1258,RIaebf1b8_1259,
        RIaebf230_1260,RIaebf2a8_1261,RIaebf320_1262,RIaebf398_1263,RIaebf410_1264,RIaebf488_1265,RIaebf500_1266,RIaebf578_1267,RIaebf5f0_1268,RIaebf668_1269,
        RIaebf6e0_1270,RIaebf758_1271,RIaebf7d0_1272,RIaebf848_1273,RIaebf8c0_1274,RIaebf938_1275,RIaebf9b0_1276,RIaebfa28_1277,RIaebfaa0_1278,RIaebfb18_1279,
        RIaebfb90_1280,RIaebfc08_1281,RIaebfc80_1282,RIaebfcf8_1283,RIaebfd70_1284,RIaebfde8_1285,RIaebfe60_1286,RIaebfed8_1287,RIaebff50_1288,RIaebffc8_1289,
        RIaec0040_1290,RIaec00b8_1291,RIaec0130_1292,RIaec01a8_1293,RIaec0220_1294,RIaec0298_1295,RIaec0310_1296,RIaec0388_1297,RIaec0400_1298,RIaec0478_1299,
        RIaec04f0_1300,RIaec0568_1301,RIaec05e0_1302,RIaec0658_1303,RIaec06d0_1304,RIaec0748_1305,RIaec07c0_1306,RIaec0838_1307,RIaec08b0_1308,RIaec0928_1309,
        RIaec09a0_1310,RIaec0a18_1311,RIaec0a90_1312,RIaec0b08_1313,RIaec0b80_1314,RIaec0bf8_1315,RIaec0c70_1316,RIaec0ce8_1317,RIaec0d60_1318,RIaec0dd8_1319,
        RIaec0e50_1320,RIaec0ec8_1321,RIaec0f40_1322,RIaec0fb8_1323,RIaec1030_1324,RIaec10a8_1325,RIaec1120_1326,RIaec1198_1327,RIaec1210_1328,RIaec1288_1329,
        RIaec1300_1330,RIaec1378_1331,RIaec13f0_1332,RIaec1468_1333,RIaec14e0_1334,RIaec1558_1335,RIaec15d0_1336,RIaec1648_1337,RIaec16c0_1338,RIaec1738_1339,
        RIaec17b0_1340,RIaec1828_1341,RIaec18a0_1342,RIaec1918_1343,RIaec1990_1344,RIaec1a08_1345,RIaec1a80_1346,RIaec1af8_1347,RIaec1b70_1348,RIaec1be8_1349,
        RIaec1c60_1350,RIaec1cd8_1351,RIaec1d50_1352,RIaec1dc8_1353,RIaec1e40_1354,RIaec1eb8_1355,RIaec1f30_1356,RIaec1fa8_1357,RIaec2020_1358,RIaec2098_1359,
        RIaec2110_1360,RIaec2188_1361,RIaec2200_1362,RIaec2278_1363,RIaec22f0_1364,RIaec2368_1365,RIaec23e0_1366,RIaec2458_1367,RIaec24d0_1368,RIaec2548_1369,
        RIaec25c0_1370,RIaec2638_1371,RIaec26b0_1372,RIaec2728_1373,RIaec27a0_1374,RIaec2818_1375,RIaec2890_1376,RIaec2908_1377,RIaec2980_1378,RIaec29f8_1379,
        RIaec2a70_1380,RIaec2ae8_1381,RIaec2b60_1382,RIaec2bd8_1383,RIaec2c50_1384,RIaec2cc8_1385,RIaec2d40_1386,RIaec2db8_1387,RIaec2e30_1388,RIaec2ea8_1389,
        RIaec2f20_1390,RIaec2f98_1391,RIaec3010_1392,RIaec3088_1393,RIaec3100_1394,RIaec3178_1395,RIaec31f0_1396,RIaec3268_1397,RIaec32e0_1398,RIaec3358_1399,
        RIaec33d0_1400,RIaec3448_1401,RIaec34c0_1402,RIaec3538_1403,RIaec35b0_1404,RIaec3628_1405,RIaec36a0_1406,RIaec3718_1407,RIaec3790_1408,RIaec3808_1409,
        RIaec3880_1410,RIaec38f8_1411,RIaec3970_1412,RIaec39e8_1413,RIaec3a60_1414,RIaec3ad8_1415,RIaec3b50_1416,RIaec3bc8_1417,RIaec3c40_1418,RIaec3cb8_1419,
        RIaec3d30_1420,RIaec3da8_1421,RIaec3e20_1422,RIaec3e98_1423,RIaec3f10_1424,RIaec3f88_1425,RIaec4000_1426,RIaec4078_1427,RIaec40f0_1428,RIaec4168_1429,
        RIaec41e0_1430,RIaec4258_1431,RIaec42d0_1432,RIaec4348_1433,RIaec43c0_1434,RIaec4438_1435,RIaec44b0_1436,RIaec4528_1437,RIaec45a0_1438,RIaec4618_1439,
        RIaec4690_1440,RIaec4708_1441,RIaec4780_1442,RIaec47f8_1443,RIaec4870_1444,RIaec48e8_1445,RIaec4960_1446,RIaec49d8_1447,RIaec4a50_1448,RIaec4ac8_1449,
        RIaec4b40_1450,RIaec4bb8_1451,RIaec4c30_1452,RIaec4ca8_1453,RIaec4d20_1454,RIaec4d98_1455,RIaec4e10_1456,RIaec4e88_1457,RIaec4f00_1458,RIaec4f78_1459,
        RIaec4ff0_1460,RIaec5068_1461,RIaec50e0_1462,RIaec5158_1463,RIaec51d0_1464,RIaec5248_1465,RIaec52c0_1466,RIaec5338_1467,RIaec53b0_1468,RIaec5428_1469,
        RIaec54a0_1470,RIaec5518_1471,RIaec5590_1472,RIaec5608_1473,RIaec5680_1474,RIaec56f8_1475,RIaec5770_1476,RIaec57e8_1477,RIaec5860_1478,RIaec58d8_1479,
        RIaec5950_1480,RIaec59c8_1481,RIaec5a40_1482,RIaec5ab8_1483,RIaec5b30_1484,RIaec5ba8_1485,RIaec5c20_1486,RIaec5c98_1487,RIaec5d10_1488,RIaec5d88_1489,
        RIaec5e00_1490,RIaec5e78_1491,RIaec5ef0_1492,RIaec5f68_1493,RIaec5fe0_1494,RIaec6058_1495,RIaec60d0_1496,RIaec6148_1497,RIaec61c0_1498,RIaec6238_1499,
        RIaec62b0_1500,RIaec6328_1501,RIaec63a0_1502,RIaec6418_1503,RIaec6490_1504,RIaec6508_1505,RIaec6580_1506,RIaec65f8_1507,RIaec6670_1508,RIaec66e8_1509,
        RIaec6760_1510,RIaec67d8_1511,RIaec6850_1512,RIaec68c8_1513,RIaec6940_1514,RIaec69b8_1515,RIaec6a30_1516,RIaec6aa8_1517,RIaec6b20_1518,RIaec6b98_1519,
        RIaec6c10_1520,RIaec6c88_1521,RIaec6d00_1522,RIaec6d78_1523,RIaec6df0_1524,RIaec6e68_1525,RIaec6ee0_1526,RIaec6f58_1527,RIaec6fd0_1528,RIaec7048_1529,
        RIaec70c0_1530,RIaec7138_1531,RIaec71b0_1532,RIaec7228_1533,RIaec72a0_1534,RIaec7318_1535,RIaec7390_1536,RIaec7408_1537,RIaec7480_1538,RIaec74f8_1539,
        RIaec7570_1540,RIaec75e8_1541,RIaec7660_1542,RIaec76d8_1543,RIaec7750_1544,RIaec77c8_1545,RIaec7840_1546,RIaec78b8_1547,RIaec7930_1548,RIaec79a8_1549,
        RIaec7a20_1550,RIaec7a98_1551,RIaec7b10_1552,RIaec7b88_1553,RIaec7c00_1554,RIaec7c78_1555,RIaec7cf0_1556,RIaec7d68_1557,RIaec7de0_1558,RIaec7e58_1559,
        RIaec7ed0_1560,RIaec7f48_1561,RIaec7fc0_1562,RIaec8038_1563,RIaec80b0_1564,RIaec8128_1565,RIaec81a0_1566,RIaec8218_1567,RIaec8290_1568,RIaec8308_1569,
        RIaec8380_1570,RIaec83f8_1571,RIaec8470_1572,RIaec84e8_1573,RIaec8560_1574,RIaec85d8_1575,RIaec8650_1576,RIaec86c8_1577,RIaec8740_1578,RIaec87b8_1579,
        RIaec8830_1580,RIaec88a8_1581,RIaec8920_1582,RIaec8998_1583,RIaec8a10_1584,RIaec8a88_1585,RIaec8b00_1586,RIaec8b78_1587,RIaec8bf0_1588,RIaec8c68_1589,
        RIaec8ce0_1590,RIaec8d58_1591,RIaec8dd0_1592,RIaec8e48_1593,RIaec8ec0_1594,RIaec8f38_1595,RIaec8fb0_1596,RIaec9028_1597,RIaec90a0_1598,RIaec9118_1599,
        RIaec9190_1600,RIaec9208_1601,RIaec9280_1602,RIaec92f8_1603,RIaec9370_1604,RIaec93e8_1605,RIaec9460_1606,RIaec94d8_1607,RIaec9550_1608,RIaec95c8_1609,
        RIaec9640_1610,RIaec96b8_1611,RIaec9730_1612,RIaec97a8_1613,RIaec9820_1614,RIaec9898_1615,RIaec9910_1616,RIaec9988_1617,RIaec9a00_1618,RIaec9a78_1619,
        RIaec9af0_1620,RIaec9b68_1621,RIaec9be0_1622,RIaec9c58_1623,RIaec9cd0_1624,RIaec9d48_1625,RIaec9dc0_1626,RIaec9e38_1627,RIaec9eb0_1628,RIaec9f28_1629,
        RIaec9fa0_1630,RIaeca018_1631,RIaeca090_1632,RIaeca108_1633,RIaeca180_1634,RIaeca1f8_1635,RIaeca270_1636,RIaeca2e8_1637,RIaeca360_1638,RIaeca3d8_1639,
        RIaeca450_1640,RIaeca4c8_1641,RIaeca540_1642,RIaeca5b8_1643,RIaeca630_1644,RIaeca6a8_1645,RIaeca720_1646,RIaeca798_1647,RIaeca810_1648,RIaeca888_1649,
        RIaeca900_1650,RIaeca978_1651,RIaeca9f0_1652,RIaecaa68_1653,RIaecaae0_1654,RIaecab58_1655,RIaecabd0_1656,RIaecac48_1657,RIaecacc0_1658,RIaecad38_1659,
        RIaecadb0_1660,RIaecae28_1661,RIaecaea0_1662,RIaecaf18_1663,RIaecaf90_1664,RIaecb008_1665,RIaecb080_1666,RIaecb0f8_1667,RIaecb170_1668,RIaecb1e8_1669,
        RIaecb260_1670,RIaecb2d8_1671,RIaecb350_1672,RIaecb3c8_1673,RIaecb440_1674,RIaecb4b8_1675,RIaecb530_1676,RIaecb5a8_1677,RIaecb620_1678,RIaecb698_1679,
        RIaecb710_1680,RIaecb788_1681,RIaecb800_1682,RIaecb878_1683,RIaecb8f0_1684,RIaecb968_1685,RIaecb9e0_1686,RIaecba58_1687,RIaecbad0_1688,RIaecbb48_1689,
        RIaecbbc0_1690,RIaecbc38_1691,RIaecbcb0_1692,RIaecbd28_1693,RIaecbda0_1694,RIaecbe18_1695,RIaecbe90_1696,RIaecbf08_1697,RIaecbf80_1698,RIaecbff8_1699,
        RIaecc070_1700,RIaecc0e8_1701,RIaecc160_1702,RIaecc1d8_1703,RIaecc250_1704,RIaecc2c8_1705,RIaecc340_1706,RIaecc3b8_1707,RIaecc430_1708,RIaecc4a8_1709,
        RIaecc520_1710,RIaecc598_1711,RIaecc610_1712,RIaecc688_1713,RIaecc700_1714,RIaecc778_1715,RIaecc7f0_1716,RIaecc868_1717,RIaecc8e0_1718,RIaecc958_1719,
        RIaecc9d0_1720,RIaecca48_1721,RIaeccac0_1722,RIaeccb38_1723,RIaeccbb0_1724,RIaeccc28_1725,RIaeccca0_1726,RIaeccd18_1727,RIaeccd90_1728,RIaecce08_1729,
        RIaecce80_1730,RIaeccef8_1731,RIaeccf70_1732,RIaeccfe8_1733,RIaecd060_1734,RIaecd0d8_1735,RIaecd150_1736,RIaecd1c8_1737,RIaecd240_1738,RIaecd2b8_1739,
        RIaecd330_1740,RIaecd3a8_1741,RIaecd420_1742,RIaecd498_1743,RIaecd510_1744,RIaecd588_1745,RIaecd600_1746,RIaecd678_1747,RIaecd6f0_1748,RIaecd768_1749,
        RIaecd7e0_1750,RIaecd858_1751,RIaecd8d0_1752,RIaecd948_1753,RIaecd9c0_1754,RIaecda38_1755,RIaecdab0_1756,RIaecdb28_1757,RIaecdba0_1758,RIaecdc18_1759,
        RIaecdc90_1760,RIaecdd08_1761,RIaecdd80_1762,RIaecddf8_1763,RIaecde70_1764,RIaecdee8_1765,RIaecdf60_1766,RIaecdfd8_1767,RIaece050_1768,RIaece0c8_1769,
        RIaece140_1770,RIaece1b8_1771,RIaece230_1772,RIaece2a8_1773,RIaece320_1774,RIaece398_1775,RIaece410_1776,RIaece488_1777,RIaece500_1778,RIaece578_1779,
        RIaece5f0_1780,RIaece668_1781,RIaece6e0_1782,RIaece758_1783,RIaece7d0_1784,RIaece848_1785,RIaece8c0_1786,RIaece938_1787,RIaece9b0_1788,RIaecea28_1789,
        RIaeceaa0_1790,RIaeceb18_1791,RIaeceb90_1792,RIaecec08_1793,RIaecec80_1794,RIaececf8_1795,RIaeced70_1796,RIaecede8_1797,RIaecee60_1798,RIaeceed8_1799,
        RIaecef50_1800,RIaecefc8_1801,RIaecf040_1802,RIaecf0b8_1803,RIaecf130_1804,RIaecf1a8_1805,RIaecf220_1806,RIaecf298_1807,RIaecf310_1808,RIaecf388_1809,
        RIaecf400_1810,RIaecf478_1811,RIaecf4f0_1812,RIaecf568_1813,RIaecf5e0_1814,RIaecf658_1815,RIaecf6d0_1816,RIaecf748_1817,RIaecf7c0_1818,RIaecf838_1819,
        RIaecf8b0_1820,RIaecf928_1821,RIaecf9a0_1822,RIaecfa18_1823,RIaecfa90_1824,RIaecfb08_1825,RIaecfb80_1826,RIaecfbf8_1827,RIaecfc70_1828,RIaecfce8_1829,
        RIaecfd60_1830,RIaecfdd8_1831,RIaecfe50_1832,RIaecfec8_1833,RIaecff40_1834,RIaecffb8_1835,RIaed0030_1836,RIaed00a8_1837,RIaed0120_1838,RIaed0198_1839,
        RIaed0210_1840,RIaed0288_1841,RIaed0300_1842,RIaed0378_1843,RIaed03f0_1844,RIaed0468_1845,RIaed04e0_1846,RIaed0558_1847,RIaed05d0_1848,RIaed0648_1849,
        RIaed06c0_1850,RIaed0738_1851,RIaed07b0_1852,RIaed0828_1853,RIaed08a0_1854,RIaed0918_1855,RIaed0990_1856,RIaed0a08_1857,RIaed0a80_1858,RIaed0af8_1859,
        RIaed0b70_1860,RIaed0be8_1861,RIaed0c60_1862,RIaed0cd8_1863,RIaed0d50_1864,RIaed0dc8_1865,RIaed0e40_1866,RIaed0eb8_1867,RIaed0f30_1868,RIaed0fa8_1869,
        RIaed1020_1870,RIaed1098_1871,RIaed1110_1872,RIaed1188_1873,RIaed1200_1874,RIaed1278_1875,RIaed12f0_1876,RIaed1368_1877,RIaed13e0_1878,RIaed1458_1879,
        RIaed14d0_1880,RIaed1548_1881,RIaed15c0_1882,RIaed1638_1883,RIaed16b0_1884,RIaed1728_1885,RIaed17a0_1886,RIaed1818_1887,RIaed1890_1888,RIaed1908_1889,
        RIaed1980_1890,RIaed19f8_1891,RIaed1a70_1892,RIaed1ae8_1893,RIaed1b60_1894,RIaed1bd8_1895,RIaed1c50_1896,RIaed1cc8_1897,RIaed1d40_1898,RIaed1db8_1899,
        RIaed1e30_1900,RIaed1ea8_1901,RIaed1f20_1902,RIaed1f98_1903,RIaed2010_1904,RIaed2088_1905,RIaed2100_1906,RIaed2178_1907,RIaed21f0_1908,RIaed2268_1909,
        RIaed22e0_1910,RIaed2358_1911,RIaed23d0_1912,RIaed2448_1913,RIaed24c0_1914,RIaed2538_1915,RIaed25b0_1916,RIaed2628_1917,RIaed26a0_1918,RIaed2718_1919,
        RIaed2790_1920,RIaed2808_1921,RIaed2880_1922,RIaed28f8_1923,RIaed2970_1924,RIaed29e8_1925,RIaed2a60_1926,RIaed2ad8_1927,RIaed2b50_1928,RIaed2bc8_1929,
        RIaed2c40_1930,RIaed2cb8_1931,RIaed2d30_1932,RIaed2da8_1933,RIaed2e20_1934,RIaed2e98_1935,RIaed2f10_1936,RIaed2f88_1937,RIaed3000_1938,RIaed3078_1939,
        RIaed30f0_1940,RIaed3168_1941,RIaed31e0_1942,RIaed3258_1943,RIaed32d0_1944,RIaed3348_1945,RIaed33c0_1946,RIaed3438_1947,RIaed34b0_1948,RIaed3528_1949,
        RIaed35a0_1950,RIaed3618_1951,RIaed3690_1952,RIaed3708_1953,RIaed3780_1954,RIaed37f8_1955,RIaed3870_1956,RIaed38e8_1957,RIaed3960_1958,RIaed39d8_1959,
        RIaed3a50_1960,RIaed3ac8_1961,RIaed3b40_1962,RIaed3bb8_1963,RIaed3c30_1964,RIaed3ca8_1965,RIaed3d20_1966,RIaed3d98_1967,RIaed3e10_1968,RIaed3e88_1969,
        RIaed3f00_1970,RIaed3f78_1971,RIaed3ff0_1972,RIaed4068_1973,RIaed40e0_1974,RIaed4158_1975,RIaed41d0_1976,RIaed4248_1977,RIaed42c0_1978,RIaed4338_1979,
        RIaed43b0_1980,RIaed4428_1981,RIaed44a0_1982,RIaed4518_1983,RIaed4590_1984,RIaed4608_1985,RIaed4680_1986,RIaed46f8_1987,RIaed4770_1988,RIaed47e8_1989,
        RIaed4860_1990,RIaed48d8_1991,RIaed4950_1992,RIaed49c8_1993,RIaed4a40_1994,RIaed4ab8_1995,RIaed4b30_1996,RIaed4ba8_1997,RIaed4c20_1998,RIaed4c98_1999,
        RIaed4d10_2000,RIaed4d88_2001,RIaed4e00_2002,RIaed4e78_2003,RIaed4ef0_2004,RIaed4f68_2005,RIaed4fe0_2006,RIaed5058_2007,RIaed50d0_2008,RIaed5148_2009,
        RIaed51c0_2010,RIaed5238_2011,RIaed52b0_2012,RIaed5328_2013,RIaed53a0_2014,RIaed5418_2015,RIaed5490_2016,RIaed5508_2017,RIaed5580_2018,RIaed55f8_2019,
        RIaed5670_2020,RIaed56e8_2021,RIaed5760_2022,RIaed57d8_2023,RIaed5850_2024,RIaed58c8_2025,RIaed5940_2026,RIaed59b8_2027,RIaed5a30_2028,RIaed5aa8_2029,
        RIaed5b20_2030,RIaed5b98_2031,RIaed5c10_2032,RIaed5c88_2033,RIaed5d00_2034,RIaed5d78_2035,RIaed5df0_2036,RIaed5e68_2037,RIaed5ee0_2038,RIaed5f58_2039,
        RIaed5fd0_2040,RIaed6048_2041,RIaed60c0_2042,RIaed6138_2043,RIaed61b0_2044,RIaed6228_2045,RIaed62a0_2046,RIaed6318_2047,RIaed6390_2048,RIaed6408_2049,
        RIaed6480_2050,RIaed64f8_2051,RIaed6570_2052,RIaed65e8_2053,RIaed6660_2054,RIaed66d8_2055,RIaed6750_2056,RIaed67c8_2057,RIaed6840_2058,RIaed68b8_2059,
        RIaed6930_2060,RIaed69a8_2061,RIaed6a20_2062,RIaed6a98_2063,RIaed6b10_2064,RIaed6b88_2065,RIaed6c00_2066,RIaed6c78_2067,RIaed6cf0_2068,RIaed6d68_2069,
        RIaed6de0_2070,RIaed6e58_2071,RIaed6ed0_2072,RIaed6f48_2073,RIaed6fc0_2074,RIaed7038_2075,RIaed70b0_2076,RIaed7128_2077,RIaed71a0_2078,RIaed7218_2079,
        RIaed7290_2080,RIaed7308_2081,RIaed7380_2082,RIaed73f8_2083,RIaed7470_2084,RIaed74e8_2085,RIaed7560_2086,RIaed75d8_2087,RIaed7650_2088,RIaed76c8_2089,
        RIaed7740_2090,RIaed77b8_2091,RIaed7830_2092,RIaed78a8_2093,RIaed7920_2094,RIaed7998_2095,RIaed7a10_2096,RIaed7a88_2097,RIaed7b00_2098,RIaed7b78_2099,
        RIaed7bf0_2100,RIaed7c68_2101,RIaed7ce0_2102,RIaed7d58_2103,RIaed7dd0_2104,RIaed7e48_2105,RIaed7ec0_2106,RIaed7f38_2107,RIaed7fb0_2108,RIaed8028_2109,
        RIaed80a0_2110,RIaed8118_2111,RIaed8190_2112,RIaed8208_2113,RIaed8280_2114,RIaed82f8_2115,RIaed8370_2116,RIaed83e8_2117,RIaed8460_2118,RIaed84d8_2119,
        RIaed8550_2120,RIaed85c8_2121,RIaed8640_2122,RIaed86b8_2123,RIaed8730_2124,RIaed87a8_2125,RIaed8820_2126,RIaed8898_2127,RIaed8910_2128,RIaed8988_2129,
        RIaed8a00_2130,RIaed8a78_2131,RIaed8af0_2132,RIaed8b68_2133,RIaed8be0_2134,RIaed8c58_2135,RIaed8cd0_2136,RIaed8d48_2137,RIaed8dc0_2138,RIaed8e38_2139,
        RIaed8eb0_2140,RIaed8f28_2141,RIaed8fa0_2142,RIaed9018_2143,RIaed9090_2144,RIaed9108_2145,RIaed9180_2146,RIaed91f8_2147,RIaed9270_2148,RIaed92e8_2149,
        RIaed9360_2150,RIaed93d8_2151,RIaed9450_2152,RIaed94c8_2153,RIaed9540_2154,RIaed95b8_2155,RIaed9630_2156,RIaed96a8_2157,RIaed9720_2158,RIaed9798_2159,
        RIaed9810_2160,RIaed9888_2161,RIaed9900_2162,RIaed9978_2163,RIaed99f0_2164,RIaed9a68_2165,RIaed9ae0_2166,RIaed9b58_2167,RIaed9bd0_2168,RIaed9c48_2169,
        RIaed9cc0_2170,RIaed9d38_2171,RIaed9db0_2172,RIaed9e28_2173,RIaed9ea0_2174,RIaed9f18_2175,RIaed9f90_2176,RIaeda008_2177,RIaeda080_2178,RIaeda0f8_2179,
        RIaeda170_2180,RIaeda1e8_2181,RIaeda260_2182,RIaeda2d8_2183,RIaeda350_2184,RIaeda3c8_2185,RIaeda440_2186,RIaeda4b8_2187,RIaeda530_2188,RIaeda5a8_2189,
        RIaeda620_2190,RIaeda698_2191,RIaeda710_2192,RIaeda788_2193,RIaeda800_2194,RIaeda878_2195,RIaeda8f0_2196,RIaeda968_2197,RIaeda9e0_2198,RIaedaa58_2199,
        RIaedaad0_2200,RIaedab48_2201,RIaedabc0_2202,RIaedac38_2203,RIaedacb0_2204,RIaedad28_2205,RIaedada0_2206,RIaedae18_2207,RIaedae90_2208,RIaedaf08_2209,
        RIaedaf80_2210,RIaedaff8_2211,RIaedb070_2212,RIaedb0e8_2213,RIaedb160_2214,RIaedb1d8_2215,RIaedb250_2216,RIaedb2c8_2217,RIaedb340_2218,RIaedb3b8_2219,
        RIaedb430_2220,RIaedb4a8_2221,RIaedb520_2222,RIaedb598_2223,RIaedb610_2224,RIaedb688_2225,RIaedb700_2226,RIaedb778_2227,RIaedb7f0_2228,RIaedb868_2229,
        RIaedb8e0_2230,RIaedb958_2231,RIaedb9d0_2232,RIaedba48_2233,RIaedbac0_2234,RIaedbb38_2235,RIaedbbb0_2236,RIaedbc28_2237,RIaedbca0_2238,RIaedbd18_2239,
        RIaedbd90_2240,RIaedbe08_2241,RIaedbe80_2242,RIaedbef8_2243,RIaedbf70_2244,RIaedbfe8_2245,RIaedc060_2246,RIaedc0d8_2247,RIaedc150_2248,RIaedc1c8_2249,
        RIaedc240_2250,RIaedc2b8_2251,RIaedc330_2252,RIaedc3a8_2253,RIaedc420_2254,RIaedc498_2255,RIaedc510_2256,RIaedc588_2257,RIaedc600_2258,RIaedc678_2259,
        RIaedc6f0_2260,RIaedc768_2261,RIaedc7e0_2262,RIaedc858_2263,RIaedc8d0_2264,RIaedc948_2265,RIaedc9c0_2266,RIaedca38_2267,RIaedcab0_2268,RIaedcb28_2269,
        RIaedcba0_2270,RIaedcc18_2271,RIaedcc90_2272,RIaedcd08_2273,RIaedcd80_2274,RIaedcdf8_2275,RIaedce70_2276,RIaedcee8_2277,RIaedcf60_2278,RIaedcfd8_2279,
        RIaedd050_2280,RIaedd0c8_2281,RIaedd140_2282,RIaedd1b8_2283,RIaedd230_2284,RIaedd2a8_2285,RIaedd320_2286,RIaedd398_2287,RIaedd410_2288,RIaedd488_2289,
        RIaedd500_2290,RIaedd578_2291,RIaedd5f0_2292,RIaedd668_2293,RIaedd6e0_2294,RIaedd758_2295,RIaedd7d0_2296,RIaedd848_2297,RIaedd8c0_2298,RIaedd938_2299,
        RIaedd9b0_2300,RIaedda28_2301,RIaeddaa0_2302,RIaeddb18_2303,RIaeddb90_2304,RIaeddc08_2305,RIaeddc80_2306,RIaeddcf8_2307,RIaeddd70_2308,RIaeddde8_2309,
        RIaedde60_2310,RIaedded8_2311,RIaeddf50_2312,RIaeddfc8_2313,RIaede040_2314,RIaede0b8_2315,RIaede130_2316,RIaede1a8_2317,RIaede220_2318,RIaede298_2319,
        RIaede310_2320,RIaede388_2321,RIaede400_2322,RIaede478_2323,RIaede4f0_2324,RIaede568_2325,RIaede5e0_2326,RIaede658_2327,RIaede6d0_2328,RIaede748_2329,
        RIaede7c0_2330,RIaede838_2331,RIaede8b0_2332,RIaede928_2333,RIaede9a0_2334,RIaedea18_2335,RIaedea90_2336,RIaedeb08_2337,RIaedeb80_2338,RIaedebf8_2339,
        RIaedec70_2340,RIaedece8_2341,RIaeded60_2342,RIaededd8_2343,RIaedee50_2344,RIaedeec8_2345,RIaedef40_2346,RIaedefb8_2347,RIaedf030_2348,RIaedf0a8_2349,
        RIaedf120_2350,RIaedf198_2351,RIaedf210_2352,RIaedf288_2353,RIaedf300_2354,RIaedf378_2355,RIaedf3f0_2356,RIaedf468_2357,RIaedf4e0_2358,RIaedf558_2359,
        RIaedf5d0_2360,RIaedf648_2361,RIaedf6c0_2362,RIaedf738_2363,RIaedf7b0_2364,RIaedf828_2365,RIaedf8a0_2366,RIaedf918_2367,RIaedf990_2368,RIaedfa08_2369,
        RIaedfa80_2370,RIaedfaf8_2371,RIaedfb70_2372,RIaedfbe8_2373,RIaedfc60_2374,RIaedfcd8_2375,RIaedfd50_2376,RIaedfdc8_2377,RIaedfe40_2378,RIaedfeb8_2379,
        RIaedff30_2380,RIaedffa8_2381,RIaee0020_2382,RIaee0098_2383,RIaee0110_2384,RIaee0188_2385,RIaee0200_2386,RIaee0278_2387,RIaee02f0_2388,RIaee0368_2389,
        RIaee03e0_2390,RIaee0458_2391,RIaee04d0_2392,RIaee0548_2393,RIaee05c0_2394,RIaee0638_2395,RIaee06b0_2396,RIaee0728_2397,RIaee07a0_2398,RIaee0818_2399,
        RIaee0890_2400,RIaee0908_2401,RIaee0980_2402,RIaee09f8_2403,RIaee0a70_2404,RIaee0ae8_2405,RIaee0b60_2406,RIaee0bd8_2407,RIaee0c50_2408,RIaee0cc8_2409,
        RIaee0d40_2410,RIaee0db8_2411,RIaee0e30_2412,RIaee0ea8_2413,RIaee0f20_2414,RIaee0f98_2415,RIaee1010_2416,RIaee1088_2417,RIaee1100_2418,RIaee1178_2419,
        RIaee11f0_2420,RIaee1268_2421,RIaee12e0_2422,RIaee1358_2423,RIaee13d0_2424,RIaee1448_2425,RIaee14c0_2426,RIaee1538_2427,RIaee15b0_2428,RIaee1628_2429,
        RIaee16a0_2430,RIaee1718_2431,RIaee1790_2432,RIaee1808_2433,RIaee1880_2434,RIaee18f8_2435,RIaee1970_2436,RIaee19e8_2437,RIaee1a60_2438,RIaee1ad8_2439,
        RIaee1b50_2440,RIaee1bc8_2441,RIaee1c40_2442,RIaee1cb8_2443,RIaee1d30_2444,RIaee1da8_2445,RIaee1e20_2446,RIaee1e98_2447,RIaee1f10_2448,RIaee1f88_2449,
        RIaee2000_2450,RIaee2078_2451,RIaee20f0_2452,RIaee2168_2453,RIaee21e0_2454,RIaee2258_2455,RIaee22d0_2456,RIaee2348_2457,RIaee23c0_2458,RIaee2438_2459,
        RIaee24b0_2460,RIaee2528_2461,RIaee25a0_2462,RIaee2618_2463,RIaee2690_2464,RIaee2708_2465,RIaee2780_2466,RIaee27f8_2467,RIaee2870_2468,RIaee28e8_2469,
        RIaee2960_2470,RIaee29d8_2471,RIaee2a50_2472,RIaee2ac8_2473,RIaee2b40_2474,RIaee2bb8_2475,RIaee2c30_2476,RIaee2ca8_2477,RIaee2d20_2478,RIaee2d98_2479,
        RIaee2e10_2480,RIaee2e88_2481,RIaee2f00_2482,RIaee2f78_2483,RIaee2ff0_2484,RIaee3068_2485,RIaee30e0_2486,RIaee3158_2487,RIaee31d0_2488,RIaee3248_2489,
        RIaee32c0_2490,RIaee3338_2491,RIaee33b0_2492,RIaee3428_2493,RIaee34a0_2494,RIaee3518_2495,RIaee3590_2496,RIaee3608_2497,RIaee3680_2498,RIaee36f8_2499,
        RIaee3770_2500,RIaee37e8_2501,RIaee3860_2502,RIaee38d8_2503,RIaee3950_2504,RIaee39c8_2505,RIaee3a40_2506,RIaee3ab8_2507,RIaee3b30_2508,RIaee3ba8_2509,
        RIaee3c20_2510,RIaee3c98_2511,RIaee3d10_2512,RIaee3d88_2513,RIaee3e00_2514,RIaee3e78_2515,RIaee3ef0_2516,RIaee3f68_2517,RIaee3fe0_2518,RIaee4058_2519,
        RIaee40d0_2520,RIaee4148_2521,RIaee41c0_2522,RIaee4238_2523,RIaee42b0_2524,RIaee4328_2525,RIaee43a0_2526,RIaee4418_2527,RIaee4490_2528,RIaee4508_2529,
        RIaee4580_2530,RIaee45f8_2531,RIaee4670_2532,RIaee46e8_2533,RIaee4760_2534,RIaee47d8_2535,RIaee4850_2536,RIaee48c8_2537,RIaee4940_2538,RIaee49b8_2539,
        RIaee4a30_2540,RIaee4aa8_2541,RIaee4b20_2542,RIaee4b98_2543,RIaee4c10_2544,RIaee4c88_2545,RIaee4d00_2546,RIaee4d78_2547,RIaee4df0_2548,RIaee4e68_2549,
        RIaee4ee0_2550,RIaee4f58_2551,RIaee4fd0_2552,RIaee5048_2553,RIaee50c0_2554,RIaee5138_2555,RIaee51b0_2556,RIaee5228_2557,RIaee52a0_2558,RIaee5318_2559,
        RIaee5390_2560,RIaee5408_2561,RIaee5480_2562,RIaee54f8_2563,RIaee5570_2564,RIaee55e8_2565,RIaee5660_2566,RIaee56d8_2567,RIaee5750_2568,RIaee57c8_2569,
        RIaee5840_2570,RIaee58b8_2571,RIaee5930_2572,RIaee59a8_2573,RIaee5a20_2574,RIaee5a98_2575,RIaee5b10_2576,RIaee5b88_2577,RIaee5c00_2578,RIaee5c78_2579,
        RIaee5cf0_2580,RIaee5d68_2581,RIaee5de0_2582,RIaee5e58_2583,RIaee5ed0_2584,RIaee5f48_2585,RIaee5fc0_2586,RIaee6038_2587,RIaee60b0_2588,RIaee6128_2589,
        RIaee61a0_2590,RIaee6218_2591,RIaee6290_2592,RIaee6308_2593,RIaee6380_2594,RIaee63f8_2595,RIaee6470_2596,RIaee64e8_2597,RIaee6560_2598,RIaee65d8_2599,
        RIaee6650_2600,RIaee66c8_2601,RIaee6740_2602,RIaee67b8_2603,RIaee6830_2604,RIaee68a8_2605,RIaee6920_2606,RIaee6998_2607,RIaee6a10_2608,RIaee6a88_2609,
        RIaee6b00_2610,RIaee6b78_2611,RIaee6bf0_2612,RIaee6c68_2613,RIaee6ce0_2614,RIaee6d58_2615,RIaee6dd0_2616,RIaee6e48_2617,RIaee6ec0_2618,RIaee6f38_2619,
        RIaee6fb0_2620,RIaee7028_2621,RIaee70a0_2622,RIaee7118_2623,RIaee7190_2624,RIaee7208_2625,RIaee7280_2626,RIaee72f8_2627,RIaee7370_2628,RIaee73e8_2629,
        RIaee7460_2630,RIaee74d8_2631,RIaee7550_2632,RIaee75c8_2633,RIaee7640_2634,RIaee76b8_2635,RIaee7730_2636,RIaee77a8_2637,RIaee7820_2638,RIaee7898_2639,
        RIaee7910_2640,RIaee7988_2641,RIaee7a00_2642,RIaee7a78_2643,RIaee7af0_2644,RIaee7b68_2645,RIaee7be0_2646,RIaee7c58_2647,RIaee7cd0_2648,RIaee7d48_2649,
        RIaee7dc0_2650,RIaee7e38_2651,RIaee7eb0_2652,RIaee7f28_2653,RIaee7fa0_2654,RIaee8018_2655,RIaee8090_2656,RIaee8108_2657,RIaee8180_2658,RIaee81f8_2659,
        RIaee8270_2660,RIaee82e8_2661,RIaee8360_2662,RIaee83d8_2663,RIaee8450_2664,RIaee84c8_2665,RIaee8540_2666,RIaee85b8_2667,RIaee8630_2668,RIaee86a8_2669,
        RIaee8720_2670,RIaee8798_2671,RIaee8810_2672,RIaee8888_2673,RIaee8900_2674,RIaee8978_2675,RIaee89f0_2676,RIaee8a68_2677,RIaee8ae0_2678,RIaee8b58_2679,
        RIaee8bd0_2680,RIaee8c48_2681,RIaee8cc0_2682,RIaee8d38_2683,RIaee8db0_2684,RIaee8e28_2685,RIaee8ea0_2686,RIaee8f18_2687,RIaee8f90_2688,RIaee9008_2689,
        RIaee9080_2690,RIaee90f8_2691,RIaee9170_2692,RIaee91e8_2693,RIaee9260_2694,RIaee92d8_2695,RIaee9350_2696,RIaee93c8_2697,RIaee9440_2698,RIaee94b8_2699,
        RIaee9530_2700,RIaee95a8_2701,RIaee9620_2702,RIaee9698_2703,RIaee9710_2704,RIaee9788_2705,RIaee9800_2706,RIaee9878_2707,RIaee98f0_2708,RIaee9968_2709,
        RIaee99e0_2710,RIaee9a58_2711,RIaee9ad0_2712,RIaee9b48_2713,RIaee9bc0_2714,RIaee9c38_2715,RIaee9cb0_2716,RIaee9d28_2717,RIaee9da0_2718,RIaee9e18_2719,
        RIaee9e90_2720,RIaee9f08_2721,RIaee9f80_2722,RIaee9ff8_2723,RIaeea070_2724,RIaeea0e8_2725,RIaeea160_2726,RIaeea1d8_2727,RIaeea250_2728,RIaeea2c8_2729,
        RIaeea340_2730,RIaeea3b8_2731,RIaeea430_2732,RIaeea4a8_2733,RIaeea520_2734,RIaeea598_2735,RIaeea610_2736,RIaeea688_2737,RIaeea700_2738,RIaeea778_2739,
        RIaeea7f0_2740,RIaeea868_2741,RIaeea8e0_2742,RIaeea958_2743,RIaeea9d0_2744,RIaeeaa48_2745,RIaeeaac0_2746,RIaeeab38_2747,RIaeeabb0_2748,RIaeeac28_2749,
        RIaeeaca0_2750,RIaeead18_2751,RIaeead90_2752,RIaeeae08_2753,RIaeeae80_2754,RIaeeaef8_2755,RIaeeaf70_2756,RIaeeafe8_2757,RIaeeb060_2758,RIaeeb0d8_2759,
        RIaeeb150_2760,RIaeeb1c8_2761,RIaeeb240_2762,RIaeeb2b8_2763,RIaeeb330_2764,RIaeeb3a8_2765,RIaeeb420_2766,RIaeeb498_2767,RIaeeb510_2768,RIaeeb588_2769,
        RIaeeb600_2770,RIaeeb678_2771,RIaeeb6f0_2772,RIaeeb768_2773,RIaeeb7e0_2774,RIaeeb858_2775,RIaeeb8d0_2776,RIaeeb948_2777,RIaeeb9c0_2778,RIaeeba38_2779,
        RIaeebab0_2780,RIaeebb28_2781,RIaeebba0_2782,RIaeebc18_2783,RIaeebc90_2784,RIaeebd08_2785,RIaeebd80_2786,RIaeebdf8_2787,RIaeebe70_2788,RIaeebee8_2789,
        RIaeebf60_2790,RIaeebfd8_2791,RIaeec050_2792,RIaeec0c8_2793,RIaeec140_2794,RIaeec1b8_2795,RIaeec230_2796,RIaeec2a8_2797,RIaeec320_2798,RIaeec398_2799,
        RIaeec410_2800,RIaeec488_2801,RIaeec500_2802,RIaeec578_2803,RIaeec5f0_2804,RIaeec668_2805,RIaeec6e0_2806,RIaeec758_2807,RIaeec7d0_2808,RIaeec848_2809,
        RIaeec8c0_2810,RIaeec938_2811,RIaeec9b0_2812,RIaeeca28_2813,RIaeecaa0_2814,RIaeecb18_2815,RIaeecb90_2816,RIaeecc08_2817,RIaeecc80_2818,RIaeeccf8_2819,
        RIaeecd70_2820,RIaeecde8_2821,RIaeece60_2822,RIaeeced8_2823,RIaeecf50_2824,RIaeecfc8_2825,RIaeed040_2826,RIaeed0b8_2827,RIaeed130_2828,RIaeed1a8_2829,
        RIaeed220_2830,RIaeed298_2831,RIaeed310_2832,RIaeed388_2833,RIaeed400_2834,RIaeed478_2835,RIaeed4f0_2836,RIaeed568_2837,RIaeed5e0_2838,RIaeed658_2839,
        RIaeed6d0_2840,RIaeed748_2841,RIaeed7c0_2842,RIaeed838_2843,RIaeed8b0_2844,RIaeed928_2845,RIaeed9a0_2846,RIaeeda18_2847,RIaeeda90_2848,RIaeedb08_2849,
        RIaeedb80_2850,RIaeedbf8_2851,RIaeedc70_2852,RIaeedce8_2853,RIaeedd60_2854,RIaeeddd8_2855,RIaeede50_2856,RIaeedec8_2857,RIaeedf40_2858,RIaeedfb8_2859,
        RIaeee030_2860,RIaeee0a8_2861,RIaeee120_2862,RIaeee198_2863,RIaeee210_2864,RIaeee288_2865,RIaeee300_2866,RIaeee378_2867,RIaeee3f0_2868,RIaeee468_2869,
        RIaeee4e0_2870,RIaeee558_2871,RIaeee5d0_2872,RIaeee648_2873,RIaeee6c0_2874,RIaeee738_2875,RIaeee7b0_2876,RIaeee828_2877,RIaeee8a0_2878,RIaeee918_2879,
        RIaeee990_2880,RIaeeea08_2881,RIaeeea80_2882,RIaeeeaf8_2883,RIaeeeb70_2884,RIaeeebe8_2885,RIaeeec60_2886,RIaeeecd8_2887,RIaeeed50_2888,RIaeeedc8_2889,
        RIaeeee40_2890,RIaeeeeb8_2891,RIaeeef30_2892,RIaeeefa8_2893,RIaeef020_2894,RIaeef098_2895,RIaeef110_2896,RIaeef188_2897,RIaeef200_2898,RIaeef278_2899,
        RIaeef2f0_2900,RIaeef368_2901,RIaeef3e0_2902,RIaeef458_2903,RIaeef4d0_2904,RIaeef548_2905,RIaeef5c0_2906,RIaeef638_2907,RIaeef6b0_2908,RIaeef728_2909,
        RIaeef7a0_2910,RIaeef818_2911,RIaeef890_2912,RIaeef908_2913,RIaeef980_2914,RIaeef9f8_2915,RIaeefa70_2916,RIaeefae8_2917,RIaeefb60_2918,RIaeefbd8_2919,
        RIaeefc50_2920,RIaeefcc8_2921,RIaeefd40_2922,RIaeefdb8_2923,RIaeefe30_2924,RIaeefea8_2925,RIaeeff20_2926,RIaeeff98_2927,RIaef0010_2928,RIaef0088_2929,
        RIaef0100_2930,RIaef0178_2931,RIaef01f0_2932,RIaef0268_2933,RIaef02e0_2934,RIaef0358_2935,RIaef03d0_2936,RIaef0448_2937,RIaef04c0_2938,RIaef0538_2939,
        RIaef05b0_2940,RIaef0628_2941,RIaef06a0_2942,RIaef0718_2943,RIaef0790_2944,RIaef0808_2945,RIaef0880_2946,RIaef08f8_2947,RIaef0970_2948,RIaef09e8_2949,
        RIaef0a60_2950,RIaef0ad8_2951,RIaef0b50_2952,RIaef0bc8_2953,RIaef0c40_2954,RIaef0cb8_2955,RIaef0d30_2956,RIaef0da8_2957,RIaef0e20_2958,RIaef0e98_2959,
        RIaef0f10_2960,RIaef0f88_2961,RIaef1000_2962,RIaef1078_2963,RIaef10f0_2964,RIaef1168_2965,RIaef11e0_2966,RIaef1258_2967,RIaef12d0_2968,RIaef1348_2969,
        RIaef13c0_2970,RIaef1438_2971,RIaef14b0_2972,RIaef1528_2973,RIaef15a0_2974,RIaef1618_2975,RIaef1690_2976,RIaef1708_2977,RIaef1780_2978,RIaef17f8_2979,
        RIaef1870_2980,RIaef18e8_2981,RIaef1960_2982,RIaef19d8_2983,RIaef1a50_2984,RIaef1ac8_2985,RIaef1b40_2986,RIaef1bb8_2987,RIaef1c30_2988,RIaef1ca8_2989,
        RIaef1d20_2990,RIaef1d98_2991,RIaef1e10_2992,RIaef1e88_2993,RIaef1f00_2994,RIaef1f78_2995,RIaef1ff0_2996,RIaef2068_2997,RIaef20e0_2998,RIaef2158_2999,
        RIaef21d0_3000,RIaef2248_3001,RIaef22c0_3002,RIaef2338_3003,RIaef23b0_3004,RIaef2428_3005,RIaef24a0_3006,RIaef2518_3007,RIaef2590_3008,RIaef2608_3009,
        RIaef2680_3010,RIaef26f8_3011,RIaef2770_3012,RIaef27e8_3013,RIaef2860_3014,RIaef28d8_3015,RIaef2950_3016,RIaef29c8_3017,RIaef2a40_3018,RIaef2ab8_3019,
        RIaef2b30_3020,RIaef2ba8_3021,RIaef2c20_3022,RIaef2c98_3023,RIaef2d10_3024,RIaef2d88_3025,RIaef2e00_3026,RIaef2e78_3027,RIaef2ef0_3028,RIaef2f68_3029,
        RIaef2fe0_3030,RIaef3058_3031,RIaef30d0_3032,RIaef3148_3033,RIaef31c0_3034,RIaef3238_3035,RIaef32b0_3036,RIaef3328_3037,RIaef33a0_3038,RIaef3418_3039,
        RIaef3490_3040,RIaef3508_3041,RIaef3580_3042,RIaef35f8_3043,RIaef3670_3044,RIaef36e8_3045,RIaef3760_3046,RIaef37d8_3047,RIaef3850_3048,RIaef38c8_3049,
        RIaef3940_3050,RIaef39b8_3051,RIaef3a30_3052,RIaef3aa8_3053,RIaef3b20_3054,RIaef3b98_3055,RIaef3c10_3056,RIaef3c88_3057,RIaef3d00_3058,RIaef3d78_3059,
        RIaef3df0_3060,RIaef3e68_3061,RIaef3ee0_3062,RIaef3f58_3063,RIaef3fd0_3064,RIaef4048_3065,RIaef40c0_3066,RIaef4138_3067,RIaef41b0_3068,RIaef4228_3069,
        RIaef42a0_3070,RIaef4318_3071,RIaef4390_3072,RIaef4408_3073,RIaef4480_3074,RIaef44f8_3075,RIaef4570_3076,RIaef45e8_3077,RIaef4660_3078,RIaef46d8_3079,
        RIaef4750_3080,RIaef47c8_3081,RIaef4840_3082,RIaef48b8_3083,RIaef4930_3084,RIaef49a8_3085,RIaef4a20_3086,RIaef4a98_3087,RIaef4b10_3088,RIaef4b88_3089,
        RIaef4c00_3090,RIaef4c78_3091,RIaef4cf0_3092,RIaef4d68_3093,RIaef4de0_3094,RIaef4e58_3095,RIaef4ed0_3096,RIaef4f48_3097,RIaef4fc0_3098,RIaef5038_3099,
        RIaef50b0_3100,RIaef5128_3101,RIaef51a0_3102,RIaef5218_3103,RIaef5290_3104,RIaef5308_3105,RIaef5380_3106,RIaef53f8_3107,RIaef5470_3108,RIaef54e8_3109,
        RIaef5560_3110,RIaef55d8_3111,RIaef5650_3112,RIaef56c8_3113,RIaef5740_3114,RIaef57b8_3115,RIaef5830_3116,RIaef58a8_3117,RIaef5920_3118,RIaef5998_3119,
        RIaef5a10_3120,RIaef5a88_3121,RIaef5b00_3122,RIaef5b78_3123,RIaef5bf0_3124,RIaef5c68_3125,RIaef5ce0_3126,RIaef5d58_3127,RIaef5dd0_3128,RIaef5e48_3129,
        RIaef5ec0_3130,RIaef5f38_3131,RIaef5fb0_3132,RIaef6028_3133,RIaef60a0_3134,RIaef6118_3135,RIaef6190_3136,RIaef6208_3137,RIaef6280_3138,RIaef62f8_3139,
        RIaef6370_3140,RIaef63e8_3141,RIaef6460_3142,RIaef64d8_3143,RIaef6550_3144,RIaef65c8_3145,RIaef6640_3146,RIaef66b8_3147,RIaef6730_3148,RIaef67a8_3149,
        RIaef6820_3150,RIaef6898_3151,RIaef6910_3152,RIaef6988_3153,RIaef6a00_3154,RIaef6a78_3155,RIaef6af0_3156,RIaef6b68_3157,RIaef6be0_3158,RIaef6c58_3159,
        RIaef6cd0_3160,RIaef6d48_3161,RIaef6dc0_3162,RIaef6e38_3163,RIaef6eb0_3164,RIaef6f28_3165,RIaef6fa0_3166,RIaef7018_3167,RIaef7090_3168,RIaef7108_3169,
        RIaef7180_3170,RIaef71f8_3171,RIaef7270_3172,RIaef72e8_3173,RIaef7360_3174,RIaef73d8_3175,RIaef7450_3176,RIaef74c8_3177,RIaef7540_3178,RIaef75b8_3179,
        RIaef7630_3180,RIaef76a8_3181,RIaef7720_3182,RIaef7798_3183,RIaef7810_3184,RIaef7888_3185,RIaef7900_3186,RIaef7978_3187,RIaef79f0_3188,RIaef7a68_3189,
        RIaef7ae0_3190,RIaef7b58_3191,RIaef7bd0_3192,RIaef7c48_3193,RIaef7cc0_3194,RIaef7d38_3195,RIaef7db0_3196,RIaef7e28_3197,RIaef7ea0_3198,RIaef7f18_3199,
        RIaef7f90_3200,RIaef8008_3201,RIaef8080_3202,RIaef80f8_3203,RIaef8170_3204,RIaef81e8_3205,RIaef8260_3206,RIaef82d8_3207,RIaef8350_3208,RIaef83c8_3209,
        RIaef8440_3210,RIaef84b8_3211,RIaef8530_3212,RIaef85a8_3213,RIaef8620_3214,RIaef8698_3215,RIaef8710_3216,RIaef8788_3217,RIaef8800_3218,RIaef8878_3219,
        RIaef88f0_3220,RIaef8968_3221,RIaef89e0_3222,RIaef8a58_3223,RIaef8ad0_3224,RIaef8b48_3225,RIaef8bc0_3226,RIaef8c38_3227,RIaef8cb0_3228,RIaef8d28_3229,
        RIaef8da0_3230,RIaef8e18_3231,RIaef8e90_3232,RIaef8f08_3233,RIaef8f80_3234,RIaef8ff8_3235,RIaef9070_3236,RIaef90e8_3237,RIaef9160_3238,RIaef91d8_3239,
        RIaef9250_3240,RIaef92c8_3241,RIaef9340_3242,RIaef93b8_3243,RIaef9430_3244,RIaef94a8_3245,RIaef9520_3246,RIaef9598_3247,RIaef9610_3248,RIaef9688_3249,
        RIaef9700_3250,RIaef9778_3251,RIaef97f0_3252,RIaef9868_3253,RIaef98e0_3254,RIaef9958_3255,RIaef99d0_3256,RIaef9a48_3257,RIaef9ac0_3258,RIaef9b38_3259,
        RIaef9bb0_3260,RIaef9c28_3261,RIaef9ca0_3262,RIaef9d18_3263,RIaef9d90_3264,RIaef9e08_3265,RIaef9e80_3266,RIaef9ef8_3267,RIaef9f70_3268,RIaef9fe8_3269,
        RIaefa060_3270,RIaefa0d8_3271,RIaefa150_3272,RIaefa1c8_3273,RIaefa240_3274,RIaefa2b8_3275,RIaefa330_3276,RIaefa3a8_3277,RIaefa420_3278,RIaefa498_3279,
        RIaefa510_3280,RIaefa588_3281,RIaefa600_3282,RIaefa678_3283,RIaefa6f0_3284,RIaefa768_3285,RIaefa7e0_3286,RIaefa858_3287,RIaefa8d0_3288,RIaefa948_3289,
        RIaefa9c0_3290,RIaefaa38_3291,RIaefaab0_3292,RIaefab28_3293,RIaefaba0_3294,RIaefac18_3295,RIaefac90_3296,RIaefad08_3297,RIaefad80_3298,RIaefadf8_3299,
        RIaefae70_3300,RIaefaee8_3301,RIaefaf60_3302,RIaefafd8_3303,RIaefb050_3304,RIaefb0c8_3305,RIaefb140_3306,RIaefb1b8_3307,RIaefb230_3308,RIaefb2a8_3309,
        RIaefb320_3310,RIaefb398_3311,RIaefb410_3312,RIaefb488_3313,RIaefb500_3314,RIaefb578_3315,RIaefb5f0_3316,RIaefb668_3317,RIaefb6e0_3318,RIaefb758_3319,
        RIaefb7d0_3320,RIaefb848_3321,RIaefb8c0_3322,RIaefb938_3323,RIaefb9b0_3324,RIaefba28_3325,RIaefbaa0_3326,RIaefbb18_3327,RIaefbb90_3328,RIaefbc08_3329,
        RIaefbc80_3330,RIaefbcf8_3331,RIaefbd70_3332,RIaefbde8_3333,RIaefbe60_3334,RIaefbed8_3335,RIaefbf50_3336,RIaefbfc8_3337,RIaefc040_3338,RIaefc0b8_3339,
        RIaefc130_3340,RIaefc1a8_3341,RIaefc220_3342,RIaefc298_3343,RIaefc310_3344,RIaefc388_3345,RIaefc400_3346,RIaefc478_3347,RIaefc4f0_3348,RIaefc568_3349,
        RIaefc5e0_3350,RIaefc658_3351,RIaefc6d0_3352,RIaefc748_3353,RIaefc7c0_3354,RIaefc838_3355,RIaefc8b0_3356,RIaefc928_3357,RIaefc9a0_3358,RIaefca18_3359,
        RIaefca90_3360,RIaefcb08_3361,RIaefcb80_3362,RIaefcbf8_3363,RIaefcc70_3364,RIaefcce8_3365,RIaefcd60_3366,RIaefcdd8_3367,RIaefce50_3368,RIaefcec8_3369,
        RIaefcf40_3370,RIaefcfb8_3371,RIaefd030_3372,RIaefd0a8_3373,RIaefd120_3374,RIaefd198_3375,RIaefd210_3376,RIaefd288_3377,RIaefd300_3378,RIaefd378_3379,
        RIaefd3f0_3380,RIaefd468_3381,RIaefd4e0_3382,RIaefd558_3383,RIaefd5d0_3384,RIaefd648_3385,RIaefd6c0_3386,RIaefd738_3387,RIaefd7b0_3388,RIaefd828_3389,
        RIaefd8a0_3390,RIaefd918_3391,RIaefd990_3392,RIaefda08_3393,RIaefda80_3394,RIaefdaf8_3395,RIaefdb70_3396,RIaefdbe8_3397,RIaefdc60_3398,RIaefdcd8_3399,
        RIaefdd50_3400,RIaefddc8_3401,RIaefde40_3402,RIaefdeb8_3403,RIaefdf30_3404,RIaefdfa8_3405,RIaefe020_3406,RIaefe098_3407,RIaefe110_3408,RIaefe188_3409,
        RIaefe200_3410,RIaefe278_3411,RIaefe2f0_3412,RIaefe368_3413,RIaefe3e0_3414,RIaefe458_3415,RIaefe4d0_3416,RIaefe548_3417,RIaefe5c0_3418,RIaefe638_3419,
        RIaefe6b0_3420,RIaefe728_3421,RIaefe7a0_3422,RIaefe818_3423,RIaefe890_3424,RIaefe908_3425,RIaefe980_3426,RIaefe9f8_3427,RIaefea70_3428,RIaefeae8_3429,
        RIaefeb60_3430,RIaefebd8_3431,RIaefec50_3432,RIaefecc8_3433,RIaefed40_3434,RIaefedb8_3435,RIaefee30_3436,RIaefeea8_3437,RIaefef20_3438,RIaefef98_3439,
        RIaeff010_3440,RIaeff088_3441,RIaeff100_3442,RIaeff178_3443,RIaeff1f0_3444,RIaeff268_3445,RIaeff2e0_3446,RIaeff358_3447,RIaeff3d0_3448,RIaeff448_3449,
        RIaeff4c0_3450,RIaeff538_3451,RIaeff5b0_3452,RIaeff628_3453,RIaeff6a0_3454,RIaeff718_3455,RIaeff790_3456,RIaeff808_3457,RIaeff880_3458,RIaeff8f8_3459,
        RIaeff970_3460,RIaeff9e8_3461,RIaeffa60_3462,RIaeffad8_3463,RIaeffb50_3464,RIaeffbc8_3465,RIaeffc40_3466,RIaeffcb8_3467,RIaeffd30_3468,RIaeffda8_3469,
        RIaeffe20_3470,RIaeffe98_3471,RIaefff10_3472,RIaefff88_3473,RIaf00000_3474,RIaf00078_3475,RIaf000f0_3476,RIaf00168_3477,RIaf001e0_3478,RIaf00258_3479,
        RIaf002d0_3480,RIaf00348_3481,RIaf003c0_3482,RIaf00438_3483,RIaf004b0_3484,RIaf00528_3485,RIaf005a0_3486,RIaf00618_3487,RIaf00690_3488,RIaf00708_3489,
        RIaf00780_3490,RIaf007f8_3491,RIaf00870_3492,RIaf008e8_3493,RIaf00960_3494,RIaf009d8_3495,RIaf00a50_3496,RIaf00ac8_3497,RIaf00b40_3498,RIaf00bb8_3499,
        RIaf00c30_3500,RIaf00ca8_3501,RIaf00d20_3502,RIaf00d98_3503,RIaf00e10_3504,RIaf00e88_3505,RIaf00f00_3506,RIaf00f78_3507,RIaf00ff0_3508,RIaf01068_3509,
        RIaf010e0_3510,RIaf01158_3511,RIaf011d0_3512,RIaf01248_3513,RIaf012c0_3514,RIaf01338_3515,RIaf013b0_3516,RIaf01428_3517,RIaf014a0_3518,RIaf01518_3519,
        RIaf01590_3520,RIaf01608_3521,RIaf01680_3522,RIaf016f8_3523,RIaf01770_3524,RIaf017e8_3525,RIaf01860_3526,RIaf018d8_3527,RIaf01950_3528,RIaf019c8_3529,
        RIaf01a40_3530,RIaf01ab8_3531,RIaf01b30_3532,RIaf01ba8_3533,RIaf01c20_3534,RIaf01c98_3535,RIaf01d10_3536,RIaf01d88_3537,RIaf01e00_3538,RIaf01e78_3539,
        RIaf01ef0_3540,RIaf01f68_3541,RIaf01fe0_3542,RIaf02058_3543,RIaf020d0_3544,RIaf02148_3545,RIaf021c0_3546,RIaf02238_3547,RIaf022b0_3548,RIaf02328_3549,
        RIaf023a0_3550,RIaf02418_3551,RIaf02490_3552,RIaf02508_3553,RIaf02580_3554,RIaf025f8_3555,RIaf02670_3556,RIaf026e8_3557,RIaf02760_3558,RIaf027d8_3559,
        RIaf02850_3560,RIaf028c8_3561,RIaf02940_3562,RIaf029b8_3563,RIaf02a30_3564,RIaf02aa8_3565,RIaf02b20_3566,RIaf02b98_3567,RIaf02c10_3568,RIaf02c88_3569,
        RIaf02d00_3570,RIaf02d78_3571,RIaf02df0_3572,RIaf02e68_3573,RIaf02ee0_3574,RIaf02f58_3575,RIaf02fd0_3576,RIaf03048_3577,RIaf030c0_3578,RIaf03138_3579,
        RIaf031b0_3580,RIaf03228_3581,RIaf032a0_3582,RIaf03318_3583,RIaf03390_3584,RIaf03408_3585,RIaf03480_3586,RIaf034f8_3587,RIaf03570_3588,RIaf035e8_3589,
        RIaf03660_3590,RIaf036d8_3591,RIaf03750_3592,RIaf037c8_3593,RIaf03840_3594,RIaf038b8_3595,RIaf03930_3596,RIaf039a8_3597,RIaf03a20_3598,RIaf03a98_3599,
        RIaf03b10_3600,RIaf03b88_3601,RIaf03c00_3602,RIaf03c78_3603,RIaf03cf0_3604,RIaf03d68_3605,RIaf03de0_3606,RIaf03e58_3607,RIaf03ed0_3608,RIaf03f48_3609,
        RIaf03fc0_3610,RIaf04038_3611,RIaf040b0_3612,RIaf04128_3613,RIaf041a0_3614,RIaf04218_3615,RIaf04290_3616,RIaf04308_3617,RIaf04380_3618,RIaf043f8_3619,
        RIaf04470_3620,RIaf044e8_3621,RIaf04560_3622,RIaf045d8_3623,RIaf04650_3624,RIaf046c8_3625,RIaf04740_3626,RIaf047b8_3627,RIaf04830_3628,RIaf048a8_3629,
        RIaf04920_3630,RIaf04998_3631,RIaf04a10_3632,RIaf04a88_3633,RIaf04b00_3634,RIaf04b78_3635,RIaf04bf0_3636,RIaf04c68_3637,RIaf04ce0_3638,RIaf04d58_3639,
        RIaf04dd0_3640,RIaf04e48_3641,RIaf04ec0_3642,RIaf04f38_3643,RIaf04fb0_3644,RIaf05028_3645,RIaf050a0_3646,RIaf05118_3647,RIaf05190_3648,RIaf05208_3649,
        RIaf05280_3650,RIaf052f8_3651,RIaf05370_3652,RIaf053e8_3653,RIaf05460_3654,RIaf054d8_3655,RIaf05550_3656,RIaf055c8_3657,RIaf05640_3658,RIaf056b8_3659,
        RIaf05730_3660,RIaf057a8_3661,RIaf05820_3662,RIaf05898_3663,RIaf05910_3664,RIaf05988_3665,RIaf05a00_3666,RIaf05a78_3667,RIaf05af0_3668,RIaf05b68_3669,
        RIaf05be0_3670,RIaf05c58_3671,RIaf05cd0_3672,RIaf05d48_3673,RIaf05dc0_3674,RIaf05e38_3675,RIaf05eb0_3676,RIaf05f28_3677,RIaf05fa0_3678,RIaf06018_3679,
        RIaf06090_3680,RIaf06108_3681,RIaf06180_3682,RIaf061f8_3683,RIaf06270_3684,RIaf062e8_3685,RIaf06360_3686,RIaf063d8_3687,RIaf06450_3688,RIaf064c8_3689,
        RIaf06540_3690,RIaf065b8_3691,RIaf06630_3692,RIaf066a8_3693,RIaf06720_3694,RIaf06798_3695,RIaf06810_3696,RIaf06888_3697,RIaf06900_3698,RIaf06978_3699,
        RIaf069f0_3700,RIaf06a68_3701,RIaf06ae0_3702,RIaf06b58_3703,RIaf06bd0_3704,RIaf06c48_3705,RIaf06cc0_3706,RIaf06d38_3707,RIaf06db0_3708,RIaf06e28_3709,
        RIaf06ea0_3710,RIaf06f18_3711,RIaf06f90_3712,RIaf07008_3713,RIaf07080_3714,RIaf070f8_3715,RIaf07170_3716,RIaf071e8_3717,RIaf07260_3718,RIaf072d8_3719,
        RIaf07350_3720,RIaf073c8_3721,RIaf07440_3722,RIaf074b8_3723,RIaf07530_3724,RIaf075a8_3725,RIaf07620_3726,RIaf07698_3727,RIaf07710_3728,RIaf07788_3729,
        RIaf07800_3730,RIaf07878_3731,RIaf078f0_3732,RIaf07968_3733,RIaf079e0_3734,RIaf07a58_3735,RIaf07ad0_3736,RIaf07b48_3737,RIaf07bc0_3738,RIaf07c38_3739,
        RIaf07cb0_3740,RIaf07d28_3741,RIaf07da0_3742,RIaf07e18_3743,RIaf07e90_3744,RIaf07f08_3745,RIaf07f80_3746,RIaf07ff8_3747,RIaf08070_3748,RIaf080e8_3749,
        RIaf08160_3750,RIaf081d8_3751,RIaf08250_3752,RIaf082c8_3753,RIaf08340_3754,RIaf083b8_3755,RIaf08430_3756,RIaf084a8_3757,RIaf08520_3758,RIaf08598_3759,
        RIaf08610_3760,RIaf08688_3761,RIaf08700_3762,RIaf08778_3763,RIaf087f0_3764,RIaf08868_3765,RIaf088e0_3766,RIaf08958_3767,RIaf089d0_3768,RIaf08a48_3769,
        RIaf08ac0_3770,RIaf08b38_3771,RIaf08bb0_3772,RIaf08c28_3773,RIaf08ca0_3774,RIaf08d18_3775,RIaf08d90_3776,RIaf08e08_3777,RIaf08e80_3778,RIaf08ef8_3779,
        RIaf08f70_3780,RIaf08fe8_3781,RIaf09060_3782,RIaf090d8_3783,RIaf09150_3784,RIaf091c8_3785,RIaf09240_3786,RIaf092b8_3787,RIaf09330_3788,RIaf093a8_3789,
        RIaf09420_3790,RIaf09498_3791,RIaf09510_3792,RIaf09588_3793,RIaf09600_3794,RIaf09678_3795,RIaf096f0_3796,RIaf09768_3797,RIaf097e0_3798,RIaf09858_3799,
        RIaf098d0_3800,RIaf09948_3801,RIaf099c0_3802,RIaf09a38_3803,RIaf09ab0_3804,RIaf09b28_3805,RIaf09ba0_3806,RIaf09c18_3807,RIaf09c90_3808,RIaf09d08_3809,
        RIaf09d80_3810,RIaf09df8_3811,RIaf09e70_3812,RIaf09ee8_3813,RIaf09f60_3814,RIaf09fd8_3815,RIaf0a050_3816,RIaf0a0c8_3817,RIaf0a140_3818,RIaf0a1b8_3819,
        RIaf0a230_3820,RIaf0a2a8_3821,RIaf0a320_3822,RIaf0a398_3823,RIaf0a410_3824,RIaf0a488_3825,RIaf0a500_3826,RIaf0a578_3827,RIaf0a5f0_3828,RIaf0a668_3829,
        RIaf0a6e0_3830,RIaf0a758_3831,RIaf0a7d0_3832,RIaf0a848_3833,RIaf0a8c0_3834,RIaf0a938_3835,RIaf0a9b0_3836,RIaf0aa28_3837,RIaf0aaa0_3838,RIaf0ab18_3839,
        RIaf0ab90_3840,RIaf0ac08_3841,RIaf0ac80_3842,RIaf0acf8_3843,RIaf0ad70_3844,RIaf0ade8_3845,RIaf0ae60_3846,RIaf0aed8_3847,RIaf0af50_3848,RIaf0afc8_3849,
        RIaf0b040_3850,RIaf0b0b8_3851,RIaf0b130_3852,RIaf0b1a8_3853,RIaf0b220_3854,RIaf0b298_3855,RIaf0b310_3856,RIaf0b388_3857,RIaf0b400_3858,RIaf0b478_3859,
        RIaf0b4f0_3860,RIaf0b568_3861,RIaf0b5e0_3862,RIaf0b658_3863,RIaf0b6d0_3864,RIaf0b748_3865,RIaf0b7c0_3866,RIaf0b838_3867,RIaf0b8b0_3868,RIaf0b928_3869,
        RIaf0b9a0_3870,RIaf0ba18_3871,RIaf0ba90_3872,RIaf0bb08_3873,RIaf0bb80_3874,RIaf0bbf8_3875,RIaf0bc70_3876,RIaf0bce8_3877,RIaf0bd60_3878,RIaf0bdd8_3879,
        RIaf0be50_3880,RIaf0bec8_3881,RIaf0bf40_3882,RIaf0bfb8_3883,RIaf0c030_3884,RIaf0c0a8_3885,RIaf0c120_3886,RIaf0c198_3887,RIaf0c210_3888,RIaf0c288_3889,
        RIaf0c300_3890,RIaf0c378_3891,RIaf0c3f0_3892,RIaf0c468_3893,RIaf0c4e0_3894,RIaf0c558_3895,RIaf0c5d0_3896,RIaf0c648_3897,RIaf0c6c0_3898,RIaf0c738_3899,
        RIaf0c7b0_3900,RIaf0c828_3901,RIaf0c8a0_3902,RIaf0c918_3903,RIaf0c990_3904,RIaf0ca08_3905,RIaf0ca80_3906,RIaf0caf8_3907,RIaf0cb70_3908,RIaf0cbe8_3909,
        RIaf0cc60_3910,RIaf0ccd8_3911,RIaf0cd50_3912,RIaf0cdc8_3913,RIaf0ce40_3914,RIaf0ceb8_3915,RIaf0cf30_3916,RIaf0cfa8_3917,RIaf0d020_3918,RIaf0d098_3919,
        RIaf0d110_3920,RIaf0d188_3921,RIaf0d200_3922,RIaf0d278_3923,RIaf0d2f0_3924,RIaf0d368_3925,RIaf0d3e0_3926,RIaf0d458_3927,RIaf0d4d0_3928,RIaf0d548_3929,
        RIaf0d5c0_3930,RIaf0d638_3931,RIaf0d6b0_3932,RIaf0d728_3933,RIaf0d7a0_3934,RIaf0d818_3935,RIaf0d890_3936,RIaf0d908_3937,RIaf0d980_3938,RIaf0d9f8_3939,
        RIaf0da70_3940,RIaf0dae8_3941,RIaf0db60_3942,RIaf0dbd8_3943,RIaf0dc50_3944,RIaf0dcc8_3945,RIaf0dd40_3946,RIaf0ddb8_3947,RIaf0de30_3948,RIaf0dea8_3949,
        RIaf0df20_3950,RIaf0df98_3951,RIaf0e010_3952,RIaf0e088_3953,RIaf0e100_3954,RIaf0e178_3955,RIaf0e1f0_3956,RIaf0e268_3957,RIaf0e2e0_3958,RIaf0e358_3959,
        RIaf0e3d0_3960,RIaf0e448_3961,RIaf0e4c0_3962,RIaf0e538_3963,RIaf0e5b0_3964,RIaf0e628_3965,RIaf0e6a0_3966,RIaf0e718_3967,RIaf0e790_3968,RIaf0e808_3969,
        RIaf0e880_3970,RIaf0e8f8_3971,RIaf0e970_3972,RIaf0e9e8_3973,RIaf0ea60_3974,RIaf0ead8_3975,RIaf0eb50_3976,RIaf0ebc8_3977,RIaf0ec40_3978,RIaf0ecb8_3979,
        RIaf0ed30_3980,RIaf0eda8_3981,RIaf0ee20_3982,RIaf0ee98_3983,RIaf0ef10_3984,RIaf0ef88_3985,RIaf0f000_3986,RIaf0f078_3987,RIaf0f0f0_3988,RIaf0f168_3989,
        RIaf0f1e0_3990,RIaf0f258_3991,RIaf0f2d0_3992,RIaf0f348_3993,RIaf0f3c0_3994,RIaf0f438_3995,RIaf0f4b0_3996,RIaf0f528_3997,RIaf0f5a0_3998,RIaf0f618_3999,
        RIaf0f690_4000,RIaf0f708_4001,RIaf0f780_4002,RIaf0f7f8_4003,RIaf0f870_4004,RIaf0f8e8_4005,RIaf0f960_4006,RIaf0f9d8_4007,RIaf0fa50_4008,RIaf0fac8_4009,
        RIaf0fb40_4010,RIaf0fbb8_4011,RIaf0fc30_4012,RIaf0fca8_4013,RIaf0fd20_4014,RIaf0fd98_4015,RIaf0fe10_4016,RIaf0fe88_4017,RIaf0ff00_4018,RIaf0ff78_4019,
        RIaf0fff0_4020,RIaf10068_4021,RIaf100e0_4022,RIaf10158_4023,RIaf101d0_4024,RIaf10248_4025,RIaf102c0_4026,RIaf10338_4027,RIaf103b0_4028,RIaf10428_4029,
        RIaf104a0_4030,RIaf10518_4031,RIaf10590_4032,RIaf10608_4033,RIaf10680_4034,RIaf106f8_4035,RIaf10770_4036,RIaf107e8_4037,RIaf10860_4038,RIaf108d8_4039,
        RIaf10950_4040,RIaf109c8_4041,RIaf10a40_4042,RIaf10ab8_4043,RIaf10b30_4044,RIaf10ba8_4045,RIaf10c20_4046,RIaf10c98_4047,RIaf10d10_4048,RIaf10d88_4049,
        RIaf10e00_4050,RIaf10e78_4051,RIaf10ef0_4052,RIaf10f68_4053,RIaf10fe0_4054,RIaf11058_4055,RIaf110d0_4056,RIaf11148_4057,RIaf111c0_4058,RIaf11238_4059,
        RIaf112b0_4060,RIaf11328_4061,RIaf113a0_4062,RIaf11418_4063,RIaf11490_4064,RIaf11508_4065,RIaf11580_4066,RIaf115f8_4067,RIaf11670_4068,RIaf116e8_4069,
        RIaf11760_4070,RIaf117d8_4071,RIaf11850_4072,RIaf118c8_4073,RIaf11940_4074,RIaf119b8_4075,RIaf11a30_4076,RIaf11aa8_4077,RIaf11b20_4078,RIaf11b98_4079,
        RIaf11c10_4080,RIaf11c88_4081,RIaf11d00_4082,RIaf11d78_4083,RIaf11df0_4084,RIaf11e68_4085,RIaf11ee0_4086,RIaf11f58_4087,RIaf11fd0_4088,RIaf12048_4089,
        RIaf120c0_4090,RIaf12138_4091,RIaf121b0_4092,RIaf12228_4093,RIaf122a0_4094,RIaf12318_4095,RIaf12390_4096,RIaf12408_4097,RIaf12480_4098,RIaf124f8_4099,
        RIaf12570_4100,RIaf125e8_4101,RIaf12660_4102,RIaf126d8_4103,RIaf12750_4104,RIaf127c8_4105,RIaf12840_4106,RIaf128b8_4107,RIaf12930_4108,RIaf129a8_4109,
        RIaf12a20_4110,RIaf12a98_4111,RIaf12b10_4112,RIaf12b88_4113,RIaf12c00_4114,RIaf12c78_4115,RIaf12cf0_4116,RIaf12d68_4117,RIaf12de0_4118,RIaf12e58_4119,
        RIaf12ed0_4120,RIaf12f48_4121,RIaf12fc0_4122,RIaf13038_4123,RIaf130b0_4124,RIaf13128_4125,RIaf131a0_4126,RIaf13218_4127,RIaf13290_4128,RIaf13308_4129,
        RIaf13380_4130,RIaf133f8_4131,RIaf13470_4132,RIaf134e8_4133,RIaf13560_4134,RIaf135d8_4135,RIaf13650_4136,RIaf136c8_4137,RIaf13740_4138,RIaf137b8_4139,
        RIaf13830_4140,RIaf138a8_4141,RIaf13920_4142,RIaf13998_4143,RIaf13a10_4144,RIaf13a88_4145,RIaf13b00_4146,RIaf13b78_4147,RIaf13bf0_4148,RIaf13c68_4149,
        RIaf13ce0_4150,RIaf13d58_4151,RIaf13dd0_4152,RIaf13e48_4153,RIaf13ec0_4154,RIaf13f38_4155,RIaf13fb0_4156,RIaf14028_4157,RIaf140a0_4158,RIaf14118_4159,
        RIaf14190_4160,RIaf14208_4161,RIaf14280_4162,RIaf142f8_4163,RIaf14370_4164,RIaf143e8_4165,RIaf14460_4166,RIaf144d8_4167,RIaf14550_4168,RIaf145c8_4169,
        RIaf14640_4170,RIaf146b8_4171,RIaf14730_4172,RIaf147a8_4173,RIaf14820_4174,RIaf14898_4175,RIaf14910_4176,RIaf14988_4177,RIaf14a00_4178,RIaf14a78_4179,
        RIaf14af0_4180,RIaf14b68_4181,RIaf14be0_4182,RIaf14c58_4183,RIaf14cd0_4184,RIaf14d48_4185,RIaf14dc0_4186,RIaf14e38_4187,RIaf14eb0_4188,RIaf14f28_4189,
        RIaf14fa0_4190,RIaf15018_4191,RIaf15090_4192,RIaf15108_4193,RIaf15180_4194,RIaf151f8_4195,RIaf15270_4196,RIaf152e8_4197,RIaf15360_4198,RIaf153d8_4199,
        RIaf15450_4200,RIaf154c8_4201,RIaf15540_4202,RIaf155b8_4203,RIaf15630_4204,RIaf156a8_4205,RIaf15720_4206,RIaf15798_4207,RIaf15810_4208,RIaf15888_4209,
        RIaf15900_4210,RIaf15978_4211,RIaf159f0_4212,RIaf15a68_4213,RIaf15ae0_4214,RIaf15b58_4215,RIaf15bd0_4216,RIaf15c48_4217,RIaf15cc0_4218,RIaf15d38_4219,
        RIaf15db0_4220,RIaf15e28_4221,RIaf15ea0_4222,RIaf15f18_4223,RIaf15f90_4224,RIaf16008_4225,RIaf16080_4226,RIaf160f8_4227,RIaf16170_4228,RIaf161e8_4229,
        RIaf16260_4230,RIaf162d8_4231,RIaf16350_4232,RIaf163c8_4233,RIaf16440_4234,RIaf164b8_4235,RIaf16530_4236,RIaf165a8_4237,RIaf16620_4238,RIaf16698_4239,
        RIaf16710_4240,RIaf16788_4241,RIaf16800_4242,RIaf16878_4243,RIaf168f0_4244,RIaf16968_4245,RIaf169e0_4246,RIaf16a58_4247,RIaf16ad0_4248,RIaf16b48_4249,
        RIaf16bc0_4250,RIaf16c38_4251,RIaf16cb0_4252,RIaf16d28_4253,RIaf16da0_4254,RIaf16e18_4255,RIaf16e90_4256,RIaf16f08_4257,RIaf16f80_4258,RIaf16ff8_4259,
        RIaf17070_4260,RIaf170e8_4261,RIaf17160_4262,RIaf171d8_4263,RIaf17250_4264,RIaf172c8_4265,RIaf17340_4266,RIaf173b8_4267,RIaf17430_4268,RIaf174a8_4269,
        RIaf17520_4270,RIaf17598_4271,RIaf17610_4272,RIaf17688_4273,RIaf17700_4274,RIaf17778_4275,RIaf177f0_4276,RIaf17868_4277,RIaf178e0_4278,RIaf17958_4279,
        RIaf179d0_4280,RIaf17a48_4281,RIaf17ac0_4282,RIaf17b38_4283,RIaf17bb0_4284,RIaf17c28_4285,RIaf17ca0_4286,RIaf17d18_4287,RIaf17d90_4288,RIaf17e08_4289,
        RIaf17e80_4290,RIaf17ef8_4291,RIaf17f70_4292,RIaf17fe8_4293,RIaf18060_4294,RIaf180d8_4295,RIaf18150_4296,RIaf181c8_4297,RIaf18240_4298,RIaf182b8_4299,
        RIaf18330_4300,RIaf183a8_4301,RIaf18420_4302,RIaf18498_4303,RIaf18510_4304,RIaf18588_4305,RIaf18600_4306,RIaf18678_4307,RIaf186f0_4308,RIaf18768_4309,
        RIaf187e0_4310,RIaf18858_4311,RIaf188d0_4312,RIaf18948_4313,RIaf189c0_4314,RIaf18a38_4315,RIaf18ab0_4316,RIaf18b28_4317,RIaf18ba0_4318,RIaf18c18_4319,
        RIaf18c90_4320,RIaf18d08_4321,RIaf18d80_4322,RIaf18df8_4323,RIaf18e70_4324,RIaf18ee8_4325,RIaf18f60_4326,RIaf18fd8_4327,RIaf19050_4328,RIaf190c8_4329,
        RIaf19140_4330,RIaf191b8_4331,RIaf19230_4332,RIaf192a8_4333,RIaf19320_4334,RIaf19398_4335,RIaf19410_4336,RIaf19488_4337,RIaf19500_4338,RIaf19578_4339,
        RIaf195f0_4340,RIaf19668_4341,RIaf196e0_4342,RIaf19758_4343,RIaf197d0_4344,RIaf19848_4345,RIaf198c0_4346,RIaf19938_4347,RIaf199b0_4348,RIaf19a28_4349,
        RIaf19aa0_4350,RIaf19b18_4351,RIaf19b90_4352,RIaf19c08_4353,RIaf19c80_4354,RIaf19cf8_4355,RIaf19d70_4356,RIaf19de8_4357,RIaf19e60_4358,RIaf19ed8_4359,
        RIaf19f50_4360,RIaf19fc8_4361,RIaf1a040_4362,RIaf1a0b8_4363,RIaf1a130_4364,RIaf1a1a8_4365,RIaf1a220_4366,RIaf1a298_4367,RIaf1a310_4368,RIaf1a388_4369,
        RIaf1a400_4370,RIaf1a478_4371,RIaf1a4f0_4372,RIaf1a568_4373,RIaf1a5e0_4374,RIaf1a658_4375,RIaf1a6d0_4376,RIaf1a748_4377,RIaf1a7c0_4378,RIaf1a838_4379,
        RIaf1a8b0_4380,RIaf1a928_4381,RIaf1a9a0_4382,RIaf1aa18_4383,RIaf1aa90_4384,RIaf1ab08_4385,RIaf1ab80_4386,RIaf1abf8_4387,RIaf1ac70_4388,RIaf1ace8_4389,
        RIaf1ad60_4390,RIaf1add8_4391,RIaf1ae50_4392,RIaf1aec8_4393,RIaf1af40_4394,RIaf1afb8_4395,RIaf1b030_4396,RIaf1b0a8_4397,RIaf1b120_4398,RIaf1b198_4399,
        RIaf1b210_4400,RIaf1b288_4401,RIaf1b300_4402,RIaf1b378_4403,RIaf1b3f0_4404,RIaf1b468_4405,RIaf1b4e0_4406,RIaf1b558_4407,RIaf1b5d0_4408,RIaf1b648_4409,
        RIaf1b6c0_4410,RIaf1b738_4411,RIaf1b7b0_4412,RIaf1b828_4413,RIaf1b8a0_4414,RIaf1b918_4415,RIaf1b990_4416,RIaf1ba08_4417,RIaf1ba80_4418,RIaf1baf8_4419,
        RIaf1bb70_4420,RIaf1bbe8_4421,RIaf1bc60_4422,RIaf1bcd8_4423,RIaf1bd50_4424,RIaf1bdc8_4425,RIaf1be40_4426,RIaf1beb8_4427,RIaf1bf30_4428,RIaf1bfa8_4429,
        RIaf1c020_4430,RIaf1c098_4431,RIaf1c110_4432,RIaf1c188_4433,RIaf1c200_4434,RIaf1c278_4435,RIaf1c2f0_4436,RIaf1c368_4437,RIaf1c3e0_4438,RIaf1c458_4439,
        RIaf1c4d0_4440,RIaf1c548_4441,RIaf1c5c0_4442,RIaf1c638_4443,RIaf1c6b0_4444,RIaf1c728_4445,RIaf1c7a0_4446,RIaf1c818_4447,RIaf1c890_4448,RIaf1c908_4449,
        RIaf1c980_4450,RIaf1c9f8_4451,RIaf1ca70_4452,RIaf1cae8_4453,RIaf1cb60_4454,RIaf1cbd8_4455,RIaf1cc50_4456,RIaf1ccc8_4457,RIaf1cd40_4458,RIaf1cdb8_4459,
        RIaf1ce30_4460,RIaf1cea8_4461,RIaf1cf20_4462,RIaf1cf98_4463,RIaf1d010_4464,RIaf1d088_4465,RIaf1d100_4466,RIaf1d178_4467,RIaf1d1f0_4468,RIaf1d268_4469,
        RIaf1d2e0_4470,RIaf1d358_4471,RIaf1d3d0_4472,RIaf1d448_4473,RIaf1d4c0_4474,RIaf1d538_4475,RIaf1d5b0_4476,RIaf1d628_4477,RIaf1d6a0_4478,RIaf1d718_4479,
        RIaf1d790_4480,RIaf1d808_4481,RIaf1d880_4482,RIaf1d8f8_4483,RIaf1d970_4484,RIaf1d9e8_4485,RIaf1da60_4486,RIaf1dad8_4487,RIaf1db50_4488,RIaf1dbc8_4489,
        RIaf1dc40_4490,RIaf1dcb8_4491,RIaf1dd30_4492,RIaf1dda8_4493,RIaf1de20_4494,RIaf1de98_4495,RIaf1df10_4496,RIaf1df88_4497,RIaf1e000_4498,RIaf1e078_4499,
        RIaf1e0f0_4500,RIaf1e168_4501,RIaf1e1e0_4502,RIaf1e258_4503,RIaf1e2d0_4504,RIaf1e348_4505,RIaf1e3c0_4506,RIaf1e438_4507,RIaf1e4b0_4508,RIaf1e528_4509,
        RIaf1e5a0_4510,RIaf1e618_4511,RIaf1e690_4512,RIaf1e708_4513,RIaf1e780_4514,RIaf1e7f8_4515,RIaf1e870_4516,RIaf1e8e8_4517,RIaf1e960_4518,RIaf1e9d8_4519,
        RIaf1ea50_4520,RIaf1eac8_4521,RIaf1eb40_4522,RIaf1ebb8_4523,RIaf1ec30_4524,RIaf1eca8_4525,RIaf1ed20_4526,RIaf1ed98_4527,RIaf1ee10_4528,RIaf1ee88_4529,
        RIaf1ef00_4530,RIaf1ef78_4531,RIaf1eff0_4532,RIaf1f068_4533,RIaf1f0e0_4534,RIaf1f158_4535,RIaf1f1d0_4536,RIaf1f248_4537,RIaf1f2c0_4538,RIaf1f338_4539,
        RIaf1f3b0_4540,RIaf1f428_4541,RIaf1f4a0_4542,RIaf1f518_4543,RIaf1f590_4544,RIaf1f608_4545,RIaf1f680_4546,RIaf1f6f8_4547,RIaf1f770_4548,RIaf1f7e8_4549,
        RIaf1f860_4550,RIaf1f8d8_4551,RIaf1f950_4552,RIaf1f9c8_4553,RIaf1fa40_4554,RIaf1fab8_4555,RIaf1fb30_4556,RIaf1fba8_4557,RIaf1fc20_4558,RIaf1fc98_4559,
        RIaf1fd10_4560,RIaf1fd88_4561,RIaf1fe00_4562,RIaf1fe78_4563,RIaf1fef0_4564,RIaf1ff68_4565,RIaf1ffe0_4566,RIaf20058_4567,RIaf200d0_4568,RIaf20148_4569,
        RIaf201c0_4570,RIaf20238_4571,RIaf202b0_4572,RIaf20328_4573,RIaf203a0_4574,RIaf20418_4575,RIaf20490_4576,RIaf20508_4577,RIaf20580_4578,RIaf205f8_4579,
        RIaf20670_4580,RIaf206e8_4581,RIaf20760_4582,RIaf207d8_4583,RIaf20850_4584,RIaf208c8_4585,RIaf20940_4586,RIaf209b8_4587,RIaf20a30_4588,RIaf20aa8_4589,
        RIaf20b20_4590,RIaf20b98_4591,RIaf20c10_4592,RIaf20c88_4593,RIaf20d00_4594,RIaf20d78_4595,RIaf20df0_4596,RIaf20e68_4597,RIaf20ee0_4598,RIaf20f58_4599,
        RIaf20fd0_4600,RIaf21048_4601,RIaf210c0_4602,RIaf21138_4603,RIaf211b0_4604,RIaf21228_4605,RIaf212a0_4606,RIaf21318_4607,RIaf21390_4608,RIaf21408_4609,
        RIaf21480_4610,RIaf214f8_4611,RIaf21570_4612,RIaf215e8_4613,RIaf21660_4614,RIaf216d8_4615,RIaf21750_4616,RIaf217c8_4617,RIaf21840_4618,RIaf218b8_4619,
        RIaf21930_4620,RIaf219a8_4621,RIaf21a20_4622,RIaf21a98_4623,RIaf21b10_4624,RIaf21b88_4625,RIaf21c00_4626,RIaf21c78_4627,RIaf21cf0_4628,RIaf21d68_4629,
        RIaf21de0_4630,RIaf21e58_4631,RIaf21ed0_4632,RIaf21f48_4633,RIaf21fc0_4634,RIaf22038_4635,RIaf220b0_4636,RIaf22128_4637,RIaf221a0_4638,RIaf22218_4639,
        RIaf22290_4640,RIaf22308_4641,RIaf22380_4642,RIaf223f8_4643,RIaf22470_4644,RIaf224e8_4645,RIaf22560_4646,RIaf225d8_4647,RIaf22650_4648,RIaf226c8_4649,
        RIaf22740_4650,RIaf227b8_4651,RIaf22830_4652,RIaf228a8_4653,RIaf22920_4654,RIaf22998_4655,RIaf22a10_4656,RIaf22a88_4657,RIaf22b00_4658,RIaf22b78_4659,
        RIaf22bf0_4660,RIaf22c68_4661,RIaf22ce0_4662,RIaf22d58_4663,RIaf22dd0_4664,RIaf22e48_4665,RIaf22ec0_4666,RIaf22f38_4667,RIaf22fb0_4668,RIaf23028_4669,
        RIaf230a0_4670,RIaf23118_4671,RIaf23190_4672,RIaf23208_4673,RIaf23280_4674,RIaf232f8_4675,RIaf23370_4676,RIaf233e8_4677,RIaf23460_4678,RIaf234d8_4679,
        RIaf23550_4680;
output R_1249_9a72be0,R_124a_9a72c88,R_124b_9a72d30,R_124c_9a72dd8,R_124d_9a72e80,R_124e_9a72f28,R_124f_9a72fd0,R_1250_9a73078,R_1251_9a73120;

wire \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 ,
         \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706_N$1 , \4707_N$2 , \4708_N$3 ,
         \4709_N$4 , \4710_N$5 , \4711_N$6 , \4712_N$7 , \4713_N$8 , \4714_ZERO , \4715_ONE , \4716 , \4717 , \4718 ,
         \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 ,
         \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 ,
         \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 ,
         \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 ,
         \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 ,
         \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 ,
         \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 ,
         \4789 , \4790 , \4791 , \4792 ;
buf \U$labajz955 ( R_1249_9a72be0, \4792 );
buf \U$labajz956 ( R_124a_9a72c88, 1'b0 );
buf \U$labajz957 ( R_124b_9a72d30, 1'b0 );
buf \U$labajz958 ( R_124c_9a72dd8, 1'b0 );
buf \U$labajz959 ( R_124d_9a72e80, 1'b0 );
buf \U$labajz960 ( R_124e_9a72f28, 1'b0 );
buf \U$labajz961 ( R_124f_9a72fd0, 1'b0 );
buf \U$labajz962 ( R_1250_9a73078, 1'b0 );
buf \U$labajz963 ( R_1251_9a73120, 1'b0 );
and \U$1 ( \4716 , RIae9a408_1, RIae9a480_2, RIae9a4f8_3, RIae9a570_4, RIae9a5e8_5, RIae9a660_6, RIae9a6d8_7, RIae9a750_8, RIae9a7c8_9, RIae9a840_10, RIae9a8b8_11, RIae9a930_12, RIae9a9a8_13, RIae9aa20_14, RIae9aa98_15, RIae9ab10_16, RIae9ab88_17, RIae9ac00_18, RIae9ac78_19, RIae9acf0_20, RIae9ad68_21, RIae9ade0_22, RIae9ae58_23, RIae9aed0_24, RIae9af48_25, RIae9afc0_26, RIae9b038_27, RIae9b0b0_28, RIae9b128_29, RIae9b1a0_30, RIae9b218_31, RIae9b290_32, RIae9b308_33, RIae9b380_34, RIae9b3f8_35, RIae9b470_36, RIae9b4e8_37, RIae9b560_38, RIae9b5d8_39, RIae9b650_40, RIae9b6c8_41, RIae9b740_42, RIae9b7b8_43, RIae9b830_44, RIae9b8a8_45, RIae9b920_46, RIae9b998_47, RIae9ba10_48, RIae9ba88_49, RIae9bb00_50, RIae9bb78_51, RIae9bbf0_52, RIae9bc68_53, RIae9bce0_54, RIae9bd58_55, RIae9bdd0_56, RIae9be48_57, RIae9bec0_58, RIae9bf38_59, RIae9bfb0_60, RIae9c028_61, RIae9c0a0_62, RIae9c118_63, RIae9c190_64);
and \U$2 ( \4717 , RIae9c208_65, RIae9c280_66, RIae9c2f8_67, RIae9c370_68, RIae9c3e8_69, RIae9c460_70, RIae9c4d8_71, RIae9c550_72, RIae9c5c8_73, RIae9c640_74, RIae9c6b8_75, RIae9c730_76, RIae9c7a8_77, RIae9c820_78, RIae9c898_79, RIae9c910_80, RIae9c988_81, RIae9ca00_82, RIae9ca78_83, RIae9caf0_84, RIae9cb68_85, RIae9cbe0_86, RIae9cc58_87, RIae9ccd0_88, RIae9cd48_89, RIae9cdc0_90, RIae9ce38_91, RIae9ceb0_92, RIae9cf28_93, RIae9cfa0_94, RIae9d018_95, RIae9d090_96, RIae9d108_97, RIae9d180_98, RIae9d1f8_99, RIae9d270_100, RIae9d2e8_101, RIae9d360_102, RIae9d3d8_103, RIae9d450_104, RIae9d4c8_105, RIae9d540_106, RIae9d5b8_107, RIae9d630_108, RIae9d6a8_109, RIae9d720_110, RIae9d798_111, RIae9d810_112, RIae9d888_113, RIae9d900_114, RIae9d978_115, RIae9d9f0_116, RIae9da68_117, RIae9dae0_118, RIae9db58_119, RIae9dbd0_120, RIae9dc48_121, RIae9dcc0_122, RIae9dd38_123, RIae9ddb0_124, RIae9de28_125, RIae9dea0_126, RIae9df18_127, RIae9df90_128);
and \U$3 ( \4718 , RIae9e008_129, RIae9e080_130, RIae9e0f8_131, RIae9e170_132, RIae9e1e8_133, RIae9e260_134, RIae9e2d8_135, RIae9e350_136, RIae9e3c8_137, RIae9e440_138, RIae9e4b8_139, RIae9e530_140, RIae9e5a8_141, RIae9e620_142, RIae9e698_143, RIae9e710_144, RIae9e788_145, RIae9e800_146, RIae9e878_147, RIae9e8f0_148, RIae9e968_149, RIae9e9e0_150, RIae9ea58_151, RIae9ead0_152, RIae9eb48_153, RIae9ebc0_154, RIae9ec38_155, RIae9ecb0_156, RIae9ed28_157, RIae9eda0_158, RIae9ee18_159, RIae9ee90_160, RIae9ef08_161, RIae9ef80_162, RIae9eff8_163, RIae9f070_164, RIae9f0e8_165, RIae9f160_166, RIae9f1d8_167, RIae9f250_168, RIae9f2c8_169, RIae9f340_170, RIae9f3b8_171, RIae9f430_172, RIae9f4a8_173, RIae9f520_174, RIae9f598_175, RIae9f610_176, RIae9f688_177, RIae9f700_178, RIae9f778_179, RIae9f7f0_180, RIae9f868_181, RIae9f8e0_182, RIae9f958_183, RIae9f9d0_184, RIae9fa48_185, RIae9fac0_186, RIae9fb38_187, RIae9fbb0_188, RIae9fc28_189, RIae9fca0_190, RIae9fd18_191, RIae9fd90_192);
and \U$4 ( \4719 , RIae9fe08_193, RIae9fe80_194, RIae9fef8_195, RIae9ff70_196, RIae9ffe8_197, RIaea0060_198, RIaea00d8_199, RIaea0150_200, RIaea01c8_201, RIaea0240_202, RIaea02b8_203, RIaea0330_204, RIaea03a8_205, RIaea0420_206, RIaea0498_207, RIaea0510_208, RIaea0588_209, RIaea0600_210, RIaea0678_211, RIaea06f0_212, RIaea0768_213, RIaea07e0_214, RIaea0858_215, RIaea08d0_216, RIaea0948_217, RIaea09c0_218, RIaea0a38_219, RIaea0ab0_220, RIaea0b28_221, RIaea0ba0_222, RIaea0c18_223, RIaea0c90_224, RIaea0d08_225, RIaea0d80_226, RIaea0df8_227, RIaea0e70_228, RIaea0ee8_229, RIaea0f60_230, RIaea0fd8_231, RIaea1050_232, RIaea10c8_233, RIaea1140_234, RIaea11b8_235, RIaea1230_236, RIaea12a8_237, RIaea1320_238, RIaea1398_239, RIaea1410_240, RIaea1488_241, RIaea1500_242, RIaea1578_243, RIaea15f0_244, RIaea1668_245, RIaea16e0_246, RIaea1758_247, RIaea17d0_248, RIaea1848_249, RIaea18c0_250, RIaea1938_251, RIaea19b0_252, RIaea1a28_253, RIaea1aa0_254, RIaea1b18_255, RIaea1b90_256);
and \U$5 ( \4720 , RIaea1c08_257, RIaea1c80_258, RIaea1cf8_259, RIaea1d70_260, RIaea1de8_261, RIaea1e60_262, RIaea1ed8_263, RIaea1f50_264, RIaea1fc8_265, RIaea2040_266, RIaea20b8_267, RIaea2130_268, RIaea21a8_269, RIaea2220_270, RIaea2298_271, RIaea2310_272, RIaea2388_273, RIaea2400_274, RIaea2478_275, RIaea24f0_276, RIaea2568_277, RIaea25e0_278, RIaea2658_279, RIaea26d0_280, RIaea2748_281, RIaea27c0_282, RIaea2838_283, RIaea28b0_284, RIaea2928_285, RIaea29a0_286, RIaea2a18_287, RIaea2a90_288, RIaea2b08_289, RIaea2b80_290, RIaea2bf8_291, RIaea2c70_292, RIaea2ce8_293, RIaea2d60_294, RIaea2dd8_295, RIaea2e50_296, RIaea2ec8_297, RIaea2f40_298, RIaea2fb8_299, RIaea3030_300, RIaea30a8_301, RIaea3120_302, RIaea3198_303, RIaea3210_304, RIaea3288_305, RIaea3300_306, RIaea3378_307, RIaea33f0_308, RIaea3468_309, RIaea34e0_310, RIaea3558_311, RIaea35d0_312, RIaea3648_313, RIaea36c0_314, RIaea3738_315, RIaea37b0_316, RIaea3828_317, RIaea38a0_318, RIaea3918_319, RIaea3990_320);
and \U$6 ( \4721 , RIaea3a08_321, RIaea3a80_322, RIaea3af8_323, RIaea3b70_324, RIaea3be8_325, RIaea3c60_326, RIaea3cd8_327, RIaea3d50_328, RIaea3dc8_329, RIaea3e40_330, RIaea3eb8_331, RIaea3f30_332, RIaea3fa8_333, RIaea4020_334, RIaea4098_335, RIaea4110_336, RIaea4188_337, RIaea4200_338, RIaea4278_339, RIaea42f0_340, RIaea4368_341, RIaea43e0_342, RIaea4458_343, RIaea44d0_344, RIaea4548_345, RIaea45c0_346, RIaea4638_347, RIaea46b0_348, RIaea4728_349, RIaea47a0_350, RIaea4818_351, RIaea4890_352, RIaea4908_353, RIaea4980_354, RIaea49f8_355, RIaea4a70_356, RIaea4ae8_357, RIaea4b60_358, RIaea4bd8_359, RIaea4c50_360, RIaea4cc8_361, RIaea4d40_362, RIaea4db8_363, RIaea4e30_364, RIaea4ea8_365, RIaea4f20_366, RIaea4f98_367, RIaea5010_368, RIaea5088_369, RIaea5100_370, RIaea5178_371, RIaea51f0_372, RIaea5268_373, RIaea52e0_374, RIaea5358_375, RIaea53d0_376, RIaea5448_377, RIaea54c0_378, RIaea5538_379, RIaea55b0_380, RIaea5628_381, RIaea56a0_382, RIaea5718_383, RIaea5790_384);
and \U$7 ( \4722 , RIaea5808_385, RIaea5880_386, RIaea58f8_387, RIaea5970_388, RIaea59e8_389, RIaea5a60_390, RIaea5ad8_391, RIaea5b50_392, RIaea5bc8_393, RIaea5c40_394, RIaea5cb8_395, RIaea5d30_396, RIaea5da8_397, RIaea5e20_398, RIaea5e98_399, RIaea5f10_400, RIaea5f88_401, RIaea6000_402, RIaea6078_403, RIaea60f0_404, RIaea6168_405, RIaea61e0_406, RIaea6258_407, RIaea62d0_408, RIaea6348_409, RIaea63c0_410, RIaea6438_411, RIaea64b0_412, RIaea6528_413, RIaea65a0_414, RIaea6618_415, RIaea6690_416, RIaea6708_417, RIaea6780_418, RIaea67f8_419, RIaea6870_420, RIaea68e8_421, RIaea6960_422, RIaea69d8_423, RIaea6a50_424, RIaea6ac8_425, RIaea6b40_426, RIaea6bb8_427, RIaea6c30_428, RIaea6ca8_429, RIaea6d20_430, RIaea6d98_431, RIaea6e10_432, RIaea6e88_433, RIaea6f00_434, RIaea6f78_435, RIaea6ff0_436, RIaea7068_437, RIaea70e0_438, RIaea7158_439, RIaea71d0_440, RIaea7248_441, RIaea72c0_442, RIaea7338_443, RIaea73b0_444, RIaea7428_445, RIaea74a0_446, RIaea7518_447, RIaea7590_448);
and \U$8 ( \4723 , RIaea7608_449, RIaea7680_450, RIaea76f8_451, RIaea7770_452, RIaea77e8_453, RIaea7860_454, RIaea78d8_455, RIaea7950_456, RIaea79c8_457, RIaea7a40_458, RIaea7ab8_459, RIaea7b30_460, RIaea7ba8_461, RIaea7c20_462, RIaea7c98_463, RIaea7d10_464, RIaea7d88_465, RIaea7e00_466, RIaea7e78_467, RIaea7ef0_468, RIaea7f68_469, RIaea7fe0_470, RIaea8058_471, RIaea80d0_472, RIaea8148_473, RIaea81c0_474, RIaea8238_475, RIaea82b0_476, RIaea8328_477, RIaea83a0_478, RIaea8418_479, RIaea8490_480, RIaea8508_481, RIaea8580_482, RIaea85f8_483, RIaea8670_484, RIaea86e8_485, RIaea8760_486, RIaea87d8_487, RIaea8850_488, RIaea88c8_489, RIaea8940_490, RIaea89b8_491, RIaea8a30_492, RIaea8aa8_493, RIaea8b20_494, RIaea8b98_495, RIaea8c10_496, RIaea8c88_497, RIaea8d00_498, RIaea8d78_499, RIaea8df0_500, RIaea8e68_501, RIaea8ee0_502, RIaea8f58_503, RIaea8fd0_504, RIaea9048_505, RIaea90c0_506, RIaea9138_507, RIaea91b0_508, RIaea9228_509, RIaea92a0_510, RIaea9318_511, RIaea9390_512);
and \U$9 ( \4724 , RIaea9408_513, RIaea9480_514, RIaea94f8_515, RIaea9570_516, RIaea95e8_517, RIaea9660_518, RIaea96d8_519, RIaea9750_520, RIaea97c8_521, RIaea9840_522, RIaea98b8_523, RIaea9930_524, RIaea99a8_525, RIaea9a20_526, RIaea9a98_527, RIaea9b10_528, RIaea9b88_529, RIaea9c00_530, RIaea9c78_531, RIaea9cf0_532, RIaea9d68_533, RIaea9de0_534, RIaea9e58_535, RIaea9ed0_536, RIaea9f48_537, RIaea9fc0_538, RIaeaa038_539, RIaeaa0b0_540, RIaeaa128_541, RIaeaa1a0_542, RIaeaa218_543, RIaeaa290_544, RIaeaa308_545, RIaeaa380_546, RIaeaa3f8_547, RIaeaa470_548, RIaeaa4e8_549, RIaeaa560_550, RIaeaa5d8_551, RIaeaa650_552, RIaeaa6c8_553, RIaeaa740_554, RIaeaa7b8_555, RIaeaa830_556, RIaeaa8a8_557, RIaeaa920_558, RIaeaa998_559, RIaeaaa10_560, RIaeaaa88_561, RIaeaab00_562, RIaeaab78_563, RIaeaabf0_564, RIaeaac68_565, RIaeaace0_566, RIaeaad58_567, RIaeaadd0_568, RIaeaae48_569, RIaeaaec0_570, RIaeaaf38_571, RIaeaafb0_572, RIaeab028_573, RIaeab0a0_574, RIaeab118_575, RIaeab190_576);
and \U$10 ( \4725 , RIaeab208_577, RIaeab280_578, RIaeab2f8_579, RIaeab370_580, RIaeab3e8_581, RIaeab460_582, RIaeab4d8_583, RIaeab550_584, RIaeab5c8_585, RIaeab640_586, RIaeab6b8_587, RIaeab730_588, RIaeab7a8_589, RIaeab820_590, RIaeab898_591, RIaeab910_592, RIaeab988_593, RIaeaba00_594, RIaeaba78_595, RIaeabaf0_596, RIaeabb68_597, RIaeabbe0_598, RIaeabc58_599, RIaeabcd0_600, RIaeabd48_601, RIaeabdc0_602, RIaeabe38_603, RIaeabeb0_604, RIaeabf28_605, RIaeabfa0_606, RIaeac018_607, RIaeac090_608, RIaeac108_609, RIaeac180_610, RIaeac1f8_611, RIaeac270_612, RIaeac2e8_613, RIaeac360_614, RIaeac3d8_615, RIaeac450_616, RIaeac4c8_617, RIaeac540_618, RIaeac5b8_619, RIaeac630_620, RIaeac6a8_621, RIaeac720_622, RIaeac798_623, RIaeac810_624, RIaeac888_625, RIaeac900_626, RIaeac978_627, RIaeac9f0_628, RIaeaca68_629, RIaeacae0_630, RIaeacb58_631, RIaeacbd0_632, RIaeacc48_633, RIaeaccc0_634, RIaeacd38_635, RIaeacdb0_636, RIaeace28_637, RIaeacea0_638, RIaeacf18_639, RIaeacf90_640);
and \U$11 ( \4726 , RIaead008_641, RIaead080_642, RIaead0f8_643, RIaead170_644, RIaead1e8_645, RIaead260_646, RIaead2d8_647, RIaead350_648, RIaead3c8_649, RIaead440_650, RIaead4b8_651, RIaead530_652, RIaead5a8_653, RIaead620_654, RIaead698_655, RIaead710_656, RIaead788_657, RIaead800_658, RIaead878_659, RIaead8f0_660, RIaead968_661, RIaead9e0_662, RIaeada58_663, RIaeadad0_664, RIaeadb48_665, RIaeadbc0_666, RIaeadc38_667, RIaeadcb0_668, RIaeadd28_669, RIaeadda0_670, RIaeade18_671, RIaeade90_672, RIaeadf08_673, RIaeadf80_674, RIaeadff8_675, RIaeae070_676, RIaeae0e8_677, RIaeae160_678, RIaeae1d8_679, RIaeae250_680, RIaeae2c8_681, RIaeae340_682, RIaeae3b8_683, RIaeae430_684, RIaeae4a8_685, RIaeae520_686, RIaeae598_687, RIaeae610_688, RIaeae688_689, RIaeae700_690, RIaeae778_691, RIaeae7f0_692, RIaeae868_693, RIaeae8e0_694, RIaeae958_695, RIaeae9d0_696, RIaeaea48_697, RIaeaeac0_698, RIaeaeb38_699, RIaeaebb0_700, RIaeaec28_701, RIaeaeca0_702, RIaeaed18_703, RIaeaed90_704);
and \U$12 ( \4727 , RIaeaee08_705, RIaeaee80_706, RIaeaeef8_707, RIaeaef70_708, RIaeaefe8_709, RIaeaf060_710, RIaeaf0d8_711, RIaeaf150_712, RIaeaf1c8_713, RIaeaf240_714, RIaeaf2b8_715, RIaeaf330_716, RIaeaf3a8_717, RIaeaf420_718, RIaeaf498_719, RIaeaf510_720, RIaeaf588_721, RIaeaf600_722, RIaeaf678_723, RIaeaf6f0_724, RIaeaf768_725, RIaeaf7e0_726, RIaeaf858_727, RIaeaf8d0_728, RIaeaf948_729, RIaeaf9c0_730, RIaeafa38_731, RIaeafab0_732, RIaeafb28_733, RIaeafba0_734, RIaeafc18_735, RIaeafc90_736, RIaeafd08_737, RIaeafd80_738, RIaeafdf8_739, RIaeafe70_740, RIaeafee8_741, RIaeaff60_742, RIaeaffd8_743, RIaeb0050_744, RIaeb00c8_745, RIaeb0140_746, RIaeb01b8_747, RIaeb0230_748, RIaeb02a8_749, RIaeb0320_750, RIaeb0398_751, RIaeb0410_752, RIaeb0488_753, RIaeb0500_754, RIaeb0578_755, RIaeb05f0_756, RIaeb0668_757, RIaeb06e0_758, RIaeb0758_759, RIaeb07d0_760, RIaeb0848_761, RIaeb08c0_762, RIaeb0938_763, RIaeb09b0_764, RIaeb0a28_765, RIaeb0aa0_766, RIaeb0b18_767, RIaeb0b90_768);
and \U$13 ( \4728 , RIaeb0c08_769, RIaeb0c80_770, RIaeb0cf8_771, RIaeb0d70_772, RIaeb0de8_773, RIaeb0e60_774, RIaeb0ed8_775, RIaeb0f50_776, RIaeb0fc8_777, RIaeb1040_778, RIaeb10b8_779, RIaeb1130_780, RIaeb11a8_781, RIaeb1220_782, RIaeb1298_783, RIaeb1310_784, RIaeb1388_785, RIaeb1400_786, RIaeb1478_787, RIaeb14f0_788, RIaeb1568_789, RIaeb15e0_790, RIaeb1658_791, RIaeb16d0_792, RIaeb1748_793, RIaeb17c0_794, RIaeb1838_795, RIaeb18b0_796, RIaeb1928_797, RIaeb19a0_798, RIaeb1a18_799, RIaeb1a90_800, RIaeb1b08_801, RIaeb1b80_802, RIaeb1bf8_803, RIaeb1c70_804, RIaeb1ce8_805, RIaeb1d60_806, RIaeb1dd8_807, RIaeb1e50_808, RIaeb1ec8_809, RIaeb1f40_810, RIaeb1fb8_811, RIaeb2030_812, RIaeb20a8_813, RIaeb2120_814, RIaeb2198_815, RIaeb2210_816, RIaeb2288_817, RIaeb2300_818, RIaeb2378_819, RIaeb23f0_820, RIaeb2468_821, RIaeb24e0_822, RIaeb2558_823, RIaeb25d0_824, RIaeb2648_825, RIaeb26c0_826, RIaeb2738_827, RIaeb27b0_828, RIaeb2828_829, RIaeb28a0_830, RIaeb2918_831, RIaeb2990_832);
and \U$14 ( \4729 , RIaeb2a08_833, RIaeb2a80_834, RIaeb2af8_835, RIaeb2b70_836, RIaeb2be8_837, RIaeb2c60_838, RIaeb2cd8_839, RIaeb2d50_840, RIaeb2dc8_841, RIaeb2e40_842, RIaeb2eb8_843, RIaeb2f30_844, RIaeb2fa8_845, RIaeb3020_846, RIaeb3098_847, RIaeb3110_848, RIaeb3188_849, RIaeb3200_850, RIaeb3278_851, RIaeb32f0_852, RIaeb3368_853, RIaeb33e0_854, RIaeb3458_855, RIaeb34d0_856, RIaeb3548_857, RIaeb35c0_858, RIaeb3638_859, RIaeb36b0_860, RIaeb3728_861, RIaeb37a0_862, RIaeb3818_863, RIaeb3890_864, RIaeb3908_865, RIaeb3980_866, RIaeb39f8_867, RIaeb3a70_868, RIaeb3ae8_869, RIaeb3b60_870, RIaeb3bd8_871, RIaeb3c50_872, RIaeb3cc8_873, RIaeb3d40_874, RIaeb3db8_875, RIaeb3e30_876, RIaeb3ea8_877, RIaeb3f20_878, RIaeb3f98_879, RIaeb4010_880, RIaeb4088_881, RIaeb4100_882, RIaeb4178_883, RIaeb41f0_884, RIaeb4268_885, RIaeb42e0_886, RIaeb4358_887, RIaeb43d0_888, RIaeb4448_889, RIaeb44c0_890, RIaeb4538_891, RIaeb45b0_892, RIaeb4628_893, RIaeb46a0_894, RIaeb4718_895, RIaeb4790_896);
and \U$15 ( \4730 , RIaeb4808_897, RIaeb4880_898, RIaeb48f8_899, RIaeb4970_900, RIaeb49e8_901, RIaeb4a60_902, RIaeb4ad8_903, RIaeb4b50_904, RIaeb4bc8_905, RIaeb4c40_906, RIaeb4cb8_907, RIaeb4d30_908, RIaeb4da8_909, RIaeb4e20_910, RIaeb4e98_911, RIaeb4f10_912, RIaeb4f88_913, RIaeb5000_914, RIaeb5078_915, RIaeb50f0_916, RIaeb5168_917, RIaeb51e0_918, RIaeb5258_919, RIaeb52d0_920, RIaeb5348_921, RIaeb53c0_922, RIaeb5438_923, RIaeb54b0_924, RIaeb5528_925, RIaeb55a0_926, RIaeb5618_927, RIaeb5690_928, RIaeb5708_929, RIaeb5780_930, RIaeb57f8_931, RIaeb5870_932, RIaeb58e8_933, RIaeb5960_934, RIaeb59d8_935, RIaeb5a50_936, RIaeb5ac8_937, RIaeb5b40_938, RIaeb5bb8_939, RIaeb5c30_940, RIaeb5ca8_941, RIaeb5d20_942, RIaeb5d98_943, RIaeb5e10_944, RIaeb5e88_945, RIaeb5f00_946, RIaeb5f78_947, RIaeb5ff0_948, RIaeb6068_949, RIaeb60e0_950, RIaeb6158_951, RIaeb61d0_952, RIaeb6248_953, RIaeb62c0_954, RIaeb6338_955, RIaeb63b0_956, RIaeb6428_957, RIaeb64a0_958, RIaeb6518_959, RIaeb6590_960);
and \U$16 ( \4731 , RIaeb6608_961, RIaeb6680_962, RIaeb66f8_963, RIaeb6770_964, RIaeb67e8_965, RIaeb6860_966, RIaeb68d8_967, RIaeb6950_968, RIaeb69c8_969, RIaeb6a40_970, RIaeb6ab8_971, RIaeb6b30_972, RIaeb6ba8_973, RIaeb6c20_974, RIaeb6c98_975, RIaeb6d10_976, RIaeb6d88_977, RIaeb6e00_978, RIaeb6e78_979, RIaeb6ef0_980, RIaeb6f68_981, RIaeb6fe0_982, RIaeb7058_983, RIaeb70d0_984, RIaeb7148_985, RIaeb71c0_986, RIaeb7238_987, RIaeb72b0_988, RIaeb7328_989, RIaeb73a0_990, RIaeb7418_991, RIaeb7490_992, RIaeb7508_993, RIaeb7580_994, RIaeb75f8_995, RIaeb7670_996, RIaeb76e8_997, RIaeb7760_998, RIaeb77d8_999, RIaeb7850_1000, RIaeb78c8_1001, RIaeb7940_1002, RIaeb79b8_1003, RIaeb7a30_1004, RIaeb7aa8_1005, RIaeb7b20_1006, RIaeb7b98_1007, RIaeb7c10_1008, RIaeb7c88_1009, RIaeb7d00_1010, RIaeb7d78_1011, RIaeb7df0_1012, RIaeb7e68_1013, RIaeb7ee0_1014, RIaeb7f58_1015, RIaeb7fd0_1016, RIaeb8048_1017, RIaeb80c0_1018, RIaeb8138_1019, RIaeb81b0_1020, RIaeb8228_1021, RIaeb82a0_1022, RIaeb8318_1023, RIaeb8390_1024);
and \U$17 ( \4732 , RIaeb8408_1025, RIaeb8480_1026, RIaeb84f8_1027, RIaeb8570_1028, RIaeb85e8_1029, RIaeb8660_1030, RIaeb86d8_1031, RIaeb8750_1032, RIaeb87c8_1033, RIaeb8840_1034, RIaeb88b8_1035, RIaeb8930_1036, RIaeb89a8_1037, RIaeb8a20_1038, RIaeb8a98_1039, RIaeb8b10_1040, RIaeb8b88_1041, RIaeb8c00_1042, RIaeb8c78_1043, RIaeb8cf0_1044, RIaeb8d68_1045, RIaeb8de0_1046, RIaeb8e58_1047, RIaeb8ed0_1048, RIaeb8f48_1049, RIaeb8fc0_1050, RIaeb9038_1051, RIaeb90b0_1052, RIaeb9128_1053, RIaeb91a0_1054, RIaeb9218_1055, RIaeb9290_1056, RIaeb9308_1057, RIaeb9380_1058, RIaeb93f8_1059, RIaeb9470_1060, RIaeb94e8_1061, RIaeb9560_1062, RIaeb95d8_1063, RIaeb9650_1064, RIaeb96c8_1065, RIaeb9740_1066, RIaeb97b8_1067, RIaeb9830_1068, RIaeb98a8_1069, RIaeb9920_1070, RIaeb9998_1071, RIaeb9a10_1072, RIaeb9a88_1073, RIaeb9b00_1074, RIaeb9b78_1075, RIaeb9bf0_1076, RIaeb9c68_1077, RIaeb9ce0_1078, RIaeb9d58_1079, RIaeb9dd0_1080, RIaeb9e48_1081, RIaeb9ec0_1082, RIaeb9f38_1083, RIaeb9fb0_1084, RIaeba028_1085, RIaeba0a0_1086, RIaeba118_1087, RIaeba190_1088);
and \U$18 ( \4733 , RIaeba208_1089, RIaeba280_1090, RIaeba2f8_1091, RIaeba370_1092, RIaeba3e8_1093, RIaeba460_1094, RIaeba4d8_1095, RIaeba550_1096, RIaeba5c8_1097, RIaeba640_1098, RIaeba6b8_1099, RIaeba730_1100, RIaeba7a8_1101, RIaeba820_1102, RIaeba898_1103, RIaeba910_1104, RIaeba988_1105, RIaebaa00_1106, RIaebaa78_1107, RIaebaaf0_1108, RIaebab68_1109, RIaebabe0_1110, RIaebac58_1111, RIaebacd0_1112, RIaebad48_1113, RIaebadc0_1114, RIaebae38_1115, RIaebaeb0_1116, RIaebaf28_1117, RIaebafa0_1118, RIaebb018_1119, RIaebb090_1120, RIaebb108_1121, RIaebb180_1122, RIaebb1f8_1123, RIaebb270_1124, RIaebb2e8_1125, RIaebb360_1126, RIaebb3d8_1127, RIaebb450_1128, RIaebb4c8_1129, RIaebb540_1130, RIaebb5b8_1131, RIaebb630_1132, RIaebb6a8_1133, RIaebb720_1134, RIaebb798_1135, RIaebb810_1136, RIaebb888_1137, RIaebb900_1138, RIaebb978_1139, RIaebb9f0_1140, RIaebba68_1141, RIaebbae0_1142, RIaebbb58_1143, RIaebbbd0_1144, RIaebbc48_1145, RIaebbcc0_1146, RIaebbd38_1147, RIaebbdb0_1148, RIaebbe28_1149, RIaebbea0_1150, RIaebbf18_1151, RIaebbf90_1152);
and \U$19 ( \4734 , RIaebc008_1153, RIaebc080_1154, RIaebc0f8_1155, RIaebc170_1156, RIaebc1e8_1157, RIaebc260_1158, RIaebc2d8_1159, RIaebc350_1160, RIaebc3c8_1161, RIaebc440_1162, RIaebc4b8_1163, RIaebc530_1164, RIaebc5a8_1165, RIaebc620_1166, RIaebc698_1167, RIaebc710_1168, RIaebc788_1169, RIaebc800_1170, RIaebc878_1171, RIaebc8f0_1172, RIaebc968_1173, RIaebc9e0_1174, RIaebca58_1175, RIaebcad0_1176, RIaebcb48_1177, RIaebcbc0_1178, RIaebcc38_1179, RIaebccb0_1180, RIaebcd28_1181, RIaebcda0_1182, RIaebce18_1183, RIaebce90_1184, RIaebcf08_1185, RIaebcf80_1186, RIaebcff8_1187, RIaebd070_1188, RIaebd0e8_1189, RIaebd160_1190, RIaebd1d8_1191, RIaebd250_1192, RIaebd2c8_1193, RIaebd340_1194, RIaebd3b8_1195, RIaebd430_1196, RIaebd4a8_1197, RIaebd520_1198, RIaebd598_1199, RIaebd610_1200, RIaebd688_1201, RIaebd700_1202, RIaebd778_1203, RIaebd7f0_1204, RIaebd868_1205, RIaebd8e0_1206, RIaebd958_1207, RIaebd9d0_1208, RIaebda48_1209, RIaebdac0_1210, RIaebdb38_1211, RIaebdbb0_1212, RIaebdc28_1213, RIaebdca0_1214, RIaebdd18_1215, RIaebdd90_1216);
and \U$20 ( \4735 , RIaebde08_1217, RIaebde80_1218, RIaebdef8_1219, RIaebdf70_1220, RIaebdfe8_1221, RIaebe060_1222, RIaebe0d8_1223, RIaebe150_1224, RIaebe1c8_1225, RIaebe240_1226, RIaebe2b8_1227, RIaebe330_1228, RIaebe3a8_1229, RIaebe420_1230, RIaebe498_1231, RIaebe510_1232, RIaebe588_1233, RIaebe600_1234, RIaebe678_1235, RIaebe6f0_1236, RIaebe768_1237, RIaebe7e0_1238, RIaebe858_1239, RIaebe8d0_1240, RIaebe948_1241, RIaebe9c0_1242, RIaebea38_1243, RIaebeab0_1244, RIaebeb28_1245, RIaebeba0_1246, RIaebec18_1247, RIaebec90_1248, RIaebed08_1249, RIaebed80_1250, RIaebedf8_1251, RIaebee70_1252, RIaebeee8_1253, RIaebef60_1254, RIaebefd8_1255, RIaebf050_1256, RIaebf0c8_1257, RIaebf140_1258, RIaebf1b8_1259, RIaebf230_1260, RIaebf2a8_1261, RIaebf320_1262, RIaebf398_1263, RIaebf410_1264, RIaebf488_1265, RIaebf500_1266, RIaebf578_1267, RIaebf5f0_1268, RIaebf668_1269, RIaebf6e0_1270, RIaebf758_1271, RIaebf7d0_1272, RIaebf848_1273, RIaebf8c0_1274, RIaebf938_1275, RIaebf9b0_1276, RIaebfa28_1277, RIaebfaa0_1278, RIaebfb18_1279, RIaebfb90_1280);
and \U$21 ( \4736 , RIaebfc08_1281, RIaebfc80_1282, RIaebfcf8_1283, RIaebfd70_1284, RIaebfde8_1285, RIaebfe60_1286, RIaebfed8_1287, RIaebff50_1288, RIaebffc8_1289, RIaec0040_1290, RIaec00b8_1291, RIaec0130_1292, RIaec01a8_1293, RIaec0220_1294, RIaec0298_1295, RIaec0310_1296, RIaec0388_1297, RIaec0400_1298, RIaec0478_1299, RIaec04f0_1300, RIaec0568_1301, RIaec05e0_1302, RIaec0658_1303, RIaec06d0_1304, RIaec0748_1305, RIaec07c0_1306, RIaec0838_1307, RIaec08b0_1308, RIaec0928_1309, RIaec09a0_1310, RIaec0a18_1311, RIaec0a90_1312, RIaec0b08_1313, RIaec0b80_1314, RIaec0bf8_1315, RIaec0c70_1316, RIaec0ce8_1317, RIaec0d60_1318, RIaec0dd8_1319, RIaec0e50_1320, RIaec0ec8_1321, RIaec0f40_1322, RIaec0fb8_1323, RIaec1030_1324, RIaec10a8_1325, RIaec1120_1326, RIaec1198_1327, RIaec1210_1328, RIaec1288_1329, RIaec1300_1330, RIaec1378_1331, RIaec13f0_1332, RIaec1468_1333, RIaec14e0_1334, RIaec1558_1335, RIaec15d0_1336, RIaec1648_1337, RIaec16c0_1338, RIaec1738_1339, RIaec17b0_1340, RIaec1828_1341, RIaec18a0_1342, RIaec1918_1343, RIaec1990_1344);
and \U$22 ( \4737 , RIaec1a08_1345, RIaec1a80_1346, RIaec1af8_1347, RIaec1b70_1348, RIaec1be8_1349, RIaec1c60_1350, RIaec1cd8_1351, RIaec1d50_1352, RIaec1dc8_1353, RIaec1e40_1354, RIaec1eb8_1355, RIaec1f30_1356, RIaec1fa8_1357, RIaec2020_1358, RIaec2098_1359, RIaec2110_1360, RIaec2188_1361, RIaec2200_1362, RIaec2278_1363, RIaec22f0_1364, RIaec2368_1365, RIaec23e0_1366, RIaec2458_1367, RIaec24d0_1368, RIaec2548_1369, RIaec25c0_1370, RIaec2638_1371, RIaec26b0_1372, RIaec2728_1373, RIaec27a0_1374, RIaec2818_1375, RIaec2890_1376, RIaec2908_1377, RIaec2980_1378, RIaec29f8_1379, RIaec2a70_1380, RIaec2ae8_1381, RIaec2b60_1382, RIaec2bd8_1383, RIaec2c50_1384, RIaec2cc8_1385, RIaec2d40_1386, RIaec2db8_1387, RIaec2e30_1388, RIaec2ea8_1389, RIaec2f20_1390, RIaec2f98_1391, RIaec3010_1392, RIaec3088_1393, RIaec3100_1394, RIaec3178_1395, RIaec31f0_1396, RIaec3268_1397, RIaec32e0_1398, RIaec3358_1399, RIaec33d0_1400, RIaec3448_1401, RIaec34c0_1402, RIaec3538_1403, RIaec35b0_1404, RIaec3628_1405, RIaec36a0_1406, RIaec3718_1407, RIaec3790_1408);
and \U$23 ( \4738 , RIaec3808_1409, RIaec3880_1410, RIaec38f8_1411, RIaec3970_1412, RIaec39e8_1413, RIaec3a60_1414, RIaec3ad8_1415, RIaec3b50_1416, RIaec3bc8_1417, RIaec3c40_1418, RIaec3cb8_1419, RIaec3d30_1420, RIaec3da8_1421, RIaec3e20_1422, RIaec3e98_1423, RIaec3f10_1424, RIaec3f88_1425, RIaec4000_1426, RIaec4078_1427, RIaec40f0_1428, RIaec4168_1429, RIaec41e0_1430, RIaec4258_1431, RIaec42d0_1432, RIaec4348_1433, RIaec43c0_1434, RIaec4438_1435, RIaec44b0_1436, RIaec4528_1437, RIaec45a0_1438, RIaec4618_1439, RIaec4690_1440, RIaec4708_1441, RIaec4780_1442, RIaec47f8_1443, RIaec4870_1444, RIaec48e8_1445, RIaec4960_1446, RIaec49d8_1447, RIaec4a50_1448, RIaec4ac8_1449, RIaec4b40_1450, RIaec4bb8_1451, RIaec4c30_1452, RIaec4ca8_1453, RIaec4d20_1454, RIaec4d98_1455, RIaec4e10_1456, RIaec4e88_1457, RIaec4f00_1458, RIaec4f78_1459, RIaec4ff0_1460, RIaec5068_1461, RIaec50e0_1462, RIaec5158_1463, RIaec51d0_1464, RIaec5248_1465, RIaec52c0_1466, RIaec5338_1467, RIaec53b0_1468, RIaec5428_1469, RIaec54a0_1470, RIaec5518_1471, RIaec5590_1472);
and \U$24 ( \4739 , RIaec5608_1473, RIaec5680_1474, RIaec56f8_1475, RIaec5770_1476, RIaec57e8_1477, RIaec5860_1478, RIaec58d8_1479, RIaec5950_1480, RIaec59c8_1481, RIaec5a40_1482, RIaec5ab8_1483, RIaec5b30_1484, RIaec5ba8_1485, RIaec5c20_1486, RIaec5c98_1487, RIaec5d10_1488, RIaec5d88_1489, RIaec5e00_1490, RIaec5e78_1491, RIaec5ef0_1492, RIaec5f68_1493, RIaec5fe0_1494, RIaec6058_1495, RIaec60d0_1496, RIaec6148_1497, RIaec61c0_1498, RIaec6238_1499, RIaec62b0_1500, RIaec6328_1501, RIaec63a0_1502, RIaec6418_1503, RIaec6490_1504, RIaec6508_1505, RIaec6580_1506, RIaec65f8_1507, RIaec6670_1508, RIaec66e8_1509, RIaec6760_1510, RIaec67d8_1511, RIaec6850_1512, RIaec68c8_1513, RIaec6940_1514, RIaec69b8_1515, RIaec6a30_1516, RIaec6aa8_1517, RIaec6b20_1518, RIaec6b98_1519, RIaec6c10_1520, RIaec6c88_1521, RIaec6d00_1522, RIaec6d78_1523, RIaec6df0_1524, RIaec6e68_1525, RIaec6ee0_1526, RIaec6f58_1527, RIaec6fd0_1528, RIaec7048_1529, RIaec70c0_1530, RIaec7138_1531, RIaec71b0_1532, RIaec7228_1533, RIaec72a0_1534, RIaec7318_1535, RIaec7390_1536);
and \U$25 ( \4740 , RIaec7408_1537, RIaec7480_1538, RIaec74f8_1539, RIaec7570_1540, RIaec75e8_1541, RIaec7660_1542, RIaec76d8_1543, RIaec7750_1544, RIaec77c8_1545, RIaec7840_1546, RIaec78b8_1547, RIaec7930_1548, RIaec79a8_1549, RIaec7a20_1550, RIaec7a98_1551, RIaec7b10_1552, RIaec7b88_1553, RIaec7c00_1554, RIaec7c78_1555, RIaec7cf0_1556, RIaec7d68_1557, RIaec7de0_1558, RIaec7e58_1559, RIaec7ed0_1560, RIaec7f48_1561, RIaec7fc0_1562, RIaec8038_1563, RIaec80b0_1564, RIaec8128_1565, RIaec81a0_1566, RIaec8218_1567, RIaec8290_1568, RIaec8308_1569, RIaec8380_1570, RIaec83f8_1571, RIaec8470_1572, RIaec84e8_1573, RIaec8560_1574, RIaec85d8_1575, RIaec8650_1576, RIaec86c8_1577, RIaec8740_1578, RIaec87b8_1579, RIaec8830_1580, RIaec88a8_1581, RIaec8920_1582, RIaec8998_1583, RIaec8a10_1584, RIaec8a88_1585, RIaec8b00_1586, RIaec8b78_1587, RIaec8bf0_1588, RIaec8c68_1589, RIaec8ce0_1590, RIaec8d58_1591, RIaec8dd0_1592, RIaec8e48_1593, RIaec8ec0_1594, RIaec8f38_1595, RIaec8fb0_1596, RIaec9028_1597, RIaec90a0_1598, RIaec9118_1599, RIaec9190_1600);
and \U$26 ( \4741 , RIaec9208_1601, RIaec9280_1602, RIaec92f8_1603, RIaec9370_1604, RIaec93e8_1605, RIaec9460_1606, RIaec94d8_1607, RIaec9550_1608, RIaec95c8_1609, RIaec9640_1610, RIaec96b8_1611, RIaec9730_1612, RIaec97a8_1613, RIaec9820_1614, RIaec9898_1615, RIaec9910_1616, RIaec9988_1617, RIaec9a00_1618, RIaec9a78_1619, RIaec9af0_1620, RIaec9b68_1621, RIaec9be0_1622, RIaec9c58_1623, RIaec9cd0_1624, RIaec9d48_1625, RIaec9dc0_1626, RIaec9e38_1627, RIaec9eb0_1628, RIaec9f28_1629, RIaec9fa0_1630, RIaeca018_1631, RIaeca090_1632, RIaeca108_1633, RIaeca180_1634, RIaeca1f8_1635, RIaeca270_1636, RIaeca2e8_1637, RIaeca360_1638, RIaeca3d8_1639, RIaeca450_1640, RIaeca4c8_1641, RIaeca540_1642, RIaeca5b8_1643, RIaeca630_1644, RIaeca6a8_1645, RIaeca720_1646, RIaeca798_1647, RIaeca810_1648, RIaeca888_1649, RIaeca900_1650, RIaeca978_1651, RIaeca9f0_1652, RIaecaa68_1653, RIaecaae0_1654, RIaecab58_1655, RIaecabd0_1656, RIaecac48_1657, RIaecacc0_1658, RIaecad38_1659, RIaecadb0_1660, RIaecae28_1661, RIaecaea0_1662, RIaecaf18_1663, RIaecaf90_1664);
and \U$27 ( \4742 , RIaecb008_1665, RIaecb080_1666, RIaecb0f8_1667, RIaecb170_1668, RIaecb1e8_1669, RIaecb260_1670, RIaecb2d8_1671, RIaecb350_1672, RIaecb3c8_1673, RIaecb440_1674, RIaecb4b8_1675, RIaecb530_1676, RIaecb5a8_1677, RIaecb620_1678, RIaecb698_1679, RIaecb710_1680, RIaecb788_1681, RIaecb800_1682, RIaecb878_1683, RIaecb8f0_1684, RIaecb968_1685, RIaecb9e0_1686, RIaecba58_1687, RIaecbad0_1688, RIaecbb48_1689, RIaecbbc0_1690, RIaecbc38_1691, RIaecbcb0_1692, RIaecbd28_1693, RIaecbda0_1694, RIaecbe18_1695, RIaecbe90_1696, RIaecbf08_1697, RIaecbf80_1698, RIaecbff8_1699, RIaecc070_1700, RIaecc0e8_1701, RIaecc160_1702, RIaecc1d8_1703, RIaecc250_1704, RIaecc2c8_1705, RIaecc340_1706, RIaecc3b8_1707, RIaecc430_1708, RIaecc4a8_1709, RIaecc520_1710, RIaecc598_1711, RIaecc610_1712, RIaecc688_1713, RIaecc700_1714, RIaecc778_1715, RIaecc7f0_1716, RIaecc868_1717, RIaecc8e0_1718, RIaecc958_1719, RIaecc9d0_1720, RIaecca48_1721, RIaeccac0_1722, RIaeccb38_1723, RIaeccbb0_1724, RIaeccc28_1725, RIaeccca0_1726, RIaeccd18_1727, RIaeccd90_1728);
and \U$28 ( \4743 , RIaecce08_1729, RIaecce80_1730, RIaeccef8_1731, RIaeccf70_1732, RIaeccfe8_1733, RIaecd060_1734, RIaecd0d8_1735, RIaecd150_1736, RIaecd1c8_1737, RIaecd240_1738, RIaecd2b8_1739, RIaecd330_1740, RIaecd3a8_1741, RIaecd420_1742, RIaecd498_1743, RIaecd510_1744, RIaecd588_1745, RIaecd600_1746, RIaecd678_1747, RIaecd6f0_1748, RIaecd768_1749, RIaecd7e0_1750, RIaecd858_1751, RIaecd8d0_1752, RIaecd948_1753, RIaecd9c0_1754, RIaecda38_1755, RIaecdab0_1756, RIaecdb28_1757, RIaecdba0_1758, RIaecdc18_1759, RIaecdc90_1760, RIaecdd08_1761, RIaecdd80_1762, RIaecddf8_1763, RIaecde70_1764, RIaecdee8_1765, RIaecdf60_1766, RIaecdfd8_1767, RIaece050_1768, RIaece0c8_1769, RIaece140_1770, RIaece1b8_1771, RIaece230_1772, RIaece2a8_1773, RIaece320_1774, RIaece398_1775, RIaece410_1776, RIaece488_1777, RIaece500_1778, RIaece578_1779, RIaece5f0_1780, RIaece668_1781, RIaece6e0_1782, RIaece758_1783, RIaece7d0_1784, RIaece848_1785, RIaece8c0_1786, RIaece938_1787, RIaece9b0_1788, RIaecea28_1789, RIaeceaa0_1790, RIaeceb18_1791, RIaeceb90_1792);
and \U$29 ( \4744 , RIaecec08_1793, RIaecec80_1794, RIaececf8_1795, RIaeced70_1796, RIaecede8_1797, RIaecee60_1798, RIaeceed8_1799, RIaecef50_1800, RIaecefc8_1801, RIaecf040_1802, RIaecf0b8_1803, RIaecf130_1804, RIaecf1a8_1805, RIaecf220_1806, RIaecf298_1807, RIaecf310_1808, RIaecf388_1809, RIaecf400_1810, RIaecf478_1811, RIaecf4f0_1812, RIaecf568_1813, RIaecf5e0_1814, RIaecf658_1815, RIaecf6d0_1816, RIaecf748_1817, RIaecf7c0_1818, RIaecf838_1819, RIaecf8b0_1820, RIaecf928_1821, RIaecf9a0_1822, RIaecfa18_1823, RIaecfa90_1824, RIaecfb08_1825, RIaecfb80_1826, RIaecfbf8_1827, RIaecfc70_1828, RIaecfce8_1829, RIaecfd60_1830, RIaecfdd8_1831, RIaecfe50_1832, RIaecfec8_1833, RIaecff40_1834, RIaecffb8_1835, RIaed0030_1836, RIaed00a8_1837, RIaed0120_1838, RIaed0198_1839, RIaed0210_1840, RIaed0288_1841, RIaed0300_1842, RIaed0378_1843, RIaed03f0_1844, RIaed0468_1845, RIaed04e0_1846, RIaed0558_1847, RIaed05d0_1848, RIaed0648_1849, RIaed06c0_1850, RIaed0738_1851, RIaed07b0_1852, RIaed0828_1853, RIaed08a0_1854, RIaed0918_1855, RIaed0990_1856);
and \U$30 ( \4745 , RIaed0a08_1857, RIaed0a80_1858, RIaed0af8_1859, RIaed0b70_1860, RIaed0be8_1861, RIaed0c60_1862, RIaed0cd8_1863, RIaed0d50_1864, RIaed0dc8_1865, RIaed0e40_1866, RIaed0eb8_1867, RIaed0f30_1868, RIaed0fa8_1869, RIaed1020_1870, RIaed1098_1871, RIaed1110_1872, RIaed1188_1873, RIaed1200_1874, RIaed1278_1875, RIaed12f0_1876, RIaed1368_1877, RIaed13e0_1878, RIaed1458_1879, RIaed14d0_1880, RIaed1548_1881, RIaed15c0_1882, RIaed1638_1883, RIaed16b0_1884, RIaed1728_1885, RIaed17a0_1886, RIaed1818_1887, RIaed1890_1888, RIaed1908_1889, RIaed1980_1890, RIaed19f8_1891, RIaed1a70_1892, RIaed1ae8_1893, RIaed1b60_1894, RIaed1bd8_1895, RIaed1c50_1896, RIaed1cc8_1897, RIaed1d40_1898, RIaed1db8_1899, RIaed1e30_1900, RIaed1ea8_1901, RIaed1f20_1902, RIaed1f98_1903, RIaed2010_1904, RIaed2088_1905, RIaed2100_1906, RIaed2178_1907, RIaed21f0_1908, RIaed2268_1909, RIaed22e0_1910, RIaed2358_1911, RIaed23d0_1912, RIaed2448_1913, RIaed24c0_1914, RIaed2538_1915, RIaed25b0_1916, RIaed2628_1917, RIaed26a0_1918, RIaed2718_1919, RIaed2790_1920);
and \U$31 ( \4746 , RIaed2808_1921, RIaed2880_1922, RIaed28f8_1923, RIaed2970_1924, RIaed29e8_1925, RIaed2a60_1926, RIaed2ad8_1927, RIaed2b50_1928, RIaed2bc8_1929, RIaed2c40_1930, RIaed2cb8_1931, RIaed2d30_1932, RIaed2da8_1933, RIaed2e20_1934, RIaed2e98_1935, RIaed2f10_1936, RIaed2f88_1937, RIaed3000_1938, RIaed3078_1939, RIaed30f0_1940, RIaed3168_1941, RIaed31e0_1942, RIaed3258_1943, RIaed32d0_1944, RIaed3348_1945, RIaed33c0_1946, RIaed3438_1947, RIaed34b0_1948, RIaed3528_1949, RIaed35a0_1950, RIaed3618_1951, RIaed3690_1952, RIaed3708_1953, RIaed3780_1954, RIaed37f8_1955, RIaed3870_1956, RIaed38e8_1957, RIaed3960_1958, RIaed39d8_1959, RIaed3a50_1960, RIaed3ac8_1961, RIaed3b40_1962, RIaed3bb8_1963, RIaed3c30_1964, RIaed3ca8_1965, RIaed3d20_1966, RIaed3d98_1967, RIaed3e10_1968, RIaed3e88_1969, RIaed3f00_1970, RIaed3f78_1971, RIaed3ff0_1972, RIaed4068_1973, RIaed40e0_1974, RIaed4158_1975, RIaed41d0_1976, RIaed4248_1977, RIaed42c0_1978, RIaed4338_1979, RIaed43b0_1980, RIaed4428_1981, RIaed44a0_1982, RIaed4518_1983, RIaed4590_1984);
and \U$32 ( \4747 , RIaed4608_1985, RIaed4680_1986, RIaed46f8_1987, RIaed4770_1988, RIaed47e8_1989, RIaed4860_1990, RIaed48d8_1991, RIaed4950_1992, RIaed49c8_1993, RIaed4a40_1994, RIaed4ab8_1995, RIaed4b30_1996, RIaed4ba8_1997, RIaed4c20_1998, RIaed4c98_1999, RIaed4d10_2000, RIaed4d88_2001, RIaed4e00_2002, RIaed4e78_2003, RIaed4ef0_2004, RIaed4f68_2005, RIaed4fe0_2006, RIaed5058_2007, RIaed50d0_2008, RIaed5148_2009, RIaed51c0_2010, RIaed5238_2011, RIaed52b0_2012, RIaed5328_2013, RIaed53a0_2014, RIaed5418_2015, RIaed5490_2016, RIaed5508_2017, RIaed5580_2018, RIaed55f8_2019, RIaed5670_2020, RIaed56e8_2021, RIaed5760_2022, RIaed57d8_2023, RIaed5850_2024, RIaed58c8_2025, RIaed5940_2026, RIaed59b8_2027, RIaed5a30_2028, RIaed5aa8_2029, RIaed5b20_2030, RIaed5b98_2031, RIaed5c10_2032, RIaed5c88_2033, RIaed5d00_2034, RIaed5d78_2035, RIaed5df0_2036, RIaed5e68_2037, RIaed5ee0_2038, RIaed5f58_2039, RIaed5fd0_2040, RIaed6048_2041, RIaed60c0_2042, RIaed6138_2043, RIaed61b0_2044, RIaed6228_2045, RIaed62a0_2046, RIaed6318_2047, RIaed6390_2048);
and \U$33 ( \4748 , RIaed6408_2049, RIaed6480_2050, RIaed64f8_2051, RIaed6570_2052, RIaed65e8_2053, RIaed6660_2054, RIaed66d8_2055, RIaed6750_2056, RIaed67c8_2057, RIaed6840_2058, RIaed68b8_2059, RIaed6930_2060, RIaed69a8_2061, RIaed6a20_2062, RIaed6a98_2063, RIaed6b10_2064, RIaed6b88_2065, RIaed6c00_2066, RIaed6c78_2067, RIaed6cf0_2068, RIaed6d68_2069, RIaed6de0_2070, RIaed6e58_2071, RIaed6ed0_2072, RIaed6f48_2073, RIaed6fc0_2074, RIaed7038_2075, RIaed70b0_2076, RIaed7128_2077, RIaed71a0_2078, RIaed7218_2079, RIaed7290_2080, RIaed7308_2081, RIaed7380_2082, RIaed73f8_2083, RIaed7470_2084, RIaed74e8_2085, RIaed7560_2086, RIaed75d8_2087, RIaed7650_2088, RIaed76c8_2089, RIaed7740_2090, RIaed77b8_2091, RIaed7830_2092, RIaed78a8_2093, RIaed7920_2094, RIaed7998_2095, RIaed7a10_2096, RIaed7a88_2097, RIaed7b00_2098, RIaed7b78_2099, RIaed7bf0_2100, RIaed7c68_2101, RIaed7ce0_2102, RIaed7d58_2103, RIaed7dd0_2104, RIaed7e48_2105, RIaed7ec0_2106, RIaed7f38_2107, RIaed7fb0_2108, RIaed8028_2109, RIaed80a0_2110, RIaed8118_2111, RIaed8190_2112);
and \U$34 ( \4749 , RIaed8208_2113, RIaed8280_2114, RIaed82f8_2115, RIaed8370_2116, RIaed83e8_2117, RIaed8460_2118, RIaed84d8_2119, RIaed8550_2120, RIaed85c8_2121, RIaed8640_2122, RIaed86b8_2123, RIaed8730_2124, RIaed87a8_2125, RIaed8820_2126, RIaed8898_2127, RIaed8910_2128, RIaed8988_2129, RIaed8a00_2130, RIaed8a78_2131, RIaed8af0_2132, RIaed8b68_2133, RIaed8be0_2134, RIaed8c58_2135, RIaed8cd0_2136, RIaed8d48_2137, RIaed8dc0_2138, RIaed8e38_2139, RIaed8eb0_2140, RIaed8f28_2141, RIaed8fa0_2142, RIaed9018_2143, RIaed9090_2144, RIaed9108_2145, RIaed9180_2146, RIaed91f8_2147, RIaed9270_2148, RIaed92e8_2149, RIaed9360_2150, RIaed93d8_2151, RIaed9450_2152, RIaed94c8_2153, RIaed9540_2154, RIaed95b8_2155, RIaed9630_2156, RIaed96a8_2157, RIaed9720_2158, RIaed9798_2159, RIaed9810_2160, RIaed9888_2161, RIaed9900_2162, RIaed9978_2163, RIaed99f0_2164, RIaed9a68_2165, RIaed9ae0_2166, RIaed9b58_2167, RIaed9bd0_2168, RIaed9c48_2169, RIaed9cc0_2170, RIaed9d38_2171, RIaed9db0_2172, RIaed9e28_2173, RIaed9ea0_2174, RIaed9f18_2175, RIaed9f90_2176);
and \U$35 ( \4750 , RIaeda008_2177, RIaeda080_2178, RIaeda0f8_2179, RIaeda170_2180, RIaeda1e8_2181, RIaeda260_2182, RIaeda2d8_2183, RIaeda350_2184, RIaeda3c8_2185, RIaeda440_2186, RIaeda4b8_2187, RIaeda530_2188, RIaeda5a8_2189, RIaeda620_2190, RIaeda698_2191, RIaeda710_2192, RIaeda788_2193, RIaeda800_2194, RIaeda878_2195, RIaeda8f0_2196, RIaeda968_2197, RIaeda9e0_2198, RIaedaa58_2199, RIaedaad0_2200, RIaedab48_2201, RIaedabc0_2202, RIaedac38_2203, RIaedacb0_2204, RIaedad28_2205, RIaedada0_2206, RIaedae18_2207, RIaedae90_2208, RIaedaf08_2209, RIaedaf80_2210, RIaedaff8_2211, RIaedb070_2212, RIaedb0e8_2213, RIaedb160_2214, RIaedb1d8_2215, RIaedb250_2216, RIaedb2c8_2217, RIaedb340_2218, RIaedb3b8_2219, RIaedb430_2220, RIaedb4a8_2221, RIaedb520_2222, RIaedb598_2223, RIaedb610_2224, RIaedb688_2225, RIaedb700_2226, RIaedb778_2227, RIaedb7f0_2228, RIaedb868_2229, RIaedb8e0_2230, RIaedb958_2231, RIaedb9d0_2232, RIaedba48_2233, RIaedbac0_2234, RIaedbb38_2235, RIaedbbb0_2236, RIaedbc28_2237, RIaedbca0_2238, RIaedbd18_2239, RIaedbd90_2240);
and \U$36 ( \4751 , RIaedbe08_2241, RIaedbe80_2242, RIaedbef8_2243, RIaedbf70_2244, RIaedbfe8_2245, RIaedc060_2246, RIaedc0d8_2247, RIaedc150_2248, RIaedc1c8_2249, RIaedc240_2250, RIaedc2b8_2251, RIaedc330_2252, RIaedc3a8_2253, RIaedc420_2254, RIaedc498_2255, RIaedc510_2256, RIaedc588_2257, RIaedc600_2258, RIaedc678_2259, RIaedc6f0_2260, RIaedc768_2261, RIaedc7e0_2262, RIaedc858_2263, RIaedc8d0_2264, RIaedc948_2265, RIaedc9c0_2266, RIaedca38_2267, RIaedcab0_2268, RIaedcb28_2269, RIaedcba0_2270, RIaedcc18_2271, RIaedcc90_2272, RIaedcd08_2273, RIaedcd80_2274, RIaedcdf8_2275, RIaedce70_2276, RIaedcee8_2277, RIaedcf60_2278, RIaedcfd8_2279, RIaedd050_2280, RIaedd0c8_2281, RIaedd140_2282, RIaedd1b8_2283, RIaedd230_2284, RIaedd2a8_2285, RIaedd320_2286, RIaedd398_2287, RIaedd410_2288, RIaedd488_2289, RIaedd500_2290, RIaedd578_2291, RIaedd5f0_2292, RIaedd668_2293, RIaedd6e0_2294, RIaedd758_2295, RIaedd7d0_2296, RIaedd848_2297, RIaedd8c0_2298, RIaedd938_2299, RIaedd9b0_2300, RIaedda28_2301, RIaeddaa0_2302, RIaeddb18_2303, RIaeddb90_2304);
and \U$37 ( \4752 , RIaeddc08_2305, RIaeddc80_2306, RIaeddcf8_2307, RIaeddd70_2308, RIaeddde8_2309, RIaedde60_2310, RIaedded8_2311, RIaeddf50_2312, RIaeddfc8_2313, RIaede040_2314, RIaede0b8_2315, RIaede130_2316, RIaede1a8_2317, RIaede220_2318, RIaede298_2319, RIaede310_2320, RIaede388_2321, RIaede400_2322, RIaede478_2323, RIaede4f0_2324, RIaede568_2325, RIaede5e0_2326, RIaede658_2327, RIaede6d0_2328, RIaede748_2329, RIaede7c0_2330, RIaede838_2331, RIaede8b0_2332, RIaede928_2333, RIaede9a0_2334, RIaedea18_2335, RIaedea90_2336, RIaedeb08_2337, RIaedeb80_2338, RIaedebf8_2339, RIaedec70_2340, RIaedece8_2341, RIaeded60_2342, RIaededd8_2343, RIaedee50_2344, RIaedeec8_2345, RIaedef40_2346, RIaedefb8_2347, RIaedf030_2348, RIaedf0a8_2349, RIaedf120_2350, RIaedf198_2351, RIaedf210_2352, RIaedf288_2353, RIaedf300_2354, RIaedf378_2355, RIaedf3f0_2356, RIaedf468_2357, RIaedf4e0_2358, RIaedf558_2359, RIaedf5d0_2360, RIaedf648_2361, RIaedf6c0_2362, RIaedf738_2363, RIaedf7b0_2364, RIaedf828_2365, RIaedf8a0_2366, RIaedf918_2367, RIaedf990_2368);
and \U$38 ( \4753 , RIaedfa08_2369, RIaedfa80_2370, RIaedfaf8_2371, RIaedfb70_2372, RIaedfbe8_2373, RIaedfc60_2374, RIaedfcd8_2375, RIaedfd50_2376, RIaedfdc8_2377, RIaedfe40_2378, RIaedfeb8_2379, RIaedff30_2380, RIaedffa8_2381, RIaee0020_2382, RIaee0098_2383, RIaee0110_2384, RIaee0188_2385, RIaee0200_2386, RIaee0278_2387, RIaee02f0_2388, RIaee0368_2389, RIaee03e0_2390, RIaee0458_2391, RIaee04d0_2392, RIaee0548_2393, RIaee05c0_2394, RIaee0638_2395, RIaee06b0_2396, RIaee0728_2397, RIaee07a0_2398, RIaee0818_2399, RIaee0890_2400, RIaee0908_2401, RIaee0980_2402, RIaee09f8_2403, RIaee0a70_2404, RIaee0ae8_2405, RIaee0b60_2406, RIaee0bd8_2407, RIaee0c50_2408, RIaee0cc8_2409, RIaee0d40_2410, RIaee0db8_2411, RIaee0e30_2412, RIaee0ea8_2413, RIaee0f20_2414, RIaee0f98_2415, RIaee1010_2416, RIaee1088_2417, RIaee1100_2418, RIaee1178_2419, RIaee11f0_2420, RIaee1268_2421, RIaee12e0_2422, RIaee1358_2423, RIaee13d0_2424, RIaee1448_2425, RIaee14c0_2426, RIaee1538_2427, RIaee15b0_2428, RIaee1628_2429, RIaee16a0_2430, RIaee1718_2431, RIaee1790_2432);
and \U$39 ( \4754 , RIaee1808_2433, RIaee1880_2434, RIaee18f8_2435, RIaee1970_2436, RIaee19e8_2437, RIaee1a60_2438, RIaee1ad8_2439, RIaee1b50_2440, RIaee1bc8_2441, RIaee1c40_2442, RIaee1cb8_2443, RIaee1d30_2444, RIaee1da8_2445, RIaee1e20_2446, RIaee1e98_2447, RIaee1f10_2448, RIaee1f88_2449, RIaee2000_2450, RIaee2078_2451, RIaee20f0_2452, RIaee2168_2453, RIaee21e0_2454, RIaee2258_2455, RIaee22d0_2456, RIaee2348_2457, RIaee23c0_2458, RIaee2438_2459, RIaee24b0_2460, RIaee2528_2461, RIaee25a0_2462, RIaee2618_2463, RIaee2690_2464, RIaee2708_2465, RIaee2780_2466, RIaee27f8_2467, RIaee2870_2468, RIaee28e8_2469, RIaee2960_2470, RIaee29d8_2471, RIaee2a50_2472, RIaee2ac8_2473, RIaee2b40_2474, RIaee2bb8_2475, RIaee2c30_2476, RIaee2ca8_2477, RIaee2d20_2478, RIaee2d98_2479, RIaee2e10_2480, RIaee2e88_2481, RIaee2f00_2482, RIaee2f78_2483, RIaee2ff0_2484, RIaee3068_2485, RIaee30e0_2486, RIaee3158_2487, RIaee31d0_2488, RIaee3248_2489, RIaee32c0_2490, RIaee3338_2491, RIaee33b0_2492, RIaee3428_2493, RIaee34a0_2494, RIaee3518_2495, RIaee3590_2496);
and \U$40 ( \4755 , RIaee3608_2497, RIaee3680_2498, RIaee36f8_2499, RIaee3770_2500, RIaee37e8_2501, RIaee3860_2502, RIaee38d8_2503, RIaee3950_2504, RIaee39c8_2505, RIaee3a40_2506, RIaee3ab8_2507, RIaee3b30_2508, RIaee3ba8_2509, RIaee3c20_2510, RIaee3c98_2511, RIaee3d10_2512, RIaee3d88_2513, RIaee3e00_2514, RIaee3e78_2515, RIaee3ef0_2516, RIaee3f68_2517, RIaee3fe0_2518, RIaee4058_2519, RIaee40d0_2520, RIaee4148_2521, RIaee41c0_2522, RIaee4238_2523, RIaee42b0_2524, RIaee4328_2525, RIaee43a0_2526, RIaee4418_2527, RIaee4490_2528, RIaee4508_2529, RIaee4580_2530, RIaee45f8_2531, RIaee4670_2532, RIaee46e8_2533, RIaee4760_2534, RIaee47d8_2535, RIaee4850_2536, RIaee48c8_2537, RIaee4940_2538, RIaee49b8_2539, RIaee4a30_2540, RIaee4aa8_2541, RIaee4b20_2542, RIaee4b98_2543, RIaee4c10_2544, RIaee4c88_2545, RIaee4d00_2546, RIaee4d78_2547, RIaee4df0_2548, RIaee4e68_2549, RIaee4ee0_2550, RIaee4f58_2551, RIaee4fd0_2552, RIaee5048_2553, RIaee50c0_2554, RIaee5138_2555, RIaee51b0_2556, RIaee5228_2557, RIaee52a0_2558, RIaee5318_2559, RIaee5390_2560);
and \U$41 ( \4756 , RIaee5408_2561, RIaee5480_2562, RIaee54f8_2563, RIaee5570_2564, RIaee55e8_2565, RIaee5660_2566, RIaee56d8_2567, RIaee5750_2568, RIaee57c8_2569, RIaee5840_2570, RIaee58b8_2571, RIaee5930_2572, RIaee59a8_2573, RIaee5a20_2574, RIaee5a98_2575, RIaee5b10_2576, RIaee5b88_2577, RIaee5c00_2578, RIaee5c78_2579, RIaee5cf0_2580, RIaee5d68_2581, RIaee5de0_2582, RIaee5e58_2583, RIaee5ed0_2584, RIaee5f48_2585, RIaee5fc0_2586, RIaee6038_2587, RIaee60b0_2588, RIaee6128_2589, RIaee61a0_2590, RIaee6218_2591, RIaee6290_2592, RIaee6308_2593, RIaee6380_2594, RIaee63f8_2595, RIaee6470_2596, RIaee64e8_2597, RIaee6560_2598, RIaee65d8_2599, RIaee6650_2600, RIaee66c8_2601, RIaee6740_2602, RIaee67b8_2603, RIaee6830_2604, RIaee68a8_2605, RIaee6920_2606, RIaee6998_2607, RIaee6a10_2608, RIaee6a88_2609, RIaee6b00_2610, RIaee6b78_2611, RIaee6bf0_2612, RIaee6c68_2613, RIaee6ce0_2614, RIaee6d58_2615, RIaee6dd0_2616, RIaee6e48_2617, RIaee6ec0_2618, RIaee6f38_2619, RIaee6fb0_2620, RIaee7028_2621, RIaee70a0_2622, RIaee7118_2623, RIaee7190_2624);
and \U$42 ( \4757 , RIaee7208_2625, RIaee7280_2626, RIaee72f8_2627, RIaee7370_2628, RIaee73e8_2629, RIaee7460_2630, RIaee74d8_2631, RIaee7550_2632, RIaee75c8_2633, RIaee7640_2634, RIaee76b8_2635, RIaee7730_2636, RIaee77a8_2637, RIaee7820_2638, RIaee7898_2639, RIaee7910_2640, RIaee7988_2641, RIaee7a00_2642, RIaee7a78_2643, RIaee7af0_2644, RIaee7b68_2645, RIaee7be0_2646, RIaee7c58_2647, RIaee7cd0_2648, RIaee7d48_2649, RIaee7dc0_2650, RIaee7e38_2651, RIaee7eb0_2652, RIaee7f28_2653, RIaee7fa0_2654, RIaee8018_2655, RIaee8090_2656, RIaee8108_2657, RIaee8180_2658, RIaee81f8_2659, RIaee8270_2660, RIaee82e8_2661, RIaee8360_2662, RIaee83d8_2663, RIaee8450_2664, RIaee84c8_2665, RIaee8540_2666, RIaee85b8_2667, RIaee8630_2668, RIaee86a8_2669, RIaee8720_2670, RIaee8798_2671, RIaee8810_2672, RIaee8888_2673, RIaee8900_2674, RIaee8978_2675, RIaee89f0_2676, RIaee8a68_2677, RIaee8ae0_2678, RIaee8b58_2679, RIaee8bd0_2680, RIaee8c48_2681, RIaee8cc0_2682, RIaee8d38_2683, RIaee8db0_2684, RIaee8e28_2685, RIaee8ea0_2686, RIaee8f18_2687, RIaee8f90_2688);
and \U$43 ( \4758 , RIaee9008_2689, RIaee9080_2690, RIaee90f8_2691, RIaee9170_2692, RIaee91e8_2693, RIaee9260_2694, RIaee92d8_2695, RIaee9350_2696, RIaee93c8_2697, RIaee9440_2698, RIaee94b8_2699, RIaee9530_2700, RIaee95a8_2701, RIaee9620_2702, RIaee9698_2703, RIaee9710_2704, RIaee9788_2705, RIaee9800_2706, RIaee9878_2707, RIaee98f0_2708, RIaee9968_2709, RIaee99e0_2710, RIaee9a58_2711, RIaee9ad0_2712, RIaee9b48_2713, RIaee9bc0_2714, RIaee9c38_2715, RIaee9cb0_2716, RIaee9d28_2717, RIaee9da0_2718, RIaee9e18_2719, RIaee9e90_2720, RIaee9f08_2721, RIaee9f80_2722, RIaee9ff8_2723, RIaeea070_2724, RIaeea0e8_2725, RIaeea160_2726, RIaeea1d8_2727, RIaeea250_2728, RIaeea2c8_2729, RIaeea340_2730, RIaeea3b8_2731, RIaeea430_2732, RIaeea4a8_2733, RIaeea520_2734, RIaeea598_2735, RIaeea610_2736, RIaeea688_2737, RIaeea700_2738, RIaeea778_2739, RIaeea7f0_2740, RIaeea868_2741, RIaeea8e0_2742, RIaeea958_2743, RIaeea9d0_2744, RIaeeaa48_2745, RIaeeaac0_2746, RIaeeab38_2747, RIaeeabb0_2748, RIaeeac28_2749, RIaeeaca0_2750, RIaeead18_2751, RIaeead90_2752);
and \U$44 ( \4759 , RIaeeae08_2753, RIaeeae80_2754, RIaeeaef8_2755, RIaeeaf70_2756, RIaeeafe8_2757, RIaeeb060_2758, RIaeeb0d8_2759, RIaeeb150_2760, RIaeeb1c8_2761, RIaeeb240_2762, RIaeeb2b8_2763, RIaeeb330_2764, RIaeeb3a8_2765, RIaeeb420_2766, RIaeeb498_2767, RIaeeb510_2768, RIaeeb588_2769, RIaeeb600_2770, RIaeeb678_2771, RIaeeb6f0_2772, RIaeeb768_2773, RIaeeb7e0_2774, RIaeeb858_2775, RIaeeb8d0_2776, RIaeeb948_2777, RIaeeb9c0_2778, RIaeeba38_2779, RIaeebab0_2780, RIaeebb28_2781, RIaeebba0_2782, RIaeebc18_2783, RIaeebc90_2784, RIaeebd08_2785, RIaeebd80_2786, RIaeebdf8_2787, RIaeebe70_2788, RIaeebee8_2789, RIaeebf60_2790, RIaeebfd8_2791, RIaeec050_2792, RIaeec0c8_2793, RIaeec140_2794, RIaeec1b8_2795, RIaeec230_2796, RIaeec2a8_2797, RIaeec320_2798, RIaeec398_2799, RIaeec410_2800, RIaeec488_2801, RIaeec500_2802, RIaeec578_2803, RIaeec5f0_2804, RIaeec668_2805, RIaeec6e0_2806, RIaeec758_2807, RIaeec7d0_2808, RIaeec848_2809, RIaeec8c0_2810, RIaeec938_2811, RIaeec9b0_2812, RIaeeca28_2813, RIaeecaa0_2814, RIaeecb18_2815, RIaeecb90_2816);
and \U$45 ( \4760 , RIaeecc08_2817, RIaeecc80_2818, RIaeeccf8_2819, RIaeecd70_2820, RIaeecde8_2821, RIaeece60_2822, RIaeeced8_2823, RIaeecf50_2824, RIaeecfc8_2825, RIaeed040_2826, RIaeed0b8_2827, RIaeed130_2828, RIaeed1a8_2829, RIaeed220_2830, RIaeed298_2831, RIaeed310_2832, RIaeed388_2833, RIaeed400_2834, RIaeed478_2835, RIaeed4f0_2836, RIaeed568_2837, RIaeed5e0_2838, RIaeed658_2839, RIaeed6d0_2840, RIaeed748_2841, RIaeed7c0_2842, RIaeed838_2843, RIaeed8b0_2844, RIaeed928_2845, RIaeed9a0_2846, RIaeeda18_2847, RIaeeda90_2848, RIaeedb08_2849, RIaeedb80_2850, RIaeedbf8_2851, RIaeedc70_2852, RIaeedce8_2853, RIaeedd60_2854, RIaeeddd8_2855, RIaeede50_2856, RIaeedec8_2857, RIaeedf40_2858, RIaeedfb8_2859, RIaeee030_2860, RIaeee0a8_2861, RIaeee120_2862, RIaeee198_2863, RIaeee210_2864, RIaeee288_2865, RIaeee300_2866, RIaeee378_2867, RIaeee3f0_2868, RIaeee468_2869, RIaeee4e0_2870, RIaeee558_2871, RIaeee5d0_2872, RIaeee648_2873, RIaeee6c0_2874, RIaeee738_2875, RIaeee7b0_2876, RIaeee828_2877, RIaeee8a0_2878, RIaeee918_2879, RIaeee990_2880);
and \U$46 ( \4761 , RIaeeea08_2881, RIaeeea80_2882, RIaeeeaf8_2883, RIaeeeb70_2884, RIaeeebe8_2885, RIaeeec60_2886, RIaeeecd8_2887, RIaeeed50_2888, RIaeeedc8_2889, RIaeeee40_2890, RIaeeeeb8_2891, RIaeeef30_2892, RIaeeefa8_2893, RIaeef020_2894, RIaeef098_2895, RIaeef110_2896, RIaeef188_2897, RIaeef200_2898, RIaeef278_2899, RIaeef2f0_2900, RIaeef368_2901, RIaeef3e0_2902, RIaeef458_2903, RIaeef4d0_2904, RIaeef548_2905, RIaeef5c0_2906, RIaeef638_2907, RIaeef6b0_2908, RIaeef728_2909, RIaeef7a0_2910, RIaeef818_2911, RIaeef890_2912, RIaeef908_2913, RIaeef980_2914, RIaeef9f8_2915, RIaeefa70_2916, RIaeefae8_2917, RIaeefb60_2918, RIaeefbd8_2919, RIaeefc50_2920, RIaeefcc8_2921, RIaeefd40_2922, RIaeefdb8_2923, RIaeefe30_2924, RIaeefea8_2925, RIaeeff20_2926, RIaeeff98_2927, RIaef0010_2928, RIaef0088_2929, RIaef0100_2930, RIaef0178_2931, RIaef01f0_2932, RIaef0268_2933, RIaef02e0_2934, RIaef0358_2935, RIaef03d0_2936, RIaef0448_2937, RIaef04c0_2938, RIaef0538_2939, RIaef05b0_2940, RIaef0628_2941, RIaef06a0_2942, RIaef0718_2943, RIaef0790_2944);
and \U$47 ( \4762 , RIaef0808_2945, RIaef0880_2946, RIaef08f8_2947, RIaef0970_2948, RIaef09e8_2949, RIaef0a60_2950, RIaef0ad8_2951, RIaef0b50_2952, RIaef0bc8_2953, RIaef0c40_2954, RIaef0cb8_2955, RIaef0d30_2956, RIaef0da8_2957, RIaef0e20_2958, RIaef0e98_2959, RIaef0f10_2960, RIaef0f88_2961, RIaef1000_2962, RIaef1078_2963, RIaef10f0_2964, RIaef1168_2965, RIaef11e0_2966, RIaef1258_2967, RIaef12d0_2968, RIaef1348_2969, RIaef13c0_2970, RIaef1438_2971, RIaef14b0_2972, RIaef1528_2973, RIaef15a0_2974, RIaef1618_2975, RIaef1690_2976, RIaef1708_2977, RIaef1780_2978, RIaef17f8_2979, RIaef1870_2980, RIaef18e8_2981, RIaef1960_2982, RIaef19d8_2983, RIaef1a50_2984, RIaef1ac8_2985, RIaef1b40_2986, RIaef1bb8_2987, RIaef1c30_2988, RIaef1ca8_2989, RIaef1d20_2990, RIaef1d98_2991, RIaef1e10_2992, RIaef1e88_2993, RIaef1f00_2994, RIaef1f78_2995, RIaef1ff0_2996, RIaef2068_2997, RIaef20e0_2998, RIaef2158_2999, RIaef21d0_3000, RIaef2248_3001, RIaef22c0_3002, RIaef2338_3003, RIaef23b0_3004, RIaef2428_3005, RIaef24a0_3006, RIaef2518_3007, RIaef2590_3008);
and \U$48 ( \4763 , RIaef2608_3009, RIaef2680_3010, RIaef26f8_3011, RIaef2770_3012, RIaef27e8_3013, RIaef2860_3014, RIaef28d8_3015, RIaef2950_3016, RIaef29c8_3017, RIaef2a40_3018, RIaef2ab8_3019, RIaef2b30_3020, RIaef2ba8_3021, RIaef2c20_3022, RIaef2c98_3023, RIaef2d10_3024, RIaef2d88_3025, RIaef2e00_3026, RIaef2e78_3027, RIaef2ef0_3028, RIaef2f68_3029, RIaef2fe0_3030, RIaef3058_3031, RIaef30d0_3032, RIaef3148_3033, RIaef31c0_3034, RIaef3238_3035, RIaef32b0_3036, RIaef3328_3037, RIaef33a0_3038, RIaef3418_3039, RIaef3490_3040, RIaef3508_3041, RIaef3580_3042, RIaef35f8_3043, RIaef3670_3044, RIaef36e8_3045, RIaef3760_3046, RIaef37d8_3047, RIaef3850_3048, RIaef38c8_3049, RIaef3940_3050, RIaef39b8_3051, RIaef3a30_3052, RIaef3aa8_3053, RIaef3b20_3054, RIaef3b98_3055, RIaef3c10_3056, RIaef3c88_3057, RIaef3d00_3058, RIaef3d78_3059, RIaef3df0_3060, RIaef3e68_3061, RIaef3ee0_3062, RIaef3f58_3063, RIaef3fd0_3064, RIaef4048_3065, RIaef40c0_3066, RIaef4138_3067, RIaef41b0_3068, RIaef4228_3069, RIaef42a0_3070, RIaef4318_3071, RIaef4390_3072);
and \U$49 ( \4764 , RIaef4408_3073, RIaef4480_3074, RIaef44f8_3075, RIaef4570_3076, RIaef45e8_3077, RIaef4660_3078, RIaef46d8_3079, RIaef4750_3080, RIaef47c8_3081, RIaef4840_3082, RIaef48b8_3083, RIaef4930_3084, RIaef49a8_3085, RIaef4a20_3086, RIaef4a98_3087, RIaef4b10_3088, RIaef4b88_3089, RIaef4c00_3090, RIaef4c78_3091, RIaef4cf0_3092, RIaef4d68_3093, RIaef4de0_3094, RIaef4e58_3095, RIaef4ed0_3096, RIaef4f48_3097, RIaef4fc0_3098, RIaef5038_3099, RIaef50b0_3100, RIaef5128_3101, RIaef51a0_3102, RIaef5218_3103, RIaef5290_3104, RIaef5308_3105, RIaef5380_3106, RIaef53f8_3107, RIaef5470_3108, RIaef54e8_3109, RIaef5560_3110, RIaef55d8_3111, RIaef5650_3112, RIaef56c8_3113, RIaef5740_3114, RIaef57b8_3115, RIaef5830_3116, RIaef58a8_3117, RIaef5920_3118, RIaef5998_3119, RIaef5a10_3120, RIaef5a88_3121, RIaef5b00_3122, RIaef5b78_3123, RIaef5bf0_3124, RIaef5c68_3125, RIaef5ce0_3126, RIaef5d58_3127, RIaef5dd0_3128, RIaef5e48_3129, RIaef5ec0_3130, RIaef5f38_3131, RIaef5fb0_3132, RIaef6028_3133, RIaef60a0_3134, RIaef6118_3135, RIaef6190_3136);
and \U$50 ( \4765 , RIaef6208_3137, RIaef6280_3138, RIaef62f8_3139, RIaef6370_3140, RIaef63e8_3141, RIaef6460_3142, RIaef64d8_3143, RIaef6550_3144, RIaef65c8_3145, RIaef6640_3146, RIaef66b8_3147, RIaef6730_3148, RIaef67a8_3149, RIaef6820_3150, RIaef6898_3151, RIaef6910_3152, RIaef6988_3153, RIaef6a00_3154, RIaef6a78_3155, RIaef6af0_3156, RIaef6b68_3157, RIaef6be0_3158, RIaef6c58_3159, RIaef6cd0_3160, RIaef6d48_3161, RIaef6dc0_3162, RIaef6e38_3163, RIaef6eb0_3164, RIaef6f28_3165, RIaef6fa0_3166, RIaef7018_3167, RIaef7090_3168, RIaef7108_3169, RIaef7180_3170, RIaef71f8_3171, RIaef7270_3172, RIaef72e8_3173, RIaef7360_3174, RIaef73d8_3175, RIaef7450_3176, RIaef74c8_3177, RIaef7540_3178, RIaef75b8_3179, RIaef7630_3180, RIaef76a8_3181, RIaef7720_3182, RIaef7798_3183, RIaef7810_3184, RIaef7888_3185, RIaef7900_3186, RIaef7978_3187, RIaef79f0_3188, RIaef7a68_3189, RIaef7ae0_3190, RIaef7b58_3191, RIaef7bd0_3192, RIaef7c48_3193, RIaef7cc0_3194, RIaef7d38_3195, RIaef7db0_3196, RIaef7e28_3197, RIaef7ea0_3198, RIaef7f18_3199, RIaef7f90_3200);
and \U$51 ( \4766 , RIaef8008_3201, RIaef8080_3202, RIaef80f8_3203, RIaef8170_3204, RIaef81e8_3205, RIaef8260_3206, RIaef82d8_3207, RIaef8350_3208, RIaef83c8_3209, RIaef8440_3210, RIaef84b8_3211, RIaef8530_3212, RIaef85a8_3213, RIaef8620_3214, RIaef8698_3215, RIaef8710_3216, RIaef8788_3217, RIaef8800_3218, RIaef8878_3219, RIaef88f0_3220, RIaef8968_3221, RIaef89e0_3222, RIaef8a58_3223, RIaef8ad0_3224, RIaef8b48_3225, RIaef8bc0_3226, RIaef8c38_3227, RIaef8cb0_3228, RIaef8d28_3229, RIaef8da0_3230, RIaef8e18_3231, RIaef8e90_3232, RIaef8f08_3233, RIaef8f80_3234, RIaef8ff8_3235, RIaef9070_3236, RIaef90e8_3237, RIaef9160_3238, RIaef91d8_3239, RIaef9250_3240, RIaef92c8_3241, RIaef9340_3242, RIaef93b8_3243, RIaef9430_3244, RIaef94a8_3245, RIaef9520_3246, RIaef9598_3247, RIaef9610_3248, RIaef9688_3249, RIaef9700_3250, RIaef9778_3251, RIaef97f0_3252, RIaef9868_3253, RIaef98e0_3254, RIaef9958_3255, RIaef99d0_3256, RIaef9a48_3257, RIaef9ac0_3258, RIaef9b38_3259, RIaef9bb0_3260, RIaef9c28_3261, RIaef9ca0_3262, RIaef9d18_3263, RIaef9d90_3264);
and \U$52 ( \4767 , RIaef9e08_3265, RIaef9e80_3266, RIaef9ef8_3267, RIaef9f70_3268, RIaef9fe8_3269, RIaefa060_3270, RIaefa0d8_3271, RIaefa150_3272, RIaefa1c8_3273, RIaefa240_3274, RIaefa2b8_3275, RIaefa330_3276, RIaefa3a8_3277, RIaefa420_3278, RIaefa498_3279, RIaefa510_3280, RIaefa588_3281, RIaefa600_3282, RIaefa678_3283, RIaefa6f0_3284, RIaefa768_3285, RIaefa7e0_3286, RIaefa858_3287, RIaefa8d0_3288, RIaefa948_3289, RIaefa9c0_3290, RIaefaa38_3291, RIaefaab0_3292, RIaefab28_3293, RIaefaba0_3294, RIaefac18_3295, RIaefac90_3296, RIaefad08_3297, RIaefad80_3298, RIaefadf8_3299, RIaefae70_3300, RIaefaee8_3301, RIaefaf60_3302, RIaefafd8_3303, RIaefb050_3304, RIaefb0c8_3305, RIaefb140_3306, RIaefb1b8_3307, RIaefb230_3308, RIaefb2a8_3309, RIaefb320_3310, RIaefb398_3311, RIaefb410_3312, RIaefb488_3313, RIaefb500_3314, RIaefb578_3315, RIaefb5f0_3316, RIaefb668_3317, RIaefb6e0_3318, RIaefb758_3319, RIaefb7d0_3320, RIaefb848_3321, RIaefb8c0_3322, RIaefb938_3323, RIaefb9b0_3324, RIaefba28_3325, RIaefbaa0_3326, RIaefbb18_3327, RIaefbb90_3328);
and \U$53 ( \4768 , RIaefbc08_3329, RIaefbc80_3330, RIaefbcf8_3331, RIaefbd70_3332, RIaefbde8_3333, RIaefbe60_3334, RIaefbed8_3335, RIaefbf50_3336, RIaefbfc8_3337, RIaefc040_3338, RIaefc0b8_3339, RIaefc130_3340, RIaefc1a8_3341, RIaefc220_3342, RIaefc298_3343, RIaefc310_3344, RIaefc388_3345, RIaefc400_3346, RIaefc478_3347, RIaefc4f0_3348, RIaefc568_3349, RIaefc5e0_3350, RIaefc658_3351, RIaefc6d0_3352, RIaefc748_3353, RIaefc7c0_3354, RIaefc838_3355, RIaefc8b0_3356, RIaefc928_3357, RIaefc9a0_3358, RIaefca18_3359, RIaefca90_3360, RIaefcb08_3361, RIaefcb80_3362, RIaefcbf8_3363, RIaefcc70_3364, RIaefcce8_3365, RIaefcd60_3366, RIaefcdd8_3367, RIaefce50_3368, RIaefcec8_3369, RIaefcf40_3370, RIaefcfb8_3371, RIaefd030_3372, RIaefd0a8_3373, RIaefd120_3374, RIaefd198_3375, RIaefd210_3376, RIaefd288_3377, RIaefd300_3378, RIaefd378_3379, RIaefd3f0_3380, RIaefd468_3381, RIaefd4e0_3382, RIaefd558_3383, RIaefd5d0_3384, RIaefd648_3385, RIaefd6c0_3386, RIaefd738_3387, RIaefd7b0_3388, RIaefd828_3389, RIaefd8a0_3390, RIaefd918_3391, RIaefd990_3392);
and \U$54 ( \4769 , RIaefda08_3393, RIaefda80_3394, RIaefdaf8_3395, RIaefdb70_3396, RIaefdbe8_3397, RIaefdc60_3398, RIaefdcd8_3399, RIaefdd50_3400, RIaefddc8_3401, RIaefde40_3402, RIaefdeb8_3403, RIaefdf30_3404, RIaefdfa8_3405, RIaefe020_3406, RIaefe098_3407, RIaefe110_3408, RIaefe188_3409, RIaefe200_3410, RIaefe278_3411, RIaefe2f0_3412, RIaefe368_3413, RIaefe3e0_3414, RIaefe458_3415, RIaefe4d0_3416, RIaefe548_3417, RIaefe5c0_3418, RIaefe638_3419, RIaefe6b0_3420, RIaefe728_3421, RIaefe7a0_3422, RIaefe818_3423, RIaefe890_3424, RIaefe908_3425, RIaefe980_3426, RIaefe9f8_3427, RIaefea70_3428, RIaefeae8_3429, RIaefeb60_3430, RIaefebd8_3431, RIaefec50_3432, RIaefecc8_3433, RIaefed40_3434, RIaefedb8_3435, RIaefee30_3436, RIaefeea8_3437, RIaefef20_3438, RIaefef98_3439, RIaeff010_3440, RIaeff088_3441, RIaeff100_3442, RIaeff178_3443, RIaeff1f0_3444, RIaeff268_3445, RIaeff2e0_3446, RIaeff358_3447, RIaeff3d0_3448, RIaeff448_3449, RIaeff4c0_3450, RIaeff538_3451, RIaeff5b0_3452, RIaeff628_3453, RIaeff6a0_3454, RIaeff718_3455, RIaeff790_3456);
and \U$55 ( \4770 , RIaeff808_3457, RIaeff880_3458, RIaeff8f8_3459, RIaeff970_3460, RIaeff9e8_3461, RIaeffa60_3462, RIaeffad8_3463, RIaeffb50_3464, RIaeffbc8_3465, RIaeffc40_3466, RIaeffcb8_3467, RIaeffd30_3468, RIaeffda8_3469, RIaeffe20_3470, RIaeffe98_3471, RIaefff10_3472, RIaefff88_3473, RIaf00000_3474, RIaf00078_3475, RIaf000f0_3476, RIaf00168_3477, RIaf001e0_3478, RIaf00258_3479, RIaf002d0_3480, RIaf00348_3481, RIaf003c0_3482, RIaf00438_3483, RIaf004b0_3484, RIaf00528_3485, RIaf005a0_3486, RIaf00618_3487, RIaf00690_3488, RIaf00708_3489, RIaf00780_3490, RIaf007f8_3491, RIaf00870_3492, RIaf008e8_3493, RIaf00960_3494, RIaf009d8_3495, RIaf00a50_3496, RIaf00ac8_3497, RIaf00b40_3498, RIaf00bb8_3499, RIaf00c30_3500, RIaf00ca8_3501, RIaf00d20_3502, RIaf00d98_3503, RIaf00e10_3504, RIaf00e88_3505, RIaf00f00_3506, RIaf00f78_3507, RIaf00ff0_3508, RIaf01068_3509, RIaf010e0_3510, RIaf01158_3511, RIaf011d0_3512, RIaf01248_3513, RIaf012c0_3514, RIaf01338_3515, RIaf013b0_3516, RIaf01428_3517, RIaf014a0_3518, RIaf01518_3519, RIaf01590_3520);
and \U$56 ( \4771 , RIaf01608_3521, RIaf01680_3522, RIaf016f8_3523, RIaf01770_3524, RIaf017e8_3525, RIaf01860_3526, RIaf018d8_3527, RIaf01950_3528, RIaf019c8_3529, RIaf01a40_3530, RIaf01ab8_3531, RIaf01b30_3532, RIaf01ba8_3533, RIaf01c20_3534, RIaf01c98_3535, RIaf01d10_3536, RIaf01d88_3537, RIaf01e00_3538, RIaf01e78_3539, RIaf01ef0_3540, RIaf01f68_3541, RIaf01fe0_3542, RIaf02058_3543, RIaf020d0_3544, RIaf02148_3545, RIaf021c0_3546, RIaf02238_3547, RIaf022b0_3548, RIaf02328_3549, RIaf023a0_3550, RIaf02418_3551, RIaf02490_3552, RIaf02508_3553, RIaf02580_3554, RIaf025f8_3555, RIaf02670_3556, RIaf026e8_3557, RIaf02760_3558, RIaf027d8_3559, RIaf02850_3560, RIaf028c8_3561, RIaf02940_3562, RIaf029b8_3563, RIaf02a30_3564, RIaf02aa8_3565, RIaf02b20_3566, RIaf02b98_3567, RIaf02c10_3568, RIaf02c88_3569, RIaf02d00_3570, RIaf02d78_3571, RIaf02df0_3572, RIaf02e68_3573, RIaf02ee0_3574, RIaf02f58_3575, RIaf02fd0_3576, RIaf03048_3577, RIaf030c0_3578, RIaf03138_3579, RIaf031b0_3580, RIaf03228_3581, RIaf032a0_3582, RIaf03318_3583, RIaf03390_3584);
and \U$57 ( \4772 , RIaf03408_3585, RIaf03480_3586, RIaf034f8_3587, RIaf03570_3588, RIaf035e8_3589, RIaf03660_3590, RIaf036d8_3591, RIaf03750_3592, RIaf037c8_3593, RIaf03840_3594, RIaf038b8_3595, RIaf03930_3596, RIaf039a8_3597, RIaf03a20_3598, RIaf03a98_3599, RIaf03b10_3600, RIaf03b88_3601, RIaf03c00_3602, RIaf03c78_3603, RIaf03cf0_3604, RIaf03d68_3605, RIaf03de0_3606, RIaf03e58_3607, RIaf03ed0_3608, RIaf03f48_3609, RIaf03fc0_3610, RIaf04038_3611, RIaf040b0_3612, RIaf04128_3613, RIaf041a0_3614, RIaf04218_3615, RIaf04290_3616, RIaf04308_3617, RIaf04380_3618, RIaf043f8_3619, RIaf04470_3620, RIaf044e8_3621, RIaf04560_3622, RIaf045d8_3623, RIaf04650_3624, RIaf046c8_3625, RIaf04740_3626, RIaf047b8_3627, RIaf04830_3628, RIaf048a8_3629, RIaf04920_3630, RIaf04998_3631, RIaf04a10_3632, RIaf04a88_3633, RIaf04b00_3634, RIaf04b78_3635, RIaf04bf0_3636, RIaf04c68_3637, RIaf04ce0_3638, RIaf04d58_3639, RIaf04dd0_3640, RIaf04e48_3641, RIaf04ec0_3642, RIaf04f38_3643, RIaf04fb0_3644, RIaf05028_3645, RIaf050a0_3646, RIaf05118_3647, RIaf05190_3648);
and \U$58 ( \4773 , RIaf05208_3649, RIaf05280_3650, RIaf052f8_3651, RIaf05370_3652, RIaf053e8_3653, RIaf05460_3654, RIaf054d8_3655, RIaf05550_3656, RIaf055c8_3657, RIaf05640_3658, RIaf056b8_3659, RIaf05730_3660, RIaf057a8_3661, RIaf05820_3662, RIaf05898_3663, RIaf05910_3664, RIaf05988_3665, RIaf05a00_3666, RIaf05a78_3667, RIaf05af0_3668, RIaf05b68_3669, RIaf05be0_3670, RIaf05c58_3671, RIaf05cd0_3672, RIaf05d48_3673, RIaf05dc0_3674, RIaf05e38_3675, RIaf05eb0_3676, RIaf05f28_3677, RIaf05fa0_3678, RIaf06018_3679, RIaf06090_3680, RIaf06108_3681, RIaf06180_3682, RIaf061f8_3683, RIaf06270_3684, RIaf062e8_3685, RIaf06360_3686, RIaf063d8_3687, RIaf06450_3688, RIaf064c8_3689, RIaf06540_3690, RIaf065b8_3691, RIaf06630_3692, RIaf066a8_3693, RIaf06720_3694, RIaf06798_3695, RIaf06810_3696, RIaf06888_3697, RIaf06900_3698, RIaf06978_3699, RIaf069f0_3700, RIaf06a68_3701, RIaf06ae0_3702, RIaf06b58_3703, RIaf06bd0_3704, RIaf06c48_3705, RIaf06cc0_3706, RIaf06d38_3707, RIaf06db0_3708, RIaf06e28_3709, RIaf06ea0_3710, RIaf06f18_3711, RIaf06f90_3712);
and \U$59 ( \4774 , RIaf07008_3713, RIaf07080_3714, RIaf070f8_3715, RIaf07170_3716, RIaf071e8_3717, RIaf07260_3718, RIaf072d8_3719, RIaf07350_3720, RIaf073c8_3721, RIaf07440_3722, RIaf074b8_3723, RIaf07530_3724, RIaf075a8_3725, RIaf07620_3726, RIaf07698_3727, RIaf07710_3728, RIaf07788_3729, RIaf07800_3730, RIaf07878_3731, RIaf078f0_3732, RIaf07968_3733, RIaf079e0_3734, RIaf07a58_3735, RIaf07ad0_3736, RIaf07b48_3737, RIaf07bc0_3738, RIaf07c38_3739, RIaf07cb0_3740, RIaf07d28_3741, RIaf07da0_3742, RIaf07e18_3743, RIaf07e90_3744, RIaf07f08_3745, RIaf07f80_3746, RIaf07ff8_3747, RIaf08070_3748, RIaf080e8_3749, RIaf08160_3750, RIaf081d8_3751, RIaf08250_3752, RIaf082c8_3753, RIaf08340_3754, RIaf083b8_3755, RIaf08430_3756, RIaf084a8_3757, RIaf08520_3758, RIaf08598_3759, RIaf08610_3760, RIaf08688_3761, RIaf08700_3762, RIaf08778_3763, RIaf087f0_3764, RIaf08868_3765, RIaf088e0_3766, RIaf08958_3767, RIaf089d0_3768, RIaf08a48_3769, RIaf08ac0_3770, RIaf08b38_3771, RIaf08bb0_3772, RIaf08c28_3773, RIaf08ca0_3774, RIaf08d18_3775, RIaf08d90_3776);
and \U$60 ( \4775 , RIaf08e08_3777, RIaf08e80_3778, RIaf08ef8_3779, RIaf08f70_3780, RIaf08fe8_3781, RIaf09060_3782, RIaf090d8_3783, RIaf09150_3784, RIaf091c8_3785, RIaf09240_3786, RIaf092b8_3787, RIaf09330_3788, RIaf093a8_3789, RIaf09420_3790, RIaf09498_3791, RIaf09510_3792, RIaf09588_3793, RIaf09600_3794, RIaf09678_3795, RIaf096f0_3796, RIaf09768_3797, RIaf097e0_3798, RIaf09858_3799, RIaf098d0_3800, RIaf09948_3801, RIaf099c0_3802, RIaf09a38_3803, RIaf09ab0_3804, RIaf09b28_3805, RIaf09ba0_3806, RIaf09c18_3807, RIaf09c90_3808, RIaf09d08_3809, RIaf09d80_3810, RIaf09df8_3811, RIaf09e70_3812, RIaf09ee8_3813, RIaf09f60_3814, RIaf09fd8_3815, RIaf0a050_3816, RIaf0a0c8_3817, RIaf0a140_3818, RIaf0a1b8_3819, RIaf0a230_3820, RIaf0a2a8_3821, RIaf0a320_3822, RIaf0a398_3823, RIaf0a410_3824, RIaf0a488_3825, RIaf0a500_3826, RIaf0a578_3827, RIaf0a5f0_3828, RIaf0a668_3829, RIaf0a6e0_3830, RIaf0a758_3831, RIaf0a7d0_3832, RIaf0a848_3833, RIaf0a8c0_3834, RIaf0a938_3835, RIaf0a9b0_3836, RIaf0aa28_3837, RIaf0aaa0_3838, RIaf0ab18_3839, RIaf0ab90_3840);
and \U$61 ( \4776 , RIaf0ac08_3841, RIaf0ac80_3842, RIaf0acf8_3843, RIaf0ad70_3844, RIaf0ade8_3845, RIaf0ae60_3846, RIaf0aed8_3847, RIaf0af50_3848, RIaf0afc8_3849, RIaf0b040_3850, RIaf0b0b8_3851, RIaf0b130_3852, RIaf0b1a8_3853, RIaf0b220_3854, RIaf0b298_3855, RIaf0b310_3856, RIaf0b388_3857, RIaf0b400_3858, RIaf0b478_3859, RIaf0b4f0_3860, RIaf0b568_3861, RIaf0b5e0_3862, RIaf0b658_3863, RIaf0b6d0_3864, RIaf0b748_3865, RIaf0b7c0_3866, RIaf0b838_3867, RIaf0b8b0_3868, RIaf0b928_3869, RIaf0b9a0_3870, RIaf0ba18_3871, RIaf0ba90_3872, RIaf0bb08_3873, RIaf0bb80_3874, RIaf0bbf8_3875, RIaf0bc70_3876, RIaf0bce8_3877, RIaf0bd60_3878, RIaf0bdd8_3879, RIaf0be50_3880, RIaf0bec8_3881, RIaf0bf40_3882, RIaf0bfb8_3883, RIaf0c030_3884, RIaf0c0a8_3885, RIaf0c120_3886, RIaf0c198_3887, RIaf0c210_3888, RIaf0c288_3889, RIaf0c300_3890, RIaf0c378_3891, RIaf0c3f0_3892, RIaf0c468_3893, RIaf0c4e0_3894, RIaf0c558_3895, RIaf0c5d0_3896, RIaf0c648_3897, RIaf0c6c0_3898, RIaf0c738_3899, RIaf0c7b0_3900, RIaf0c828_3901, RIaf0c8a0_3902, RIaf0c918_3903, RIaf0c990_3904);
and \U$62 ( \4777 , RIaf0ca08_3905, RIaf0ca80_3906, RIaf0caf8_3907, RIaf0cb70_3908, RIaf0cbe8_3909, RIaf0cc60_3910, RIaf0ccd8_3911, RIaf0cd50_3912, RIaf0cdc8_3913, RIaf0ce40_3914, RIaf0ceb8_3915, RIaf0cf30_3916, RIaf0cfa8_3917, RIaf0d020_3918, RIaf0d098_3919, RIaf0d110_3920, RIaf0d188_3921, RIaf0d200_3922, RIaf0d278_3923, RIaf0d2f0_3924, RIaf0d368_3925, RIaf0d3e0_3926, RIaf0d458_3927, RIaf0d4d0_3928, RIaf0d548_3929, RIaf0d5c0_3930, RIaf0d638_3931, RIaf0d6b0_3932, RIaf0d728_3933, RIaf0d7a0_3934, RIaf0d818_3935, RIaf0d890_3936, RIaf0d908_3937, RIaf0d980_3938, RIaf0d9f8_3939, RIaf0da70_3940, RIaf0dae8_3941, RIaf0db60_3942, RIaf0dbd8_3943, RIaf0dc50_3944, RIaf0dcc8_3945, RIaf0dd40_3946, RIaf0ddb8_3947, RIaf0de30_3948, RIaf0dea8_3949, RIaf0df20_3950, RIaf0df98_3951, RIaf0e010_3952, RIaf0e088_3953, RIaf0e100_3954, RIaf0e178_3955, RIaf0e1f0_3956, RIaf0e268_3957, RIaf0e2e0_3958, RIaf0e358_3959, RIaf0e3d0_3960, RIaf0e448_3961, RIaf0e4c0_3962, RIaf0e538_3963, RIaf0e5b0_3964, RIaf0e628_3965, RIaf0e6a0_3966, RIaf0e718_3967, RIaf0e790_3968);
and \U$63 ( \4778 , RIaf0e808_3969, RIaf0e880_3970, RIaf0e8f8_3971, RIaf0e970_3972, RIaf0e9e8_3973, RIaf0ea60_3974, RIaf0ead8_3975, RIaf0eb50_3976, RIaf0ebc8_3977, RIaf0ec40_3978, RIaf0ecb8_3979, RIaf0ed30_3980, RIaf0eda8_3981, RIaf0ee20_3982, RIaf0ee98_3983, RIaf0ef10_3984, RIaf0ef88_3985, RIaf0f000_3986, RIaf0f078_3987, RIaf0f0f0_3988, RIaf0f168_3989, RIaf0f1e0_3990, RIaf0f258_3991, RIaf0f2d0_3992, RIaf0f348_3993, RIaf0f3c0_3994, RIaf0f438_3995, RIaf0f4b0_3996, RIaf0f528_3997, RIaf0f5a0_3998, RIaf0f618_3999, RIaf0f690_4000, RIaf0f708_4001, RIaf0f780_4002, RIaf0f7f8_4003, RIaf0f870_4004, RIaf0f8e8_4005, RIaf0f960_4006, RIaf0f9d8_4007, RIaf0fa50_4008, RIaf0fac8_4009, RIaf0fb40_4010, RIaf0fbb8_4011, RIaf0fc30_4012, RIaf0fca8_4013, RIaf0fd20_4014, RIaf0fd98_4015, RIaf0fe10_4016, RIaf0fe88_4017, RIaf0ff00_4018, RIaf0ff78_4019, RIaf0fff0_4020, RIaf10068_4021, RIaf100e0_4022, RIaf10158_4023, RIaf101d0_4024, RIaf10248_4025, RIaf102c0_4026, RIaf10338_4027, RIaf103b0_4028, RIaf10428_4029, RIaf104a0_4030, RIaf10518_4031, RIaf10590_4032);
and \U$64 ( \4779 , RIaf10608_4033, RIaf10680_4034, RIaf106f8_4035, RIaf10770_4036, RIaf107e8_4037, RIaf10860_4038, RIaf108d8_4039, RIaf10950_4040, RIaf109c8_4041, RIaf10a40_4042, RIaf10ab8_4043, RIaf10b30_4044, RIaf10ba8_4045, RIaf10c20_4046, RIaf10c98_4047, RIaf10d10_4048, RIaf10d88_4049, RIaf10e00_4050, RIaf10e78_4051, RIaf10ef0_4052, RIaf10f68_4053, RIaf10fe0_4054, RIaf11058_4055, RIaf110d0_4056, RIaf11148_4057, RIaf111c0_4058, RIaf11238_4059, RIaf112b0_4060, RIaf11328_4061, RIaf113a0_4062, RIaf11418_4063, RIaf11490_4064, RIaf11508_4065, RIaf11580_4066, RIaf115f8_4067, RIaf11670_4068, RIaf116e8_4069, RIaf11760_4070, RIaf117d8_4071, RIaf11850_4072, RIaf118c8_4073, RIaf11940_4074, RIaf119b8_4075, RIaf11a30_4076, RIaf11aa8_4077, RIaf11b20_4078, RIaf11b98_4079, RIaf11c10_4080, RIaf11c88_4081, RIaf11d00_4082, RIaf11d78_4083, RIaf11df0_4084, RIaf11e68_4085, RIaf11ee0_4086, RIaf11f58_4087, RIaf11fd0_4088, RIaf12048_4089, RIaf120c0_4090, RIaf12138_4091, RIaf121b0_4092, RIaf12228_4093, RIaf122a0_4094, RIaf12318_4095, RIaf12390_4096);
and \U$65 ( \4780 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 );
and \U$66 ( \4781 , RIaf12408_4097, RIaf12480_4098, RIaf124f8_4099, RIaf12570_4100, RIaf125e8_4101, RIaf12660_4102, RIaf126d8_4103, RIaf12750_4104, RIaf127c8_4105, RIaf12840_4106, RIaf128b8_4107, RIaf12930_4108, RIaf129a8_4109, RIaf12a20_4110, RIaf12a98_4111, RIaf12b10_4112, RIaf12b88_4113, RIaf12c00_4114, RIaf12c78_4115, RIaf12cf0_4116, RIaf12d68_4117, RIaf12de0_4118, RIaf12e58_4119, RIaf12ed0_4120, RIaf12f48_4121, RIaf12fc0_4122, RIaf13038_4123, RIaf130b0_4124, RIaf13128_4125, RIaf131a0_4126, RIaf13218_4127, RIaf13290_4128, RIaf13308_4129, RIaf13380_4130, RIaf133f8_4131, RIaf13470_4132, RIaf134e8_4133, RIaf13560_4134, RIaf135d8_4135, RIaf13650_4136, RIaf136c8_4137, RIaf13740_4138, RIaf137b8_4139, RIaf13830_4140, RIaf138a8_4141, RIaf13920_4142, RIaf13998_4143, RIaf13a10_4144, RIaf13a88_4145, RIaf13b00_4146, RIaf13b78_4147, RIaf13bf0_4148, RIaf13c68_4149, RIaf13ce0_4150, RIaf13d58_4151, RIaf13dd0_4152, RIaf13e48_4153, RIaf13ec0_4154, RIaf13f38_4155, RIaf13fb0_4156, RIaf14028_4157, RIaf140a0_4158, RIaf14118_4159, RIaf14190_4160);
and \U$67 ( \4782 , RIaf14208_4161, RIaf14280_4162, RIaf142f8_4163, RIaf14370_4164, RIaf143e8_4165, RIaf14460_4166, RIaf144d8_4167, RIaf14550_4168, RIaf145c8_4169, RIaf14640_4170, RIaf146b8_4171, RIaf14730_4172, RIaf147a8_4173, RIaf14820_4174, RIaf14898_4175, RIaf14910_4176, RIaf14988_4177, RIaf14a00_4178, RIaf14a78_4179, RIaf14af0_4180, RIaf14b68_4181, RIaf14be0_4182, RIaf14c58_4183, RIaf14cd0_4184, RIaf14d48_4185, RIaf14dc0_4186, RIaf14e38_4187, RIaf14eb0_4188, RIaf14f28_4189, RIaf14fa0_4190, RIaf15018_4191, RIaf15090_4192, RIaf15108_4193, RIaf15180_4194, RIaf151f8_4195, RIaf15270_4196, RIaf152e8_4197, RIaf15360_4198, RIaf153d8_4199, RIaf15450_4200, RIaf154c8_4201, RIaf15540_4202, RIaf155b8_4203, RIaf15630_4204, RIaf156a8_4205, RIaf15720_4206, RIaf15798_4207, RIaf15810_4208, RIaf15888_4209, RIaf15900_4210, RIaf15978_4211, RIaf159f0_4212, RIaf15a68_4213, RIaf15ae0_4214, RIaf15b58_4215, RIaf15bd0_4216, RIaf15c48_4217, RIaf15cc0_4218, RIaf15d38_4219, RIaf15db0_4220, RIaf15e28_4221, RIaf15ea0_4222, RIaf15f18_4223, RIaf15f90_4224);
and \U$68 ( \4783 , RIaf16008_4225, RIaf16080_4226, RIaf160f8_4227, RIaf16170_4228, RIaf161e8_4229, RIaf16260_4230, RIaf162d8_4231, RIaf16350_4232, RIaf163c8_4233, RIaf16440_4234, RIaf164b8_4235, RIaf16530_4236, RIaf165a8_4237, RIaf16620_4238, RIaf16698_4239, RIaf16710_4240, RIaf16788_4241, RIaf16800_4242, RIaf16878_4243, RIaf168f0_4244, RIaf16968_4245, RIaf169e0_4246, RIaf16a58_4247, RIaf16ad0_4248, RIaf16b48_4249, RIaf16bc0_4250, RIaf16c38_4251, RIaf16cb0_4252, RIaf16d28_4253, RIaf16da0_4254, RIaf16e18_4255, RIaf16e90_4256, RIaf16f08_4257, RIaf16f80_4258, RIaf16ff8_4259, RIaf17070_4260, RIaf170e8_4261, RIaf17160_4262, RIaf171d8_4263, RIaf17250_4264, RIaf172c8_4265, RIaf17340_4266, RIaf173b8_4267, RIaf17430_4268, RIaf174a8_4269, RIaf17520_4270, RIaf17598_4271, RIaf17610_4272, RIaf17688_4273, RIaf17700_4274, RIaf17778_4275, RIaf177f0_4276, RIaf17868_4277, RIaf178e0_4278, RIaf17958_4279, RIaf179d0_4280, RIaf17a48_4281, RIaf17ac0_4282, RIaf17b38_4283, RIaf17bb0_4284, RIaf17c28_4285, RIaf17ca0_4286, RIaf17d18_4287, RIaf17d90_4288);
and \U$69 ( \4784 , RIaf17e08_4289, RIaf17e80_4290, RIaf17ef8_4291, RIaf17f70_4292, RIaf17fe8_4293, RIaf18060_4294, RIaf180d8_4295, RIaf18150_4296, RIaf181c8_4297, RIaf18240_4298, RIaf182b8_4299, RIaf18330_4300, RIaf183a8_4301, RIaf18420_4302, RIaf18498_4303, RIaf18510_4304, RIaf18588_4305, RIaf18600_4306, RIaf18678_4307, RIaf186f0_4308, RIaf18768_4309, RIaf187e0_4310, RIaf18858_4311, RIaf188d0_4312, RIaf18948_4313, RIaf189c0_4314, RIaf18a38_4315, RIaf18ab0_4316, RIaf18b28_4317, RIaf18ba0_4318, RIaf18c18_4319, RIaf18c90_4320, RIaf18d08_4321, RIaf18d80_4322, RIaf18df8_4323, RIaf18e70_4324, RIaf18ee8_4325, RIaf18f60_4326, RIaf18fd8_4327, RIaf19050_4328, RIaf190c8_4329, RIaf19140_4330, RIaf191b8_4331, RIaf19230_4332, RIaf192a8_4333, RIaf19320_4334, RIaf19398_4335, RIaf19410_4336, RIaf19488_4337, RIaf19500_4338, RIaf19578_4339, RIaf195f0_4340, RIaf19668_4341, RIaf196e0_4342, RIaf19758_4343, RIaf197d0_4344, RIaf19848_4345, RIaf198c0_4346, RIaf19938_4347, RIaf199b0_4348, RIaf19a28_4349, RIaf19aa0_4350, RIaf19b18_4351, RIaf19b90_4352);
and \U$70 ( \4785 , RIaf19c08_4353, RIaf19c80_4354, RIaf19cf8_4355, RIaf19d70_4356, RIaf19de8_4357, RIaf19e60_4358, RIaf19ed8_4359, RIaf19f50_4360, RIaf19fc8_4361, RIaf1a040_4362, RIaf1a0b8_4363, RIaf1a130_4364, RIaf1a1a8_4365, RIaf1a220_4366, RIaf1a298_4367, RIaf1a310_4368, RIaf1a388_4369, RIaf1a400_4370, RIaf1a478_4371, RIaf1a4f0_4372, RIaf1a568_4373, RIaf1a5e0_4374, RIaf1a658_4375, RIaf1a6d0_4376, RIaf1a748_4377, RIaf1a7c0_4378, RIaf1a838_4379, RIaf1a8b0_4380, RIaf1a928_4381, RIaf1a9a0_4382, RIaf1aa18_4383, RIaf1aa90_4384, RIaf1ab08_4385, RIaf1ab80_4386, RIaf1abf8_4387, RIaf1ac70_4388, RIaf1ace8_4389, RIaf1ad60_4390, RIaf1add8_4391, RIaf1ae50_4392, RIaf1aec8_4393, RIaf1af40_4394, RIaf1afb8_4395, RIaf1b030_4396, RIaf1b0a8_4397, RIaf1b120_4398, RIaf1b198_4399, RIaf1b210_4400, RIaf1b288_4401, RIaf1b300_4402, RIaf1b378_4403, RIaf1b3f0_4404, RIaf1b468_4405, RIaf1b4e0_4406, RIaf1b558_4407, RIaf1b5d0_4408, RIaf1b648_4409, RIaf1b6c0_4410, RIaf1b738_4411, RIaf1b7b0_4412, RIaf1b828_4413, RIaf1b8a0_4414, RIaf1b918_4415, RIaf1b990_4416);
and \U$71 ( \4786 , RIaf1ba08_4417, RIaf1ba80_4418, RIaf1baf8_4419, RIaf1bb70_4420, RIaf1bbe8_4421, RIaf1bc60_4422, RIaf1bcd8_4423, RIaf1bd50_4424, RIaf1bdc8_4425, RIaf1be40_4426, RIaf1beb8_4427, RIaf1bf30_4428, RIaf1bfa8_4429, RIaf1c020_4430, RIaf1c098_4431, RIaf1c110_4432, RIaf1c188_4433, RIaf1c200_4434, RIaf1c278_4435, RIaf1c2f0_4436, RIaf1c368_4437, RIaf1c3e0_4438, RIaf1c458_4439, RIaf1c4d0_4440, RIaf1c548_4441, RIaf1c5c0_4442, RIaf1c638_4443, RIaf1c6b0_4444, RIaf1c728_4445, RIaf1c7a0_4446, RIaf1c818_4447, RIaf1c890_4448, RIaf1c908_4449, RIaf1c980_4450, RIaf1c9f8_4451, RIaf1ca70_4452, RIaf1cae8_4453, RIaf1cb60_4454, RIaf1cbd8_4455, RIaf1cc50_4456, RIaf1ccc8_4457, RIaf1cd40_4458, RIaf1cdb8_4459, RIaf1ce30_4460, RIaf1cea8_4461, RIaf1cf20_4462, RIaf1cf98_4463, RIaf1d010_4464, RIaf1d088_4465, RIaf1d100_4466, RIaf1d178_4467, RIaf1d1f0_4468, RIaf1d268_4469, RIaf1d2e0_4470, RIaf1d358_4471, RIaf1d3d0_4472, RIaf1d448_4473, RIaf1d4c0_4474, RIaf1d538_4475, RIaf1d5b0_4476, RIaf1d628_4477, RIaf1d6a0_4478, RIaf1d718_4479, RIaf1d790_4480);
and \U$72 ( \4787 , RIaf1d808_4481, RIaf1d880_4482, RIaf1d8f8_4483, RIaf1d970_4484, RIaf1d9e8_4485, RIaf1da60_4486, RIaf1dad8_4487, RIaf1db50_4488, RIaf1dbc8_4489, RIaf1dc40_4490, RIaf1dcb8_4491, RIaf1dd30_4492, RIaf1dda8_4493, RIaf1de20_4494, RIaf1de98_4495, RIaf1df10_4496, RIaf1df88_4497, RIaf1e000_4498, RIaf1e078_4499, RIaf1e0f0_4500, RIaf1e168_4501, RIaf1e1e0_4502, RIaf1e258_4503, RIaf1e2d0_4504, RIaf1e348_4505, RIaf1e3c0_4506, RIaf1e438_4507, RIaf1e4b0_4508, RIaf1e528_4509, RIaf1e5a0_4510, RIaf1e618_4511, RIaf1e690_4512, RIaf1e708_4513, RIaf1e780_4514, RIaf1e7f8_4515, RIaf1e870_4516, RIaf1e8e8_4517, RIaf1e960_4518, RIaf1e9d8_4519, RIaf1ea50_4520, RIaf1eac8_4521, RIaf1eb40_4522, RIaf1ebb8_4523, RIaf1ec30_4524, RIaf1eca8_4525, RIaf1ed20_4526, RIaf1ed98_4527, RIaf1ee10_4528, RIaf1ee88_4529, RIaf1ef00_4530, RIaf1ef78_4531, RIaf1eff0_4532, RIaf1f068_4533, RIaf1f0e0_4534, RIaf1f158_4535, RIaf1f1d0_4536, RIaf1f248_4537, RIaf1f2c0_4538, RIaf1f338_4539, RIaf1f3b0_4540, RIaf1f428_4541, RIaf1f4a0_4542, RIaf1f518_4543, RIaf1f590_4544);
and \U$73 ( \4788 , RIaf1f608_4545, RIaf1f680_4546, RIaf1f6f8_4547, RIaf1f770_4548, RIaf1f7e8_4549, RIaf1f860_4550, RIaf1f8d8_4551, RIaf1f950_4552, RIaf1f9c8_4553, RIaf1fa40_4554, RIaf1fab8_4555, RIaf1fb30_4556, RIaf1fba8_4557, RIaf1fc20_4558, RIaf1fc98_4559, RIaf1fd10_4560, RIaf1fd88_4561, RIaf1fe00_4562, RIaf1fe78_4563, RIaf1fef0_4564, RIaf1ff68_4565, RIaf1ffe0_4566, RIaf20058_4567, RIaf200d0_4568, RIaf20148_4569, RIaf201c0_4570, RIaf20238_4571, RIaf202b0_4572, RIaf20328_4573, RIaf203a0_4574, RIaf20418_4575, RIaf20490_4576, RIaf20508_4577, RIaf20580_4578, RIaf205f8_4579, RIaf20670_4580, RIaf206e8_4581, RIaf20760_4582, RIaf207d8_4583, RIaf20850_4584, RIaf208c8_4585, RIaf20940_4586, RIaf209b8_4587, RIaf20a30_4588, RIaf20aa8_4589, RIaf20b20_4590, RIaf20b98_4591, RIaf20c10_4592, RIaf20c88_4593, RIaf20d00_4594, RIaf20d78_4595, RIaf20df0_4596, RIaf20e68_4597, RIaf20ee0_4598, RIaf20f58_4599, RIaf20fd0_4600, RIaf21048_4601, RIaf210c0_4602, RIaf21138_4603, RIaf211b0_4604, RIaf21228_4605, RIaf212a0_4606, RIaf21318_4607, RIaf21390_4608);
and \U$74 ( \4789 , RIaf21408_4609, RIaf21480_4610, RIaf214f8_4611, RIaf21570_4612, RIaf215e8_4613, RIaf21660_4614, RIaf216d8_4615, RIaf21750_4616, RIaf217c8_4617, RIaf21840_4618, RIaf218b8_4619, RIaf21930_4620, RIaf219a8_4621, RIaf21a20_4622, RIaf21a98_4623, RIaf21b10_4624, RIaf21b88_4625, RIaf21c00_4626, RIaf21c78_4627, RIaf21cf0_4628, RIaf21d68_4629, RIaf21de0_4630, RIaf21e58_4631, RIaf21ed0_4632, RIaf21f48_4633, RIaf21fc0_4634, RIaf22038_4635, RIaf220b0_4636, RIaf22128_4637, RIaf221a0_4638, RIaf22218_4639, RIaf22290_4640, RIaf22308_4641, RIaf22380_4642, RIaf223f8_4643, RIaf22470_4644, RIaf224e8_4645, RIaf22560_4646, RIaf225d8_4647, RIaf22650_4648, RIaf226c8_4649, RIaf22740_4650, RIaf227b8_4651, RIaf22830_4652, RIaf228a8_4653, RIaf22920_4654, RIaf22998_4655, RIaf22a10_4656, RIaf22a88_4657, RIaf22b00_4658, RIaf22b78_4659, RIaf22bf0_4660, RIaf22c68_4661, RIaf22ce0_4662, RIaf22d58_4663, RIaf22dd0_4664, RIaf22e48_4665, RIaf22ec0_4666, RIaf22f38_4667, RIaf22fb0_4668, RIaf23028_4669, RIaf230a0_4670, RIaf23118_4671, RIaf23190_4672);
and \U$75 ( \4790 , RIaf23208_4673, RIaf23280_4674, RIaf232f8_4675, RIaf23370_4676, RIaf233e8_4677, RIaf23460_4678, RIaf234d8_4679, RIaf23550_4680);
and \U$76 ( \4791 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 );
buf \U$77 ( \4792 , \4791 );
endmodule

