//
// Conformal-LEC Version 20.10-d213 (02-Sep-2020)
//
module top(RI986e350_15,RI986e3c8_16,RI986e260_13,RI986e2d8_14,RI986e080_9,RI986e0f8_10,RI986e170_11,RI986e1e8_12,RI986dcc0_1,
        RI986dd38_2,RI986dea0_5,RI986df18_6,RI986df90_7,RI986e008_8,RI986de28_4,RI986ddb0_3,RI986ef80_41,RI986eff8_42,RI986f070_43,
        RI986f0e8_44,RI986f250_47,RI986f2c8_48,RI986f160_45,RI986f1d8_46,RI986e878_26,RI986e800_25,RI986e9e0_29,RI986ea58_30,RI986ead0_31,
        RI986eb48_32,RI986e8f0_27,RI986e968_28,RI986ebc0_33,RI986ec38_34,RI986ecb0_35,RI986ed28_36,RI986eda0_37,RI986ee18_38,RI986ee90_39,
        RI986ef08_40,RI986e710_23,RI986e788_24,RI986e620_21,RI986e698_22,RI986e530_19,RI986e5a8_20,RI986e440_17,RI986e4b8_18,RI986ffe8_76,
        RI986ff70_75,RI9870060_77,RI98700d8_78,RI986fe80_73,RI986fef8_74,RI9870150_79,RI98701c8_80,RI986fca0_69,RI986fd18_70,RI986fd90_71,
        RI986fe08_72,RI986fbb0_67,RI986fc28_68,RI986fac0_65,RI986fb38_66,RI9870240_81,RI98702b8_82,RI9870330_83,RI98703a8_84,RI9870420_85,
        RI9870498_86,RI9870510_87,RI9870588_88,RI98707e0_93,RI9870858_94,RI9870600_89,RI9870678_90,RI98708d0_95,RI9870948_96,RI9870768_92,
        RI98706f0_91,RI9871050_111,RI98710c8_112,RI9870e70_107,RI9870ee8_108,RI9870ba0_101,RI9870c18_102,RI9870f60_109,RI9870fd8_110,RI9870ab0_99,
        RI9870b28_100,RI98709c0_97,RI9870a38_98,RI9870d80_105,RI9870df8_106,RI9870c90_103,RI9870d08_104,RI9871398_118,RI9871320_117,RI9871230_115,
        RI98712a8_116,RI9871140_113,RI98711b8_114,RI9871410_119,RI9871488_120,RI98716e0_125,RI9871758_126,RI98717d0_127,RI9871848_128,RI98715f0_123,
        RI9871668_124,RI9871500_121,RI9871578_122,RI986f700_57,RI986f778_58,RI986f868_60,RI986f7f0_59,RI986f9d0_63,RI986fa48_64,RI986f340_49,
        RI986f3b8_50,RI986f430_51,RI986f4a8_52,RI986f598_54,RI986f520_53,RI986f688_56,RI986f610_55,RI986f8e0_61,RI986f958_62,RI98719b0_131,
        RI9871aa0_133,RI9871a28_132,RI9871d70_139,RI9872130_147,RI9872220_149,RI9871c80_137,RI98721a8_148,RI9871ed8_142,RI9871f50_143,RI9871e60_141,
        RI98718c0_129,RI9871938_130,RI9872040_145,RI9871fc8_144,RI9871b18_134,RI9871b90_135,RI9871c08_136,RI9871de8_140,RI9872298_150,RI9872310_151,
        RI98720b8_146,RI9871cf8_138,RI98726d0_159,RI9872748_160,RI98725e0_157,RI9872658_158,RI9872388_152,RI98727c0_161,RI9872400_153,RI9872478_154,
        RI98724f0_155,RI9872568_156,RI9872838_162,RI98728b0_163,RI9872928_164,RI98729a0_165,RI9872a18_166,RI9872a90_167,RI9872b08_168,RI9872b80_169,
        RI9872f40_177,RI9872fb8_178,RI9873030_179,RI9872e50_175,RI9872dd8_174,RI9872d60_173,RI9872bf8_170,RI9872c70_171,RI9872ce8_172,RI9872ec8_176,
        RI98730a8_180,RI9873120_181,RI9873210_183,RI9873198_182,RI9873288_184,RI9873300_185,RI9873378_186,RI98733f0_187,RI9873558_190,RI98735d0_191,
        RI98734e0_189,RI9873468_188,RI9873648_192,RI9874020_213,RI9874098_214,RI9875100_249,RI9875178_250,RI98751f0_251,RI9875268_252,RI9874200_217,
        RI9874278_218,RI9874b60_237,RI9874bd8_238,RI9874c50_239,RI9874cc8_240,RI9874110_215,RI9874188_216,RI98736c0_193,RI9873738_194,RI9873a08_200,
        RI9873990_199,RI98738a0_197,RI9873918_198,RI9873c60_205,RI9873cd8_206,RI9873dc8_208,RI9873d50_207,RI9874f20_245,RI9874f98_246,RI9875010_247,
        RI9875088_248,RI9874d40_241,RI9874db8_242,RI9874e30_243,RI9874ea8_244,RI98742f0_219,RI9874368_220,RI9874890_231,RI9874908_232,RI98752e0_253,
        RI9875358_254,RI98747a0_229,RI9874818_230,RI98743e0_221,RI9874458_222,RI9874548_224,RI98744d0_223,RI9873fa8_212,RI9873f30_211,RI9873e40_209,
        RI9873eb8_210,RI98737b0_195,RI9873828_196,RI98753d0_255,RI9875448_256,RI9873a80_201,RI9873af8_202,RI9873b70_203,RI9873be8_204,RI9874980_233,
        RI98749f8_234,RI9874ae8_236,RI9874a70_235,RI98746b0_227,RI9874728_228,RI98745c0_225,RI9874638_226,R_101_8a8e950,R_102_8a8f868,R_103_8a8f910,
        R_104_8a8f9b8,R_105_8a8fa60,R_106_8a8fb08,R_107_8a8fbb0,R_108_8a8fc58,R_109_8a8fd00,R_10a_8a8fda8,R_10b_8a8fe50,R_10c_8a8fef8,R_10d_8a8ffa0,
        R_10e_8a90048,R_10f_8a900f0,R_110_8a90198,R_111_8a90240,R_112_8a902e8,R_113_8a90390,R_114_8a90438,R_115_8a904e0,R_116_8a90588,R_117_8a90630,
        R_118_8a906d8,R_119_8a90780,R_11a_8a90828,R_11b_8a908d0,R_11c_8a90978,R_11d_8a90a20,R_11e_8a90ac8,R_11f_8a90b70,R_120_8a90c18,R_121_8a90cc0,
        R_122_8a90d68,R_123_8a90e10,R_124_8a90eb8,R_125_8a90f60,R_126_8a91008,R_127_8a910b0,R_128_8a91158,R_129_8a91200,R_12a_8a912a8,R_12b_8a91350,
        R_12c_8a913f8,R_12d_8a914a0,R_12e_8a91548,R_12f_8a915f0,R_130_8a91698,R_131_8a91740,R_132_8a917e8,R_133_8a91890,R_134_8a91938,R_135_8a919e0,
        R_136_8a91a88,R_137_8a91b30,R_138_8a91bd8,R_139_8a91c80,R_13a_8a91d28,R_13b_8a91dd0,R_13c_8a91e78,R_13d_8a91f20,R_13e_8a91fc8,R_13f_8a92070,
        R_140_8a92118,R_141_8a921c0,R_142_8a92268,R_143_8a92310,R_144_8a923b8,R_145_8a92460,R_146_8a92508,R_147_8a925b0,R_148_8a92658,R_149_8a92700,
        R_14a_8a927a8,R_14b_8a92850,R_14c_8a928f8,R_14d_8a929a0,R_14e_8a92a48,R_14f_8a92af0,R_150_8a92b98,R_151_8a92c40,R_152_8a92ce8,R_153_8a92d90,
        R_154_8a92e38,R_155_8a92ee0);
input RI986e350_15,RI986e3c8_16,RI986e260_13,RI986e2d8_14,RI986e080_9,RI986e0f8_10,RI986e170_11,RI986e1e8_12,RI986dcc0_1,
        RI986dd38_2,RI986dea0_5,RI986df18_6,RI986df90_7,RI986e008_8,RI986de28_4,RI986ddb0_3,RI986ef80_41,RI986eff8_42,RI986f070_43,
        RI986f0e8_44,RI986f250_47,RI986f2c8_48,RI986f160_45,RI986f1d8_46,RI986e878_26,RI986e800_25,RI986e9e0_29,RI986ea58_30,RI986ead0_31,
        RI986eb48_32,RI986e8f0_27,RI986e968_28,RI986ebc0_33,RI986ec38_34,RI986ecb0_35,RI986ed28_36,RI986eda0_37,RI986ee18_38,RI986ee90_39,
        RI986ef08_40,RI986e710_23,RI986e788_24,RI986e620_21,RI986e698_22,RI986e530_19,RI986e5a8_20,RI986e440_17,RI986e4b8_18,RI986ffe8_76,
        RI986ff70_75,RI9870060_77,RI98700d8_78,RI986fe80_73,RI986fef8_74,RI9870150_79,RI98701c8_80,RI986fca0_69,RI986fd18_70,RI986fd90_71,
        RI986fe08_72,RI986fbb0_67,RI986fc28_68,RI986fac0_65,RI986fb38_66,RI9870240_81,RI98702b8_82,RI9870330_83,RI98703a8_84,RI9870420_85,
        RI9870498_86,RI9870510_87,RI9870588_88,RI98707e0_93,RI9870858_94,RI9870600_89,RI9870678_90,RI98708d0_95,RI9870948_96,RI9870768_92,
        RI98706f0_91,RI9871050_111,RI98710c8_112,RI9870e70_107,RI9870ee8_108,RI9870ba0_101,RI9870c18_102,RI9870f60_109,RI9870fd8_110,RI9870ab0_99,
        RI9870b28_100,RI98709c0_97,RI9870a38_98,RI9870d80_105,RI9870df8_106,RI9870c90_103,RI9870d08_104,RI9871398_118,RI9871320_117,RI9871230_115,
        RI98712a8_116,RI9871140_113,RI98711b8_114,RI9871410_119,RI9871488_120,RI98716e0_125,RI9871758_126,RI98717d0_127,RI9871848_128,RI98715f0_123,
        RI9871668_124,RI9871500_121,RI9871578_122,RI986f700_57,RI986f778_58,RI986f868_60,RI986f7f0_59,RI986f9d0_63,RI986fa48_64,RI986f340_49,
        RI986f3b8_50,RI986f430_51,RI986f4a8_52,RI986f598_54,RI986f520_53,RI986f688_56,RI986f610_55,RI986f8e0_61,RI986f958_62,RI98719b0_131,
        RI9871aa0_133,RI9871a28_132,RI9871d70_139,RI9872130_147,RI9872220_149,RI9871c80_137,RI98721a8_148,RI9871ed8_142,RI9871f50_143,RI9871e60_141,
        RI98718c0_129,RI9871938_130,RI9872040_145,RI9871fc8_144,RI9871b18_134,RI9871b90_135,RI9871c08_136,RI9871de8_140,RI9872298_150,RI9872310_151,
        RI98720b8_146,RI9871cf8_138,RI98726d0_159,RI9872748_160,RI98725e0_157,RI9872658_158,RI9872388_152,RI98727c0_161,RI9872400_153,RI9872478_154,
        RI98724f0_155,RI9872568_156,RI9872838_162,RI98728b0_163,RI9872928_164,RI98729a0_165,RI9872a18_166,RI9872a90_167,RI9872b08_168,RI9872b80_169,
        RI9872f40_177,RI9872fb8_178,RI9873030_179,RI9872e50_175,RI9872dd8_174,RI9872d60_173,RI9872bf8_170,RI9872c70_171,RI9872ce8_172,RI9872ec8_176,
        RI98730a8_180,RI9873120_181,RI9873210_183,RI9873198_182,RI9873288_184,RI9873300_185,RI9873378_186,RI98733f0_187,RI9873558_190,RI98735d0_191,
        RI98734e0_189,RI9873468_188,RI9873648_192,RI9874020_213,RI9874098_214,RI9875100_249,RI9875178_250,RI98751f0_251,RI9875268_252,RI9874200_217,
        RI9874278_218,RI9874b60_237,RI9874bd8_238,RI9874c50_239,RI9874cc8_240,RI9874110_215,RI9874188_216,RI98736c0_193,RI9873738_194,RI9873a08_200,
        RI9873990_199,RI98738a0_197,RI9873918_198,RI9873c60_205,RI9873cd8_206,RI9873dc8_208,RI9873d50_207,RI9874f20_245,RI9874f98_246,RI9875010_247,
        RI9875088_248,RI9874d40_241,RI9874db8_242,RI9874e30_243,RI9874ea8_244,RI98742f0_219,RI9874368_220,RI9874890_231,RI9874908_232,RI98752e0_253,
        RI9875358_254,RI98747a0_229,RI9874818_230,RI98743e0_221,RI9874458_222,RI9874548_224,RI98744d0_223,RI9873fa8_212,RI9873f30_211,RI9873e40_209,
        RI9873eb8_210,RI98737b0_195,RI9873828_196,RI98753d0_255,RI9875448_256,RI9873a80_201,RI9873af8_202,RI9873b70_203,RI9873be8_204,RI9874980_233,
        RI98749f8_234,RI9874ae8_236,RI9874a70_235,RI98746b0_227,RI9874728_228,RI98745c0_225,RI9874638_226;
output R_101_8a8e950,R_102_8a8f868,R_103_8a8f910,R_104_8a8f9b8,R_105_8a8fa60,R_106_8a8fb08,R_107_8a8fbb0,R_108_8a8fc58,R_109_8a8fd00,
        R_10a_8a8fda8,R_10b_8a8fe50,R_10c_8a8fef8,R_10d_8a8ffa0,R_10e_8a90048,R_10f_8a900f0,R_110_8a90198,R_111_8a90240,R_112_8a902e8,R_113_8a90390,
        R_114_8a90438,R_115_8a904e0,R_116_8a90588,R_117_8a90630,R_118_8a906d8,R_119_8a90780,R_11a_8a90828,R_11b_8a908d0,R_11c_8a90978,R_11d_8a90a20,
        R_11e_8a90ac8,R_11f_8a90b70,R_120_8a90c18,R_121_8a90cc0,R_122_8a90d68,R_123_8a90e10,R_124_8a90eb8,R_125_8a90f60,R_126_8a91008,R_127_8a910b0,
        R_128_8a91158,R_129_8a91200,R_12a_8a912a8,R_12b_8a91350,R_12c_8a913f8,R_12d_8a914a0,R_12e_8a91548,R_12f_8a915f0,R_130_8a91698,R_131_8a91740,
        R_132_8a917e8,R_133_8a91890,R_134_8a91938,R_135_8a919e0,R_136_8a91a88,R_137_8a91b30,R_138_8a91bd8,R_139_8a91c80,R_13a_8a91d28,R_13b_8a91dd0,
        R_13c_8a91e78,R_13d_8a91f20,R_13e_8a91fc8,R_13f_8a92070,R_140_8a92118,R_141_8a921c0,R_142_8a92268,R_143_8a92310,R_144_8a923b8,R_145_8a92460,
        R_146_8a92508,R_147_8a925b0,R_148_8a92658,R_149_8a92700,R_14a_8a927a8,R_14b_8a92850,R_14c_8a928f8,R_14d_8a929a0,R_14e_8a92a48,R_14f_8a92af0,
        R_150_8a92b98,R_151_8a92c40,R_152_8a92ce8,R_153_8a92d90,R_154_8a92e38,R_155_8a92ee0;

wire \342_ZERO , \343_ONE , \344 , \345 , \346 , \347 , \348 , \349 , \350 ,
         \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 ,
         \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 ,
         \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 ,
         \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 ,
         \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 ,
         \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 ,
         \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 ,
         \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 ,
         \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 ,
         \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 ,
         \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 ,
         \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 ,
         \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 ,
         \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 ,
         \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 ,
         \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 ,
         \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 ,
         \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 ,
         \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 ,
         \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 ,
         \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 ,
         \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 ,
         \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 ,
         \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 ,
         \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 ,
         \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 ,
         \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 ,
         \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 ,
         \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 ,
         \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 ,
         \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 ,
         \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 ,
         \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 ,
         \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 ,
         \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 ,
         \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 ,
         \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 ,
         \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 ,
         \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 ,
         \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 ,
         \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 ,
         \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 ,
         \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 ,
         \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 ,
         \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 ,
         \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 ,
         \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 ,
         \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 ,
         \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 ,
         \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 ,
         \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 ,
         \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 ,
         \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 ,
         \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 ,
         \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 ,
         \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 ,
         \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 ,
         \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 ,
         \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 ,
         \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 ,
         \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 ,
         \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 ,
         \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 ,
         \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 ,
         \991 , \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 ,
         \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 ,
         \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 ,
         \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 ,
         \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 ,
         \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 ,
         \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 ,
         \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 ,
         \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 ,
         \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 ,
         \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 ,
         \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 ,
         \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 ,
         \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 ,
         \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 ,
         \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 ,
         \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 ,
         \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 ,
         \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 ,
         \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 ,
         \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 ,
         \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 ,
         \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 ,
         \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 ,
         \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 ,
         \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 ,
         \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 ,
         \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 ,
         \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 ,
         \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 ,
         \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 ,
         \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 ,
         \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 ,
         \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 ,
         \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 ,
         \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 ,
         \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 ,
         \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 ,
         \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 ,
         \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 ,
         \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 ,
         \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 ,
         \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 ,
         \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 ,
         \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 ,
         \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 ,
         \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 ,
         \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 ,
         \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 ,
         \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 ,
         \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 ,
         \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 ,
         \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 ,
         \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 ,
         \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 ,
         \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 ,
         \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 ,
         \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 ,
         \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 ,
         \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 ,
         \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 ,
         \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 ,
         \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 ,
         \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 ,
         \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 ,
         \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 ,
         \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 ,
         \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 ,
         \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 ,
         \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 ,
         \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 ,
         \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 ,
         \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 ,
         \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 ,
         \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 ,
         \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 ,
         \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 ,
         \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 ,
         \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 ,
         \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 ,
         \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 ,
         \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 ,
         \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 ,
         \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 ,
         \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 ,
         \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 ,
         \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 ,
         \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 ,
         \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 ,
         \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 ,
         \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 ,
         \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 ,
         \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 ,
         \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 ,
         \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 ,
         \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 ,
         \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 ,
         \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 ,
         \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 ,
         \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 ,
         \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 ,
         \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 ,
         \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 ,
         \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 ,
         \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 ,
         \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 ,
         \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 ,
         \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 ,
         \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 ,
         \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 ,
         \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 ,
         \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 ,
         \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 ,
         \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 ,
         \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 ,
         \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 ,
         \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 ,
         \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 ,
         \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 ,
         \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 ,
         \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 ,
         \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 ,
         \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 ,
         \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 ,
         \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 ,
         \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 ,
         \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 ,
         \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 ,
         \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 ,
         \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 ,
         \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 ,
         \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 ,
         \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 ,
         \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 ,
         \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 ,
         \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 ,
         \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 ,
         \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 ,
         \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 ,
         \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 ,
         \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 ,
         \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 ,
         \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 ,
         \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 ,
         \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 ,
         \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 ,
         \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 ,
         \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 ,
         \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 ,
         \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 ,
         \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 ,
         \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 ,
         \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 ,
         \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 ,
         \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 ,
         \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 ,
         \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 ,
         \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 ,
         \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 ,
         \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 ,
         \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 ,
         \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 ,
         \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 ,
         \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 ,
         \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 ,
         \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 ,
         \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 ,
         \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 ,
         \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 ,
         \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 ,
         \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 ,
         \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 ,
         \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 ,
         \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 ,
         \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 ,
         \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 ,
         \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 ,
         \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 ,
         \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 ,
         \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 ,
         \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 ,
         \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 ,
         \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 ,
         \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 ,
         \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 ,
         \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 ,
         \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 ,
         \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 ,
         \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 ,
         \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 ,
         \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 ,
         \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 ,
         \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 ,
         \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 ,
         \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 ,
         \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 ,
         \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 ,
         \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 ,
         \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 ,
         \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 ,
         \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 ,
         \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 ,
         \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 ,
         \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 ,
         \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 ,
         \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 ,
         \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 ,
         \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 ,
         \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 ,
         \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 ,
         \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 ,
         \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 ,
         \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 ,
         \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 ,
         \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 ,
         \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 ,
         \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 ,
         \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 ,
         \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 ,
         \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 ,
         \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 ,
         \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 ,
         \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 ,
         \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 ,
         \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 ,
         \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 ,
         \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 ,
         \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 ,
         \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 ,
         \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 ,
         \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 ,
         \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 ,
         \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 ,
         \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 ,
         \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 ,
         \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 ,
         \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 ,
         \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 ,
         \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 ,
         \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 ,
         \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 ,
         \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 ,
         \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 ,
         \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 ,
         \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 ,
         \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 ,
         \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 ,
         \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 ,
         \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 ,
         \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 ,
         \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 ,
         \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 ,
         \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 ,
         \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 ,
         \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 ,
         \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 ,
         \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 ,
         \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 ,
         \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 ,
         \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 ,
         \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 ,
         \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 ,
         \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 ,
         \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 ,
         \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 ,
         \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 ,
         \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 ,
         \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 ,
         \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 ,
         \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 ,
         \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 ,
         \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 ,
         \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 ,
         \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 ,
         \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 ,
         \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 ,
         \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 ,
         \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 ,
         \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 ,
         \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 ,
         \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 ,
         \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 ,
         \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 ,
         \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 ,
         \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 ,
         \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 ,
         \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 ,
         \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 ,
         \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 ,
         \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 ,
         \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 ,
         \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 ,
         \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 ,
         \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 ,
         \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 ,
         \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 ,
         \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 ,
         \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 ,
         \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 ,
         \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 ,
         \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 ,
         \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 ,
         \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 ,
         \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 ,
         \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 ,
         \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 ,
         \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 ,
         \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 ,
         \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 ,
         \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 ,
         \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 ,
         \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 ,
         \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 ,
         \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 ,
         \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 ,
         \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 ,
         \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 ,
         \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 ,
         \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 ,
         \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 ,
         \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 ,
         \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 ,
         \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 ,
         \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 ,
         \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 ,
         \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 ,
         \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 ,
         \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 ,
         \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 ,
         \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 ,
         \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 ,
         \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 ,
         \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 ,
         \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 ,
         \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 ,
         \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 ,
         \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 ,
         \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 ,
         \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 ,
         \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 ,
         \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 ,
         \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 ,
         \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 ,
         \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 ,
         \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 ,
         \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 ,
         \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 ,
         \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 ,
         \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 ,
         \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 ,
         \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 ,
         \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 ,
         \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 ,
         \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 ,
         \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 ,
         \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 ,
         \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 ,
         \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 ,
         \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 ,
         \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 ,
         \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 ,
         \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 ,
         \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 ,
         \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 ,
         \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 ,
         \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 ,
         \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 ,
         \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 ,
         \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 ,
         \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 ,
         \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 ,
         \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 ,
         \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 ,
         \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 ,
         \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 ,
         \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 ,
         \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 ,
         \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 ,
         \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 ,
         \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 ,
         \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 ,
         \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 ,
         \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 ,
         \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 ,
         \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 ,
         \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 ,
         \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 ,
         \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 ,
         \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 ,
         \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 ,
         \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 ,
         \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 ,
         \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 ,
         \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 ,
         \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 ,
         \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 ,
         \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 ,
         \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 ,
         \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 ,
         \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 ,
         \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 ,
         \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 ,
         \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 ,
         \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 ,
         \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 ,
         \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 ,
         \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 ,
         \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 ,
         \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 ,
         \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 ,
         \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 ,
         \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 ,
         \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 ,
         \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 ,
         \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 ,
         \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 ,
         \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 ,
         \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 ,
         \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 ,
         \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 ,
         \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 ,
         \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 ,
         \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 ,
         \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 ,
         \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 ,
         \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 ,
         \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 ,
         \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 ,
         \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 ,
         \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 ,
         \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 ,
         \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 ,
         \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 ,
         \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 ,
         \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 ,
         \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 ,
         \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 ,
         \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 ,
         \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 ,
         \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 ,
         \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 ,
         \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 ,
         \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 ,
         \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 ,
         \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 ,
         \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 ,
         \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 ,
         \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 ,
         \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 ,
         \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 ,
         \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 ,
         \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 ,
         \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 ,
         \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 ,
         \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 ,
         \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 ,
         \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 ,
         \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 ,
         \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 ,
         \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 ,
         \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 ,
         \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 ,
         \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 ,
         \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 ,
         \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 ,
         \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 ,
         \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 ,
         \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 ,
         \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 ,
         \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 ,
         \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 ,
         \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 ,
         \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 ,
         \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 ,
         \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 ,
         \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 ,
         \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 ,
         \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 ,
         \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 ,
         \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 ,
         \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 ,
         \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 ,
         \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 ,
         \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 ,
         \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 ,
         \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 ,
         \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 ,
         \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 ,
         \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 ,
         \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 ,
         \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 ,
         \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 ,
         \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 ,
         \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 ,
         \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 ,
         \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 ,
         \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 ,
         \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 ,
         \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 ,
         \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 ,
         \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 ,
         \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 ,
         \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 ,
         \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 ,
         \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 ,
         \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 ,
         \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 ,
         \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 ,
         \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 ,
         \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 ,
         \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 ,
         \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 ,
         \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 ,
         \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 ,
         \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 ,
         \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 ,
         \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 ,
         \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 ,
         \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 ,
         \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 ,
         \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 ,
         \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 ,
         \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 ,
         \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 ,
         \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 ,
         \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 ,
         \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 ,
         \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 ,
         \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 ,
         \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 ,
         \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 ,
         \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 ,
         \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 ,
         \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 ,
         \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 ,
         \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 ,
         \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 ,
         \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 ,
         \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 ,
         \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 ,
         \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 ,
         \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 ,
         \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 ,
         \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 ,
         \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 ,
         \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 ,
         \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 ,
         \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 ,
         \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 ,
         \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 ,
         \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 ,
         \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 ,
         \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 ,
         \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 ,
         \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 ,
         \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 ,
         \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 ,
         \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 ,
         \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 ,
         \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 ,
         \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 ,
         \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 ,
         \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 ,
         \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 ,
         \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 ,
         \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 ,
         \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 ,
         \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 ,
         \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 ,
         \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 ,
         \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 ,
         \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 ,
         \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 ,
         \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 ,
         \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 ,
         \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 ,
         \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 ,
         \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 ,
         \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 ,
         \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 ,
         \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 ,
         \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 ,
         \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 ,
         \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 ,
         \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 ,
         \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 ,
         \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 ,
         \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 ,
         \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 ,
         \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 ,
         \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 ,
         \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 ,
         \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 ,
         \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 ,
         \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 ,
         \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 ,
         \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 ,
         \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 ,
         \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 ,
         \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 ,
         \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 ,
         \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 ,
         \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 ,
         \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 ,
         \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 ,
         \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 ,
         \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 ,
         \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 ,
         \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 ,
         \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 ,
         \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 ,
         \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 ,
         \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 ,
         \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 ,
         \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 ,
         \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 ,
         \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 ,
         \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 ,
         \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 ,
         \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 ,
         \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 ,
         \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 ,
         \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 ,
         \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 ,
         \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 ,
         \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 ,
         \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 ,
         \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 ,
         \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 ,
         \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 ,
         \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 ,
         \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 ,
         \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 ,
         \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 ,
         \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 ,
         \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 ,
         \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 ,
         \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 ,
         \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 ,
         \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 ,
         \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 ,
         \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 ,
         \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 ,
         \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 ,
         \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 ,
         \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 ,
         \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 ,
         \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 ,
         \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 ,
         \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 ,
         \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 ,
         \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 ,
         \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 ,
         \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 ,
         \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 ,
         \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 ,
         \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 ,
         \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 ,
         \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 ,
         \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 ,
         \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 ,
         \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 ,
         \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 ,
         \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 ,
         \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 ,
         \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 ,
         \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 ,
         \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 ,
         \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 ,
         \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 ,
         \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 ,
         \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 ,
         \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 ,
         \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 ,
         \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 ,
         \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 ,
         \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 ,
         \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 ,
         \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 ,
         \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 ,
         \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 ,
         \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 ,
         \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 ,
         \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 ,
         \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 ,
         \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 ,
         \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 ,
         \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 ,
         \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 ,
         \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 ,
         \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 ,
         \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 ,
         \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 ,
         \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 ,
         \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 ,
         \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 ,
         \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 ,
         \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 ,
         \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 ,
         \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 ,
         \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 ,
         \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 ,
         \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 ,
         \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 ,
         \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 ,
         \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 ,
         \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 ,
         \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 ,
         \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 ,
         \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 ,
         \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 ,
         \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 ,
         \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 ,
         \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 ,
         \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 ,
         \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 ,
         \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 ,
         \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 ,
         \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 ,
         \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 ,
         \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 ,
         \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 ,
         \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 ,
         \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 ,
         \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 ,
         \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 ,
         \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 ,
         \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 ,
         \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 ,
         \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 ,
         \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 ,
         \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 ,
         \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 ,
         \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 ,
         \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 ,
         \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 ,
         \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 ,
         \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 ,
         \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 ,
         \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 ,
         \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 ,
         \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 ,
         \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 ,
         \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 ,
         \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 ,
         \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 ,
         \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 ,
         \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 ,
         \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 ,
         \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 ,
         \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 ,
         \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 ,
         \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 ,
         \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 ,
         \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 ,
         \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 ,
         \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 ,
         \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 ,
         \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 ,
         \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 ,
         \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 ,
         \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 ,
         \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 ,
         \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 ,
         \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 ,
         \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 ,
         \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 ,
         \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 ,
         \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 ,
         \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 ,
         \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 ,
         \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 ,
         \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 ,
         \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 ,
         \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 ,
         \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 ,
         \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 ,
         \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 ,
         \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 ,
         \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 ,
         \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 ,
         \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 ,
         \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 ,
         \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 ,
         \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 ,
         \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 ,
         \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 ,
         \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 ,
         \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 ,
         \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 ,
         \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 ,
         \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 ,
         \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 ,
         \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 ,
         \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 ,
         \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 ,
         \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 ,
         \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 ,
         \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 ,
         \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 ,
         \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 ,
         \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 ,
         \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 ,
         \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 ,
         \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 ,
         \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 ,
         \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 ,
         \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 ,
         \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 ,
         \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 ,
         \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 ,
         \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 ,
         \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 ,
         \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 ,
         \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 ,
         \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 ,
         \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 ,
         \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 ,
         \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 ,
         \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 ,
         \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 ,
         \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 ,
         \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 ,
         \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 ,
         \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 ,
         \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 ,
         \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 ,
         \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 ,
         \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 ,
         \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 ,
         \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 ,
         \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 ,
         \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 ,
         \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 ,
         \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 ,
         \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 ,
         \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 ,
         \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 ,
         \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 ,
         \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 ,
         \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 ,
         \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 ,
         \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 ,
         \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 ,
         \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 ,
         \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 ,
         \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 ,
         \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 ,
         \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 ,
         \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 ,
         \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 ,
         \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 ,
         \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 ,
         \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 ,
         \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 ,
         \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 ,
         \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 ,
         \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 ,
         \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 ,
         \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 ,
         \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 ,
         \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 ,
         \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 ,
         \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 ,
         \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 ,
         \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 ,
         \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 ,
         \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 ,
         \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 ,
         \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 ,
         \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 ,
         \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 ,
         \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 ,
         \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 ,
         \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 ,
         \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 ,
         \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 ,
         \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 ,
         \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 ,
         \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 ,
         \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 ,
         \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 ,
         \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 ,
         \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 ,
         \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 ,
         \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 ,
         \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 ,
         \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 ,
         \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 ,
         \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 ,
         \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 ,
         \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 ,
         \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 ,
         \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 ,
         \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 ,
         \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 ,
         \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 ,
         \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 ,
         \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 ,
         \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 ,
         \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 ,
         \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 ,
         \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 ,
         \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 ,
         \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 ,
         \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 ,
         \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 ,
         \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 ,
         \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 ,
         \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 ,
         \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 ,
         \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 ,
         \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 ,
         \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 ,
         \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 ,
         \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 ,
         \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 ,
         \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 ,
         \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 ,
         \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 ,
         \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 ,
         \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 ,
         \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 ,
         \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 ,
         \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 ,
         \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 ,
         \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 ,
         \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 ,
         \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 ,
         \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 ,
         \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 ,
         \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 ,
         \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 ,
         \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 ,
         \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 ,
         \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 ,
         \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 ,
         \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 ,
         \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 ,
         \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 ,
         \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 ,
         \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 ,
         \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 ,
         \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 ,
         \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 ,
         \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 ,
         \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 ,
         \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 ,
         \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 ,
         \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 ,
         \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 ,
         \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 ,
         \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 ,
         \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 ,
         \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 ,
         \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 ,
         \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 ,
         \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 ,
         \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 ,
         \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 ,
         \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 ,
         \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 ,
         \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 ,
         \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 ,
         \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 ,
         \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 ,
         \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 ,
         \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 ,
         \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 ,
         \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 ,
         \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 ,
         \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 ,
         \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 ,
         \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 ,
         \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 ,
         \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 ,
         \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 ,
         \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 ,
         \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 ,
         \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 ,
         \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 ,
         \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 ,
         \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 ,
         \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 ,
         \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 ,
         \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 ,
         \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 ,
         \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 ,
         \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 ,
         \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 ,
         \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 ,
         \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 ,
         \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 ,
         \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 ,
         \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 ,
         \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 , \10948 , \10949 , \10950 ,
         \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 , \10958 , \10959 , \10960 ,
         \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 , \10968 , \10969 , \10970 ,
         \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 , \10978 , \10979 , \10980 ,
         \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 , \10988 , \10989 , \10990 ,
         \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 , \10998 , \10999 , \11000 ,
         \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 , \11008 , \11009 , \11010 ,
         \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 , \11018 , \11019 , \11020 ,
         \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 , \11028 , \11029 , \11030 ,
         \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 , \11038 , \11039 , \11040 ,
         \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 , \11048 , \11049 , \11050 ,
         \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 , \11058 , \11059 , \11060 ,
         \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 , \11068 , \11069 , \11070 ,
         \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 , \11078 , \11079 , \11080 ,
         \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 , \11088 , \11089 , \11090 ,
         \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 , \11098 , \11099 , \11100 ,
         \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 , \11108 , \11109 , \11110 ,
         \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 , \11118 , \11119 , \11120 ,
         \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 , \11128 , \11129 , \11130 ,
         \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 , \11138 , \11139 , \11140 ,
         \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 , \11148 , \11149 , \11150 ,
         \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 , \11158 , \11159 , \11160 ,
         \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 , \11168 , \11169 , \11170 ,
         \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 , \11178 , \11179 , \11180 ,
         \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 , \11188 , \11189 , \11190 ,
         \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 , \11198 , \11199 , \11200 ,
         \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 , \11208 , \11209 , \11210 ,
         \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 , \11218 , \11219 , \11220 ,
         \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 , \11228 , \11229 , \11230 ,
         \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 , \11238 , \11239 , \11240 ,
         \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 , \11248 , \11249 , \11250 ,
         \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 , \11258 , \11259 , \11260 ,
         \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 , \11268 , \11269 , \11270 ,
         \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 , \11278 , \11279 , \11280 ,
         \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 , \11288 , \11289 , \11290 ,
         \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 , \11298 , \11299 , \11300 ,
         \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 , \11308 , \11309 , \11310 ,
         \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 , \11318 , \11319 , \11320 ,
         \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 , \11328 , \11329 , \11330 ,
         \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 , \11338 , \11339 , \11340 ,
         \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 , \11348 , \11349 , \11350 ,
         \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 , \11358 , \11359 , \11360 ,
         \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 , \11368 , \11369 , \11370 ,
         \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 , \11378 , \11379 , \11380 ,
         \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 , \11388 , \11389 , \11390 ,
         \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 , \11398 , \11399 , \11400 ,
         \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 , \11408 , \11409 , \11410 ,
         \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 , \11418 , \11419 , \11420 ,
         \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 , \11428 , \11429 , \11430 ,
         \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 , \11438 , \11439 , \11440 ,
         \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 , \11448 , \11449 , \11450 ,
         \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 , \11458 , \11459 , \11460 ,
         \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 , \11468 , \11469 , \11470 ,
         \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 , \11478 , \11479 , \11480 ,
         \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 , \11488 , \11489 , \11490 ,
         \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 , \11498 , \11499 , \11500 ,
         \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 , \11508 , \11509 , \11510 ,
         \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 , \11518 , \11519 , \11520 ,
         \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 , \11528 , \11529 , \11530 ,
         \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 , \11538 , \11539 , \11540 ,
         \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 , \11548 , \11549 , \11550 ,
         \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 , \11558 , \11559 , \11560 ,
         \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 , \11568 , \11569 , \11570 ,
         \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 , \11578 , \11579 , \11580 ,
         \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 , \11588 , \11589 , \11590 ,
         \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 , \11598 , \11599 , \11600 ,
         \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 , \11608 , \11609 , \11610 ,
         \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 , \11618 , \11619 , \11620 ,
         \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 , \11628 , \11629 , \11630 ,
         \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 , \11638 , \11639 , \11640 ,
         \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 , \11648 , \11649 , \11650 ,
         \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 , \11658 , \11659 , \11660 ,
         \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 , \11668 , \11669 , \11670 ,
         \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 , \11678 , \11679 , \11680 ,
         \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 , \11688 , \11689 , \11690 ,
         \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 , \11698 , \11699 , \11700 ,
         \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 , \11708 , \11709 , \11710 ,
         \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 , \11718 , \11719 , \11720 ,
         \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 , \11728 , \11729 , \11730 ,
         \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 , \11738 , \11739 , \11740 ,
         \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 , \11748 , \11749 , \11750 ,
         \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 , \11758 , \11759 , \11760 ,
         \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 , \11768 , \11769 , \11770 ,
         \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 , \11778 , \11779 , \11780 ,
         \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 , \11788 , \11789 , \11790 ,
         \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 , \11798 , \11799 , \11800 ,
         \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 , \11808 , \11809 , \11810 ,
         \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 , \11818 , \11819 , \11820 ,
         \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 , \11828 , \11829 , \11830 ,
         \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 , \11838 , \11839 , \11840 ,
         \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 , \11848 , \11849 , \11850 ,
         \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 , \11858 , \11859 , \11860 ,
         \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 , \11868 , \11869 , \11870 ,
         \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 , \11878 , \11879 , \11880 ,
         \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 , \11888 , \11889 , \11890 ,
         \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 , \11898 , \11899 , \11900 ,
         \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 , \11908 , \11909 , \11910 ,
         \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 , \11918 , \11919 , \11920 ,
         \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 , \11928 , \11929 , \11930 ,
         \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 , \11938 , \11939 , \11940 ,
         \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 , \11948 , \11949 , \11950 ,
         \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 , \11958 , \11959 , \11960 ,
         \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 , \11968 , \11969 , \11970 ,
         \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 , \11978 , \11979 , \11980 ,
         \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 , \11988 , \11989 , \11990 ,
         \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 , \11998 , \11999 , \12000 ,
         \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 , \12008 , \12009 , \12010 ,
         \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 , \12018 , \12019 , \12020 ,
         \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 , \12028 , \12029 , \12030 ,
         \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 , \12038 , \12039 , \12040 ,
         \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 , \12048 , \12049 , \12050 ,
         \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 , \12058 , \12059 , \12060 ,
         \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 , \12068 , \12069 , \12070 ,
         \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 , \12078 , \12079 , \12080 ,
         \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 , \12088 , \12089 , \12090 ,
         \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 , \12098 , \12099 , \12100 ,
         \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 , \12108 , \12109 , \12110 ,
         \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 , \12118 , \12119 , \12120 ,
         \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 , \12128 , \12129 , \12130 ,
         \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 , \12138 , \12139 , \12140 ,
         \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 , \12148 , \12149 , \12150 ,
         \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 , \12158 , \12159 , \12160 ,
         \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 , \12168 , \12169 , \12170 ,
         \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 , \12178 , \12179 , \12180 ,
         \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 , \12188 , \12189 , \12190 ,
         \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 , \12198 , \12199 , \12200 ,
         \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 , \12208 , \12209 , \12210 ,
         \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 , \12218 , \12219 , \12220 ,
         \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 , \12228 , \12229 , \12230 ,
         \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 , \12238 , \12239 , \12240 ,
         \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 , \12248 , \12249 , \12250 ,
         \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 , \12258 , \12259 , \12260 ,
         \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 , \12268 , \12269 , \12270 ,
         \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 , \12278 , \12279 , \12280 ,
         \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 , \12288 , \12289 , \12290 ,
         \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 , \12298 , \12299 , \12300 ,
         \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 , \12308 , \12309 , \12310 ,
         \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 , \12318 , \12319 , \12320 ,
         \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 , \12328 , \12329 , \12330 ,
         \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 , \12338 , \12339 , \12340 ,
         \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 , \12348 , \12349 , \12350 ,
         \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 , \12358 , \12359 , \12360 ,
         \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 , \12368 , \12369 , \12370 ,
         \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 , \12378 , \12379 , \12380 ,
         \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 , \12388 , \12389 , \12390 ,
         \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 , \12398 , \12399 , \12400 ,
         \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 , \12408 , \12409 , \12410 ,
         \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 , \12418 , \12419 , \12420 ,
         \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 , \12428 , \12429 , \12430 ,
         \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 , \12438 , \12439 , \12440 ,
         \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 , \12448 , \12449 , \12450 ,
         \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 , \12458 , \12459 , \12460 ,
         \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 , \12468 , \12469 , \12470 ,
         \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 , \12478 , \12479 , \12480 ,
         \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 , \12488 , \12489 , \12490 ,
         \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 , \12498 , \12499 , \12500 ,
         \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 , \12508 , \12509 , \12510 ,
         \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 , \12518 , \12519 , \12520 ,
         \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 , \12528 , \12529 , \12530 ,
         \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 , \12538 , \12539 , \12540 ,
         \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 , \12548 , \12549 , \12550 ,
         \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 , \12558 , \12559 , \12560 ,
         \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 , \12568 , \12569 , \12570 ,
         \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 , \12578 , \12579 , \12580 ,
         \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 , \12588 , \12589 , \12590 ,
         \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 , \12598 , \12599 , \12600 ,
         \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 , \12608 , \12609 , \12610 ,
         \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 , \12618 , \12619 , \12620 ,
         \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 , \12628 , \12629 , \12630 ,
         \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 , \12638 , \12639 , \12640 ,
         \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 , \12648 , \12649 , \12650 ,
         \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 , \12658 , \12659 , \12660 ,
         \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 , \12668 , \12669 , \12670 ,
         \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 , \12678 , \12679 , \12680 ,
         \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 , \12688 , \12689 , \12690 ,
         \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 , \12698 , \12699 , \12700 ,
         \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 , \12708 , \12709 , \12710 ,
         \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 , \12718 , \12719 , \12720 ,
         \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 , \12728 , \12729 , \12730 ,
         \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 , \12738 , \12739 , \12740 ,
         \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 , \12748 , \12749 , \12750 ,
         \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 , \12758 , \12759 , \12760 ,
         \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 , \12768 , \12769 , \12770 ,
         \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 , \12778 , \12779 , \12780 ,
         \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 , \12788 , \12789 , \12790 ,
         \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 , \12798 , \12799 , \12800 ,
         \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 , \12808 , \12809 , \12810 ,
         \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 , \12818 , \12819 , \12820 ,
         \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 , \12828 , \12829 , \12830 ,
         \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 , \12838 , \12839 , \12840 ,
         \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 , \12848 , \12849 , \12850 ,
         \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 , \12858 , \12859 , \12860 ,
         \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 , \12868 , \12869 , \12870 ,
         \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 , \12878 , \12879 , \12880 ,
         \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 , \12888 , \12889 , \12890 ,
         \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 , \12898 , \12899 , \12900 ,
         \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 , \12908 , \12909 , \12910 ,
         \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 , \12918 , \12919 , \12920 ,
         \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 , \12928 , \12929 , \12930 ,
         \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 , \12938 , \12939 , \12940 ,
         \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 , \12948 , \12949 , \12950 ,
         \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 , \12958 , \12959 , \12960 ,
         \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 , \12968 , \12969 , \12970 ,
         \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 , \12978 , \12979 , \12980 ,
         \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 , \12988 , \12989 , \12990 ,
         \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 , \12998 , \12999 , \13000 ,
         \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 , \13008 , \13009 , \13010 ,
         \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 , \13018 , \13019 , \13020 ,
         \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 , \13028 , \13029 , \13030 ,
         \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 , \13038 , \13039 , \13040 ,
         \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 , \13048 , \13049 , \13050 ,
         \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 , \13058 , \13059 , \13060 ,
         \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 , \13068 , \13069 , \13070 ,
         \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 , \13078 , \13079 , \13080 ,
         \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 , \13088 , \13089 , \13090 ,
         \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 , \13098 , \13099 , \13100 ,
         \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 , \13108 , \13109 , \13110 ,
         \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 , \13118 , \13119 , \13120 ,
         \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 , \13128 , \13129 , \13130 ,
         \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 , \13138 , \13139 , \13140 ,
         \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 , \13148 , \13149 , \13150 ,
         \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 , \13158 , \13159 , \13160 ,
         \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 , \13168 , \13169 , \13170 ,
         \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 , \13178 , \13179 , \13180 ,
         \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 , \13188 , \13189 , \13190 ,
         \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 , \13198 , \13199 , \13200 ,
         \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 , \13208 , \13209 , \13210 ,
         \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 , \13218 , \13219 , \13220 ,
         \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 , \13228 , \13229 , \13230 ,
         \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 , \13238 , \13239 , \13240 ,
         \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 , \13248 , \13249 , \13250 ,
         \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 , \13258 , \13259 , \13260 ,
         \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 , \13268 , \13269 , \13270 ,
         \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 , \13278 , \13279 , \13280 ,
         \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 , \13288 , \13289 , \13290 ,
         \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 , \13298 , \13299 , \13300 ,
         \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 , \13308 , \13309 , \13310 ,
         \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 , \13318 , \13319 , \13320 ,
         \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 , \13328 , \13329 , \13330 ,
         \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 , \13338 , \13339 , \13340 ,
         \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 , \13348 , \13349 , \13350 ,
         \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 , \13358 , \13359 , \13360 ,
         \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 , \13368 , \13369 , \13370 ,
         \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 , \13378 , \13379 , \13380 ,
         \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 , \13388 , \13389 , \13390 ,
         \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 , \13398 , \13399 , \13400 ,
         \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 , \13408 , \13409 , \13410 ,
         \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 , \13418 , \13419 , \13420 ,
         \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 , \13428 , \13429 , \13430 ,
         \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 , \13438 , \13439 , \13440 ,
         \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 , \13448 , \13449 , \13450 ,
         \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 , \13458 , \13459 , \13460 ,
         \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 , \13468 , \13469 , \13470 ,
         \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 , \13478 , \13479 , \13480 ,
         \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 , \13488 , \13489 , \13490 ,
         \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 , \13498 , \13499 , \13500 ,
         \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 , \13508 , \13509 , \13510 ,
         \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 , \13518 , \13519 , \13520 ,
         \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 , \13528 , \13529 , \13530 ,
         \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 , \13538 , \13539 , \13540 ,
         \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 , \13548 , \13549 , \13550 ,
         \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 , \13558 , \13559 , \13560 ,
         \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 , \13568 , \13569 , \13570 ,
         \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 , \13578 , \13579 , \13580 ,
         \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 , \13588 , \13589 , \13590 ,
         \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 , \13598 , \13599 , \13600 ,
         \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 , \13608 , \13609 , \13610 ,
         \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 , \13618 , \13619 , \13620 ,
         \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 , \13628 , \13629 , \13630 ,
         \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 , \13638 , \13639 , \13640 ,
         \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 , \13648 , \13649 , \13650 ,
         \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 , \13658 , \13659 , \13660 ,
         \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 , \13668 , \13669 , \13670 ,
         \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 , \13678 , \13679 , \13680 ,
         \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 , \13688 , \13689 , \13690 ,
         \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 , \13698 , \13699 , \13700 ,
         \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 , \13708 , \13709 , \13710 ,
         \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 , \13718 , \13719 , \13720 ,
         \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 , \13728 , \13729 , \13730 ,
         \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 , \13738 , \13739 , \13740 ,
         \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 , \13748 , \13749 , \13750 ,
         \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 , \13758 , \13759 , \13760 ,
         \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 , \13768 , \13769 , \13770 ,
         \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 , \13778 , \13779 , \13780 ,
         \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 , \13788 , \13789 , \13790 ,
         \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 , \13798 , \13799 , \13800 ,
         \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 , \13808 , \13809 , \13810 ,
         \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 , \13818 , \13819 , \13820 ,
         \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 , \13828 , \13829 , \13830 ,
         \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 , \13838 , \13839 , \13840 ,
         \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 , \13848 , \13849 , \13850 ,
         \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 , \13858 , \13859 , \13860 ,
         \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 , \13868 , \13869 , \13870 ,
         \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 , \13878 , \13879 , \13880 ,
         \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 , \13888 , \13889 , \13890 ,
         \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 , \13898 , \13899 , \13900 ,
         \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 , \13908 , \13909 , \13910 ,
         \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 , \13918 , \13919 , \13920 ,
         \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 , \13928 , \13929 , \13930 ,
         \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 , \13938 , \13939 , \13940 ,
         \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 , \13948 , \13949 , \13950 ,
         \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 , \13958 , \13959 , \13960 ,
         \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 , \13968 , \13969 , \13970 ,
         \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 , \13978 , \13979 , \13980 ,
         \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 , \13988 , \13989 , \13990 ,
         \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 , \13998 , \13999 , \14000 ,
         \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 , \14008 , \14009 , \14010 ,
         \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 , \14018 , \14019 , \14020 ,
         \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 , \14028 , \14029 , \14030 ,
         \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 , \14038 , \14039 , \14040 ,
         \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 , \14048 , \14049 , \14050 ,
         \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 , \14058 , \14059 , \14060 ,
         \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 , \14068 , \14069 , \14070 ,
         \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 , \14078 , \14079 , \14080 ,
         \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 , \14088 , \14089 , \14090 ,
         \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 , \14098 , \14099 , \14100 ,
         \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 , \14108 , \14109 , \14110 ,
         \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 , \14118 , \14119 , \14120 ,
         \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 , \14128 , \14129 , \14130 ,
         \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 , \14138 , \14139 , \14140 ,
         \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 , \14148 , \14149 , \14150 ,
         \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 , \14158 , \14159 , \14160 ,
         \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 , \14168 , \14169 , \14170 ,
         \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 , \14178 , \14179 , \14180 ,
         \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 , \14188 , \14189 , \14190 ,
         \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 , \14198 , \14199 , \14200 ,
         \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 , \14208 , \14209 , \14210 ,
         \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 , \14218 , \14219 , \14220 ,
         \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 , \14228 , \14229 , \14230 ,
         \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 , \14238 , \14239 , \14240 ,
         \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 , \14248 , \14249 , \14250 ,
         \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 , \14258 , \14259 , \14260 ,
         \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 , \14268 , \14269 , \14270 ,
         \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 , \14278 , \14279 , \14280 ,
         \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 , \14288 , \14289 , \14290 ,
         \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 , \14298 , \14299 , \14300 ,
         \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 , \14308 , \14309 , \14310 ,
         \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 , \14318 , \14319 , \14320 ,
         \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 , \14328 , \14329 , \14330 ,
         \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 , \14338 , \14339 , \14340 ,
         \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 , \14348 , \14349 , \14350 ,
         \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 , \14358 , \14359 , \14360 ,
         \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 , \14368 , \14369 , \14370 ,
         \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 , \14378 , \14379 , \14380 ,
         \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 , \14388 , \14389 , \14390 ,
         \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 , \14398 , \14399 , \14400 ,
         \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 , \14408 , \14409 , \14410 ,
         \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 , \14418 , \14419 , \14420 ,
         \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 , \14428 , \14429 , \14430 ,
         \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 , \14438 , \14439 , \14440 ,
         \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 , \14448 , \14449 , \14450 ,
         \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 , \14458 , \14459 , \14460 ,
         \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 , \14468 , \14469 , \14470 ,
         \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 , \14478 , \14479 , \14480 ,
         \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 , \14488 , \14489 , \14490 ,
         \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 , \14498 , \14499 , \14500 ,
         \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 , \14508 , \14509 , \14510 ,
         \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 , \14518 , \14519 , \14520 ,
         \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 , \14528 , \14529 , \14530 ,
         \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 , \14538 , \14539 , \14540 ,
         \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 , \14548 , \14549 , \14550 ,
         \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 , \14558 , \14559 , \14560 ,
         \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 , \14568 , \14569 , \14570 ,
         \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 , \14578 , \14579 , \14580 ,
         \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 , \14588 , \14589 , \14590 ,
         \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 , \14598 , \14599 , \14600 ,
         \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 , \14608 , \14609 , \14610 ,
         \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 , \14618 , \14619 , \14620 ,
         \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 , \14628 , \14629 , \14630 ,
         \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 , \14638 , \14639 , \14640 ,
         \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 , \14648 , \14649 , \14650 ,
         \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 , \14658 , \14659 , \14660 ,
         \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 , \14668 , \14669 , \14670 ,
         \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 , \14678 , \14679 , \14680 ,
         \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 , \14688 , \14689 , \14690 ,
         \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 , \14698 , \14699 , \14700 ,
         \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 , \14708 , \14709 , \14710 ,
         \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 , \14718 , \14719 , \14720 ,
         \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 , \14728 , \14729 , \14730 ,
         \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 , \14738 , \14739 , \14740 ,
         \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 , \14748 , \14749 , \14750 ,
         \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 , \14758 , \14759 , \14760 ,
         \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 , \14768 , \14769 , \14770 ,
         \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 , \14778 , \14779 , \14780 ,
         \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 , \14788 , \14789 , \14790 ,
         \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 , \14798 , \14799 , \14800 ,
         \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 , \14808 , \14809 , \14810 ,
         \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 , \14818 , \14819 , \14820 ,
         \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 , \14828 , \14829 , \14830 ,
         \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 , \14838 , \14839 , \14840 ,
         \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 , \14848 , \14849 , \14850 ,
         \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 , \14858 , \14859 , \14860 ,
         \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 , \14868 , \14869 , \14870 ,
         \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 , \14878 , \14879 , \14880 ,
         \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 , \14888 , \14889 , \14890 ,
         \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 , \14898 , \14899 , \14900 ,
         \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 , \14908 , \14909 , \14910 ,
         \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 , \14918 , \14919 , \14920 ,
         \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 , \14928 , \14929 , \14930 ,
         \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 , \14938 , \14939 , \14940 ,
         \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 , \14948 , \14949 , \14950 ,
         \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 , \14958 , \14959 , \14960 ,
         \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 , \14968 , \14969 , \14970 ,
         \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 , \14978 , \14979 , \14980 ,
         \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 , \14988 , \14989 , \14990 ,
         \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 , \14998 , \14999 , \15000 ,
         \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 , \15008 , \15009 , \15010 ,
         \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 , \15018 , \15019 , \15020 ,
         \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 , \15028 , \15029 , \15030 ,
         \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 , \15038 , \15039 , \15040 ,
         \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 , \15048 , \15049 , \15050 ,
         \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 , \15058 , \15059 , \15060 ,
         \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 , \15068 , \15069 , \15070 ,
         \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 , \15078 , \15079 , \15080 ,
         \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 , \15088 , \15089 , \15090 ,
         \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 , \15098 , \15099 , \15100 ,
         \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 , \15108 , \15109 , \15110 ,
         \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 , \15118 , \15119 , \15120 ,
         \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 , \15128 , \15129 , \15130 ,
         \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 , \15138 , \15139 , \15140 ,
         \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 , \15148 , \15149 , \15150 ,
         \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 , \15158 , \15159 , \15160 ,
         \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 , \15168 , \15169 , \15170 ,
         \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 , \15178 , \15179 , \15180 ,
         \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 , \15188 , \15189 , \15190 ,
         \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 , \15198 , \15199 , \15200 ,
         \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 , \15208 , \15209 , \15210 ,
         \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 , \15218 , \15219 , \15220 ,
         \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 , \15228 , \15229 , \15230 ,
         \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 , \15238 , \15239 , \15240 ,
         \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 , \15248 , \15249 , \15250 ,
         \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 , \15258 , \15259 , \15260 ,
         \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 , \15268 , \15269 , \15270 ,
         \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 , \15278 , \15279 , \15280 ,
         \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 , \15288 , \15289 , \15290 ,
         \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 , \15298 , \15299 , \15300 ,
         \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 , \15308 , \15309 , \15310 ,
         \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 , \15318 , \15319 , \15320 ,
         \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 , \15328 , \15329 , \15330 ,
         \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 , \15338 , \15339 , \15340 ,
         \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 , \15348 , \15349 , \15350 ,
         \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 , \15358 , \15359 , \15360 ,
         \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 , \15368 , \15369 , \15370 ,
         \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 , \15378 , \15379 , \15380 ,
         \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 , \15388 , \15389 , \15390 ,
         \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 , \15398 , \15399 , \15400 ,
         \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 , \15408 , \15409 , \15410 ,
         \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 , \15418 , \15419 , \15420 ,
         \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 , \15428 , \15429 , \15430 ,
         \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 , \15438 , \15439 , \15440 ,
         \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 , \15448 , \15449 , \15450 ,
         \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 , \15458 , \15459 , \15460 ,
         \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 , \15468 , \15469 , \15470 ,
         \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 , \15478 , \15479 , \15480 ,
         \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 , \15488 , \15489 , \15490 ,
         \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 , \15498 , \15499 , \15500 ,
         \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 , \15508 , \15509 , \15510 ,
         \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 , \15518 , \15519 , \15520 ,
         \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 , \15528 , \15529 , \15530 ,
         \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 , \15538 , \15539 , \15540 ,
         \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 , \15548 , \15549 , \15550 ,
         \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 , \15558 , \15559 , \15560 ,
         \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 , \15568 , \15569 , \15570 ,
         \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 , \15578 , \15579 , \15580 ,
         \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 , \15588 , \15589 , \15590 ,
         \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 , \15598 , \15599 , \15600 ,
         \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 , \15608 , \15609 , \15610 ,
         \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 , \15618 , \15619 , \15620 ,
         \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 , \15628 , \15629 , \15630 ,
         \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 , \15638 , \15639 , \15640 ,
         \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 , \15648 , \15649 , \15650 ,
         \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 , \15658 , \15659 , \15660 ,
         \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 , \15668 , \15669 , \15670 ,
         \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 , \15678 , \15679 , \15680 ,
         \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 , \15688 , \15689 , \15690 ,
         \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 , \15698 , \15699 , \15700 ,
         \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 , \15708 , \15709 , \15710 ,
         \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 , \15718 , \15719 , \15720 ,
         \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 , \15728 , \15729 , \15730 ,
         \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 , \15738 , \15739 , \15740 ,
         \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 , \15748 , \15749 , \15750 ,
         \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 , \15758 , \15759 , \15760 ,
         \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 , \15768 , \15769 , \15770 ,
         \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 , \15778 , \15779 , \15780 ,
         \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 , \15788 , \15789 , \15790 ,
         \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 , \15798 , \15799 , \15800 ,
         \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 , \15808 , \15809 , \15810 ,
         \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 , \15818 , \15819 , \15820 ,
         \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 , \15828 , \15829 , \15830 ,
         \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 , \15838 , \15839 , \15840 ,
         \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 , \15848 , \15849 , \15850 ,
         \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 , \15858 , \15859 , \15860 ,
         \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 , \15868 , \15869 , \15870 ,
         \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 , \15878 , \15879 , \15880 ,
         \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 , \15888 , \15889 , \15890 ,
         \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 , \15898 , \15899 , \15900 ,
         \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 , \15908 , \15909 , \15910 ,
         \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 , \15918 , \15919 , \15920 ,
         \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 , \15928 , \15929 , \15930 ,
         \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 , \15938 , \15939 , \15940 ,
         \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 , \15948 , \15949 , \15950 ,
         \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 , \15958 , \15959 , \15960 ,
         \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 , \15968 , \15969 , \15970 ,
         \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 , \15978 , \15979 , \15980 ,
         \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 , \15988 , \15989 , \15990 ,
         \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 , \15998 , \15999 , \16000 ,
         \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 , \16008 , \16009 , \16010 ,
         \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 , \16018 , \16019 , \16020 ,
         \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 , \16028 , \16029 , \16030 ,
         \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 , \16038 , \16039 , \16040 ,
         \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 , \16048 , \16049 , \16050 ,
         \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 , \16058 , \16059 , \16060 ,
         \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 , \16068 , \16069 , \16070 ,
         \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 , \16078 , \16079 , \16080 ,
         \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 , \16088 , \16089 , \16090 ,
         \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 , \16098 , \16099 , \16100 ,
         \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 , \16108 , \16109 , \16110 ,
         \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 , \16118 , \16119 , \16120 ,
         \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 , \16128 , \16129 , \16130 ,
         \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 , \16138 , \16139 , \16140 ,
         \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 , \16148 , \16149 , \16150 ,
         \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 , \16158 , \16159 , \16160 ,
         \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 , \16168 , \16169 , \16170 ,
         \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 , \16178 , \16179 , \16180 ,
         \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 , \16188 , \16189 , \16190 ,
         \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 , \16198 , \16199 , \16200 ,
         \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 , \16208 , \16209 , \16210 ,
         \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 , \16218 , \16219 , \16220 ,
         \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 , \16228 , \16229 , \16230 ,
         \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 , \16238 , \16239 , \16240 ,
         \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 , \16248 , \16249 , \16250 ,
         \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 , \16258 , \16259 , \16260 ,
         \16261 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 , \16268 , \16269 , \16270 ,
         \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 , \16278 , \16279 , \16280 ,
         \16281 , \16282 , \16283 , \16284 , \16285 , \16286 , \16287 , \16288 , \16289 , \16290 ,
         \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 , \16298 , \16299 , \16300 ,
         \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 , \16308 , \16309 , \16310 ,
         \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 , \16318 , \16319 , \16320 ,
         \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 , \16328 , \16329 , \16330 ,
         \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 , \16338 , \16339 , \16340 ,
         \16341 , \16342 , \16343 , \16344 , \16345 , \16346 , \16347 , \16348 , \16349 , \16350 ,
         \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 , \16358 , \16359 , \16360 ,
         \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 , \16368 , \16369 , \16370 ,
         \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 , \16378 , \16379 , \16380 ,
         \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 , \16388 , \16389 , \16390 ,
         \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 , \16398 , \16399 , \16400 ,
         \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 , \16408 , \16409 , \16410 ,
         \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 , \16418 , \16419 , \16420 ,
         \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 , \16428 , \16429 , \16430 ,
         \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 , \16438 , \16439 , \16440 ,
         \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 , \16448 , \16449 , \16450 ,
         \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 , \16458 , \16459 , \16460 ,
         \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 , \16468 , \16469 , \16470 ,
         \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 , \16478 , \16479 , \16480 ,
         \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 , \16488 , \16489 , \16490 ,
         \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 , \16498 , \16499 , \16500 ,
         \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 , \16508 , \16509 , \16510 ,
         \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 , \16518 , \16519 , \16520 ,
         \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 , \16528 , \16529 , \16530 ,
         \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 , \16538 , \16539 , \16540 ,
         \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 , \16548 , \16549 , \16550 ,
         \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 , \16558 , \16559 , \16560 ,
         \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 , \16568 , \16569 , \16570 ,
         \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 , \16578 , \16579 , \16580 ,
         \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 , \16588 , \16589 , \16590 ,
         \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 , \16598 , \16599 , \16600 ,
         \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 , \16608 , \16609 , \16610 ,
         \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 , \16618 , \16619 , \16620 ,
         \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 , \16628 , \16629 , \16630 ,
         \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 , \16638 , \16639 , \16640 ,
         \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 , \16648 , \16649 , \16650 ,
         \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 , \16658 , \16659 , \16660 ,
         \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 , \16668 , \16669 , \16670 ,
         \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 , \16678 , \16679 , \16680 ,
         \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 , \16688 , \16689 , \16690 ,
         \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 , \16698 , \16699 , \16700 ,
         \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 , \16708 , \16709 , \16710 ,
         \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 , \16718 , \16719 , \16720 ,
         \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 , \16728 , \16729 , \16730 ,
         \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 , \16738 , \16739 , \16740 ,
         \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 , \16748 , \16749 , \16750 ,
         \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 , \16758 , \16759 , \16760 ,
         \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 , \16768 , \16769 , \16770 ,
         \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 , \16778 , \16779 , \16780 ,
         \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 , \16788 , \16789 , \16790 ,
         \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 , \16798 , \16799 , \16800 ,
         \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 , \16808 , \16809 , \16810 ,
         \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 , \16818 , \16819 , \16820 ,
         \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 , \16828 , \16829 , \16830 ,
         \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 , \16838 , \16839 , \16840 ,
         \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 , \16848 , \16849 , \16850 ,
         \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 , \16858 , \16859 , \16860 ,
         \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 , \16868 , \16869 , \16870 ,
         \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 , \16878 , \16879 , \16880 ,
         \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 , \16888 , \16889 , \16890 ,
         \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 , \16898 , \16899 , \16900 ,
         \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 , \16908 , \16909 , \16910 ,
         \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 , \16918 , \16919 , \16920 ,
         \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 , \16928 , \16929 , \16930 ,
         \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 , \16938 , \16939 , \16940 ,
         \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 , \16948 , \16949 , \16950 ,
         \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 , \16958 , \16959 , \16960 ,
         \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 , \16968 , \16969 , \16970 ,
         \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 , \16978 , \16979 , \16980 ,
         \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 , \16988 , \16989 , \16990 ,
         \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 , \16998 , \16999 , \17000 ,
         \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 , \17008 , \17009 , \17010 ,
         \17011 , \17012 , \17013 , \17014 , \17015 , \17016 , \17017 , \17018 , \17019 , \17020 ,
         \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 , \17028 , \17029 , \17030 ,
         \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 , \17038 , \17039 , \17040 ,
         \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 , \17048 , \17049 , \17050 ,
         \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 , \17058 , \17059 , \17060 ,
         \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 , \17068 , \17069 , \17070 ,
         \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 , \17078 , \17079 , \17080 ,
         \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 , \17088 , \17089 , \17090 ,
         \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 , \17098 , \17099 , \17100 ,
         \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 , \17108 , \17109 , \17110 ,
         \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 , \17118 , \17119 , \17120 ,
         \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 , \17128 , \17129 , \17130 ,
         \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 , \17138 , \17139 , \17140 ,
         \17141 , \17142 , \17143 , \17144 , \17145 , \17146 , \17147 , \17148 , \17149 , \17150 ,
         \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 , \17158 , \17159 , \17160 ,
         \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 , \17168 , \17169 , \17170 ,
         \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 , \17178 , \17179 , \17180 ,
         \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 , \17188 , \17189 , \17190 ,
         \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 , \17198 , \17199 , \17200 ,
         \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 , \17208 , \17209 , \17210 ,
         \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 , \17218 , \17219 , \17220 ,
         \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 , \17228 , \17229 , \17230 ,
         \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 , \17238 , \17239 , \17240 ,
         \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 , \17248 , \17249 , \17250 ,
         \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 , \17258 , \17259 , \17260 ,
         \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 , \17268 , \17269 , \17270 ,
         \17271 , \17272 , \17273 , \17274 , \17275 , \17276 , \17277 , \17278 , \17279 , \17280 ,
         \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 , \17288 , \17289 , \17290 ,
         \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 , \17298 , \17299 , \17300 ,
         \17301 , \17302 , \17303 , \17304 , \17305 , \17306 , \17307 , \17308 , \17309 , \17310 ,
         \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 , \17318 , \17319 , \17320 ,
         \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 , \17328 , \17329 , \17330 ,
         \17331 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 , \17338 , \17339 , \17340 ,
         \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 , \17348 , \17349 , \17350 ,
         \17351 , \17352 , \17353 , \17354 , \17355 , \17356 , \17357 , \17358 , \17359 , \17360 ,
         \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 , \17368 , \17369 , \17370 ,
         \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 , \17378 , \17379 , \17380 ,
         \17381 , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 , \17388 , \17389 , \17390 ,
         \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 , \17398 , \17399 , \17400 ,
         \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 , \17408 , \17409 , \17410 ,
         \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 , \17418 , \17419 , \17420 ,
         \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 , \17428 , \17429 , \17430 ,
         \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 , \17438 , \17439 , \17440 ,
         \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 , \17448 , \17449 , \17450 ,
         \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 , \17458 , \17459 , \17460 ,
         \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 , \17468 , \17469 , \17470 ,
         \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 , \17478 , \17479 , \17480 ,
         \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 , \17488 , \17489 , \17490 ,
         \17491 , \17492 , \17493 , \17494 , \17495 , \17496 , \17497 , \17498 , \17499 , \17500 ,
         \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 , \17508 , \17509 , \17510 ,
         \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 , \17518 , \17519 , \17520 ,
         \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 , \17528 , \17529 , \17530 ,
         \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 , \17538 , \17539 , \17540 ,
         \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 , \17548 , \17549 , \17550 ,
         \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 , \17558 , \17559 , \17560 ,
         \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 , \17568 , \17569 , \17570 ,
         \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 , \17578 , \17579 , \17580 ,
         \17581 , \17582 , \17583 , \17584 , \17585 , \17586 , \17587 , \17588 , \17589 , \17590 ,
         \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 , \17598 , \17599 , \17600 ,
         \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 , \17608 , \17609 , \17610 ,
         \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 , \17618 , \17619 , \17620 ,
         \17621 , \17622 , \17623 , \17624 , \17625 , \17626 , \17627 , \17628 , \17629 , \17630 ,
         \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 , \17638 , \17639 , \17640 ,
         \17641 , \17642 , \17643 , \17644 , \17645 , \17646 , \17647 , \17648 , \17649 , \17650 ,
         \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 , \17658 , \17659 , \17660 ,
         \17661 , \17662 , \17663 , \17664 , \17665 , \17666 , \17667 , \17668 , \17669 , \17670 ,
         \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 , \17678 , \17679 , \17680 ,
         \17681 , \17682 , \17683 , \17684 , \17685 , \17686 , \17687 , \17688 , \17689 , \17690 ,
         \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 , \17698 , \17699 , \17700 ,
         \17701 , \17702 , \17703 , \17704 , \17705 , \17706 , \17707 , \17708 , \17709 , \17710 ,
         \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 , \17718 , \17719 , \17720 ,
         \17721 , \17722 , \17723 , \17724 , \17725 , \17726 , \17727 , \17728 , \17729 , \17730 ,
         \17731 , \17732 , \17733 , \17734 , \17735 , \17736 , \17737 , \17738 , \17739 , \17740 ,
         \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 , \17748 , \17749 , \17750 ,
         \17751 , \17752 , \17753 , \17754 , \17755 , \17756 , \17757 , \17758 , \17759 , \17760 ,
         \17761 , \17762 , \17763 , \17764 , \17765 , \17766 , \17767 , \17768 , \17769 , \17770 ,
         \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 , \17778 , \17779 , \17780 ,
         \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 , \17788 , \17789 , \17790 ,
         \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 , \17798 , \17799 , \17800 ,
         \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 , \17808 , \17809 , \17810 ,
         \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 , \17818 , \17819 , \17820 ,
         \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 , \17828 , \17829 , \17830 ,
         \17831 , \17832 , \17833 , \17834 , \17835 , \17836 , \17837 , \17838 , \17839 , \17840 ,
         \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 , \17848 , \17849 , \17850 ,
         \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 , \17858 , \17859 , \17860 ,
         \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 , \17868 , \17869 , \17870 ,
         \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 , \17878 , \17879 , \17880 ,
         \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 , \17888 , \17889 , \17890 ,
         \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 , \17898 , \17899 , \17900 ,
         \17901 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 , \17908 , \17909 , \17910 ,
         \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 , \17918 , \17919 , \17920 ,
         \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 , \17928 , \17929 , \17930 ,
         \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 , \17938 , \17939 , \17940 ,
         \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 , \17948 , \17949 , \17950 ,
         \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 , \17958 , \17959 , \17960 ,
         \17961 , \17962 , \17963 , \17964 , \17965 , \17966 , \17967 , \17968 , \17969 , \17970 ,
         \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 , \17978 , \17979 , \17980 ,
         \17981 , \17982 , \17983 , \17984 , \17985 , \17986 , \17987 , \17988 , \17989 , \17990 ,
         \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 , \17998 , \17999 , \18000 ,
         \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 , \18008 , \18009 , \18010 ,
         \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 , \18018 , \18019 , \18020 ,
         \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 , \18028 , \18029 , \18030 ,
         \18031 , \18032 , \18033 , \18034 , \18035 , \18036 , \18037 , \18038 , \18039 , \18040 ,
         \18041 , \18042 , \18043 , \18044 , \18045 , \18046 , \18047 , \18048 , \18049 , \18050 ,
         \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 , \18058 , \18059 , \18060 ,
         \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 , \18068 , \18069 , \18070 ,
         \18071 , \18072 , \18073 , \18074 , \18075 , \18076 , \18077 , \18078 , \18079 , \18080 ,
         \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 , \18088 , \18089 , \18090 ,
         \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 , \18098 , \18099 , \18100 ,
         \18101 , \18102 , \18103 , \18104 , \18105 , \18106 , \18107 , \18108 , \18109 , \18110 ,
         \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 , \18118 , \18119 , \18120 ,
         \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 , \18128 , \18129 , \18130 ,
         \18131 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 , \18138 , \18139 , \18140 ,
         \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 , \18148 , \18149 , \18150 ,
         \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 , \18158 , \18159 , \18160 ,
         \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 , \18168 , \18169 , \18170 ,
         \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 , \18178 , \18179 , \18180 ,
         \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 , \18188 , \18189 , \18190 ,
         \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 , \18198 , \18199 , \18200 ,
         \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 , \18208 , \18209 , \18210 ,
         \18211 , \18212 , \18213 , \18214 , \18215 , \18216 , \18217 , \18218 , \18219 , \18220 ,
         \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 , \18228 , \18229 , \18230 ,
         \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 , \18238 , \18239 , \18240 ,
         \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 , \18248 , \18249 , \18250 ,
         \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 , \18258 , \18259 , \18260 ,
         \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 , \18268 , \18269 , \18270 ,
         \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 , \18278 , \18279 , \18280 ,
         \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 , \18288 , \18289 , \18290 ,
         \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 , \18298 , \18299 , \18300 ,
         \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 , \18308 , \18309 , \18310 ,
         \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 , \18318 , \18319 , \18320 ,
         \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 , \18328 , \18329 , \18330 ,
         \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 , \18338 , \18339 , \18340 ,
         \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 , \18348 , \18349 , \18350 ,
         \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 , \18358 , \18359 , \18360 ,
         \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 , \18368 , \18369 , \18370 ,
         \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 , \18378 , \18379 , \18380 ,
         \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 , \18388 , \18389 , \18390 ,
         \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 , \18398 , \18399 , \18400 ,
         \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 , \18408 , \18409 , \18410 ,
         \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 , \18418 , \18419 , \18420 ,
         \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 , \18428 , \18429 , \18430 ,
         \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 , \18438 , \18439 , \18440 ,
         \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 , \18448 , \18449 , \18450 ,
         \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 , \18458 , \18459 , \18460 ,
         \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 , \18468 , \18469 , \18470 ,
         \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 , \18478 , \18479 , \18480 ,
         \18481 , \18482 , \18483 , \18484 , \18485 , \18486 , \18487 , \18488 , \18489 , \18490 ,
         \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 , \18498 , \18499 , \18500 ,
         \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 , \18508 , \18509 , \18510 ,
         \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 , \18518 , \18519 , \18520 ,
         \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 , \18528 , \18529 , \18530 ,
         \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 , \18538 , \18539 , \18540 ,
         \18541 , \18542 , \18543 , \18544 , \18545 , \18546 , \18547 , \18548 , \18549 , \18550 ,
         \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 , \18558 , \18559 , \18560 ,
         \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 , \18568 , \18569 , \18570 ,
         \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 , \18578 , \18579 , \18580 ,
         \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 , \18588 , \18589 , \18590 ,
         \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 , \18598 , \18599 , \18600 ,
         \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 , \18608 , \18609 , \18610 ,
         \18611 , \18612 , \18613 , \18614 , \18615 , \18616 , \18617 , \18618 , \18619 , \18620 ,
         \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 , \18628 , \18629 , \18630 ,
         \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 , \18638 , \18639 , \18640 ,
         \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 , \18648 , \18649 , \18650 ,
         \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 , \18658 , \18659 , \18660 ,
         \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 , \18668 , \18669 , \18670 ,
         \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 , \18678 , \18679 , \18680 ,
         \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 , \18688 , \18689 , \18690 ,
         \18691 , \18692 , \18693 , \18694 , \18695 , \18696 , \18697 , \18698 , \18699 , \18700 ,
         \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 , \18708 , \18709 , \18710 ,
         \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717 , \18718 , \18719 , \18720 ,
         \18721 , \18722 , \18723 , \18724 , \18725 , \18726 , \18727 , \18728 , \18729 , \18730 ,
         \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 , \18738 , \18739 , \18740 ,
         \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 , \18748 , \18749 , \18750 ,
         \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 , \18758 , \18759 , \18760 ,
         \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 , \18768 , \18769 , \18770 ,
         \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 , \18778 , \18779 , \18780 ,
         \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 , \18788 , \18789 , \18790 ,
         \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 , \18798 , \18799 , \18800 ,
         \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 , \18808 , \18809 , \18810 ,
         \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 , \18818 , \18819 , \18820 ,
         \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 , \18828 , \18829 , \18830 ,
         \18831 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 , \18838 , \18839 , \18840 ,
         \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 , \18848 , \18849 , \18850 ,
         \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 , \18858 , \18859 , \18860 ,
         \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 , \18868 , \18869 , \18870 ,
         \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 , \18878 , \18879 , \18880 ,
         \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887 , \18888 , \18889 , \18890 ,
         \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 , \18898 , \18899 , \18900 ,
         \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 , \18908 , \18909 , \18910 ,
         \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 , \18918 , \18919 , \18920 ,
         \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 , \18928 , \18929 , \18930 ,
         \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 , \18938 , \18939 , \18940 ,
         \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 , \18948 , \18949 , \18950 ,
         \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 , \18958 , \18959 , \18960 ,
         \18961 , \18962 , \18963 , \18964 , \18965 , \18966 , \18967 , \18968 , \18969 , \18970 ,
         \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 , \18978 , \18979 , \18980 ,
         \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 , \18988 , \18989 , \18990 ,
         \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 , \18998 , \18999 , \19000 ,
         \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 , \19008 , \19009 , \19010 ,
         \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 , \19018 , \19019 , \19020 ,
         \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 , \19028 , \19029 , \19030 ,
         \19031 , \19032 , \19033 , \19034 , \19035 , \19036 , \19037 , \19038 , \19039 , \19040 ,
         \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 , \19048 , \19049 , \19050 ,
         \19051 , \19052 , \19053 , \19054 , \19055 , \19056 , \19057 , \19058 , \19059 , \19060 ,
         \19061 , \19062 , \19063 , \19064 , \19065 , \19066 , \19067 , \19068 , \19069 , \19070 ,
         \19071 , \19072 , \19073 , \19074 , \19075 , \19076 , \19077 , \19078 , \19079 , \19080 ,
         \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 , \19088 , \19089 , \19090 ,
         \19091 , \19092 , \19093 , \19094 , \19095 , \19096 , \19097 , \19098 , \19099 , \19100 ,
         \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 , \19108 , \19109 , \19110 ,
         \19111 , \19112 , \19113 , \19114 , \19115 , \19116 , \19117 , \19118 , \19119 , \19120 ,
         \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 , \19128 , \19129 , \19130 ,
         \19131 , \19132 , \19133 , \19134 , \19135 , \19136 , \19137 , \19138 , \19139 , \19140 ,
         \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 , \19148 , \19149 , \19150 ,
         \19151 , \19152 , \19153 , \19154 , \19155 , \19156 , \19157 , \19158 , \19159 , \19160 ,
         \19161 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 , \19168 , \19169 , \19170 ,
         \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 , \19178 , \19179 , \19180 ,
         \19181 , \19182 , \19183 , \19184 , \19185 , \19186 , \19187 , \19188 , \19189 , \19190 ,
         \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 , \19198 , \19199 , \19200 ,
         \19201 , \19202 , \19203 , \19204 , \19205 , \19206 , \19207 , \19208 , \19209 , \19210 ,
         \19211 , \19212 , \19213 , \19214 , \19215 , \19216 , \19217 , \19218 , \19219 , \19220 ,
         \19221 , \19222 , \19223 , \19224 , \19225 , \19226 , \19227 , \19228 , \19229 , \19230 ,
         \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 , \19238 , \19239 , \19240 ,
         \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 , \19248 , \19249 , \19250 ,
         \19251 , \19252 , \19253 , \19254 , \19255 , \19256 , \19257 , \19258 , \19259 , \19260 ,
         \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 , \19268 , \19269 , \19270 ,
         \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 , \19278 , \19279 , \19280 ,
         \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 , \19288 , \19289 , \19290 ,
         \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 , \19298 , \19299 , \19300 ,
         \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 , \19308 , \19309 , \19310 ,
         \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 , \19318 , \19319 , \19320 ,
         \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 , \19328 , \19329 , \19330 ,
         \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 , \19338 , \19339 , \19340 ,
         \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 , \19348 , \19349 , \19350 ,
         \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 , \19358 , \19359 , \19360 ,
         \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 , \19368 , \19369 , \19370 ,
         \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 , \19378 , \19379 , \19380 ,
         \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 , \19388 , \19389 , \19390 ,
         \19391 , \19392 , \19393 , \19394 , \19395 , \19396 , \19397 , \19398 , \19399 , \19400 ,
         \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 , \19408 , \19409 , \19410 ,
         \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 , \19418 , \19419 , \19420 ,
         \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 , \19428 , \19429 , \19430 ,
         \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 , \19438 , \19439 , \19440 ,
         \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 , \19448 , \19449 , \19450 ,
         \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 , \19458 , \19459 , \19460 ,
         \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 , \19468 , \19469 , \19470 ,
         \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 , \19478 , \19479 , \19480 ,
         \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 , \19488 , \19489 , \19490 ,
         \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 , \19498 , \19499 , \19500 ,
         \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 , \19508 , \19509 , \19510 ,
         \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 , \19518 , \19519 , \19520 ,
         \19521 , \19522 , \19523 , \19524 , \19525 , \19526 , \19527 , \19528 , \19529 , \19530 ,
         \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 , \19538 , \19539 , \19540 ,
         \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 , \19548 , \19549 , \19550 ,
         \19551 , \19552 , \19553 , \19554 , \19555 , \19556 , \19557 , \19558 , \19559 , \19560 ,
         \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 , \19568 , \19569 , \19570 ,
         \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 , \19578 , \19579 , \19580 ,
         \19581 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 , \19588 , \19589 , \19590 ,
         \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 , \19598 , \19599 , \19600 ,
         \19601 , \19602 , \19603 , \19604 , \19605 , \19606 , \19607 , \19608 , \19609 , \19610 ,
         \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 , \19618 , \19619 , \19620 ,
         \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 , \19628 , \19629 , \19630 ,
         \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 , \19638 , \19639 , \19640 ,
         \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 , \19648 , \19649 , \19650 ,
         \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 , \19658 , \19659 , \19660 ,
         \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 , \19668 , \19669 , \19670 ,
         \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 , \19678 , \19679 , \19680 ,
         \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 , \19688 , \19689 , \19690 ,
         \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 , \19698 , \19699 , \19700 ,
         \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 , \19708 , \19709 , \19710 ,
         \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 , \19718 , \19719 , \19720 ,
         \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 , \19728 , \19729 , \19730 ,
         \19731 , \19732 , \19733 , \19734 , \19735 , \19736 , \19737 , \19738 , \19739 , \19740 ,
         \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 , \19748 , \19749 , \19750 ,
         \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 , \19758 , \19759 , \19760 ,
         \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 , \19768 , \19769 , \19770 ,
         \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 , \19778 , \19779 , \19780 ,
         \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 , \19788 , \19789 , \19790 ,
         \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 , \19798 , \19799 , \19800 ,
         \19801 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 , \19808 , \19809 , \19810 ,
         \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 , \19818 , \19819 , \19820 ,
         \19821 , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 , \19828 , \19829 , \19830 ,
         \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 , \19838 , \19839 , \19840 ,
         \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 , \19848 , \19849 , \19850 ,
         \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 , \19858 , \19859 , \19860 ,
         \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 , \19868 , \19869 , \19870 ,
         \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 , \19878 , \19879 , \19880 ,
         \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 , \19888 , \19889 , \19890 ,
         \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 , \19898 , \19899 , \19900 ,
         \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 , \19908 , \19909 , \19910 ,
         \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 , \19918 , \19919 , \19920 ,
         \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 , \19928 , \19929 , \19930 ,
         \19931 , \19932 , \19933 , \19934 , \19935 , \19936 , \19937 , \19938 , \19939 , \19940 ,
         \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 , \19948 , \19949 , \19950 ,
         \19951 , \19952 , \19953 , \19954 , \19955 , \19956 , \19957 , \19958 , \19959 , \19960 ,
         \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 , \19968 , \19969 , \19970 ,
         \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 , \19978 , \19979 , \19980 ,
         \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 , \19988 , \19989 , \19990 ,
         \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 , \19998 , \19999 , \20000 ,
         \20001 , \20002 , \20003 , \20004 , \20005 , \20006 , \20007 , \20008 , \20009 , \20010 ,
         \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 , \20018 , \20019 , \20020 ,
         \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 , \20028 , \20029 , \20030 ,
         \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 , \20038 , \20039 , \20040 ,
         \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 , \20048 , \20049 , \20050 ,
         \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 , \20058 , \20059 , \20060 ,
         \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 , \20068 , \20069 , \20070 ,
         \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 , \20078 , \20079 , \20080 ,
         \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 , \20088 , \20089 , \20090 ,
         \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 , \20098 , \20099 , \20100 ,
         \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 , \20108 , \20109 , \20110 ,
         \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 , \20118 , \20119 , \20120 ,
         \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 , \20128 , \20129 , \20130 ,
         \20131 , \20132 , \20133 , \20134 , \20135 , \20136 , \20137 , \20138 , \20139 , \20140 ,
         \20141 , \20142 , \20143 , \20144 , \20145 , \20146 , \20147 , \20148 , \20149 , \20150 ,
         \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , \20157 , \20158 , \20159 , \20160 ,
         \20161 , \20162 , \20163 , \20164 , \20165 , \20166 , \20167 , \20168 , \20169 , \20170 ,
         \20171 , \20172 , \20173 , \20174 , \20175 , \20176 , \20177 , \20178 , \20179 , \20180 ,
         \20181 , \20182 , \20183 , \20184 , \20185 , \20186 , \20187 , \20188 , \20189 , \20190 ,
         \20191 , \20192 , \20193 , \20194 , \20195 , \20196 , \20197 , \20198 , \20199 , \20200 ,
         \20201 , \20202 , \20203 , \20204 , \20205 , \20206 , \20207 , \20208 , \20209 , \20210 ,
         \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 , \20218 , \20219 , \20220 ,
         \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 , \20228 , \20229 , \20230 ,
         \20231 , \20232 , \20233 , \20234 , \20235 , \20236 , \20237 , \20238 , \20239 , \20240 ,
         \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 , \20248 , \20249 , \20250 ,
         \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 , \20258 , \20259 , \20260 ,
         \20261 , \20262 , \20263 , \20264 , \20265 , \20266 , \20267 , \20268 , \20269 , \20270 ,
         \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 , \20278 , \20279 , \20280 ,
         \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 , \20288 , \20289 , \20290 ,
         \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 , \20298 , \20299 , \20300 ,
         \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 , \20308 , \20309 , \20310 ,
         \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 , \20318 , \20319 , \20320 ,
         \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 , \20328 , \20329 , \20330 ,
         \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 , \20338 , \20339 , \20340 ,
         \20341 , \20342 , \20343 , \20344 , \20345 , \20346 , \20347 , \20348 , \20349 , \20350 ,
         \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 , \20358 , \20359 , \20360 ,
         \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 , \20368 , \20369 , \20370 ,
         \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 , \20378 , \20379 , \20380 ,
         \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 , \20388 , \20389 , \20390 ,
         \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 , \20398 , \20399 , \20400 ,
         \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 , \20408 , \20409 , \20410 ,
         \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 , \20418 , \20419 , \20420 ,
         \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 , \20428 , \20429 , \20430 ,
         \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 , \20438 , \20439 , \20440 ,
         \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 , \20448 , \20449 , \20450 ,
         \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457 , \20458 , \20459 , \20460 ,
         \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 , \20468 , \20469 , \20470 ,
         \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 , \20478 , \20479 , \20480 ,
         \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 , \20488 , \20489 , \20490 ,
         \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 , \20498 , \20499 , \20500 ,
         \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 , \20508 , \20509 , \20510 ,
         \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 , \20518 , \20519 , \20520 ,
         \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 , \20528 , \20529 , \20530 ,
         \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 , \20538 , \20539 , \20540 ,
         \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 , \20548 , \20549 , \20550 ,
         \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 , \20558 , \20559 , \20560 ,
         \20561 , \20562 , \20563 , \20564 , \20565 , \20566 , \20567 , \20568 , \20569 , \20570 ,
         \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 , \20578 , \20579 , \20580 ,
         \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 , \20588 , \20589 , \20590 ,
         \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 , \20598 , \20599 , \20600 ,
         \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 , \20608 , \20609 , \20610 ,
         \20611 , \20612 , \20613 , \20614 , \20615 , \20616 , \20617 , \20618 , \20619 , \20620 ,
         \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 , \20628 , \20629 , \20630 ,
         \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 , \20638 , \20639 , \20640 ,
         \20641 , \20642 , \20643 , \20644 , \20645 , \20646 , \20647 , \20648 , \20649 , \20650 ,
         \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 , \20658 , \20659 , \20660 ,
         \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 , \20668 , \20669 , \20670 ,
         \20671 , \20672 , \20673 , \20674 , \20675 , \20676 , \20677 , \20678 , \20679 , \20680 ,
         \20681 , \20682 , \20683 , \20684 , \20685 , \20686 , \20687 , \20688 , \20689 , \20690 ,
         \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 , \20698 , \20699 , \20700 ,
         \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 , \20708 , \20709 , \20710 ,
         \20711 , \20712 , \20713 , \20714 , \20715 , \20716 , \20717 , \20718 , \20719 , \20720 ,
         \20721 , \20722 , \20723 , \20724 , \20725 , \20726 , \20727 , \20728 , \20729 , \20730 ,
         \20731 , \20732 , \20733 , \20734 , \20735 , \20736 , \20737 , \20738 , \20739 , \20740 ,
         \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 , \20748 , \20749 , \20750 ,
         \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 , \20758 , \20759 , \20760 ,
         \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 , \20768 , \20769 , \20770 ,
         \20771 , \20772 , \20773 , \20774 , \20775 , \20776 , \20777 , \20778 , \20779 , \20780 ,
         \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 , \20788 , \20789 , \20790 ,
         \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 , \20798 , \20799 , \20800 ,
         \20801 , \20802 , \20803 , \20804 , \20805 , \20806 , \20807 , \20808 , \20809 , \20810 ,
         \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 , \20818 , \20819 , \20820 ,
         \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 , \20828 , \20829 , \20830 ,
         \20831 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 , \20838 , \20839 , \20840 ,
         \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 , \20848 , \20849 , \20850 ,
         \20851 , \20852 , \20853 , \20854 , \20855 , \20856 , \20857 , \20858 , \20859 , \20860 ,
         \20861 , \20862 , \20863 , \20864 , \20865 , \20866 , \20867 , \20868 , \20869 , \20870 ,
         \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 , \20878 , \20879 , \20880 ,
         \20881 , \20882 , \20883 , \20884 , \20885 , \20886 , \20887 , \20888 , \20889 , \20890 ,
         \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 , \20898 , \20899 , \20900 ,
         \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 , \20908 , \20909 , \20910 ,
         \20911 , \20912 , \20913 , \20914 , \20915 , \20916 , \20917 , \20918 , \20919 , \20920 ,
         \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 , \20928 , \20929 , \20930 ,
         \20931 , \20932 , \20933 , \20934 , \20935 , \20936 , \20937 , \20938 , \20939 , \20940 ,
         \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 , \20948 , \20949 , \20950 ,
         \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 , \20958 , \20959 , \20960 ,
         \20961 , \20962 , \20963 , \20964 , \20965 , \20966 , \20967 , \20968 , \20969 , \20970 ,
         \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 , \20978 , \20979 , \20980 ,
         \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 , \20988 , \20989 , \20990 ,
         \20991 , \20992 , \20993 , \20994 , \20995 , \20996 , \20997 , \20998 , \20999 , \21000 ,
         \21001 , \21002 , \21003 , \21004 , \21005 , \21006 , \21007 , \21008 , \21009 , \21010 ,
         \21011 , \21012 , \21013 , \21014 , \21015 , \21016 , \21017 , \21018 , \21019 , \21020 ,
         \21021 , \21022 , \21023 , \21024 , \21025 , \21026 , \21027 , \21028 , \21029 , \21030 ,
         \21031 , \21032 , \21033 , \21034 , \21035 , \21036 , \21037 , \21038 , \21039 , \21040 ,
         \21041 , \21042 , \21043 , \21044 , \21045 , \21046 , \21047 , \21048 , \21049 , \21050 ,
         \21051 , \21052 , \21053 , \21054 , \21055 , \21056 , \21057 , \21058 , \21059 , \21060 ,
         \21061 , \21062 , \21063 , \21064 , \21065 , \21066 , \21067 , \21068 , \21069 , \21070 ,
         \21071 , \21072 , \21073 , \21074 , \21075 , \21076 , \21077 , \21078 , \21079 , \21080 ,
         \21081 , \21082 , \21083 , \21084 , \21085 , \21086 , \21087 , \21088 , \21089 , \21090 ,
         \21091 , \21092 , \21093 , \21094 , \21095 , \21096 , \21097 , \21098 , \21099 , \21100 ,
         \21101 , \21102 , \21103 , \21104 , \21105 , \21106 , \21107 , \21108 , \21109 , \21110 ,
         \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 , \21118 , \21119 , \21120 ,
         \21121 , \21122 , \21123 , \21124 , \21125 , \21126 , \21127 , \21128 , \21129 , \21130 ,
         \21131 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 , \21138 , \21139 , \21140 ,
         \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 , \21148 , \21149 , \21150 ,
         \21151 , \21152 , \21153 , \21154 , \21155 , \21156 , \21157 , \21158 , \21159 , \21160 ,
         \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 , \21168 , \21169 , \21170 ,
         \21171 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 , \21178 , \21179 , \21180 ,
         \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 , \21188 , \21189 , \21190 ,
         \21191 , \21192 , \21193 , \21194 , \21195 , \21196 , \21197 , \21198 , \21199 , \21200 ,
         \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207 , \21208 , \21209 , \21210 ,
         \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 , \21218 , \21219 , \21220 ,
         \21221 , \21222 , \21223 , \21224 , \21225 , \21226 , \21227 , \21228 , \21229 , \21230 ,
         \21231 , \21232 , \21233 , \21234 , \21235 , \21236 , \21237 , \21238 , \21239 , \21240 ,
         \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 , \21248 , \21249 , \21250 ,
         \21251 , \21252 , \21253 , \21254 , \21255 , \21256 , \21257 , \21258 , \21259 , \21260 ,
         \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 , \21268 , \21269 , \21270 ,
         \21271 , \21272 , \21273 , \21274 , \21275 , \21276 , \21277 , \21278 , \21279 , \21280 ,
         \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 , \21288 , \21289 , \21290 ,
         \21291 , \21292 , \21293 , \21294 , \21295 , \21296 , \21297 , \21298 , \21299 , \21300 ,
         \21301 , \21302 , \21303 , \21304 , \21305 , \21306 , \21307 , \21308 , \21309 , \21310 ,
         \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 , \21318 , \21319 , \21320 ,
         \21321 , \21322 , \21323 , \21324 , \21325 , \21326 , \21327 , \21328 , \21329 , \21330 ,
         \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 , \21338 , \21339 , \21340 ,
         \21341 , \21342 , \21343 , \21344 , \21345 , \21346 , \21347 , \21348 , \21349 , \21350 ,
         \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 , \21358 , \21359 , \21360 ,
         \21361 , \21362 , \21363 , \21364 , \21365 , \21366 , \21367 , \21368 , \21369 , \21370 ,
         \21371 , \21372 , \21373 , \21374 , \21375 , \21376 , \21377 , \21378 , \21379 , \21380 ,
         \21381 , \21382 , \21383 , \21384 , \21385 , \21386 , \21387 , \21388 , \21389 , \21390 ,
         \21391 , \21392 , \21393 , \21394 , \21395 , \21396 , \21397 , \21398 , \21399 , \21400 ,
         \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 , \21408 , \21409 , \21410 ,
         \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 , \21418 , \21419 , \21420 ,
         \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 , \21428 , \21429 , \21430 ,
         \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 , \21438 , \21439 , \21440 ,
         \21441 , \21442 , \21443 , \21444 , \21445 , \21446 , \21447 , \21448 , \21449 , \21450 ,
         \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 , \21458 , \21459 , \21460 ,
         \21461 , \21462 , \21463 , \21464 , \21465 , \21466 , \21467 , \21468 , \21469 , \21470 ,
         \21471 , \21472 , \21473 , \21474 , \21475 , \21476 , \21477 , \21478 , \21479 , \21480 ,
         \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 , \21488 , \21489 , \21490 ,
         \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 , \21498 , \21499 , \21500 ,
         \21501 , \21502 , \21503 , \21504 , \21505 , \21506 , \21507 , \21508 , \21509 , \21510 ,
         \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517 , \21518 , \21519 , \21520 ,
         \21521 , \21522 , \21523 , \21524 , \21525 , \21526 , \21527 , \21528 , \21529 , \21530 ,
         \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 , \21538 , \21539 , \21540 ,
         \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 , \21548 , \21549 , \21550 ,
         \21551 , \21552 , \21553 , \21554 , \21555 , \21556 , \21557 , \21558 , \21559 , \21560 ,
         \21561 , \21562 , \21563 , \21564 , \21565 , \21566 , \21567 , \21568 , \21569 , \21570 ,
         \21571 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 , \21578 , \21579 , \21580 ,
         \21581 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 , \21588 , \21589 , \21590 ,
         \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 , \21598 , \21599 , \21600 ,
         \21601 , \21602 , \21603 , \21604 , \21605 , \21606 , \21607 , \21608 , \21609 , \21610 ,
         \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 , \21618 , \21619 , \21620 ,
         \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 , \21628 , \21629 , \21630 ,
         \21631 , \21632 , \21633 , \21634 , \21635 , \21636 , \21637 , \21638 , \21639 , \21640 ,
         \21641 , \21642 , \21643 , \21644 , \21645 , \21646 , \21647 , \21648 , \21649 , \21650 ,
         \21651 , \21652 , \21653 , \21654 , \21655 , \21656 , \21657 , \21658 , \21659 , \21660 ,
         \21661 , \21662 , \21663 , \21664 , \21665 , \21666 , \21667 , \21668 , \21669 , \21670 ,
         \21671 , \21672 , \21673 , \21674 , \21675 , \21676 , \21677 , \21678 , \21679 , \21680 ,
         \21681 , \21682 , \21683 , \21684 , \21685 , \21686 , \21687 , \21688 , \21689 , \21690 ,
         \21691 , \21692 , \21693 , \21694 , \21695 , \21696 , \21697 , \21698 , \21699 , \21700 ,
         \21701 , \21702 , \21703 , \21704 , \21705 , \21706 , \21707 , \21708 , \21709 , \21710 ,
         \21711 , \21712 , \21713 , \21714 , \21715 , \21716 , \21717 , \21718 , \21719 , \21720 ,
         \21721 , \21722 , \21723 , \21724 , \21725 , \21726 , \21727 , \21728 , \21729 , \21730 ,
         \21731 , \21732 , \21733 , \21734 , \21735 , \21736 , \21737 , \21738 , \21739 , \21740 ,
         \21741 , \21742 , \21743 , \21744 , \21745 , \21746 , \21747 , \21748 , \21749 , \21750 ,
         \21751 , \21752 , \21753 , \21754 , \21755 , \21756 , \21757 , \21758 , \21759 , \21760 ,
         \21761 , \21762 , \21763 , \21764 , \21765 , \21766 , \21767 , \21768 , \21769 , \21770 ,
         \21771 , \21772 , \21773 , \21774 , \21775 , \21776 , \21777 , \21778 , \21779 , \21780 ,
         \21781 , \21782 , \21783 , \21784 , \21785 , \21786 , \21787 , \21788 , \21789 , \21790 ,
         \21791 , \21792 , \21793 , \21794 , \21795 , \21796 , \21797 , \21798 , \21799 , \21800 ,
         \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 , \21808 , \21809 , \21810 ,
         \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 , \21818 , \21819 , \21820 ,
         \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 , \21828 , \21829 , \21830 ,
         \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 , \21838 , \21839 , \21840 ,
         \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 , \21848 , \21849 , \21850 ,
         \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 , \21858 , \21859 , \21860 ,
         \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 , \21868 , \21869 , \21870 ,
         \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 , \21878 , \21879 , \21880 ,
         \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 , \21888 , \21889 , \21890 ,
         \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 , \21898 , \21899 , \21900 ,
         \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 , \21908 , \21909 , \21910 ,
         \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 , \21918 , \21919 , \21920 ,
         \21921 , \21922 , \21923 , \21924 , \21925 , \21926 , \21927 , \21928 , \21929 , \21930 ,
         \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937 , \21938 , \21939 , \21940 ,
         \21941 , \21942 , \21943 , \21944 , \21945 , \21946 , \21947 , \21948 , \21949 , \21950 ,
         \21951 , \21952 , \21953 , \21954 , \21955 , \21956 , \21957 , \21958 , \21959 , \21960 ,
         \21961 , \21962 , \21963 , \21964 , \21965 , \21966 , \21967 , \21968 , \21969 , \21970 ,
         \21971 , \21972 , \21973 , \21974 , \21975 , \21976 , \21977 , \21978 , \21979 , \21980 ,
         \21981 , \21982 , \21983 , \21984 , \21985 , \21986 , \21987 , \21988 , \21989 , \21990 ,
         \21991 , \21992 , \21993 , \21994 , \21995 , \21996 , \21997 , \21998 , \21999 , \22000 ,
         \22001 , \22002 , \22003 , \22004 , \22005 , \22006 , \22007 , \22008 , \22009 , \22010 ,
         \22011 , \22012 , \22013 , \22014 , \22015 , \22016 , \22017 , \22018 , \22019 , \22020 ,
         \22021 , \22022 , \22023 , \22024 , \22025 , \22026 , \22027 , \22028 , \22029 , \22030 ,
         \22031 , \22032 , \22033 , \22034 , \22035 , \22036 , \22037 , \22038 , \22039 , \22040 ,
         \22041 , \22042 , \22043 , \22044 , \22045 , \22046 , \22047 , \22048 , \22049 , \22050 ,
         \22051 , \22052 , \22053 , \22054 , \22055 , \22056 , \22057 , \22058 , \22059 , \22060 ,
         \22061 , \22062 , \22063 , \22064 , \22065 , \22066 , \22067 , \22068 , \22069 , \22070 ,
         \22071 , \22072 , \22073 , \22074 , \22075 , \22076 , \22077 , \22078 , \22079 , \22080 ,
         \22081 , \22082 , \22083 , \22084 , \22085 , \22086 , \22087 , \22088 , \22089 , \22090 ,
         \22091 , \22092 , \22093 , \22094 , \22095 , \22096 , \22097 , \22098 , \22099 , \22100 ,
         \22101 , \22102 , \22103 , \22104 , \22105 , \22106 , \22107 , \22108 , \22109 , \22110 ,
         \22111 , \22112 , \22113 , \22114 , \22115 , \22116 , \22117 , \22118 , \22119 , \22120 ,
         \22121 , \22122 , \22123 , \22124 , \22125 , \22126 , \22127 , \22128 , \22129 , \22130 ,
         \22131 , \22132 , \22133 , \22134 , \22135 , \22136 , \22137 , \22138 , \22139 , \22140 ,
         \22141 , \22142 , \22143 , \22144 , \22145 , \22146 , \22147 , \22148 , \22149 , \22150 ,
         \22151 , \22152 , \22153 , \22154 , \22155 , \22156 , \22157 , \22158 , \22159 , \22160 ,
         \22161 , \22162 , \22163 , \22164 , \22165 , \22166 , \22167 , \22168 , \22169 , \22170 ,
         \22171 , \22172 , \22173 , \22174 , \22175 , \22176 , \22177 , \22178 , \22179 , \22180 ,
         \22181 , \22182 , \22183 , \22184 , \22185 , \22186 , \22187 , \22188 , \22189 , \22190 ,
         \22191 , \22192 , \22193 , \22194 , \22195 , \22196 , \22197 , \22198 , \22199 , \22200 ,
         \22201 , \22202 , \22203 , \22204 , \22205 , \22206 , \22207 , \22208 , \22209 , \22210 ,
         \22211 , \22212 , \22213 , \22214 , \22215 , \22216 , \22217 , \22218 , \22219 , \22220 ,
         \22221 , \22222 , \22223 , \22224 , \22225 , \22226 , \22227 , \22228 , \22229 , \22230 ,
         \22231 , \22232 , \22233 , \22234 , \22235 , \22236 , \22237 , \22238 , \22239 , \22240 ,
         \22241 , \22242 , \22243 , \22244 , \22245 , \22246 , \22247 , \22248 , \22249 , \22250 ,
         \22251 , \22252 , \22253 , \22254 , \22255 , \22256 , \22257 , \22258 , \22259 , \22260 ,
         \22261 , \22262 , \22263 , \22264 , \22265 , \22266 , \22267 , \22268 , \22269 , \22270 ,
         \22271 , \22272 , \22273 , \22274 , \22275 , \22276 , \22277 , \22278 , \22279 , \22280 ,
         \22281 , \22282 , \22283 , \22284 , \22285 , \22286 , \22287 , \22288 , \22289 , \22290 ,
         \22291 , \22292 , \22293 , \22294 , \22295 , \22296 , \22297 , \22298 , \22299 , \22300 ,
         \22301 , \22302 , \22303 , \22304 , \22305 , \22306 , \22307 , \22308 , \22309 , \22310 ,
         \22311 , \22312 , \22313 , \22314 , \22315 , \22316 , \22317 , \22318 , \22319 , \22320 ,
         \22321 , \22322 , \22323 , \22324 , \22325 , \22326 , \22327 , \22328 , \22329 , \22330 ,
         \22331 , \22332 , \22333 , \22334 , \22335 , \22336 , \22337 , \22338 , \22339 , \22340 ,
         \22341 , \22342 , \22343 , \22344 , \22345 , \22346 , \22347 , \22348 , \22349 , \22350 ,
         \22351 , \22352 , \22353 , \22354 , \22355 , \22356 , \22357 , \22358 , \22359 , \22360 ,
         \22361 , \22362 , \22363 , \22364 , \22365 , \22366 , \22367 , \22368 , \22369 , \22370 ,
         \22371 , \22372 , \22373 , \22374 , \22375 , \22376 , \22377 , \22378 , \22379 , \22380 ,
         \22381 , \22382 , \22383 , \22384 , \22385 , \22386 , \22387 , \22388 , \22389 , \22390 ,
         \22391 , \22392 , \22393 , \22394 , \22395 , \22396 , \22397 , \22398 , \22399 , \22400 ,
         \22401 , \22402 , \22403 , \22404 , \22405 , \22406 , \22407 , \22408 , \22409 , \22410 ,
         \22411 , \22412 , \22413 , \22414 , \22415 , \22416 , \22417 , \22418 , \22419 , \22420 ,
         \22421 , \22422 , \22423 , \22424 , \22425 , \22426 , \22427 , \22428 , \22429 , \22430 ,
         \22431 , \22432 , \22433 , \22434 , \22435 , \22436 , \22437 , \22438 , \22439 , \22440 ,
         \22441 , \22442 , \22443 , \22444 , \22445 , \22446 , \22447 , \22448 , \22449 , \22450 ,
         \22451 , \22452 , \22453 , \22454 , \22455 , \22456 , \22457 , \22458 , \22459 , \22460 ,
         \22461 , \22462 , \22463 , \22464 , \22465 , \22466 , \22467 , \22468 , \22469 , \22470 ,
         \22471 , \22472 , \22473 , \22474 , \22475 , \22476 , \22477 , \22478 , \22479 , \22480 ,
         \22481 , \22482 , \22483 , \22484 , \22485 , \22486 , \22487 , \22488 , \22489 , \22490 ,
         \22491 , \22492 , \22493 , \22494 , \22495 , \22496 , \22497 , \22498 , \22499 , \22500 ,
         \22501 , \22502 , \22503 , \22504 , \22505 , \22506 , \22507 , \22508 , \22509 , \22510 ,
         \22511 , \22512 , \22513 , \22514 , \22515 , \22516 , \22517 , \22518 , \22519 , \22520 ,
         \22521 , \22522 , \22523 , \22524 , \22525 , \22526 , \22527 , \22528 , \22529 , \22530 ,
         \22531 , \22532 , \22533 , \22534 , \22535 , \22536 , \22537 , \22538 , \22539 , \22540 ,
         \22541 , \22542 , \22543 , \22544 , \22545 , \22546 , \22547 , \22548 , \22549 , \22550 ,
         \22551 , \22552 , \22553 , \22554 , \22555 , \22556 , \22557 , \22558 , \22559 , \22560 ,
         \22561 , \22562 , \22563 , \22564 , \22565 , \22566 , \22567 , \22568 , \22569 , \22570 ,
         \22571 , \22572 , \22573 , \22574 , \22575 , \22576 , \22577 , \22578 , \22579 , \22580 ,
         \22581 , \22582 , \22583 , \22584 , \22585 , \22586 , \22587 , \22588 , \22589 , \22590 ,
         \22591 , \22592 , \22593 , \22594 , \22595 , \22596 , \22597 , \22598 , \22599 , \22600 ,
         \22601 , \22602 , \22603 , \22604 , \22605 , \22606 , \22607 , \22608 , \22609 , \22610 ,
         \22611 , \22612 , \22613 , \22614 , \22615 , \22616 , \22617 , \22618 , \22619 , \22620 ,
         \22621 , \22622 , \22623 , \22624 , \22625 , \22626 , \22627 , \22628 , \22629 , \22630 ,
         \22631 , \22632 , \22633 , \22634 , \22635 , \22636 , \22637 , \22638 , \22639 , \22640 ,
         \22641 , \22642 , \22643 , \22644 , \22645 , \22646 , \22647 , \22648 , \22649 , \22650 ,
         \22651 , \22652 , \22653 , \22654 , \22655 , \22656 , \22657 , \22658 , \22659 , \22660 ,
         \22661 , \22662 , \22663 , \22664 , \22665 , \22666 , \22667 , \22668 , \22669 , \22670 ,
         \22671 , \22672 , \22673 , \22674 , \22675 , \22676 , \22677 , \22678 , \22679 , \22680 ,
         \22681 , \22682 , \22683 , \22684 , \22685 , \22686 , \22687 , \22688 , \22689 , \22690 ,
         \22691 , \22692 , \22693 , \22694 , \22695 , \22696 , \22697 , \22698 , \22699 , \22700 ,
         \22701 , \22702 , \22703 , \22704 , \22705 , \22706 , \22707 , \22708 , \22709 , \22710 ,
         \22711 , \22712 , \22713 , \22714 , \22715 , \22716 , \22717 , \22718 , \22719 , \22720 ,
         \22721 , \22722 , \22723 , \22724 , \22725 , \22726 , \22727 , \22728 , \22729 , \22730 ,
         \22731 , \22732 , \22733 , \22734 , \22735 , \22736 , \22737 , \22738 , \22739 , \22740 ,
         \22741 , \22742 , \22743 , \22744 , \22745 , \22746 , \22747 , \22748 , \22749 , \22750 ,
         \22751 , \22752 , \22753 , \22754 , \22755 , \22756 , \22757 , \22758 , \22759 , \22760 ,
         \22761 , \22762 , \22763 , \22764 , \22765 , \22766 , \22767 , \22768 , \22769 , \22770 ,
         \22771 , \22772 , \22773 , \22774 , \22775 , \22776 , \22777 , \22778 , \22779 , \22780 ,
         \22781 , \22782 , \22783 , \22784 , \22785 , \22786 , \22787 , \22788 , \22789 , \22790 ,
         \22791 , \22792 , \22793 , \22794 , \22795 , \22796 , \22797 , \22798 , \22799 , \22800 ,
         \22801 , \22802 , \22803 , \22804 , \22805 , \22806 , \22807 , \22808 , \22809 , \22810 ,
         \22811 , \22812 , \22813 , \22814 , \22815 , \22816 , \22817 , \22818 , \22819 , \22820 ,
         \22821 , \22822 , \22823 , \22824 , \22825 , \22826 , \22827 , \22828 , \22829 , \22830 ,
         \22831 , \22832 , \22833 , \22834 , \22835 , \22836 , \22837 , \22838 , \22839 , \22840 ,
         \22841 , \22842 , \22843 , \22844 , \22845 , \22846 , \22847 , \22848 , \22849 , \22850 ,
         \22851 , \22852 , \22853 , \22854 , \22855 , \22856 , \22857 , \22858 , \22859 , \22860 ,
         \22861 , \22862 , \22863 , \22864 , \22865 , \22866 , \22867 , \22868 , \22869 , \22870 ,
         \22871 , \22872 , \22873 , \22874 , \22875 , \22876 , \22877 , \22878 , \22879 , \22880 ,
         \22881 , \22882 , \22883 , \22884 , \22885 , \22886 , \22887 , \22888 , \22889 , \22890 ,
         \22891 , \22892 , \22893 , \22894 , \22895 , \22896 , \22897 , \22898 , \22899 , \22900 ,
         \22901 , \22902 , \22903 , \22904 , \22905 , \22906 , \22907 , \22908 , \22909 , \22910 ,
         \22911 , \22912 , \22913 , \22914 , \22915 , \22916 , \22917 , \22918 , \22919 , \22920 ,
         \22921 , \22922 , \22923 , \22924 , \22925 , \22926 , \22927 , \22928 , \22929 , \22930 ,
         \22931 , \22932 , \22933 , \22934 , \22935 , \22936 , \22937 , \22938 , \22939 , \22940 ,
         \22941 , \22942 , \22943 , \22944 , \22945 , \22946 , \22947 , \22948 , \22949 , \22950 ,
         \22951 , \22952 , \22953 , \22954 , \22955 , \22956 , \22957 , \22958 , \22959 , \22960 ,
         \22961 , \22962 , \22963 , \22964 , \22965 , \22966 , \22967 , \22968 , \22969 , \22970 ,
         \22971 , \22972 , \22973 , \22974 , \22975 , \22976 , \22977 , \22978 , \22979 , \22980 ,
         \22981 , \22982 , \22983 , \22984 , \22985 , \22986 , \22987 , \22988 , \22989 , \22990 ,
         \22991 , \22992 , \22993 , \22994 , \22995 , \22996 , \22997 , \22998 , \22999 , \23000 ,
         \23001 , \23002 , \23003 , \23004 , \23005 , \23006 , \23007 , \23008 , \23009 , \23010 ,
         \23011 , \23012 , \23013 , \23014 , \23015 , \23016 , \23017 , \23018 , \23019 , \23020 ,
         \23021 , \23022 , \23023 , \23024 , \23025 , \23026 , \23027 , \23028 , \23029 , \23030 ,
         \23031 , \23032 , \23033 , \23034 , \23035 , \23036 , \23037 , \23038 , \23039 , \23040 ,
         \23041 , \23042 , \23043 , \23044 , \23045 , \23046 , \23047 , \23048 , \23049 , \23050 ,
         \23051 , \23052 , \23053 , \23054 , \23055 , \23056 , \23057 , \23058 , \23059 , \23060 ,
         \23061 , \23062 , \23063 , \23064 , \23065 , \23066 , \23067 , \23068 , \23069 , \23070 ,
         \23071 , \23072 , \23073 , \23074 , \23075 , \23076 , \23077 , \23078 , \23079 , \23080 ,
         \23081 , \23082 , \23083 , \23084 , \23085 , \23086 , \23087 , \23088 , \23089 , \23090 ,
         \23091 , \23092 , \23093 , \23094 , \23095 , \23096 , \23097 , \23098 , \23099 , \23100 ,
         \23101 , \23102 , \23103 , \23104 , \23105 , \23106 , \23107 , \23108 , \23109 , \23110 ,
         \23111 , \23112 , \23113 , \23114 , \23115 , \23116 , \23117 , \23118 , \23119 , \23120 ,
         \23121 , \23122 , \23123 , \23124 , \23125 , \23126 , \23127 , \23128 , \23129 , \23130 ,
         \23131 , \23132 , \23133 , \23134 , \23135 , \23136 , \23137 , \23138 , \23139 , \23140 ,
         \23141 , \23142 , \23143 , \23144 , \23145 , \23146 , \23147 , \23148 , \23149 , \23150 ,
         \23151 , \23152 , \23153 , \23154 , \23155 , \23156 , \23157 , \23158 , \23159 , \23160 ,
         \23161 , \23162 , \23163 , \23164 , \23165 , \23166 , \23167 , \23168 , \23169 , \23170 ,
         \23171 , \23172 , \23173 , \23174 , \23175 , \23176 , \23177 , \23178 , \23179 , \23180 ,
         \23181 , \23182 , \23183 , \23184 , \23185 , \23186 , \23187 , \23188 , \23189 , \23190 ,
         \23191 , \23192 , \23193 , \23194 , \23195 , \23196 , \23197 , \23198 , \23199 , \23200 ,
         \23201 , \23202 , \23203 , \23204 , \23205 , \23206 , \23207 , \23208 , \23209 , \23210 ,
         \23211 , \23212 , \23213 , \23214 , \23215 , \23216 , \23217 , \23218 , \23219 , \23220 ,
         \23221 , \23222 , \23223 , \23224 , \23225 , \23226 , \23227 , \23228 , \23229 , \23230 ,
         \23231 , \23232 , \23233 , \23234 , \23235 , \23236 , \23237 , \23238 , \23239 , \23240 ,
         \23241 , \23242 , \23243 , \23244 , \23245 , \23246 , \23247 , \23248 , \23249 , \23250 ,
         \23251 , \23252 , \23253 , \23254 , \23255 , \23256 , \23257 , \23258 , \23259 , \23260 ,
         \23261 , \23262 , \23263 , \23264 , \23265 , \23266 , \23267 , \23268 , \23269 , \23270 ,
         \23271 , \23272 , \23273 , \23274 , \23275 , \23276 , \23277 , \23278 , \23279 , \23280 ,
         \23281 , \23282 , \23283 , \23284 , \23285 , \23286 , \23287 , \23288 , \23289 , \23290 ,
         \23291 , \23292 , \23293 , \23294 , \23295 , \23296 , \23297 , \23298 , \23299 , \23300 ,
         \23301 , \23302 , \23303 , \23304 , \23305 , \23306 , \23307 , \23308 , \23309 , \23310 ,
         \23311 , \23312 , \23313 , \23314 , \23315 , \23316 , \23317 , \23318 , \23319 , \23320 ,
         \23321 , \23322 , \23323 , \23324 , \23325 , \23326 , \23327 , \23328 , \23329 , \23330 ,
         \23331 , \23332 , \23333 , \23334 , \23335 , \23336 , \23337 , \23338 , \23339 , \23340 ,
         \23341 , \23342 , \23343 , \23344 , \23345 , \23346 , \23347 , \23348 , \23349 , \23350 ,
         \23351 , \23352 , \23353 , \23354 , \23355 , \23356 , \23357 , \23358 , \23359 , \23360 ,
         \23361 , \23362 , \23363 , \23364 , \23365 , \23366 , \23367 , \23368 , \23369 , \23370 ,
         \23371 , \23372 , \23373 , \23374 , \23375 , \23376 , \23377 , \23378 , \23379 , \23380 ,
         \23381 , \23382 , \23383 , \23384 , \23385 , \23386 , \23387 , \23388 , \23389 , \23390 ,
         \23391 , \23392 , \23393 , \23394 , \23395 , \23396 , \23397 , \23398 , \23399 , \23400 ,
         \23401 , \23402 , \23403 , \23404 , \23405 , \23406 , \23407 , \23408 , \23409 , \23410 ,
         \23411 , \23412 , \23413 , \23414 , \23415 , \23416 , \23417 , \23418 , \23419 , \23420 ,
         \23421 , \23422 , \23423 , \23424 , \23425 , \23426 , \23427 , \23428 , \23429 , \23430 ,
         \23431 , \23432 , \23433 , \23434 , \23435 , \23436 , \23437 , \23438 , \23439 , \23440 ,
         \23441 , \23442 , \23443 , \23444 , \23445 , \23446 , \23447 , \23448 , \23449 , \23450 ,
         \23451 , \23452 , \23453 , \23454 , \23455 , \23456 , \23457 , \23458 , \23459 , \23460 ,
         \23461 , \23462 , \23463 , \23464 , \23465 , \23466 , \23467 , \23468 , \23469 , \23470 ,
         \23471 , \23472 , \23473 , \23474 , \23475 , \23476 , \23477 , \23478 , \23479 , \23480 ,
         \23481 , \23482 , \23483 , \23484 , \23485 , \23486 , \23487 , \23488 , \23489 , \23490 ,
         \23491 , \23492 , \23493 , \23494 , \23495 , \23496 , \23497 , \23498 , \23499 , \23500 ,
         \23501 , \23502 , \23503 , \23504 , \23505 , \23506 , \23507 , \23508 , \23509 , \23510 ,
         \23511 , \23512 , \23513 , \23514 , \23515 , \23516 , \23517 , \23518 , \23519 , \23520 ,
         \23521 , \23522 , \23523 , \23524 , \23525 , \23526 , \23527 , \23528 , \23529 , \23530 ,
         \23531 , \23532 , \23533 , \23534 , \23535 , \23536 , \23537 , \23538 , \23539 , \23540 ,
         \23541 , \23542 , \23543 , \23544 , \23545 , \23546 , \23547 , \23548 , \23549 , \23550 ,
         \23551 , \23552 , \23553 , \23554 , \23555 , \23556 , \23557 , \23558 , \23559 , \23560 ,
         \23561 , \23562 , \23563 , \23564 , \23565 , \23566 , \23567 , \23568 , \23569 , \23570 ,
         \23571 , \23572 , \23573 , \23574 , \23575 , \23576 , \23577 , \23578 , \23579 , \23580 ,
         \23581 , \23582 , \23583 , \23584 , \23585 , \23586 , \23587 , \23588 , \23589 , \23590 ,
         \23591 , \23592 , \23593 , \23594 , \23595 , \23596 , \23597 , \23598 , \23599 , \23600 ,
         \23601 , \23602 , \23603 , \23604 , \23605 , \23606 , \23607 , \23608 , \23609 , \23610 ,
         \23611 , \23612 , \23613 , \23614 , \23615 , \23616 , \23617 , \23618 , \23619 , \23620 ,
         \23621 , \23622 , \23623 , \23624 , \23625 , \23626 , \23627 , \23628 , \23629 , \23630 ,
         \23631 , \23632 , \23633 , \23634 , \23635 , \23636 , \23637 , \23638 , \23639 , \23640 ,
         \23641 , \23642 , \23643 , \23644 , \23645 , \23646 , \23647 , \23648 , \23649 , \23650 ,
         \23651 , \23652 , \23653 , \23654 , \23655 , \23656 , \23657 , \23658 , \23659 , \23660 ,
         \23661 , \23662 , \23663 , \23664 , \23665 , \23666 , \23667 , \23668 , \23669 , \23670 ,
         \23671 , \23672 , \23673 , \23674 , \23675 , \23676 , \23677 , \23678 , \23679 , \23680 ,
         \23681 , \23682 , \23683 , \23684 , \23685 , \23686 , \23687 , \23688 , \23689 , \23690 ,
         \23691 , \23692 , \23693 , \23694 , \23695 , \23696 , \23697 , \23698 , \23699 , \23700 ,
         \23701 , \23702 , \23703 , \23704 , \23705 , \23706 , \23707 , \23708 , \23709 , \23710 ,
         \23711 , \23712 , \23713 , \23714 , \23715 , \23716 , \23717 , \23718 , \23719 , \23720 ,
         \23721 , \23722 , \23723 , \23724 , \23725 , \23726 , \23727 , \23728 , \23729 , \23730 ,
         \23731 , \23732 , \23733 , \23734 , \23735 , \23736 , \23737 , \23738 , \23739 , \23740 ,
         \23741 , \23742 , \23743 , \23744 , \23745 , \23746 , \23747 , \23748 , \23749 , \23750 ,
         \23751 , \23752 , \23753 , \23754 , \23755 , \23756 , \23757 , \23758 , \23759 , \23760 ,
         \23761 , \23762 , \23763 , \23764 , \23765 , \23766 , \23767 , \23768 , \23769 , \23770 ,
         \23771 , \23772 , \23773 , \23774 , \23775 , \23776 , \23777 , \23778 , \23779 , \23780 ,
         \23781 , \23782 , \23783 , \23784 , \23785 , \23786 , \23787 , \23788 , \23789 , \23790 ,
         \23791 , \23792 , \23793 , \23794 , \23795 , \23796 , \23797 , \23798 , \23799 , \23800 ,
         \23801 , \23802 , \23803 , \23804 , \23805 , \23806 , \23807 , \23808 , \23809 , \23810 ,
         \23811 , \23812 , \23813 , \23814 , \23815 , \23816 , \23817 , \23818 , \23819 , \23820 ,
         \23821 , \23822 , \23823 , \23824 , \23825 , \23826 , \23827 , \23828 , \23829 , \23830 ,
         \23831 , \23832 , \23833 , \23834 , \23835 , \23836 , \23837 , \23838 , \23839 , \23840 ,
         \23841 , \23842 , \23843 , \23844 , \23845 , \23846 , \23847 , \23848 , \23849 , \23850 ,
         \23851 , \23852 , \23853 , \23854 , \23855 , \23856 , \23857 , \23858 , \23859 , \23860 ,
         \23861 , \23862 , \23863 , \23864 , \23865 , \23866 , \23867 , \23868 , \23869 , \23870 ,
         \23871 , \23872 , \23873 , \23874 , \23875 , \23876 , \23877 , \23878 , \23879 , \23880 ,
         \23881 , \23882 , \23883 , \23884 , \23885 , \23886 , \23887 , \23888 , \23889 , \23890 ,
         \23891 , \23892 , \23893 , \23894 , \23895 , \23896 , \23897 , \23898 , \23899 , \23900 ,
         \23901 , \23902 , \23903 , \23904 , \23905 , \23906 , \23907 , \23908 , \23909 , \23910 ,
         \23911 , \23912 , \23913 , \23914 , \23915 , \23916 , \23917 , \23918 , \23919 , \23920 ,
         \23921 , \23922 , \23923 , \23924 , \23925 , \23926 , \23927 , \23928 , \23929 , \23930 ,
         \23931 , \23932 , \23933 , \23934 , \23935 , \23936 , \23937 , \23938 , \23939 , \23940 ,
         \23941 , \23942 , \23943 , \23944 , \23945 , \23946 , \23947 , \23948 , \23949 , \23950 ,
         \23951 , \23952 , \23953 , \23954 , \23955 , \23956 , \23957 , \23958 , \23959 , \23960 ,
         \23961 , \23962 , \23963 , \23964 , \23965 , \23966 , \23967 , \23968 , \23969 , \23970 ,
         \23971 , \23972 , \23973 , \23974 , \23975 , \23976 , \23977 , \23978 , \23979 , \23980 ,
         \23981 , \23982 , \23983 , \23984 , \23985 , \23986 , \23987 , \23988 , \23989 , \23990 ,
         \23991 , \23992 , \23993 , \23994 , \23995 , \23996 , \23997 , \23998 , \23999 , \24000 ,
         \24001 , \24002 , \24003 , \24004 , \24005 , \24006 , \24007 , \24008 , \24009 , \24010 ,
         \24011 , \24012 , \24013 , \24014 , \24015 , \24016 , \24017 , \24018 , \24019 , \24020 ,
         \24021 , \24022 , \24023 , \24024 , \24025 , \24026 , \24027 , \24028 , \24029 , \24030 ,
         \24031 , \24032 , \24033 , \24034 , \24035 , \24036 , \24037 , \24038 , \24039 , \24040 ,
         \24041 , \24042 , \24043 , \24044 , \24045 , \24046 , \24047 , \24048 , \24049 , \24050 ,
         \24051 , \24052 , \24053 , \24054 , \24055 , \24056 , \24057 , \24058 , \24059 , \24060 ,
         \24061 , \24062 , \24063 , \24064 , \24065 , \24066 , \24067 , \24068 , \24069 , \24070 ,
         \24071 , \24072 , \24073 , \24074 , \24075 , \24076 , \24077 , \24078 , \24079 , \24080 ,
         \24081 , \24082 , \24083 , \24084 , \24085 , \24086 , \24087 , \24088 , \24089 , \24090 ,
         \24091 , \24092 , \24093 , \24094 , \24095 , \24096 , \24097 , \24098 , \24099 , \24100 ,
         \24101 , \24102 , \24103 , \24104 , \24105 , \24106 , \24107 , \24108 , \24109 , \24110 ,
         \24111 , \24112 , \24113 , \24114 , \24115 , \24116 , \24117 , \24118 , \24119 , \24120 ,
         \24121 , \24122 , \24123 , \24124 , \24125 , \24126 , \24127 , \24128 , \24129 , \24130 ,
         \24131 , \24132 , \24133 , \24134 , \24135 , \24136 , \24137 , \24138 , \24139 , \24140 ,
         \24141 , \24142 , \24143 , \24144 , \24145 , \24146 , \24147 , \24148 , \24149 , \24150 ,
         \24151 , \24152 , \24153 , \24154 , \24155 , \24156 , \24157 , \24158 , \24159 , \24160 ,
         \24161 , \24162 , \24163 , \24164 , \24165 , \24166 , \24167 , \24168 , \24169 , \24170 ,
         \24171 , \24172 , \24173 , \24174 , \24175 , \24176 , \24177 , \24178 , \24179 , \24180 ,
         \24181 , \24182 , \24183 , \24184 , \24185 , \24186 , \24187 , \24188 , \24189 , \24190 ,
         \24191 , \24192 , \24193 , \24194 , \24195 , \24196 , \24197 , \24198 , \24199 , \24200 ,
         \24201 , \24202 , \24203 , \24204 , \24205 , \24206 , \24207 , \24208 , \24209 , \24210 ,
         \24211 , \24212 , \24213 , \24214 , \24215 , \24216 , \24217 , \24218 , \24219 , \24220 ,
         \24221 , \24222 , \24223 , \24224 , \24225 , \24226 , \24227 , \24228 , \24229 , \24230 ,
         \24231 , \24232 , \24233 , \24234 , \24235 , \24236 , \24237 , \24238 , \24239 , \24240 ,
         \24241 , \24242 , \24243 , \24244 , \24245 , \24246 , \24247 , \24248 , \24249 , \24250 ,
         \24251 , \24252 , \24253 , \24254 , \24255 , \24256 , \24257 , \24258 , \24259 , \24260 ,
         \24261 , \24262 , \24263 , \24264 , \24265 , \24266 , \24267 , \24268 , \24269 , \24270 ,
         \24271 , \24272 , \24273 , \24274 , \24275 , \24276 , \24277 , \24278 , \24279 , \24280 ,
         \24281 , \24282 , \24283 , \24284 , \24285 , \24286 , \24287 , \24288 , \24289 , \24290 ,
         \24291 , \24292 , \24293 , \24294 , \24295 , \24296 , \24297 , \24298 , \24299 , \24300 ,
         \24301 , \24302 , \24303 , \24304 , \24305 , \24306 , \24307 , \24308 , \24309 , \24310 ,
         \24311 , \24312 , \24313 , \24314 , \24315 , \24316 , \24317 , \24318 , \24319 , \24320 ,
         \24321 , \24322 , \24323 , \24324 , \24325 , \24326 , \24327 , \24328 , \24329 , \24330 ,
         \24331 , \24332 , \24333 , \24334 , \24335 , \24336 , \24337 , \24338 , \24339 , \24340 ,
         \24341 , \24342 , \24343 , \24344 , \24345 , \24346 , \24347 , \24348 , \24349 , \24350 ,
         \24351 , \24352 , \24353 , \24354 , \24355 , \24356 , \24357 , \24358 , \24359 , \24360 ,
         \24361 , \24362 , \24363 , \24364 , \24365 , \24366 , \24367 , \24368 , \24369 , \24370 ,
         \24371 , \24372 , \24373 , \24374 , \24375 , \24376 , \24377 , \24378 , \24379 , \24380 ,
         \24381 , \24382 , \24383 , \24384 , \24385 , \24386 , \24387 , \24388 , \24389 , \24390 ,
         \24391 , \24392 , \24393 , \24394 , \24395 , \24396 , \24397 , \24398 , \24399 , \24400 ,
         \24401 , \24402 , \24403 , \24404 , \24405 , \24406 , \24407 , \24408 , \24409 , \24410 ,
         \24411 , \24412 , \24413 , \24414 , \24415 , \24416 , \24417 , \24418 , \24419 , \24420 ,
         \24421 , \24422 , \24423 , \24424 , \24425 , \24426 , \24427 , \24428 , \24429 , \24430 ,
         \24431 , \24432 , \24433 , \24434 , \24435 , \24436 , \24437 , \24438 , \24439 , \24440 ,
         \24441 , \24442 , \24443 , \24444 , \24445 , \24446 , \24447 , \24448 , \24449 , \24450 ,
         \24451 , \24452 , \24453 , \24454 , \24455 , \24456 , \24457 , \24458 , \24459 , \24460 ,
         \24461 , \24462 , \24463 , \24464 , \24465 , \24466 , \24467 , \24468 , \24469 , \24470 ,
         \24471 , \24472 , \24473 , \24474 , \24475 , \24476 , \24477 , \24478 , \24479 , \24480 ,
         \24481 , \24482 , \24483 , \24484 , \24485 , \24486 , \24487 , \24488 , \24489 , \24490 ,
         \24491 , \24492 , \24493 , \24494 , \24495 , \24496 , \24497 , \24498 , \24499 , \24500 ,
         \24501 , \24502 , \24503 , \24504 , \24505 , \24506 , \24507 , \24508 , \24509 , \24510 ,
         \24511 , \24512 , \24513 , \24514 , \24515 , \24516 , \24517 , \24518 , \24519 , \24520 ,
         \24521 , \24522 , \24523 , \24524 , \24525 , \24526 , \24527 , \24528 , \24529 , \24530 ,
         \24531 , \24532 , \24533 , \24534 , \24535 , \24536 , \24537 , \24538 , \24539 , \24540 ,
         \24541 , \24542 , \24543 , \24544 , \24545 , \24546 , \24547 , \24548 , \24549 , \24550 ,
         \24551 , \24552 , \24553 , \24554 , \24555 , \24556 , \24557 , \24558 , \24559 , \24560 ,
         \24561 , \24562 , \24563 , \24564 , \24565 , \24566 , \24567 , \24568 , \24569 , \24570 ,
         \24571 , \24572 , \24573 , \24574 , \24575 , \24576 , \24577 , \24578 , \24579 , \24580 ,
         \24581 , \24582 , \24583 , \24584 , \24585 , \24586 , \24587 , \24588 , \24589 , \24590 ,
         \24591 , \24592 , \24593 , \24594 , \24595 , \24596 , \24597 , \24598 , \24599 , \24600 ,
         \24601 , \24602 , \24603 , \24604 , \24605 , \24606 , \24607 , \24608 , \24609 , \24610 ,
         \24611 , \24612 , \24613 , \24614 , \24615 , \24616 , \24617 , \24618 , \24619 , \24620 ,
         \24621 , \24622 , \24623 , \24624 , \24625 , \24626 , \24627 , \24628 , \24629 , \24630 ,
         \24631 , \24632 , \24633 , \24634 , \24635 , \24636 , \24637 , \24638 , \24639 , \24640 ,
         \24641 , \24642 , \24643 , \24644 , \24645 , \24646 , \24647 , \24648 , \24649 , \24650 ,
         \24651 , \24652 , \24653 , \24654 , \24655 , \24656 , \24657 , \24658 , \24659 , \24660 ,
         \24661 , \24662 , \24663 , \24664 , \24665 , \24666 , \24667 , \24668 , \24669 , \24670 ,
         \24671 , \24672 , \24673 , \24674 , \24675 , \24676 , \24677 , \24678 , \24679 , \24680 ,
         \24681 , \24682 , \24683 , \24684 , \24685 , \24686 , \24687 , \24688 , \24689 , \24690 ,
         \24691 , \24692 , \24693 , \24694 , \24695 , \24696 , \24697 , \24698 , \24699 , \24700 ,
         \24701 , \24702 , \24703 , \24704 , \24705 , \24706 , \24707 , \24708 , \24709 , \24710 ,
         \24711 , \24712 , \24713 , \24714 , \24715 , \24716 , \24717 , \24718 , \24719 , \24720 ,
         \24721 , \24722 , \24723 , \24724 , \24725 , \24726 , \24727 , \24728 , \24729 , \24730 ,
         \24731 , \24732 , \24733 , \24734 , \24735 , \24736 , \24737 , \24738 , \24739 , \24740 ,
         \24741 , \24742 , \24743 , \24744 , \24745 , \24746 , \24747 , \24748 , \24749 , \24750 ,
         \24751 , \24752 , \24753 , \24754 , \24755 , \24756 , \24757 , \24758 , \24759 , \24760 ,
         \24761 , \24762 , \24763 , \24764 , \24765 , \24766 , \24767 , \24768 , \24769 , \24770 ,
         \24771 , \24772 , \24773 , \24774 , \24775 , \24776 , \24777 , \24778 , \24779 , \24780 ,
         \24781 , \24782 , \24783 , \24784 , \24785 , \24786 , \24787 , \24788 , \24789 , \24790 ,
         \24791 , \24792 , \24793 , \24794 , \24795 , \24796 , \24797 , \24798 , \24799 , \24800 ,
         \24801 , \24802 , \24803 , \24804 , \24805 , \24806 , \24807 , \24808 , \24809 , \24810 ,
         \24811 , \24812 , \24813 , \24814 , \24815 , \24816 , \24817 , \24818 , \24819 , \24820 ,
         \24821 , \24822 , \24823 , \24824 , \24825 , \24826 , \24827 , \24828 , \24829 , \24830 ,
         \24831 , \24832 , \24833 , \24834 , \24835 , \24836 , \24837 , \24838 , \24839 , \24840 ,
         \24841 , \24842 , \24843 , \24844 , \24845 , \24846 , \24847 , \24848 , \24849 , \24850 ,
         \24851 , \24852 , \24853 , \24854 , \24855 , \24856 , \24857 , \24858 , \24859 , \24860 ,
         \24861 , \24862 , \24863 , \24864 , \24865 , \24866 , \24867 , \24868 , \24869 , \24870 ,
         \24871 , \24872 , \24873 , \24874 , \24875 , \24876 , \24877 , \24878 , \24879 , \24880 ,
         \24881 , \24882 , \24883 , \24884 , \24885 , \24886 , \24887 , \24888 , \24889 , \24890 ,
         \24891 , \24892 , \24893 , \24894 , \24895 , \24896 , \24897 , \24898 , \24899 , \24900 ,
         \24901 , \24902 , \24903 , \24904 , \24905 , \24906 , \24907 , \24908 , \24909 , \24910 ,
         \24911 , \24912 , \24913 , \24914 , \24915 , \24916 , \24917 , \24918 , \24919 , \24920 ,
         \24921 , \24922 , \24923 , \24924 , \24925 , \24926 , \24927 , \24928 , \24929 , \24930 ,
         \24931 , \24932 , \24933 , \24934 , \24935 , \24936 , \24937 , \24938 , \24939 , \24940 ,
         \24941 , \24942 , \24943 , \24944 , \24945 , \24946 , \24947 , \24948 , \24949 , \24950 ,
         \24951 , \24952 , \24953 , \24954 , \24955 , \24956 , \24957 , \24958 , \24959 , \24960 ,
         \24961 , \24962 , \24963 , \24964 , \24965 , \24966 , \24967 , \24968 , \24969 , \24970 ,
         \24971 , \24972 , \24973 , \24974 , \24975 , \24976 , \24977 , \24978 , \24979 , \24980 ,
         \24981 , \24982 , \24983 , \24984 , \24985 , \24986 , \24987 , \24988 , \24989 , \24990 ,
         \24991 , \24992 , \24993 , \24994 , \24995 , \24996 , \24997 , \24998 , \24999 , \25000 ,
         \25001 , \25002 , \25003 , \25004 , \25005 , \25006 , \25007 , \25008 , \25009 , \25010 ,
         \25011 , \25012 , \25013 , \25014 , \25015 , \25016 , \25017 , \25018 , \25019 , \25020 ,
         \25021 , \25022 , \25023 , \25024 , \25025 , \25026 , \25027 , \25028 , \25029 , \25030 ,
         \25031 , \25032 , \25033 , \25034 , \25035 , \25036 , \25037 , \25038 , \25039 , \25040 ,
         \25041 , \25042 , \25043 , \25044 , \25045 , \25046 , \25047 , \25048 , \25049 , \25050 ,
         \25051 , \25052 , \25053 , \25054 , \25055 , \25056 , \25057 , \25058 , \25059 , \25060 ,
         \25061 , \25062 , \25063 , \25064 , \25065 , \25066 , \25067 , \25068 , \25069 , \25070 ,
         \25071 , \25072 , \25073 , \25074 , \25075 , \25076 , \25077 , \25078 , \25079 , \25080 ,
         \25081 , \25082 , \25083 , \25084 , \25085 , \25086 , \25087 , \25088 , \25089 , \25090 ,
         \25091 , \25092 , \25093 , \25094 , \25095 , \25096 , \25097 , \25098 , \25099 , \25100 ,
         \25101 , \25102 , \25103 , \25104 , \25105 , \25106 , \25107 , \25108 , \25109 , \25110 ,
         \25111 , \25112 , \25113 , \25114 , \25115 , \25116 , \25117 , \25118 , \25119 , \25120 ,
         \25121 , \25122 , \25123 , \25124 , \25125 , \25126 , \25127 , \25128 , \25129 , \25130 ,
         \25131 , \25132 , \25133 , \25134 , \25135 , \25136 , \25137 , \25138 , \25139 , \25140 ,
         \25141 , \25142 , \25143 , \25144 , \25145 , \25146 , \25147 , \25148 , \25149 , \25150 ,
         \25151 , \25152 , \25153 , \25154 , \25155 , \25156 , \25157 , \25158 , \25159 , \25160 ,
         \25161 , \25162 , \25163 , \25164 , \25165 , \25166 , \25167 , \25168 , \25169 , \25170 ,
         \25171 , \25172 , \25173 , \25174 , \25175 , \25176 , \25177 , \25178 , \25179 , \25180 ,
         \25181 , \25182 , \25183 , \25184 , \25185 , \25186 , \25187 , \25188 , \25189 , \25190 ,
         \25191 , \25192 , \25193 , \25194 , \25195 , \25196 , \25197 , \25198 , \25199 , \25200 ,
         \25201 , \25202 , \25203 , \25204 , \25205 , \25206 , \25207 , \25208 , \25209 , \25210 ,
         \25211 , \25212 , \25213 , \25214 , \25215 , \25216 , \25217 , \25218 , \25219 , \25220 ,
         \25221 , \25222 , \25223 , \25224 , \25225 , \25226 , \25227 , \25228 , \25229 , \25230 ,
         \25231 , \25232 , \25233 , \25234 , \25235 , \25236 , \25237 , \25238 , \25239 , \25240 ,
         \25241 , \25242 , \25243 , \25244 , \25245 , \25246 , \25247 , \25248 , \25249 , \25250 ,
         \25251 , \25252 , \25253 , \25254 , \25255 , \25256 , \25257 , \25258 , \25259 , \25260 ,
         \25261 , \25262 , \25263 , \25264 , \25265 , \25266 , \25267 , \25268 , \25269 , \25270 ,
         \25271 , \25272 , \25273 , \25274 , \25275 , \25276 , \25277 , \25278 , \25279 , \25280 ,
         \25281 , \25282 , \25283 , \25284 , \25285 , \25286 , \25287 , \25288 , \25289 , \25290 ,
         \25291 , \25292 , \25293 , \25294 , \25295 , \25296 , \25297 , \25298 , \25299 , \25300 ,
         \25301 , \25302 , \25303 , \25304 , \25305 , \25306 , \25307 , \25308 , \25309 , \25310 ,
         \25311 , \25312 , \25313 , \25314 , \25315 , \25316 , \25317 , \25318 , \25319 , \25320 ,
         \25321 , \25322 , \25323 , \25324 , \25325 , \25326 , \25327 , \25328 , \25329 , \25330 ,
         \25331 , \25332 , \25333 , \25334 , \25335 , \25336 , \25337 , \25338 , \25339 , \25340 ,
         \25341 , \25342 , \25343 , \25344 , \25345 , \25346 , \25347 , \25348 , \25349 , \25350 ,
         \25351 , \25352 , \25353 , \25354 , \25355 , \25356 , \25357 , \25358 , \25359 , \25360 ,
         \25361 , \25362 , \25363 , \25364 , \25365 , \25366 , \25367 , \25368 , \25369 , \25370 ,
         \25371 , \25372 , \25373 , \25374 , \25375 , \25376 , \25377 , \25378 , \25379 , \25380 ,
         \25381 , \25382 , \25383 , \25384 , \25385 , \25386 , \25387 , \25388 , \25389 , \25390 ,
         \25391 , \25392 , \25393 , \25394 , \25395 , \25396 , \25397 , \25398 , \25399 , \25400 ,
         \25401 , \25402 , \25403 , \25404 , \25405 , \25406 , \25407 , \25408 , \25409 , \25410 ,
         \25411 , \25412 , \25413 , \25414 , \25415 , \25416 , \25417 , \25418 , \25419 , \25420 ,
         \25421 , \25422 , \25423 , \25424 , \25425 , \25426 , \25427 , \25428 , \25429 , \25430 ,
         \25431 , \25432 , \25433 , \25434 , \25435 , \25436 , \25437 , \25438 , \25439 , \25440 ,
         \25441 , \25442 , \25443 , \25444 , \25445 , \25446 , \25447 , \25448 , \25449 , \25450 ,
         \25451 , \25452 , \25453 , \25454 , \25455 , \25456 , \25457 , \25458 , \25459 , \25460 ,
         \25461 , \25462 , \25463 , \25464 , \25465 , \25466 , \25467 , \25468 , \25469 , \25470 ,
         \25471 , \25472 , \25473 , \25474 , \25475 , \25476 , \25477 , \25478 , \25479 , \25480 ,
         \25481 , \25482 , \25483 , \25484 , \25485 , \25486 , \25487 , \25488 , \25489 , \25490 ,
         \25491 , \25492 , \25493 , \25494 , \25495 , \25496 , \25497 , \25498 , \25499 , \25500 ,
         \25501 , \25502 , \25503 , \25504 , \25505 , \25506 , \25507 , \25508 , \25509 , \25510 ,
         \25511 , \25512 , \25513 , \25514 , \25515 , \25516 , \25517 , \25518 , \25519 , \25520 ,
         \25521 , \25522 , \25523 , \25524 , \25525 , \25526 , \25527 , \25528 , \25529 , \25530 ,
         \25531 , \25532 , \25533 , \25534 , \25535 , \25536 , \25537 , \25538 , \25539 , \25540 ,
         \25541 , \25542 , \25543 , \25544 , \25545 , \25546 , \25547 , \25548 , \25549 , \25550 ,
         \25551 , \25552 , \25553 , \25554 , \25555 , \25556 , \25557 , \25558 , \25559 , \25560 ,
         \25561 , \25562 , \25563 , \25564 , \25565 , \25566 , \25567 , \25568 , \25569 , \25570 ,
         \25571 , \25572 , \25573 , \25574 , \25575 , \25576 , \25577 , \25578 , \25579 , \25580 ,
         \25581 , \25582 , \25583 , \25584 , \25585 , \25586 , \25587 , \25588 , \25589 , \25590 ,
         \25591 , \25592 , \25593 , \25594 , \25595 , \25596 , \25597 , \25598 , \25599 , \25600 ,
         \25601 , \25602 , \25603 , \25604 , \25605 , \25606 , \25607 , \25608 , \25609 , \25610 ,
         \25611 , \25612 , \25613 , \25614 , \25615 , \25616 , \25617 , \25618 , \25619 , \25620 ,
         \25621 , \25622 , \25623 , \25624 , \25625 , \25626 , \25627 , \25628 , \25629 , \25630 ,
         \25631 , \25632 , \25633 , \25634 , \25635 , \25636 , \25637 , \25638 , \25639 , \25640 ,
         \25641 , \25642 , \25643 , \25644 , \25645 , \25646 , \25647 , \25648 , \25649 , \25650 ,
         \25651 , \25652 , \25653 , \25654 , \25655 , \25656 , \25657 , \25658 , \25659 , \25660 ,
         \25661 , \25662 , \25663 , \25664 , \25665 , \25666 , \25667 , \25668 , \25669 , \25670 ,
         \25671 , \25672 , \25673 , \25674 , \25675 , \25676 , \25677 , \25678 , \25679 , \25680 ,
         \25681 , \25682 , \25683 , \25684 , \25685 , \25686 , \25687 , \25688 , \25689 , \25690 ,
         \25691 , \25692 , \25693 , \25694 , \25695 , \25696 , \25697 , \25698 , \25699 , \25700 ,
         \25701 , \25702 , \25703 , \25704 , \25705 , \25706 , \25707 , \25708 , \25709 , \25710 ,
         \25711 , \25712 , \25713 , \25714 , \25715 , \25716 , \25717 , \25718 , \25719 , \25720 ,
         \25721 , \25722 , \25723 , \25724 , \25725 , \25726 , \25727 , \25728 , \25729 , \25730 ,
         \25731 , \25732 , \25733 , \25734 , \25735 , \25736 , \25737 , \25738 , \25739 , \25740 ,
         \25741 , \25742 , \25743 , \25744 , \25745 , \25746 , \25747 , \25748 , \25749 , \25750 ,
         \25751 , \25752 , \25753 , \25754 , \25755 , \25756 , \25757 , \25758 , \25759 , \25760 ,
         \25761 , \25762 , \25763 , \25764 , \25765 , \25766 , \25767 , \25768 , \25769 , \25770 ,
         \25771 , \25772 , \25773 , \25774 , \25775 , \25776 , \25777 , \25778 , \25779 , \25780 ,
         \25781 , \25782 , \25783 , \25784 , \25785 , \25786 , \25787 , \25788 , \25789 , \25790 ,
         \25791 , \25792 , \25793 , \25794 , \25795 , \25796 , \25797 , \25798 , \25799 , \25800 ,
         \25801 , \25802 , \25803 , \25804 , \25805 , \25806 , \25807 , \25808 , \25809 , \25810 ,
         \25811 , \25812 , \25813 , \25814 , \25815 , \25816 , \25817 , \25818 , \25819 , \25820 ,
         \25821 , \25822 , \25823 , \25824 , \25825 , \25826 , \25827 , \25828 , \25829 , \25830 ,
         \25831 , \25832 , \25833 , \25834 , \25835 , \25836 , \25837 , \25838 , \25839 , \25840 ,
         \25841 , \25842 , \25843 , \25844 , \25845 , \25846 , \25847 , \25848 , \25849 , \25850 ,
         \25851 , \25852 , \25853 , \25854 , \25855 , \25856 , \25857 , \25858 , \25859 , \25860 ,
         \25861 , \25862 , \25863 , \25864 , \25865 , \25866 , \25867 , \25868 , \25869 , \25870 ,
         \25871 , \25872 , \25873 , \25874 , \25875 , \25876 , \25877 , \25878 , \25879 , \25880 ,
         \25881 , \25882 , \25883 , \25884 , \25885 , \25886 , \25887 , \25888 , \25889 , \25890 ,
         \25891 , \25892 , \25893 , \25894 , \25895 , \25896 , \25897 , \25898 , \25899 , \25900 ,
         \25901 , \25902 , \25903 , \25904 , \25905 , \25906 , \25907 , \25908 , \25909 , \25910 ,
         \25911 , \25912 , \25913 , \25914 , \25915 , \25916 , \25917 , \25918 , \25919 , \25920 ,
         \25921 , \25922 , \25923 , \25924 , \25925 , \25926 , \25927 , \25928 , \25929 , \25930 ,
         \25931 , \25932 , \25933 , \25934 , \25935 , \25936 , \25937 , \25938 , \25939 , \25940 ,
         \25941 , \25942 , \25943 , \25944 , \25945 , \25946 , \25947 , \25948 , \25949 , \25950 ,
         \25951 , \25952 , \25953 , \25954 , \25955 , \25956 , \25957 , \25958 , \25959 , \25960 ,
         \25961 , \25962 , \25963 , \25964 , \25965 , \25966 , \25967 , \25968 , \25969 , \25970 ,
         \25971 , \25972 , \25973 , \25974 , \25975 , \25976 , \25977 , \25978 , \25979 , \25980 ,
         \25981 , \25982 , \25983 , \25984 , \25985 , \25986 , \25987 , \25988 , \25989 , \25990 ,
         \25991 , \25992 , \25993 , \25994 , \25995 , \25996 , \25997 , \25998 , \25999 , \26000 ,
         \26001 , \26002 , \26003 , \26004 , \26005 , \26006 , \26007 , \26008 , \26009 , \26010 ,
         \26011 , \26012 , \26013 , \26014 , \26015 , \26016 , \26017 , \26018 , \26019 , \26020 ,
         \26021 , \26022 , \26023 , \26024 , \26025 , \26026 , \26027 , \26028 , \26029 , \26030 ,
         \26031 , \26032 , \26033 , \26034 , \26035 , \26036 , \26037 , \26038 , \26039 , \26040 ,
         \26041 , \26042 , \26043 , \26044 , \26045 , \26046 , \26047 , \26048 , \26049 , \26050 ,
         \26051 , \26052 , \26053 , \26054 , \26055 , \26056 , \26057 , \26058 , \26059 , \26060 ,
         \26061 , \26062 , \26063 , \26064 , \26065 , \26066 , \26067 , \26068 , \26069 , \26070 ,
         \26071 , \26072 , \26073 , \26074 , \26075 , \26076 , \26077 , \26078 , \26079 , \26080 ,
         \26081 , \26082 , \26083 , \26084 , \26085 , \26086 , \26087 , \26088 , \26089 , \26090 ,
         \26091 , \26092 , \26093 , \26094 , \26095 , \26096 , \26097 , \26098 , \26099 , \26100 ,
         \26101 , \26102 , \26103 , \26104 , \26105 , \26106 , \26107 , \26108 , \26109 , \26110 ,
         \26111 , \26112 , \26113 , \26114 , \26115 , \26116 , \26117 , \26118 , \26119 , \26120 ,
         \26121 , \26122 , \26123 , \26124 , \26125 , \26126 , \26127 , \26128 , \26129 , \26130 ,
         \26131 , \26132 , \26133 , \26134 , \26135 , \26136 , \26137 , \26138 , \26139 , \26140 ,
         \26141 , \26142 , \26143 , \26144 , \26145 , \26146 , \26147 , \26148 , \26149 , \26150 ,
         \26151 , \26152 , \26153 , \26154 , \26155 , \26156 , \26157 , \26158 , \26159 , \26160 ,
         \26161 , \26162 , \26163 , \26164 , \26165 , \26166 , \26167 , \26168 , \26169 , \26170 ,
         \26171 , \26172 , \26173 , \26174 , \26175 , \26176 , \26177 , \26178 , \26179 , \26180 ,
         \26181 , \26182 , \26183 , \26184 , \26185 , \26186 , \26187 , \26188 , \26189 , \26190 ,
         \26191 , \26192 , \26193 , \26194 , \26195 , \26196 , \26197 , \26198 , \26199 , \26200 ,
         \26201 , \26202 , \26203 , \26204 , \26205 , \26206 , \26207 , \26208 , \26209 , \26210 ,
         \26211 , \26212 , \26213 , \26214 , \26215 , \26216 , \26217 , \26218 , \26219 , \26220 ,
         \26221 , \26222 , \26223 , \26224 , \26225 , \26226 , \26227 , \26228 , \26229 , \26230 ,
         \26231 , \26232 , \26233 , \26234 , \26235 , \26236 , \26237 , \26238 , \26239 , \26240 ,
         \26241 , \26242 , \26243 , \26244 , \26245 , \26246 , \26247 , \26248 , \26249 , \26250 ,
         \26251 , \26252 , \26253 , \26254 , \26255 , \26256 , \26257 , \26258 , \26259 , \26260 ,
         \26261 , \26262 , \26263 , \26264 , \26265 , \26266 , \26267 , \26268 , \26269 , \26270 ,
         \26271 , \26272 , \26273 , \26274 , \26275 , \26276 , \26277 , \26278 , \26279 , \26280 ,
         \26281 , \26282 , \26283 , \26284 , \26285 , \26286 , \26287 , \26288 , \26289 , \26290 ,
         \26291 , \26292 , \26293 , \26294 , \26295 , \26296 , \26297 , \26298 , \26299 , \26300 ,
         \26301 , \26302 , \26303 , \26304 , \26305 , \26306 , \26307 , \26308 , \26309 , \26310 ,
         \26311 , \26312 , \26313 , \26314 , \26315 , \26316 , \26317 , \26318 , \26319 , \26320 ,
         \26321 , \26322 , \26323 , \26324 , \26325 , \26326 , \26327 , \26328 , \26329 , \26330 ,
         \26331 , \26332 , \26333 , \26334 , \26335 , \26336 , \26337 , \26338 , \26339 , \26340 ,
         \26341 , \26342 , \26343 , \26344 , \26345 , \26346 , \26347 , \26348 , \26349 , \26350 ,
         \26351 , \26352 , \26353 , \26354 , \26355 , \26356 , \26357 , \26358 , \26359 , \26360 ,
         \26361 , \26362 , \26363 , \26364 , \26365 , \26366 , \26367 , \26368 , \26369 , \26370 ,
         \26371 , \26372 , \26373 , \26374 , \26375 , \26376 , \26377 , \26378 , \26379 , \26380 ,
         \26381 , \26382 , \26383 , \26384 , \26385 , \26386 , \26387 , \26388 , \26389 , \26390 ,
         \26391 , \26392 , \26393 , \26394 , \26395 , \26396 , \26397 , \26398 , \26399 , \26400 ,
         \26401 , \26402 , \26403 , \26404 , \26405 , \26406 , \26407 , \26408 , \26409 , \26410 ,
         \26411 , \26412 , \26413 , \26414 , \26415 , \26416 , \26417 , \26418 , \26419 , \26420 ,
         \26421 , \26422 , \26423 , \26424 , \26425 , \26426 , \26427 , \26428 , \26429 , \26430 ,
         \26431 , \26432 , \26433 , \26434 , \26435 , \26436 , \26437 , \26438 , \26439 , \26440 ,
         \26441 , \26442 , \26443 , \26444 , \26445 , \26446 , \26447 , \26448 , \26449 , \26450 ,
         \26451 , \26452 , \26453 , \26454 , \26455 , \26456 , \26457 , \26458 , \26459 , \26460 ,
         \26461 , \26462 , \26463 , \26464 , \26465 , \26466 , \26467 , \26468 , \26469 , \26470 ,
         \26471 , \26472 , \26473 , \26474 , \26475 , \26476 , \26477 , \26478 , \26479 , \26480 ,
         \26481 , \26482 , \26483 , \26484 , \26485 , \26486 , \26487 , \26488 , \26489 , \26490 ,
         \26491 , \26492 , \26493 , \26494 , \26495 , \26496 , \26497 , \26498 , \26499 , \26500 ,
         \26501 , \26502 , \26503 , \26504 , \26505 , \26506 , \26507 , \26508 , \26509 , \26510 ,
         \26511 , \26512 , \26513 , \26514 , \26515 , \26516 , \26517 , \26518 , \26519 , \26520 ,
         \26521 , \26522 , \26523 , \26524 , \26525 , \26526 , \26527 , \26528 , \26529 , \26530 ,
         \26531 , \26532 , \26533 , \26534 , \26535 , \26536 , \26537 , \26538 , \26539 , \26540 ,
         \26541 , \26542 , \26543 , \26544 , \26545 , \26546 , \26547 , \26548 , \26549 , \26550 ,
         \26551 , \26552 , \26553 , \26554 , \26555 , \26556 , \26557 , \26558 , \26559 , \26560 ,
         \26561 , \26562 , \26563 , \26564 , \26565 , \26566 , \26567 , \26568 , \26569 , \26570 ,
         \26571 , \26572 , \26573 , \26574 , \26575 , \26576 , \26577 , \26578 , \26579 , \26580 ,
         \26581 , \26582 , \26583 , \26584 , \26585 , \26586 , \26587 , \26588 , \26589 , \26590 ,
         \26591 , \26592 , \26593 , \26594 , \26595 , \26596 , \26597 , \26598 , \26599 , \26600 ,
         \26601 , \26602 , \26603 , \26604 , \26605 , \26606 , \26607 , \26608 , \26609 , \26610 ,
         \26611 , \26612 , \26613 , \26614 , \26615 , \26616 , \26617 , \26618 , \26619 , \26620 ,
         \26621 , \26622 , \26623 , \26624 , \26625 , \26626 , \26627 , \26628 , \26629 , \26630 ,
         \26631 , \26632 , \26633 , \26634 , \26635 , \26636 , \26637 , \26638 , \26639 , \26640 ,
         \26641 , \26642 , \26643 , \26644 , \26645 , \26646 , \26647 , \26648 , \26649 , \26650 ,
         \26651 , \26652 , \26653 , \26654 , \26655 , \26656 , \26657 , \26658 , \26659 , \26660 ,
         \26661 , \26662 , \26663 , \26664 , \26665 , \26666 , \26667 , \26668 , \26669 , \26670 ,
         \26671 , \26672 , \26673 , \26674 , \26675 , \26676 , \26677 , \26678 , \26679 , \26680 ,
         \26681 , \26682 , \26683 , \26684 , \26685 , \26686 , \26687 , \26688 , \26689 , \26690 ,
         \26691 , \26692 , \26693 , \26694 , \26695 , \26696 , \26697 , \26698 , \26699 , \26700 ,
         \26701 , \26702 , \26703 , \26704 , \26705 , \26706 , \26707 , \26708 , \26709 , \26710 ,
         \26711 , \26712 , \26713 , \26714 , \26715 , \26716 , \26717 , \26718 , \26719 , \26720 ,
         \26721 , \26722 , \26723 , \26724 , \26725 , \26726 , \26727 , \26728 , \26729 , \26730 ,
         \26731 , \26732 , \26733 , \26734 , \26735 , \26736 , \26737 , \26738 , \26739 , \26740 ,
         \26741 , \26742 , \26743 , \26744 , \26745 , \26746 , \26747 , \26748 , \26749 , \26750 ,
         \26751 , \26752 , \26753 , \26754 , \26755 , \26756 , \26757 , \26758 , \26759 , \26760 ,
         \26761 , \26762 , \26763 , \26764 , \26765 , \26766 , \26767 , \26768 , \26769 , \26770 ,
         \26771 , \26772 , \26773 , \26774 , \26775 , \26776 , \26777 , \26778 , \26779 , \26780 ,
         \26781 , \26782 , \26783 , \26784 , \26785 , \26786 , \26787 , \26788 , \26789 , \26790 ,
         \26791 , \26792 , \26793 , \26794 , \26795 , \26796 , \26797 , \26798 , \26799 , \26800 ,
         \26801 , \26802 , \26803 , \26804 , \26805 , \26806 , \26807 , \26808 , \26809 , \26810 ,
         \26811 , \26812 , \26813 , \26814 , \26815 , \26816 , \26817 , \26818 , \26819 , \26820 ,
         \26821 , \26822 , \26823 , \26824 , \26825 , \26826 , \26827 , \26828 , \26829 , \26830 ,
         \26831 , \26832 , \26833 , \26834 , \26835 , \26836 , \26837 , \26838 , \26839 , \26840 ,
         \26841 , \26842 , \26843 , \26844 , \26845 , \26846 , \26847 , \26848 , \26849 , \26850 ,
         \26851 , \26852 , \26853 , \26854 , \26855 , \26856 , \26857 , \26858 , \26859 , \26860 ,
         \26861 , \26862 , \26863 , \26864 , \26865 , \26866 , \26867 , \26868 , \26869 , \26870 ,
         \26871 , \26872 , \26873 , \26874 , \26875 , \26876 , \26877 , \26878 , \26879 , \26880 ,
         \26881 , \26882 , \26883 , \26884 , \26885 , \26886 , \26887 , \26888 , \26889 , \26890 ,
         \26891 , \26892 , \26893 , \26894 , \26895 , \26896 , \26897 , \26898 , \26899 , \26900 ,
         \26901 , \26902 , \26903 , \26904 , \26905 , \26906 , \26907 , \26908 , \26909 , \26910 ,
         \26911 , \26912 , \26913 , \26914 , \26915 , \26916 , \26917 , \26918 , \26919 , \26920 ,
         \26921 , \26922 , \26923 , \26924 , \26925 , \26926 , \26927 , \26928 , \26929 , \26930 ,
         \26931 , \26932 , \26933 , \26934 , \26935 , \26936 , \26937 , \26938 , \26939 , \26940 ,
         \26941 , \26942 , \26943 , \26944 , \26945 , \26946 , \26947 , \26948 , \26949 , \26950 ,
         \26951 , \26952 , \26953 , \26954 , \26955 , \26956 , \26957 , \26958 , \26959 , \26960 ,
         \26961 , \26962 , \26963 , \26964 , \26965 , \26966 , \26967 , \26968 , \26969 , \26970 ,
         \26971 , \26972 , \26973 , \26974 , \26975 , \26976 , \26977 , \26978 , \26979 , \26980 ,
         \26981 , \26982 , \26983 , \26984 , \26985 , \26986 , \26987 , \26988 , \26989 , \26990 ,
         \26991 , \26992 , \26993 , \26994 , \26995 , \26996 , \26997 , \26998 , \26999 , \27000 ,
         \27001 , \27002 , \27003 , \27004 , \27005 , \27006 , \27007 , \27008 , \27009 , \27010 ,
         \27011 , \27012 , \27013 , \27014 , \27015 , \27016 , \27017 , \27018 , \27019 , \27020 ,
         \27021 , \27022 , \27023 , \27024 , \27025 , \27026 , \27027 , \27028 , \27029 , \27030 ,
         \27031 , \27032 , \27033 , \27034 , \27035 , \27036 , \27037 , \27038 , \27039 , \27040 ,
         \27041 , \27042 , \27043 , \27044 , \27045 , \27046 , \27047 , \27048 , \27049 , \27050 ,
         \27051 , \27052 , \27053 , \27054 , \27055 , \27056 , \27057 , \27058 , \27059 , \27060 ,
         \27061 , \27062 , \27063 , \27064 , \27065 , \27066 , \27067 , \27068 , \27069 , \27070 ,
         \27071 , \27072 , \27073 , \27074 , \27075 , \27076 , \27077 , \27078 , \27079 , \27080 ,
         \27081 , \27082 , \27083 , \27084 , \27085 , \27086 , \27087 , \27088 , \27089 , \27090 ,
         \27091 , \27092 , \27093 , \27094 , \27095 , \27096 , \27097 , \27098 , \27099 , \27100 ,
         \27101 , \27102 , \27103 , \27104 , \27105 , \27106 , \27107 , \27108 , \27109 , \27110 ,
         \27111 , \27112 , \27113 , \27114 , \27115 , \27116 , \27117 , \27118 , \27119 , \27120 ,
         \27121 , \27122 , \27123 , \27124 , \27125 , \27126 , \27127 , \27128 , \27129 , \27130 ,
         \27131 , \27132 , \27133 , \27134 , \27135 , \27136 , \27137 , \27138 , \27139 , \27140 ,
         \27141 , \27142 , \27143 , \27144 , \27145 , \27146 , \27147 , \27148 , \27149 , \27150 ,
         \27151 , \27152 , \27153 , \27154 , \27155 , \27156 , \27157 , \27158 , \27159 , \27160 ,
         \27161 , \27162 , \27163 , \27164 , \27165 , \27166 , \27167 , \27168 , \27169 , \27170 ,
         \27171 , \27172 , \27173 , \27174 , \27175 , \27176 , \27177 , \27178 , \27179 , \27180 ,
         \27181 , \27182 , \27183 , \27184 , \27185 , \27186 , \27187 , \27188 , \27189 , \27190 ,
         \27191 , \27192 , \27193 , \27194 , \27195 , \27196 , \27197 , \27198 , \27199 , \27200 ,
         \27201 , \27202 , \27203 , \27204 , \27205 , \27206 , \27207 , \27208 , \27209 , \27210 ,
         \27211 , \27212 , \27213 , \27214 , \27215 , \27216 , \27217 , \27218 , \27219 , \27220 ,
         \27221 , \27222 , \27223 , \27224 , \27225 , \27226 , \27227 , \27228 , \27229 , \27230 ,
         \27231 , \27232 , \27233 , \27234 , \27235 , \27236 , \27237 , \27238 , \27239 , \27240 ,
         \27241 , \27242 , \27243 , \27244 , \27245 , \27246 , \27247 , \27248 , \27249 , \27250 ,
         \27251 , \27252 , \27253 , \27254 , \27255 , \27256 , \27257 , \27258 , \27259 , \27260 ,
         \27261 , \27262 , \27263 , \27264 , \27265 , \27266 , \27267 , \27268 , \27269 , \27270 ,
         \27271 , \27272 , \27273 , \27274 , \27275 , \27276 , \27277 , \27278 , \27279 , \27280 ,
         \27281 , \27282 , \27283 , \27284 , \27285 , \27286 , \27287 , \27288 , \27289 , \27290 ,
         \27291 , \27292 , \27293 , \27294 , \27295 , \27296 , \27297 , \27298 , \27299 , \27300 ,
         \27301 , \27302 , \27303 , \27304 , \27305 , \27306 , \27307 , \27308 , \27309 , \27310 ,
         \27311 , \27312 , \27313 , \27314 , \27315 , \27316 , \27317 , \27318 , \27319 , \27320 ,
         \27321 , \27322 , \27323 , \27324 , \27325 , \27326 , \27327 , \27328 , \27329 , \27330 ,
         \27331 , \27332 , \27333 , \27334 , \27335 , \27336 , \27337 , \27338 , \27339 , \27340 ,
         \27341 , \27342 , \27343 , \27344 , \27345 , \27346 , \27347 , \27348 , \27349 , \27350 ,
         \27351 , \27352 , \27353 , \27354 , \27355 , \27356 , \27357 , \27358 , \27359 , \27360 ,
         \27361 , \27362 , \27363 , \27364 , \27365 , \27366 , \27367 , \27368 , \27369 , \27370 ,
         \27371 , \27372 , \27373 , \27374 , \27375 , \27376 , \27377 , \27378 , \27379 , \27380 ,
         \27381 , \27382 , \27383 , \27384 , \27385 , \27386 , \27387 , \27388 , \27389 , \27390 ,
         \27391 , \27392 , \27393 , \27394 , \27395 , \27396 , \27397 , \27398 , \27399 , \27400 ,
         \27401 , \27402 , \27403 , \27404 , \27405 , \27406 , \27407 , \27408 , \27409 , \27410 ,
         \27411 , \27412 , \27413 , \27414 , \27415 , \27416 , \27417 , \27418 , \27419 , \27420 ,
         \27421 , \27422 , \27423 , \27424 , \27425 , \27426 , \27427 , \27428 , \27429 , \27430 ,
         \27431 , \27432 , \27433 , \27434 , \27435 , \27436 , \27437 , \27438 , \27439 , \27440 ,
         \27441 , \27442 , \27443 , \27444 , \27445 , \27446 , \27447 , \27448 , \27449 , \27450 ,
         \27451 , \27452 , \27453 , \27454 , \27455 , \27456 , \27457 , \27458 , \27459 , \27460 ,
         \27461 , \27462 , \27463 , \27464 , \27465 , \27466 , \27467 , \27468 , \27469 , \27470 ,
         \27471 , \27472 , \27473 , \27474 , \27475 , \27476 , \27477 , \27478 , \27479 , \27480 ,
         \27481 , \27482 , \27483 , \27484 , \27485 , \27486 , \27487 , \27488 , \27489 , \27490 ,
         \27491 , \27492 , \27493 , \27494 , \27495 , \27496 , \27497 , \27498 , \27499 , \27500 ,
         \27501 , \27502 , \27503 , \27504 , \27505 , \27506 , \27507 , \27508 , \27509 , \27510 ,
         \27511 , \27512 , \27513 , \27514 , \27515 , \27516 , \27517 , \27518 , \27519 , \27520 ,
         \27521 , \27522 , \27523 , \27524 , \27525 , \27526 , \27527 , \27528 , \27529 , \27530 ,
         \27531 , \27532 , \27533 , \27534 , \27535 , \27536 , \27537 , \27538 , \27539 , \27540 ,
         \27541 , \27542 , \27543 , \27544 , \27545 , \27546 , \27547 , \27548 , \27549 , \27550 ,
         \27551 , \27552 , \27553 , \27554 , \27555 , \27556 , \27557 , \27558 , \27559 , \27560 ,
         \27561 , \27562 , \27563 , \27564 , \27565 , \27566 , \27567 , \27568 , \27569 , \27570 ,
         \27571 , \27572 , \27573 , \27574 , \27575 , \27576 , \27577 , \27578 , \27579 , \27580 ,
         \27581 , \27582 , \27583 , \27584 , \27585 , \27586 , \27587 , \27588 , \27589 , \27590 ,
         \27591 , \27592 , \27593 , \27594 , \27595 , \27596 , \27597 , \27598 , \27599 , \27600 ,
         \27601 , \27602 , \27603 , \27604 , \27605 , \27606 , \27607 , \27608 , \27609 , \27610 ,
         \27611 , \27612 , \27613 , \27614 , \27615 , \27616 , \27617 , \27618 , \27619 , \27620 ,
         \27621 , \27622 , \27623 , \27624 , \27625 , \27626 , \27627 , \27628 , \27629 , \27630 ,
         \27631 , \27632 , \27633 , \27634 , \27635 , \27636 , \27637 , \27638 , \27639 , \27640 ,
         \27641 , \27642 , \27643 , \27644 , \27645 , \27646 , \27647 , \27648 , \27649 , \27650 ,
         \27651 , \27652 , \27653 , \27654 , \27655 , \27656 , \27657 , \27658 , \27659 , \27660 ,
         \27661 , \27662 , \27663 , \27664 , \27665 , \27666 , \27667 , \27668 , \27669 , \27670 ,
         \27671 , \27672 , \27673 , \27674 , \27675 , \27676 , \27677 , \27678 , \27679 , \27680 ,
         \27681 , \27682 , \27683 , \27684 , \27685 , \27686 , \27687 , \27688 , \27689 , \27690 ,
         \27691 , \27692 , \27693 , \27694 , \27695 , \27696 , \27697 , \27698 , \27699 , \27700 ,
         \27701 , \27702 , \27703 , \27704 , \27705 , \27706 , \27707 , \27708 , \27709 , \27710 ,
         \27711 , \27712 , \27713 , \27714 , \27715 , \27716 , \27717 , \27718 , \27719 , \27720 ,
         \27721 , \27722 , \27723 , \27724 , \27725 , \27726 , \27727 , \27728 , \27729 , \27730 ,
         \27731 , \27732 , \27733 , \27734 , \27735 , \27736 , \27737 , \27738 , \27739 , \27740 ,
         \27741 , \27742 , \27743 , \27744 , \27745 , \27746 , \27747 , \27748 , \27749 , \27750 ,
         \27751 , \27752 , \27753 , \27754 , \27755 , \27756 , \27757 , \27758 , \27759 , \27760 ,
         \27761 , \27762 , \27763 , \27764 , \27765 , \27766 , \27767 , \27768 , \27769 , \27770 ,
         \27771 , \27772 , \27773 , \27774 , \27775 , \27776 , \27777 , \27778 , \27779 , \27780 ,
         \27781 , \27782 , \27783 , \27784 , \27785 , \27786 , \27787 , \27788 , \27789 , \27790 ,
         \27791 , \27792 , \27793 , \27794 , \27795 , \27796 , \27797 , \27798 , \27799 , \27800 ,
         \27801 , \27802 , \27803 , \27804 , \27805 , \27806 , \27807 , \27808 , \27809 , \27810 ,
         \27811 , \27812 , \27813 , \27814 , \27815 , \27816 , \27817 , \27818 , \27819 , \27820 ,
         \27821 , \27822 , \27823 , \27824 , \27825 , \27826 , \27827 , \27828 , \27829 , \27830 ,
         \27831 , \27832 , \27833 , \27834 , \27835 , \27836 , \27837 , \27838 , \27839 , \27840 ,
         \27841 , \27842 , \27843 , \27844 , \27845 , \27846 , \27847 , \27848 , \27849 , \27850 ,
         \27851 , \27852 , \27853 , \27854 , \27855 , \27856 , \27857 , \27858 , \27859 , \27860 ,
         \27861 , \27862 , \27863 , \27864 , \27865 , \27866 , \27867 , \27868 , \27869 , \27870 ,
         \27871 , \27872 , \27873 , \27874 , \27875 , \27876 , \27877 , \27878 , \27879 , \27880 ,
         \27881 , \27882 , \27883 , \27884 , \27885 , \27886 , \27887 , \27888 , \27889 , \27890 ,
         \27891 , \27892 , \27893 , \27894 , \27895 , \27896 , \27897 , \27898 , \27899 , \27900 ,
         \27901 , \27902 , \27903 , \27904 , \27905 , \27906 , \27907 , \27908 , \27909 , \27910 ,
         \27911 , \27912 , \27913 , \27914 , \27915 , \27916 , \27917 , \27918 , \27919 , \27920 ,
         \27921 , \27922 , \27923 , \27924 , \27925 , \27926 , \27927 , \27928 , \27929 , \27930 ,
         \27931 , \27932 , \27933 , \27934 , \27935 , \27936 , \27937 , \27938 , \27939 , \27940 ,
         \27941 , \27942 , \27943 , \27944 , \27945 , \27946 , \27947 , \27948 , \27949 , \27950 ,
         \27951 , \27952 , \27953 , \27954 , \27955 , \27956 , \27957 , \27958 , \27959 , \27960 ,
         \27961 , \27962 , \27963 , \27964 , \27965 , \27966 , \27967 , \27968 , \27969 , \27970 ,
         \27971 , \27972 , \27973 , \27974 , \27975 , \27976 , \27977 , \27978 , \27979 , \27980 ,
         \27981 , \27982 , \27983 , \27984 , \27985 , \27986 , \27987 , \27988 , \27989 , \27990 ,
         \27991 , \27992 , \27993 , \27994 , \27995 , \27996 , \27997 , \27998 , \27999 , \28000 ,
         \28001 , \28002 , \28003 , \28004 , \28005 , \28006 , \28007 , \28008 , \28009 , \28010 ,
         \28011 , \28012 , \28013 , \28014 , \28015 , \28016 , \28017 , \28018 , \28019 , \28020 ,
         \28021 , \28022 , \28023 , \28024 , \28025 , \28026 , \28027 , \28028 , \28029 , \28030 ,
         \28031 , \28032 , \28033 , \28034 , \28035 , \28036 , \28037 , \28038 , \28039 , \28040 ,
         \28041 , \28042 , \28043 , \28044 , \28045 , \28046 , \28047 , \28048 , \28049 , \28050 ,
         \28051 , \28052 , \28053 , \28054 , \28055 , \28056 , \28057 , \28058 , \28059 , \28060 ,
         \28061 , \28062 , \28063 , \28064 , \28065 , \28066 , \28067 , \28068 , \28069 , \28070 ,
         \28071 , \28072 , \28073 , \28074 , \28075 , \28076 , \28077 , \28078 , \28079 , \28080 ,
         \28081 , \28082 , \28083 , \28084 , \28085 , \28086 , \28087 , \28088 , \28089 , \28090 ,
         \28091 , \28092 , \28093 , \28094 , \28095 , \28096 , \28097 , \28098 , \28099 , \28100 ,
         \28101 , \28102 , \28103 , \28104 , \28105 , \28106 , \28107 , \28108 , \28109 , \28110 ,
         \28111 , \28112 , \28113 , \28114 , \28115 , \28116 , \28117 , \28118 , \28119 , \28120 ,
         \28121 , \28122 , \28123 , \28124 , \28125 , \28126 , \28127 , \28128 , \28129 , \28130 ,
         \28131 , \28132 , \28133 , \28134 , \28135 , \28136 , \28137 , \28138 , \28139 , \28140 ,
         \28141 , \28142 , \28143 , \28144 , \28145 , \28146 , \28147 , \28148 , \28149 , \28150 ,
         \28151 , \28152 , \28153 , \28154 , \28155 , \28156 , \28157 , \28158 , \28159 , \28160 ,
         \28161 , \28162 , \28163 , \28164 , \28165 , \28166 , \28167 , \28168 , \28169 , \28170 ,
         \28171 , \28172 , \28173 , \28174 , \28175 , \28176 , \28177 , \28178 , \28179 , \28180 ,
         \28181 , \28182 , \28183 , \28184 , \28185 , \28186 , \28187 , \28188 , \28189 , \28190 ,
         \28191 , \28192 , \28193 , \28194 , \28195 , \28196 , \28197 , \28198 , \28199 , \28200 ,
         \28201 , \28202 , \28203 , \28204 , \28205 , \28206 , \28207 , \28208 , \28209 , \28210 ,
         \28211 , \28212 , \28213 , \28214 , \28215 , \28216 , \28217 , \28218 , \28219 , \28220 ,
         \28221 , \28222 , \28223 , \28224 , \28225 , \28226 , \28227 , \28228 , \28229 , \28230 ,
         \28231 , \28232 , \28233 , \28234 , \28235 , \28236 , \28237 , \28238 , \28239 , \28240 ,
         \28241 , \28242 , \28243 , \28244 , \28245 , \28246 , \28247 , \28248 , \28249 , \28250 ,
         \28251 , \28252 , \28253 , \28254 , \28255 , \28256 , \28257 , \28258 , \28259 , \28260 ,
         \28261 , \28262 , \28263 , \28264 , \28265 , \28266 , \28267 , \28268 , \28269 , \28270 ,
         \28271 , \28272 , \28273 , \28274 , \28275 , \28276 , \28277 , \28278 , \28279 , \28280 ,
         \28281 , \28282 , \28283 , \28284 , \28285 , \28286 , \28287 , \28288 , \28289 , \28290 ,
         \28291 , \28292 , \28293 , \28294 , \28295 , \28296 , \28297 , \28298 , \28299 , \28300 ,
         \28301 , \28302 , \28303 , \28304 , \28305 , \28306 , \28307 , \28308 , \28309 , \28310 ,
         \28311 , \28312 , \28313 , \28314 , \28315 , \28316 , \28317 , \28318 , \28319 , \28320 ,
         \28321 , \28322 , \28323 , \28324 , \28325 , \28326 , \28327 , \28328 , \28329 , \28330 ,
         \28331 , \28332 , \28333 , \28334 , \28335 , \28336 , \28337 , \28338 , \28339 , \28340 ,
         \28341 , \28342 , \28343 , \28344 , \28345 , \28346 , \28347 , \28348 , \28349 , \28350 ,
         \28351 , \28352 , \28353 , \28354 , \28355 , \28356 , \28357 , \28358 , \28359 , \28360 ,
         \28361 , \28362 , \28363 , \28364 , \28365 , \28366 , \28367 , \28368 , \28369 , \28370 ,
         \28371 , \28372 , \28373 , \28374 , \28375 , \28376 , \28377 , \28378 , \28379 , \28380 ,
         \28381 , \28382 , \28383 , \28384 , \28385 , \28386 , \28387 , \28388 , \28389 , \28390 ,
         \28391 , \28392 , \28393 , \28394 , \28395 , \28396 , \28397 , \28398 , \28399 , \28400 ,
         \28401 , \28402 , \28403 , \28404 , \28405 , \28406 , \28407 , \28408 , \28409 , \28410 ,
         \28411 , \28412 , \28413 , \28414 , \28415 , \28416 , \28417 , \28418 , \28419 , \28420 ,
         \28421 , \28422 , \28423 , \28424 , \28425 , \28426 , \28427 , \28428 , \28429 , \28430 ,
         \28431 , \28432 , \28433 , \28434 , \28435 , \28436 , \28437 , \28438 , \28439 , \28440 ,
         \28441 , \28442 , \28443 , \28444 , \28445 , \28446 , \28447 , \28448 , \28449 , \28450 ,
         \28451 , \28452 , \28453 , \28454 , \28455 , \28456 , \28457 , \28458 , \28459 , \28460 ,
         \28461 , \28462 , \28463 , \28464 , \28465 , \28466 , \28467 , \28468 , \28469 , \28470 ,
         \28471 , \28472 , \28473 , \28474 , \28475 , \28476 , \28477 , \28478 , \28479 , \28480 ,
         \28481 , \28482 , \28483 , \28484 , \28485 , \28486 , \28487 , \28488 , \28489 , \28490 ,
         \28491 , \28492 , \28493 , \28494 , \28495 , \28496 , \28497 , \28498 , \28499 , \28500 ,
         \28501 , \28502 , \28503 , \28504 , \28505 , \28506 , \28507 , \28508 , \28509 , \28510 ,
         \28511 , \28512 , \28513 , \28514 , \28515 , \28516 , \28517 , \28518 , \28519 , \28520 ,
         \28521 , \28522 , \28523 , \28524 , \28525 , \28526 , \28527 , \28528 , \28529 , \28530 ,
         \28531 , \28532 , \28533 , \28534 , \28535 , \28536 , \28537 , \28538 , \28539 , \28540 ,
         \28541 , \28542 , \28543 , \28544 , \28545 , \28546 , \28547 , \28548 , \28549 , \28550 ,
         \28551 , \28552 , \28553 , \28554 , \28555 , \28556 , \28557 , \28558 , \28559 , \28560 ,
         \28561 , \28562 , \28563 , \28564 , \28565 , \28566 , \28567 , \28568 , \28569 , \28570 ,
         \28571 , \28572 , \28573 , \28574 , \28575 , \28576 , \28577 , \28578 , \28579 , \28580 ,
         \28581 , \28582 , \28583 , \28584 , \28585 , \28586 , \28587 , \28588 , \28589 , \28590 ,
         \28591 , \28592 , \28593 , \28594 , \28595 , \28596 , \28597 , \28598 , \28599 , \28600 ,
         \28601 , \28602 , \28603 , \28604 , \28605 , \28606 , \28607 , \28608 , \28609 , \28610 ,
         \28611 , \28612 , \28613 , \28614 , \28615 , \28616 , \28617 , \28618 , \28619 , \28620 ,
         \28621 , \28622 , \28623 , \28624 , \28625 , \28626 , \28627 , \28628 , \28629 , \28630 ,
         \28631 , \28632 , \28633 , \28634 , \28635 , \28636 , \28637 , \28638 , \28639 , \28640 ,
         \28641 , \28642 , \28643 , \28644 , \28645 , \28646 , \28647 , \28648 , \28649 , \28650 ,
         \28651 , \28652 , \28653 , \28654 , \28655 , \28656 , \28657 , \28658 , \28659 , \28660 ,
         \28661 , \28662 , \28663 , \28664 , \28665 , \28666 , \28667 , \28668 , \28669 , \28670 ,
         \28671 , \28672 , \28673 , \28674 , \28675 , \28676 , \28677 , \28678 , \28679 , \28680 ,
         \28681 , \28682 , \28683 , \28684 , \28685 , \28686 , \28687 , \28688 , \28689 , \28690 ,
         \28691 , \28692 , \28693 , \28694 , \28695 , \28696 , \28697 , \28698 , \28699 , \28700 ,
         \28701 , \28702 , \28703 , \28704 , \28705 , \28706 , \28707 , \28708 , \28709 , \28710 ,
         \28711 , \28712 , \28713 , \28714 , \28715 , \28716 , \28717 , \28718 , \28719 , \28720 ,
         \28721 , \28722 , \28723 , \28724 , \28725 , \28726 , \28727 , \28728 , \28729 , \28730 ,
         \28731 , \28732 , \28733 , \28734 , \28735 , \28736 , \28737 , \28738 , \28739 , \28740 ,
         \28741 , \28742 , \28743 , \28744 , \28745 , \28746 , \28747 , \28748 , \28749 , \28750 ,
         \28751 , \28752 , \28753 , \28754 , \28755 , \28756 , \28757 , \28758 , \28759 , \28760 ,
         \28761 , \28762 , \28763 , \28764 , \28765 , \28766 , \28767 , \28768 , \28769 , \28770 ,
         \28771 , \28772 , \28773 , \28774 , \28775 , \28776 , \28777 , \28778 , \28779 , \28780 ,
         \28781 , \28782 , \28783 , \28784 , \28785 , \28786 , \28787 , \28788 , \28789 , \28790 ,
         \28791 , \28792 , \28793 , \28794 , \28795 , \28796 , \28797 , \28798 , \28799 , \28800 ,
         \28801 , \28802 , \28803 , \28804 , \28805 , \28806 , \28807 , \28808 , \28809 , \28810 ,
         \28811 , \28812 , \28813 , \28814 , \28815 , \28816 , \28817 , \28818 , \28819 , \28820 ,
         \28821 , \28822 , \28823 , \28824 , \28825 , \28826 , \28827 , \28828 , \28829 , \28830 ,
         \28831 , \28832 , \28833 , \28834 , \28835 , \28836 , \28837 , \28838 , \28839 , \28840 ,
         \28841 , \28842 , \28843 , \28844 , \28845 , \28846 , \28847 , \28848 , \28849 , \28850 ,
         \28851 , \28852 , \28853 , \28854 , \28855 , \28856 , \28857 , \28858 , \28859 , \28860 ,
         \28861 , \28862 , \28863 , \28864 , \28865 , \28866 , \28867 , \28868 , \28869 , \28870 ,
         \28871 , \28872 , \28873 , \28874 , \28875 , \28876 , \28877 , \28878 , \28879 , \28880 ,
         \28881 , \28882 , \28883 , \28884 , \28885 , \28886 , \28887 , \28888 , \28889 , \28890 ,
         \28891 , \28892 , \28893 , \28894 , \28895 , \28896 , \28897 , \28898 , \28899 , \28900 ,
         \28901 , \28902 , \28903 , \28904 , \28905 , \28906 , \28907 , \28908 , \28909 , \28910 ,
         \28911 , \28912 , \28913 , \28914 , \28915 , \28916 , \28917 , \28918 , \28919 , \28920 ,
         \28921 , \28922 , \28923 , \28924 , \28925 , \28926 , \28927 , \28928 , \28929 , \28930 ,
         \28931 , \28932 , \28933 , \28934 , \28935 , \28936 , \28937 , \28938 , \28939 , \28940 ,
         \28941 , \28942 , \28943 , \28944 , \28945 , \28946 , \28947 , \28948 , \28949 , \28950 ,
         \28951 , \28952 , \28953 , \28954 , \28955 , \28956 , \28957 , \28958 , \28959 , \28960 ,
         \28961 , \28962 , \28963 , \28964 , \28965 , \28966 , \28967 , \28968 , \28969 , \28970 ,
         \28971 , \28972 , \28973 , \28974 , \28975 , \28976 , \28977 , \28978 , \28979 , \28980 ,
         \28981 , \28982 , \28983 , \28984 , \28985 , \28986 , \28987 , \28988 , \28989 , \28990 ,
         \28991 , \28992 , \28993 , \28994 , \28995 , \28996 , \28997 , \28998 , \28999 , \29000 ,
         \29001 , \29002 , \29003 , \29004 , \29005 , \29006 , \29007 , \29008 , \29009 , \29010 ,
         \29011 , \29012 , \29013 , \29014 , \29015 , \29016 , \29017 , \29018 , \29019 , \29020 ,
         \29021 , \29022 , \29023 , \29024 , \29025 , \29026 , \29027 , \29028 , \29029 , \29030 ,
         \29031 , \29032 , \29033 , \29034 , \29035 , \29036 , \29037 , \29038 , \29039 , \29040 ,
         \29041 , \29042 , \29043 , \29044 , \29045 , \29046 , \29047 , \29048 , \29049 , \29050 ,
         \29051 , \29052 , \29053 , \29054 , \29055 , \29056 , \29057 , \29058 , \29059 , \29060 ,
         \29061 , \29062 , \29063 , \29064 , \29065 , \29066 , \29067 , \29068 , \29069 , \29070 ,
         \29071 , \29072 , \29073 , \29074 , \29075 , \29076 , \29077 , \29078 , \29079 , \29080 ,
         \29081 , \29082 , \29083 , \29084 , \29085 , \29086 , \29087 , \29088 , \29089 , \29090 ,
         \29091 , \29092 , \29093 , \29094 , \29095 , \29096 , \29097 , \29098 , \29099 , \29100 ,
         \29101 , \29102 , \29103 , \29104 , \29105 , \29106 , \29107 , \29108 , \29109 , \29110 ,
         \29111 , \29112 , \29113 , \29114 , \29115 , \29116 , \29117 , \29118 , \29119 , \29120 ,
         \29121 , \29122 , \29123 , \29124 , \29125 , \29126 , \29127 , \29128 , \29129 , \29130 ,
         \29131 , \29132 , \29133 , \29134 , \29135 , \29136 , \29137 , \29138 , \29139 , \29140 ,
         \29141 , \29142 , \29143 , \29144 , \29145 , \29146 , \29147 , \29148 , \29149 , \29150 ,
         \29151 , \29152 , \29153 , \29154 , \29155 , \29156 , \29157 , \29158 , \29159 , \29160 ,
         \29161 , \29162 , \29163 , \29164 , \29165 , \29166 , \29167 , \29168 , \29169 , \29170 ,
         \29171 , \29172 , \29173 , \29174 , \29175 , \29176 , \29177 , \29178 , \29179 , \29180 ,
         \29181 , \29182 , \29183 , \29184 , \29185 , \29186 , \29187 , \29188 , \29189 , \29190 ,
         \29191 , \29192 , \29193 , \29194 , \29195 , \29196 , \29197 , \29198 , \29199 , \29200 ,
         \29201 , \29202 , \29203 , \29204 , \29205 , \29206 , \29207 , \29208 , \29209 , \29210 ,
         \29211 , \29212 , \29213 , \29214 , \29215 , \29216 , \29217 , \29218 , \29219 , \29220 ,
         \29221 , \29222 , \29223 , \29224 , \29225 , \29226 , \29227 , \29228 , \29229 , \29230 ,
         \29231 , \29232 , \29233 , \29234 , \29235 , \29236 , \29237 , \29238 , \29239 , \29240 ,
         \29241 , \29242 , \29243 , \29244 , \29245 , \29246 , \29247 , \29248 , \29249 , \29250 ,
         \29251 , \29252 , \29253 , \29254 , \29255 , \29256 , \29257 , \29258 , \29259 , \29260 ,
         \29261 , \29262 , \29263 , \29264 , \29265 , \29266 , \29267 , \29268 , \29269 , \29270 ,
         \29271 , \29272 , \29273 , \29274 , \29275 , \29276 , \29277 , \29278 , \29279 , \29280 ,
         \29281 , \29282 , \29283 , \29284 , \29285 , \29286 , \29287 , \29288 , \29289 , \29290 ,
         \29291 , \29292 , \29293 , \29294 , \29295 , \29296 , \29297 , \29298 , \29299 , \29300 ,
         \29301 , \29302 , \29303 , \29304 , \29305 , \29306 , \29307 , \29308 , \29309 , \29310 ,
         \29311 , \29312 , \29313 , \29314 , \29315 , \29316 , \29317 , \29318 , \29319 , \29320 ,
         \29321 , \29322 , \29323 , \29324 , \29325 , \29326 , \29327 , \29328 , \29329 , \29330 ,
         \29331 , \29332 , \29333 , \29334 , \29335 , \29336 , \29337 , \29338 , \29339 , \29340 ,
         \29341 , \29342 , \29343 , \29344 , \29345 , \29346 , \29347 , \29348 , \29349 , \29350 ,
         \29351 , \29352 , \29353 , \29354 , \29355 , \29356 , \29357 , \29358 , \29359 , \29360 ,
         \29361 , \29362 , \29363 , \29364 , \29365 , \29366 , \29367 , \29368 , \29369 , \29370 ,
         \29371 , \29372 , \29373 , \29374 , \29375 , \29376 , \29377 , \29378 , \29379 , \29380 ,
         \29381 , \29382 , \29383 , \29384 , \29385 , \29386 , \29387 , \29388 , \29389 , \29390 ,
         \29391 , \29392 , \29393 , \29394 , \29395 , \29396 , \29397 , \29398 , \29399 , \29400 ,
         \29401 , \29402 , \29403 , \29404 , \29405 , \29406 , \29407 , \29408 , \29409 , \29410 ,
         \29411 , \29412 , \29413 , \29414 , \29415 , \29416 , \29417 , \29418 , \29419 , \29420 ,
         \29421 , \29422 , \29423 , \29424 , \29425 , \29426 , \29427 , \29428 , \29429 , \29430 ,
         \29431 , \29432 , \29433 , \29434 , \29435 , \29436 , \29437 , \29438 , \29439 , \29440 ,
         \29441 , \29442 , \29443 , \29444 , \29445 , \29446 , \29447 , \29448 , \29449 , \29450 ,
         \29451 , \29452 , \29453 , \29454 , \29455 , \29456 , \29457 , \29458 , \29459 , \29460 ,
         \29461 , \29462 , \29463 , \29464 , \29465 , \29466 , \29467 , \29468 , \29469 , \29470 ,
         \29471 , \29472 , \29473 , \29474 , \29475 , \29476 , \29477 , \29478 , \29479 , \29480 ,
         \29481 , \29482 , \29483 , \29484 , \29485 , \29486 , \29487 , \29488 , \29489 , \29490 ,
         \29491 , \29492 , \29493 , \29494 , \29495 , \29496 , \29497 , \29498 , \29499 , \29500 ,
         \29501 , \29502 , \29503 , \29504 , \29505 , \29506 , \29507 , \29508 , \29509 , \29510 ,
         \29511 , \29512 , \29513 , \29514 , \29515 , \29516 , \29517 , \29518 , \29519 , \29520 ,
         \29521 , \29522 , \29523 , \29524 , \29525 , \29526 , \29527 , \29528 , \29529 , \29530 ,
         \29531 , \29532 , \29533 , \29534 , \29535 , \29536 , \29537 , \29538 , \29539 , \29540 ,
         \29541 , \29542 , \29543 , \29544 , \29545 , \29546 , \29547 , \29548 , \29549 , \29550 ,
         \29551 , \29552 , \29553 , \29554 , \29555 , \29556 , \29557 , \29558 , \29559 , \29560 ,
         \29561 , \29562 , \29563 , \29564 , \29565 , \29566 , \29567 , \29568 , \29569 , \29570 ,
         \29571 , \29572 , \29573 , \29574 , \29575 , \29576 , \29577 , \29578 , \29579 , \29580 ,
         \29581 , \29582 , \29583 , \29584 , \29585 , \29586 , \29587 , \29588 , \29589 , \29590 ,
         \29591 , \29592 , \29593 , \29594 , \29595 , \29596 , \29597 , \29598 , \29599 , \29600 ,
         \29601 , \29602 , \29603 , \29604 , \29605 , \29606 , \29607 , \29608 , \29609 , \29610 ,
         \29611 , \29612 , \29613 , \29614 , \29615 , \29616 , \29617 , \29618 , \29619 , \29620 ,
         \29621 , \29622 , \29623 , \29624 , \29625 , \29626 , \29627 , \29628 , \29629 , \29630 ,
         \29631 , \29632 , \29633 , \29634 , \29635 , \29636 , \29637 , \29638 , \29639 , \29640 ,
         \29641 , \29642 , \29643 , \29644 , \29645 , \29646 , \29647 , \29648 , \29649 , \29650 ,
         \29651 , \29652 , \29653 , \29654 , \29655 , \29656 , \29657 , \29658 , \29659 , \29660 ,
         \29661 , \29662 , \29663 , \29664 , \29665 , \29666 , \29667 , \29668 , \29669 , \29670 ,
         \29671 , \29672 , \29673 , \29674 , \29675 , \29676 , \29677 , \29678 , \29679 , \29680 ,
         \29681 , \29682 , \29683 , \29684 , \29685 , \29686 , \29687 , \29688 , \29689 , \29690 ,
         \29691 , \29692 , \29693 , \29694 , \29695 , \29696 , \29697 , \29698 , \29699 , \29700 ,
         \29701 , \29702 , \29703 , \29704 , \29705 , \29706 , \29707 , \29708 , \29709 , \29710 ,
         \29711 , \29712 , \29713 , \29714 , \29715 , \29716 , \29717 , \29718 , \29719 , \29720 ,
         \29721 , \29722 , \29723 , \29724 , \29725 , \29726 , \29727 , \29728 , \29729 , \29730 ,
         \29731 , \29732 , \29733 , \29734 , \29735 , \29736 , \29737 , \29738 , \29739 , \29740 ,
         \29741 , \29742 , \29743 , \29744 , \29745 , \29746 , \29747 , \29748 , \29749 , \29750 ,
         \29751 , \29752 , \29753 , \29754 , \29755 , \29756 , \29757 , \29758 , \29759 , \29760 ,
         \29761 , \29762 , \29763 , \29764 , \29765 , \29766 , \29767 , \29768 , \29769 , \29770 ,
         \29771 , \29772 , \29773 , \29774 , \29775 , \29776 , \29777 , \29778 , \29779 , \29780 ,
         \29781 , \29782 , \29783 , \29784 , \29785 , \29786 , \29787 , \29788 , \29789 , \29790 ,
         \29791 , \29792 , \29793 , \29794 , \29795 , \29796 , \29797 , \29798 , \29799 , \29800 ,
         \29801 , \29802 , \29803 , \29804 , \29805 , \29806 , \29807 , \29808 , \29809 , \29810 ,
         \29811 , \29812 , \29813 , \29814 , \29815 , \29816 , \29817 , \29818 , \29819 , \29820 ,
         \29821 , \29822 , \29823 , \29824 , \29825 , \29826 , \29827 , \29828 , \29829 , \29830 ,
         \29831 , \29832 , \29833 , \29834 , \29835 , \29836 , \29837 , \29838 , \29839 , \29840 ,
         \29841 , \29842 , \29843 , \29844 , \29845 , \29846 , \29847 , \29848 , \29849 , \29850 ,
         \29851 , \29852 , \29853 , \29854 , \29855 , \29856 , \29857 , \29858 , \29859 , \29860 ,
         \29861 , \29862 , \29863 , \29864 , \29865 , \29866 , \29867 , \29868 , \29869 , \29870 ,
         \29871 , \29872 , \29873 , \29874 , \29875 , \29876 , \29877 , \29878 , \29879 , \29880 ,
         \29881 , \29882 , \29883 , \29884 , \29885 , \29886 , \29887 , \29888 , \29889 , \29890 ,
         \29891 , \29892 , \29893 , \29894 , \29895 , \29896 , \29897 , \29898 , \29899 , \29900 ,
         \29901 , \29902 , \29903 , \29904 , \29905 , \29906 , \29907 , \29908 , \29909 , \29910 ,
         \29911 , \29912 , \29913 , \29914 , \29915 , \29916 , \29917 , \29918 , \29919 , \29920 ,
         \29921 , \29922 , \29923 , \29924 , \29925 , \29926 , \29927 , \29928 , \29929 , \29930 ,
         \29931 , \29932 , \29933 , \29934 , \29935 , \29936 , \29937 , \29938 , \29939 , \29940 ,
         \29941 , \29942 , \29943 , \29944 , \29945 , \29946 , \29947 , \29948 , \29949 , \29950 ,
         \29951 , \29952 , \29953 , \29954 , \29955 , \29956 , \29957 , \29958 , \29959 , \29960 ,
         \29961 , \29962 , \29963 , \29964 , \29965 , \29966 , \29967 , \29968 , \29969 , \29970 ,
         \29971 , \29972 , \29973 , \29974 , \29975 , \29976 , \29977 , \29978 , \29979 , \29980 ,
         \29981 , \29982 , \29983 , \29984 , \29985 , \29986 , \29987 , \29988 , \29989 , \29990 ,
         \29991 , \29992 , \29993 , \29994 , \29995 , \29996 , \29997 , \29998 , \29999 , \30000 ,
         \30001 , \30002 , \30003 , \30004 , \30005 , \30006 , \30007 , \30008 , \30009 , \30010 ,
         \30011 , \30012 , \30013 , \30014 , \30015 , \30016 , \30017 , \30018 , \30019 , \30020 ,
         \30021 , \30022 , \30023 , \30024 , \30025 , \30026 , \30027 , \30028 , \30029 , \30030 ,
         \30031 , \30032 , \30033 , \30034 , \30035 , \30036 , \30037 , \30038 , \30039 , \30040 ,
         \30041 , \30042 , \30043 , \30044 , \30045 , \30046 , \30047 , \30048 , \30049 , \30050 ,
         \30051 , \30052 , \30053 , \30054 , \30055 , \30056 , \30057 , \30058 , \30059 , \30060 ,
         \30061 , \30062 , \30063 , \30064 , \30065 , \30066 , \30067 , \30068 , \30069 , \30070 ,
         \30071 , \30072 , \30073 , \30074 , \30075 , \30076 , \30077 , \30078 , \30079 , \30080 ,
         \30081 , \30082 , \30083 , \30084 , \30085 , \30086 , \30087 , \30088 , \30089 , \30090 ,
         \30091 , \30092 , \30093 , \30094 , \30095 , \30096 , \30097 , \30098 , \30099 , \30100 ,
         \30101 , \30102 , \30103 , \30104 , \30105 , \30106 , \30107 , \30108 , \30109 , \30110 ,
         \30111 , \30112 , \30113 , \30114 , \30115 , \30116 , \30117 , \30118 , \30119 , \30120 ,
         \30121 , \30122 , \30123 , \30124 , \30125 , \30126 , \30127 , \30128 , \30129 , \30130 ,
         \30131 , \30132 , \30133 , \30134 , \30135 , \30136 , \30137 , \30138 , \30139 , \30140 ,
         \30141 , \30142 , \30143 , \30144 , \30145 , \30146 , \30147 , \30148 , \30149 , \30150 ,
         \30151 , \30152 , \30153 , \30154 , \30155 , \30156 , \30157 , \30158 , \30159 , \30160 ,
         \30161 , \30162 , \30163 , \30164 , \30165 , \30166 , \30167 , \30168 , \30169 , \30170 ,
         \30171 , \30172 , \30173 , \30174 , \30175 , \30176 , \30177 , \30178 , \30179 , \30180 ,
         \30181 , \30182 , \30183 , \30184 , \30185 , \30186 , \30187 , \30188 , \30189 , \30190 ,
         \30191 , \30192 , \30193 , \30194 , \30195 , \30196 , \30197 , \30198 , \30199 , \30200 ,
         \30201 , \30202 , \30203 , \30204 , \30205 , \30206 , \30207 , \30208 , \30209 , \30210 ,
         \30211 , \30212 , \30213 , \30214 , \30215 , \30216 , \30217 , \30218 , \30219 , \30220 ,
         \30221 , \30222 , \30223 , \30224 , \30225 , \30226 , \30227 , \30228 , \30229 , \30230 ,
         \30231 , \30232 , \30233 , \30234 , \30235 , \30236 , \30237 , \30238 , \30239 , \30240 ,
         \30241 , \30242 , \30243 , \30244 , \30245 , \30246 , \30247 , \30248 , \30249 , \30250 ,
         \30251 , \30252 , \30253 , \30254 , \30255 , \30256 , \30257 , \30258 , \30259 , \30260 ,
         \30261 , \30262 , \30263 , \30264 , \30265 , \30266 , \30267 , \30268 , \30269 , \30270 ,
         \30271 , \30272 , \30273 , \30274 , \30275 , \30276 , \30277 , \30278 , \30279 , \30280 ,
         \30281 , \30282 , \30283 , \30284 , \30285 , \30286 , \30287 , \30288 , \30289 , \30290 ,
         \30291 , \30292 , \30293 , \30294 , \30295 , \30296 , \30297 , \30298 , \30299 , \30300 ,
         \30301 , \30302 , \30303 , \30304 , \30305 , \30306 , \30307 , \30308 , \30309 , \30310 ,
         \30311 , \30312 , \30313 , \30314 , \30315 , \30316 , \30317 , \30318 , \30319 , \30320 ,
         \30321 , \30322 , \30323 , \30324 , \30325 , \30326 , \30327 , \30328 , \30329 , \30330 ,
         \30331 , \30332 , \30333 , \30334 , \30335 , \30336 , \30337 , \30338 , \30339 , \30340 ,
         \30341 , \30342 , \30343 , \30344 , \30345 , \30346 , \30347 , \30348 , \30349 , \30350 ,
         \30351 , \30352 , \30353 , \30354 , \30355 , \30356 , \30357 , \30358 , \30359 , \30360 ,
         \30361 , \30362 , \30363 , \30364 , \30365 , \30366 , \30367 , \30368 , \30369 , \30370 ,
         \30371 , \30372 , \30373 , \30374 , \30375 , \30376 , \30377 , \30378 , \30379 , \30380 ,
         \30381 , \30382 , \30383 , \30384 , \30385 , \30386 , \30387 , \30388 , \30389 , \30390 ,
         \30391 , \30392 , \30393 , \30394 , \30395 , \30396 , \30397 , \30398 , \30399 , \30400 ,
         \30401 , \30402 , \30403 , \30404 , \30405 , \30406 , \30407 , \30408 , \30409 , \30410 ,
         \30411 , \30412 , \30413 , \30414 , \30415 , \30416 , \30417 , \30418 , \30419 , \30420 ,
         \30421 , \30422 , \30423 , \30424 , \30425 , \30426 , \30427 , \30428 , \30429 , \30430 ,
         \30431 , \30432 , \30433 , \30434 , \30435 , \30436 , \30437 , \30438 , \30439 , \30440 ,
         \30441 , \30442 , \30443 , \30444 , \30445 , \30446 , \30447 , \30448 , \30449 , \30450 ,
         \30451 , \30452 , \30453 , \30454 , \30455 , \30456 , \30457 , \30458 , \30459 , \30460 ,
         \30461 , \30462 , \30463 , \30464 , \30465 , \30466 , \30467 , \30468 , \30469 , \30470 ,
         \30471 , \30472 , \30473 , \30474 , \30475 , \30476 , \30477 , \30478 , \30479 , \30480 ,
         \30481 , \30482 , \30483 , \30484 , \30485 , \30486 , \30487 , \30488 , \30489 , \30490 ,
         \30491 , \30492 , \30493 , \30494 , \30495 , \30496 , \30497 , \30498 , \30499 , \30500 ,
         \30501 , \30502 , \30503 , \30504 , \30505 , \30506 , \30507 , \30508 , \30509 , \30510 ,
         \30511 , \30512 , \30513 , \30514 , \30515 , \30516 , \30517 , \30518 , \30519 , \30520 ,
         \30521 , \30522 , \30523 , \30524 , \30525 , \30526 , \30527 , \30528 , \30529 , \30530 ,
         \30531 , \30532 , \30533 , \30534 , \30535 , \30536 , \30537 , \30538 , \30539 , \30540 ,
         \30541 , \30542 , \30543 , \30544 , \30545 , \30546 , \30547 , \30548 , \30549 , \30550 ,
         \30551 , \30552 , \30553 , \30554 , \30555 , \30556 , \30557 , \30558 , \30559 , \30560 ,
         \30561 , \30562 , \30563 , \30564 , \30565 , \30566 , \30567 , \30568 , \30569 , \30570 ,
         \30571 , \30572 , \30573 , \30574 , \30575 , \30576 , \30577 , \30578 , \30579 , \30580 ,
         \30581 , \30582 , \30583 , \30584 , \30585 , \30586 , \30587 , \30588 , \30589 , \30590 ,
         \30591 , \30592 , \30593 , \30594 , \30595 , \30596 , \30597 , \30598 , \30599 , \30600 ,
         \30601 , \30602 , \30603 , \30604 , \30605 , \30606 , \30607 , \30608 , \30609 , \30610 ,
         \30611 , \30612 , \30613 , \30614 , \30615 , \30616 , \30617 , \30618 , \30619 , \30620 ,
         \30621 , \30622 , \30623 , \30624 , \30625 , \30626 , \30627 , \30628 , \30629 , \30630 ,
         \30631 , \30632 , \30633 , \30634 , \30635 , \30636 , \30637 , \30638 , \30639 , \30640 ,
         \30641 , \30642 , \30643 , \30644 , \30645 , \30646 , \30647 , \30648 , \30649 , \30650 ,
         \30651 , \30652 , \30653 , \30654 , \30655 , \30656 , \30657 , \30658 , \30659 , \30660 ,
         \30661 , \30662 , \30663 , \30664 , \30665 , \30666 , \30667 , \30668 , \30669 , \30670 ,
         \30671 , \30672 , \30673 , \30674 , \30675 , \30676 , \30677 , \30678 , \30679 , \30680 ,
         \30681 , \30682 , \30683 , \30684 , \30685 , \30686 , \30687 , \30688 , \30689 , \30690 ,
         \30691 , \30692 , \30693 , \30694 , \30695 , \30696 , \30697 , \30698 , \30699 , \30700 ,
         \30701 , \30702 , \30703 , \30704 , \30705 , \30706 , \30707 , \30708 , \30709 , \30710 ,
         \30711 , \30712 , \30713 , \30714 , \30715 , \30716 , \30717 , \30718 , \30719 , \30720 ,
         \30721 , \30722 , \30723 , \30724 , \30725 , \30726 , \30727 , \30728 , \30729 , \30730 ,
         \30731 , \30732 , \30733 , \30734 , \30735 , \30736 , \30737 , \30738 , \30739 , \30740 ,
         \30741 , \30742 , \30743 , \30744 , \30745 , \30746 , \30747 , \30748 , \30749 , \30750 ,
         \30751 , \30752 , \30753 , \30754 , \30755 , \30756 , \30757 , \30758 , \30759 , \30760 ,
         \30761 , \30762 , \30763 , \30764 , \30765 , \30766 , \30767 , \30768 , \30769 , \30770 ,
         \30771 , \30772 , \30773 , \30774 , \30775 , \30776 , \30777 , \30778 , \30779 , \30780 ,
         \30781 , \30782 , \30783 , \30784 , \30785 , \30786 , \30787 , \30788 , \30789 , \30790 ,
         \30791 , \30792 , \30793 , \30794 , \30795 , \30796 , \30797 , \30798 , \30799 , \30800 ,
         \30801 , \30802 , \30803 , \30804 , \30805 , \30806 , \30807 , \30808 , \30809 , \30810 ,
         \30811 , \30812 , \30813 , \30814 , \30815 , \30816 , \30817 , \30818 , \30819 , \30820 ,
         \30821 , \30822 , \30823 , \30824 , \30825 , \30826 , \30827 , \30828 , \30829 , \30830 ,
         \30831 , \30832 , \30833 , \30834 , \30835 , \30836 , \30837 , \30838 , \30839 , \30840 ,
         \30841 , \30842 , \30843 , \30844 , \30845 , \30846 , \30847 , \30848 , \30849 , \30850 ,
         \30851 , \30852 , \30853 , \30854 , \30855 , \30856 , \30857 , \30858 , \30859 , \30860 ,
         \30861 , \30862 , \30863 , \30864 , \30865 , \30866 , \30867 , \30868 , \30869 , \30870 ,
         \30871 , \30872 , \30873 , \30874 , \30875 , \30876 , \30877 , \30878 , \30879 , \30880 ,
         \30881 , \30882 , \30883 , \30884 , \30885 , \30886 , \30887 , \30888 , \30889 , \30890 ,
         \30891 , \30892 , \30893 , \30894 , \30895 , \30896 , \30897 , \30898 , \30899 , \30900 ,
         \30901 , \30902 , \30903 , \30904 , \30905 , \30906 , \30907 , \30908 , \30909 , \30910 ,
         \30911 , \30912 , \30913 , \30914 , \30915 , \30916 , \30917 , \30918 , \30919 , \30920 ,
         \30921 , \30922 , \30923 , \30924 , \30925 , \30926 , \30927 , \30928 , \30929 , \30930 ,
         \30931 , \30932 , \30933 , \30934 , \30935 , \30936 , \30937 , \30938 , \30939 , \30940 ,
         \30941 , \30942 , \30943 , \30944 , \30945 , \30946 , \30947 , \30948 , \30949 , \30950 ,
         \30951 , \30952 , \30953 , \30954 , \30955 , \30956 , \30957 , \30958 , \30959 , \30960 ,
         \30961 , \30962 , \30963 , \30964 , \30965 , \30966 , \30967 , \30968 , \30969 , \30970 ,
         \30971 , \30972 , \30973 , \30974 , \30975 , \30976 , \30977 , \30978 , \30979 , \30980 ,
         \30981 , \30982 , \30983 , \30984 , \30985 , \30986 , \30987 , \30988 , \30989 , \30990 ,
         \30991 , \30992 , \30993 , \30994 , \30995 , \30996 , \30997 , \30998 , \30999 , \31000 ,
         \31001 , \31002 , \31003 , \31004 , \31005 , \31006 , \31007 , \31008 , \31009 , \31010 ,
         \31011 , \31012 , \31013 , \31014 , \31015 , \31016 , \31017 , \31018 , \31019 , \31020 ,
         \31021 , \31022 , \31023 , \31024 , \31025 , \31026 , \31027 , \31028 , \31029 , \31030 ,
         \31031 , \31032 , \31033 , \31034 , \31035 , \31036 , \31037 , \31038 , \31039 , \31040 ,
         \31041 , \31042 , \31043 , \31044 , \31045 , \31046 , \31047 , \31048 , \31049 , \31050 ,
         \31051 , \31052 , \31053 , \31054 , \31055 , \31056 , \31057 , \31058 , \31059 , \31060 ,
         \31061 , \31062 , \31063 , \31064 , \31065 , \31066 , \31067 , \31068 , \31069 , \31070 ,
         \31071 , \31072 , \31073 , \31074 , \31075 , \31076 , \31077 , \31078 , \31079 , \31080 ,
         \31081 , \31082 , \31083 , \31084 , \31085 , \31086 , \31087 , \31088 , \31089 , \31090 ,
         \31091 , \31092 , \31093 , \31094 , \31095 , \31096 , \31097 , \31098 , \31099 , \31100 ,
         \31101 , \31102 , \31103 , \31104 , \31105 , \31106 , \31107 , \31108 , \31109 , \31110 ,
         \31111 , \31112 , \31113 , \31114 , \31115 , \31116 , \31117 , \31118 , \31119 , \31120 ,
         \31121 , \31122 , \31123 , \31124 , \31125 , \31126 , \31127 , \31128 , \31129 , \31130 ,
         \31131 , \31132 , \31133 , \31134 , \31135 , \31136 , \31137 , \31138 , \31139 , \31140 ,
         \31141 , \31142 , \31143 , \31144 , \31145 , \31146 , \31147 , \31148 , \31149 , \31150 ,
         \31151 , \31152 , \31153 , \31154 , \31155 , \31156 , \31157 , \31158 , \31159 , \31160 ,
         \31161 , \31162 , \31163 , \31164 , \31165 , \31166 , \31167 , \31168 , \31169 , \31170 ,
         \31171 , \31172 , \31173 , \31174 , \31175 , \31176 , \31177 , \31178 , \31179 , \31180 ,
         \31181 , \31182 , \31183 , \31184 , \31185 , \31186 , \31187 , \31188 , \31189 , \31190 ,
         \31191 , \31192 , \31193 , \31194 , \31195 , \31196 , \31197 , \31198 , \31199 , \31200 ,
         \31201 , \31202 , \31203 , \31204 , \31205 , \31206 , \31207 , \31208 , \31209 , \31210 ,
         \31211 , \31212 , \31213 , \31214 , \31215 , \31216 , \31217 , \31218 , \31219 , \31220 ,
         \31221 , \31222 , \31223 , \31224 , \31225 , \31226 , \31227 , \31228 , \31229 , \31230 ,
         \31231 , \31232 , \31233 , \31234 , \31235 , \31236 , \31237 , \31238 , \31239 , \31240 ,
         \31241 , \31242 , \31243 , \31244 , \31245 , \31246 , \31247 , \31248 , \31249 , \31250 ,
         \31251 , \31252 , \31253 , \31254 , \31255 , \31256 , \31257 , \31258 , \31259 , \31260 ,
         \31261 , \31262 , \31263 , \31264 , \31265 , \31266 , \31267 , \31268 , \31269 , \31270 ,
         \31271 , \31272 , \31273 , \31274 , \31275 , \31276 , \31277 , \31278 , \31279 , \31280 ,
         \31281 , \31282 , \31283 , \31284 , \31285 , \31286 , \31287 , \31288 , \31289 , \31290 ,
         \31291 , \31292 , \31293 , \31294 , \31295 , \31296 , \31297 , \31298 , \31299 , \31300 ,
         \31301 , \31302 , \31303 , \31304 , \31305 , \31306 , \31307 , \31308 , \31309 , \31310 ,
         \31311 , \31312 , \31313 , \31314 , \31315 , \31316 , \31317 , \31318 , \31319 , \31320 ,
         \31321 , \31322 , \31323 , \31324 , \31325 , \31326 , \31327 , \31328 , \31329 , \31330 ,
         \31331 , \31332 , \31333 , \31334 , \31335 , \31336 , \31337 , \31338 , \31339 , \31340 ,
         \31341 , \31342 , \31343 , \31344 , \31345 , \31346 , \31347 , \31348 , \31349 , \31350 ,
         \31351 , \31352 , \31353 , \31354 , \31355 , \31356 , \31357 , \31358 , \31359 , \31360 ,
         \31361 , \31362 , \31363 , \31364 , \31365 , \31366 , \31367 , \31368 , \31369 , \31370 ,
         \31371 , \31372 , \31373 , \31374 , \31375 , \31376 , \31377 , \31378 , \31379 , \31380 ,
         \31381 , \31382 , \31383 , \31384 , \31385 , \31386 , \31387 , \31388 , \31389 , \31390 ,
         \31391 , \31392 , \31393 , \31394 , \31395 , \31396 , \31397 , \31398 , \31399 , \31400 ,
         \31401 , \31402 , \31403 , \31404 , \31405 , \31406 , \31407 , \31408 , \31409 , \31410 ,
         \31411 , \31412 , \31413 , \31414 , \31415 , \31416 , \31417 , \31418 , \31419 , \31420 ,
         \31421 , \31422 , \31423 , \31424 , \31425 , \31426 , \31427 , \31428 , \31429 , \31430 ,
         \31431 , \31432 , \31433 , \31434 , \31435 , \31436 , \31437 , \31438 , \31439 , \31440 ,
         \31441 , \31442 , \31443 , \31444 , \31445 , \31446 , \31447 , \31448 , \31449 , \31450 ,
         \31451 , \31452 , \31453 , \31454 , \31455 , \31456 , \31457 , \31458 , \31459 , \31460 ,
         \31461 , \31462 , \31463 , \31464 , \31465 , \31466 , \31467 , \31468 , \31469 , \31470 ,
         \31471 , \31472 , \31473 , \31474 , \31475 , \31476 , \31477 , \31478 , \31479 , \31480 ,
         \31481 , \31482 , \31483 , \31484 , \31485 , \31486 , \31487 , \31488 , \31489 , \31490 ,
         \31491 , \31492 , \31493 , \31494 , \31495 , \31496 , \31497 , \31498 , \31499 , \31500 ,
         \31501 , \31502 , \31503 , \31504 , \31505 , \31506 , \31507 , \31508 , \31509 , \31510 ,
         \31511 , \31512 , \31513 , \31514 , \31515 , \31516 , \31517 , \31518 , \31519 , \31520 ,
         \31521 , \31522 , \31523 , \31524 , \31525 , \31526 , \31527 , \31528 , \31529 , \31530 ,
         \31531 , \31532 , \31533 , \31534 , \31535 , \31536 , \31537 , \31538 , \31539 , \31540 ,
         \31541 , \31542 , \31543 , \31544 , \31545 , \31546 , \31547 , \31548 , \31549 , \31550 ,
         \31551 , \31552 , \31553 , \31554 , \31555 , \31556 , \31557 , \31558 , \31559 , \31560 ,
         \31561 , \31562 , \31563 , \31564 , \31565 , \31566 , \31567 , \31568 , \31569 , \31570 ,
         \31571 , \31572 , \31573 , \31574 , \31575 , \31576 , \31577 , \31578 , \31579 , \31580 ,
         \31581 , \31582 , \31583 , \31584 , \31585 , \31586 , \31587 , \31588 , \31589 , \31590 ,
         \31591 , \31592 , \31593 , \31594 , \31595 , \31596 , \31597 , \31598 , \31599 , \31600 ,
         \31601 , \31602 , \31603 , \31604 , \31605 , \31606 , \31607 , \31608 , \31609 , \31610 ,
         \31611 , \31612 , \31613 , \31614 , \31615 , \31616 , \31617 , \31618 , \31619 , \31620 ,
         \31621 , \31622 , \31623 , \31624 , \31625 , \31626 , \31627 , \31628 , \31629 , \31630 ,
         \31631 , \31632 , \31633 , \31634 , \31635 , \31636 , \31637 , \31638 , \31639 , \31640 ,
         \31641 , \31642 , \31643 , \31644 , \31645 , \31646 , \31647 , \31648 , \31649 , \31650 ,
         \31651 , \31652 , \31653 , \31654 , \31655 , \31656 , \31657 , \31658 , \31659 , \31660 ,
         \31661 , \31662 , \31663 , \31664 , \31665 , \31666 , \31667 , \31668 , \31669 , \31670 ,
         \31671 , \31672 , \31673 , \31674 , \31675 , \31676 , \31677 , \31678 , \31679 , \31680 ,
         \31681 , \31682 , \31683 , \31684 , \31685 , \31686 , \31687 , \31688 , \31689 , \31690 ,
         \31691 , \31692 , \31693 , \31694 , \31695 , \31696 , \31697 , \31698 , \31699 , \31700 ,
         \31701 , \31702 , \31703 , \31704 , \31705 , \31706 , \31707 , \31708 , \31709 , \31710 ,
         \31711 , \31712 , \31713 , \31714 , \31715 , \31716 , \31717 , \31718 , \31719 , \31720 ,
         \31721 , \31722 , \31723 , \31724 , \31725 , \31726 , \31727 , \31728 , \31729 , \31730 ,
         \31731 , \31732 , \31733 , \31734 , \31735 , \31736 , \31737 , \31738 , \31739 , \31740 ,
         \31741 , \31742 , \31743 , \31744 , \31745 , \31746 , \31747 , \31748 , \31749 , \31750 ,
         \31751 , \31752 , \31753 , \31754 , \31755 , \31756 , \31757 , \31758 , \31759 , \31760 ,
         \31761 , \31762 , \31763 , \31764 , \31765 , \31766 , \31767 , \31768 , \31769 , \31770 ,
         \31771 , \31772 , \31773 , \31774 , \31775 , \31776 , \31777 , \31778 , \31779 , \31780 ,
         \31781 , \31782 , \31783 , \31784 , \31785 , \31786 , \31787 , \31788 , \31789 , \31790 ,
         \31791 , \31792 , \31793 , \31794 , \31795 , \31796 , \31797 , \31798 , \31799 , \31800 ,
         \31801 , \31802 , \31803 , \31804 , \31805 , \31806 , \31807 , \31808 , \31809 , \31810 ,
         \31811 , \31812 , \31813 , \31814 , \31815 , \31816 , \31817 , \31818 , \31819 , \31820 ,
         \31821 , \31822 , \31823 , \31824 , \31825 , \31826 , \31827 , \31828 , \31829 , \31830 ,
         \31831 , \31832 , \31833 , \31834 , \31835 , \31836 , \31837 , \31838 , \31839 , \31840 ,
         \31841 , \31842 , \31843 , \31844 , \31845 , \31846 , \31847 , \31848 , \31849 , \31850 ,
         \31851 , \31852 , \31853 , \31854 , \31855 , \31856 , \31857 , \31858 , \31859 , \31860 ,
         \31861 , \31862 , \31863 , \31864 , \31865 , \31866 , \31867 , \31868 , \31869 , \31870 ,
         \31871 , \31872 , \31873 , \31874 , \31875 , \31876 , \31877 , \31878 , \31879 , \31880 ,
         \31881 , \31882 , \31883 , \31884 , \31885 , \31886 , \31887 , \31888 , \31889 , \31890 ,
         \31891 , \31892 , \31893 , \31894 , \31895 , \31896 , \31897 , \31898 , \31899 , \31900 ,
         \31901 , \31902 , \31903 , \31904 , \31905 , \31906 , \31907 , \31908 , \31909 , \31910 ,
         \31911 , \31912 , \31913 , \31914 , \31915 , \31916 , \31917 , \31918 , \31919 , \31920 ,
         \31921 , \31922 , \31923 , \31924 , \31925 , \31926 , \31927 , \31928 , \31929 , \31930 ,
         \31931 , \31932 , \31933 , \31934 , \31935 , \31936 , \31937 , \31938 , \31939 , \31940 ,
         \31941 , \31942 , \31943 , \31944 , \31945 , \31946 , \31947 , \31948 , \31949 , \31950 ,
         \31951 , \31952 , \31953 , \31954 , \31955 , \31956 , \31957 , \31958 , \31959 , \31960 ,
         \31961 , \31962 , \31963 , \31964 , \31965 , \31966 , \31967 , \31968 , \31969 , \31970 ,
         \31971 , \31972 , \31973 , \31974 , \31975 , \31976 , \31977 , \31978 , \31979 , \31980 ,
         \31981 , \31982 , \31983 , \31984 , \31985 , \31986 , \31987 , \31988 , \31989 , \31990 ,
         \31991 , \31992 , \31993 , \31994 , \31995 , \31996 , \31997 , \31998 , \31999 , \32000 ,
         \32001 , \32002 , \32003 , \32004 , \32005 , \32006 , \32007 , \32008 , \32009 , \32010 ,
         \32011 , \32012 , \32013 , \32014 , \32015 , \32016 , \32017 , \32018 , \32019 , \32020 ,
         \32021 , \32022 , \32023 , \32024 , \32025 , \32026 , \32027 , \32028 , \32029 , \32030 ,
         \32031 , \32032 , \32033 , \32034 , \32035 , \32036 , \32037 , \32038 , \32039 , \32040 ,
         \32041 , \32042 , \32043 , \32044 , \32045 , \32046 , \32047 , \32048 , \32049 , \32050 ,
         \32051 , \32052 , \32053 , \32054 , \32055 , \32056 , \32057 , \32058 , \32059 , \32060 ,
         \32061 , \32062 , \32063 , \32064 , \32065 , \32066 , \32067 , \32068 , \32069 , \32070 ,
         \32071 , \32072 , \32073 , \32074 , \32075 , \32076 , \32077 , \32078 , \32079 , \32080 ,
         \32081 , \32082 , \32083 , \32084 , \32085 , \32086 , \32087 , \32088 , \32089 , \32090 ,
         \32091 , \32092 , \32093 , \32094 , \32095 , \32096 , \32097 , \32098 , \32099 , \32100 ,
         \32101 , \32102 , \32103 , \32104 , \32105 , \32106 , \32107 , \32108 , \32109 , \32110 ,
         \32111 , \32112 , \32113 , \32114 , \32115 , \32116 , \32117 , \32118 , \32119 , \32120 ,
         \32121 , \32122 , \32123 , \32124 , \32125 , \32126 , \32127 , \32128 , \32129 , \32130 ,
         \32131 , \32132 , \32133 , \32134 , \32135 , \32136 , \32137 , \32138 , \32139 , \32140 ,
         \32141 , \32142 , \32143 , \32144 , \32145 , \32146 , \32147 , \32148 , \32149 , \32150 ,
         \32151 , \32152 , \32153 , \32154 , \32155 , \32156 , \32157 , \32158 , \32159 , \32160 ,
         \32161 , \32162 , \32163 , \32164 , \32165 , \32166 , \32167 , \32168 , \32169 , \32170 ,
         \32171 , \32172 , \32173 , \32174 , \32175 , \32176 , \32177 , \32178 , \32179 , \32180 ,
         \32181 , \32182 , \32183 , \32184 , \32185 , \32186 , \32187 , \32188 , \32189 , \32190 ,
         \32191 , \32192 , \32193 , \32194 , \32195 , \32196 , \32197 , \32198 , \32199 , \32200 ,
         \32201 , \32202 , \32203 , \32204 , \32205 , \32206 , \32207 , \32208 , \32209 , \32210 ,
         \32211 , \32212 , \32213 , \32214 , \32215 , \32216 , \32217 , \32218 , \32219 , \32220 ,
         \32221 , \32222 , \32223 , \32224 , \32225 , \32226 , \32227 , \32228 , \32229 , \32230 ,
         \32231 , \32232 , \32233 , \32234 , \32235 , \32236 , \32237 , \32238 , \32239 , \32240 ,
         \32241 , \32242 , \32243 , \32244 , \32245 , \32246 , \32247 , \32248 , \32249 , \32250 ,
         \32251 , \32252 , \32253 , \32254 , \32255 , \32256 , \32257 , \32258 , \32259 , \32260 ,
         \32261 , \32262 , \32263 , \32264 , \32265 , \32266 , \32267 , \32268 , \32269 , \32270 ,
         \32271 , \32272 , \32273 , \32274 , \32275 , \32276 , \32277 , \32278 , \32279 , \32280 ,
         \32281 , \32282 , \32283 , \32284 , \32285 , \32286 , \32287 , \32288 , \32289 , \32290 ,
         \32291 , \32292 , \32293 , \32294 , \32295 , \32296 , \32297 , \32298 , \32299 , \32300 ,
         \32301 , \32302 , \32303 , \32304 , \32305 , \32306 , \32307 , \32308 , \32309 , \32310 ,
         \32311 , \32312 , \32313 , \32314 , \32315 , \32316 , \32317 , \32318 , \32319 , \32320 ,
         \32321 , \32322 , \32323 , \32324 , \32325 , \32326 , \32327 , \32328 , \32329 , \32330 ,
         \32331 , \32332 , \32333 , \32334 , \32335 , \32336 , \32337 , \32338 , \32339 , \32340 ,
         \32341 , \32342 , \32343 , \32344 , \32345 , \32346 , \32347 , \32348 , \32349 , \32350 ,
         \32351 , \32352 , \32353 , \32354 , \32355 , \32356 , \32357 , \32358 , \32359 , \32360 ,
         \32361 , \32362 , \32363 , \32364 , \32365 , \32366 , \32367 , \32368 , \32369 , \32370 ,
         \32371 , \32372 , \32373 , \32374 , \32375 , \32376 , \32377 , \32378 , \32379 , \32380 ,
         \32381 , \32382 , \32383 , \32384 , \32385 , \32386 , \32387 , \32388 , \32389 , \32390 ,
         \32391 , \32392 , \32393 , \32394 , \32395 , \32396 , \32397 , \32398 , \32399 , \32400 ,
         \32401 , \32402 , \32403 , \32404 , \32405 , \32406 , \32407 , \32408 , \32409 , \32410 ,
         \32411 , \32412 , \32413 , \32414 , \32415 , \32416 , \32417 , \32418 , \32419 , \32420 ,
         \32421 , \32422 , \32423 , \32424 , \32425 , \32426 , \32427 , \32428 , \32429 , \32430 ,
         \32431 , \32432 , \32433 , \32434 , \32435 , \32436 , \32437 , \32438 , \32439 , \32440 ,
         \32441 , \32442 , \32443 , \32444 , \32445 , \32446 , \32447 , \32448 , \32449 , \32450 ,
         \32451 , \32452 , \32453 , \32454 , \32455 , \32456 , \32457 , \32458 , \32459 , \32460 ,
         \32461 , \32462 , \32463 , \32464 , \32465 , \32466 , \32467 , \32468 , \32469 , \32470 ,
         \32471 , \32472 , \32473 , \32474 , \32475 , \32476 , \32477 , \32478 , \32479 , \32480 ,
         \32481 , \32482 , \32483 , \32484 , \32485 , \32486 , \32487 , \32488 , \32489 , \32490 ,
         \32491 , \32492 , \32493 , \32494 , \32495 , \32496 , \32497 , \32498 , \32499 , \32500 ,
         \32501 , \32502 , \32503 , \32504 , \32505 , \32506 , \32507 , \32508 , \32509 , \32510 ,
         \32511 , \32512 , \32513 , \32514 , \32515 , \32516 , \32517 , \32518 , \32519 , \32520 ,
         \32521 , \32522 , \32523 , \32524 , \32525 , \32526 , \32527 , \32528 , \32529 , \32530 ,
         \32531 , \32532 , \32533 , \32534 , \32535 , \32536 , \32537 , \32538 , \32539 , \32540 ,
         \32541 , \32542 , \32543 , \32544 , \32545 , \32546 , \32547 , \32548 , \32549 , \32550 ,
         \32551 , \32552 , \32553 , \32554 , \32555 , \32556 , \32557 , \32558 , \32559 , \32560 ,
         \32561 , \32562 , \32563 , \32564 , \32565 , \32566 , \32567 , \32568 , \32569 , \32570 ,
         \32571 , \32572 , \32573 , \32574 , \32575 , \32576 , \32577 , \32578 , \32579 , \32580 ,
         \32581 , \32582 , \32583 , \32584 , \32585 , \32586 , \32587 , \32588 , \32589 , \32590 ,
         \32591 , \32592 , \32593 , \32594 , \32595 , \32596 , \32597 , \32598 , \32599 , \32600 ,
         \32601 , \32602 , \32603 , \32604 , \32605 , \32606 , \32607 , \32608 , \32609 , \32610 ,
         \32611 , \32612 , \32613 , \32614 , \32615 , \32616 , \32617 , \32618 , \32619 , \32620 ,
         \32621 , \32622 , \32623 , \32624 , \32625 , \32626 , \32627 , \32628 , \32629 , \32630 ,
         \32631 , \32632 , \32633 , \32634 , \32635 , \32636 , \32637 , \32638 , \32639 , \32640 ,
         \32641 , \32642 , \32643 , \32644 , \32645 , \32646 , \32647 , \32648 , \32649 , \32650 ,
         \32651 , \32652 , \32653 , \32654 , \32655 , \32656 , \32657 , \32658 , \32659 , \32660 ,
         \32661 , \32662 , \32663 , \32664 , \32665 , \32666 , \32667 , \32668 , \32669 , \32670 ,
         \32671 , \32672 , \32673 , \32674 , \32675 , \32676 , \32677 , \32678 , \32679 , \32680 ,
         \32681 , \32682 , \32683 , \32684 , \32685 , \32686 , \32687 , \32688 , \32689 , \32690 ,
         \32691 , \32692 , \32693 , \32694 , \32695 , \32696 , \32697 , \32698 , \32699 , \32700 ,
         \32701 , \32702 , \32703 , \32704 , \32705 , \32706 , \32707 , \32708 , \32709 , \32710 ,
         \32711 , \32712 , \32713 , \32714 , \32715 , \32716 , \32717 , \32718 , \32719 , \32720 ,
         \32721 , \32722 , \32723 , \32724 , \32725 , \32726 , \32727 , \32728 , \32729 , \32730 ,
         \32731 , \32732 , \32733 , \32734 , \32735 , \32736 , \32737 , \32738 , \32739 , \32740 ,
         \32741 , \32742 , \32743 , \32744 , \32745 , \32746 , \32747 , \32748 , \32749 , \32750 ,
         \32751 , \32752 , \32753 , \32754 , \32755 , \32756 , \32757 , \32758 , \32759 , \32760 ,
         \32761 , \32762 , \32763 , \32764 , \32765 , \32766 , \32767 , \32768 , \32769 , \32770 ,
         \32771 , \32772 , \32773 , \32774 , \32775 , \32776 , \32777 , \32778 , \32779 , \32780 ,
         \32781 , \32782 , \32783 , \32784 , \32785 , \32786 , \32787 , \32788 , \32789 , \32790 ,
         \32791 , \32792 , \32793 , \32794 , \32795 , \32796 , \32797 , \32798 , \32799 , \32800 ,
         \32801 , \32802 , \32803 , \32804 , \32805 , \32806 , \32807 , \32808 , \32809 , \32810 ,
         \32811 , \32812 , \32813 , \32814 , \32815 , \32816 , \32817 , \32818 , \32819 , \32820 ,
         \32821 , \32822 , \32823 , \32824 , \32825 , \32826 , \32827 , \32828 , \32829 , \32830 ,
         \32831 , \32832 , \32833 , \32834 , \32835 , \32836 , \32837 , \32838 , \32839 , \32840 ,
         \32841 , \32842 , \32843 , \32844 , \32845 , \32846 , \32847 , \32848 , \32849 , \32850 ,
         \32851 , \32852 , \32853 , \32854 , \32855 , \32856 , \32857 , \32858 , \32859 , \32860 ,
         \32861 , \32862 , \32863 , \32864 , \32865 , \32866 , \32867 , \32868 , \32869 , \32870 ,
         \32871 , \32872 , \32873 , \32874 , \32875 , \32876 , \32877 , \32878 , \32879 , \32880 ,
         \32881 , \32882 , \32883 , \32884 , \32885 , \32886 , \32887 , \32888 , \32889 , \32890 ,
         \32891 , \32892 , \32893 , \32894 , \32895 , \32896 , \32897 , \32898 , \32899 , \32900 ,
         \32901 , \32902 , \32903 , \32904 , \32905 , \32906 , \32907 , \32908 , \32909 , \32910 ,
         \32911 , \32912 , \32913 , \32914 , \32915 , \32916 , \32917 , \32918 , \32919 , \32920 ,
         \32921 , \32922 , \32923 , \32924 , \32925 , \32926 , \32927 , \32928 , \32929 , \32930 ,
         \32931 , \32932 , \32933 , \32934 , \32935 , \32936 , \32937 , \32938 , \32939 , \32940 ,
         \32941 , \32942 , \32943 , \32944 , \32945 , \32946 , \32947 , \32948 , \32949 , \32950 ,
         \32951 , \32952 , \32953 , \32954 , \32955 , \32956 , \32957 , \32958 , \32959 , \32960 ,
         \32961 , \32962 , \32963 , \32964 , \32965 , \32966 , \32967 , \32968 , \32969 , \32970 ,
         \32971 , \32972 , \32973 , \32974 , \32975 , \32976 , \32977 , \32978 , \32979 , \32980 ,
         \32981 , \32982 , \32983 , \32984 , \32985 , \32986 , \32987 , \32988 , \32989 , \32990 ,
         \32991 , \32992 , \32993 , \32994 , \32995 , \32996 , \32997 , \32998 , \32999 , \33000 ,
         \33001 , \33002 , \33003 , \33004 , \33005 , \33006 , \33007 , \33008 , \33009 , \33010 ,
         \33011 , \33012 , \33013 , \33014 , \33015 , \33016 , \33017 , \33018 , \33019 , \33020 ,
         \33021 , \33022 , \33023 , \33024 , \33025 , \33026 , \33027 , \33028 , \33029 , \33030 ,
         \33031 , \33032 , \33033 , \33034 , \33035 , \33036 , \33037 , \33038 , \33039 , \33040 ,
         \33041 , \33042 , \33043 , \33044 , \33045 , \33046 , \33047 , \33048 , \33049 , \33050 ,
         \33051 , \33052 , \33053 , \33054 , \33055 , \33056 , \33057 , \33058 , \33059 , \33060 ,
         \33061 , \33062 , \33063 , \33064 , \33065 , \33066 , \33067 , \33068 , \33069 , \33070 ,
         \33071 , \33072 , \33073 , \33074 , \33075 , \33076 , \33077 , \33078 , \33079 , \33080 ,
         \33081 , \33082 , \33083 , \33084 , \33085 , \33086 , \33087 , \33088 , \33089 , \33090 ,
         \33091 , \33092 , \33093 , \33094 , \33095 , \33096 , \33097 , \33098 , \33099 , \33100 ,
         \33101 , \33102 , \33103 , \33104 , \33105 , \33106 , \33107 , \33108 , \33109 , \33110 ,
         \33111 , \33112 , \33113 , \33114 , \33115 , \33116 , \33117 , \33118 , \33119 , \33120 ,
         \33121 , \33122 , \33123 , \33124 , \33125 , \33126 , \33127 , \33128 , \33129 , \33130 ,
         \33131 , \33132 , \33133 , \33134 , \33135 , \33136 , \33137 , \33138 , \33139 , \33140 ,
         \33141 , \33142 , \33143 , \33144 , \33145 , \33146 , \33147 , \33148 , \33149 , \33150 ,
         \33151 , \33152 , \33153 , \33154 , \33155 , \33156 , \33157 , \33158 , \33159 , \33160 ,
         \33161 , \33162 , \33163 , \33164 , \33165 , \33166 , \33167 , \33168 , \33169 , \33170 ,
         \33171 , \33172 , \33173 , \33174 , \33175 , \33176 , \33177 , \33178 , \33179 , \33180 ,
         \33181 , \33182 , \33183 , \33184 , \33185 , \33186 , \33187 , \33188 , \33189 , \33190 ,
         \33191 , \33192 , \33193 , \33194 , \33195 , \33196 , \33197 , \33198 , \33199 , \33200 ,
         \33201 , \33202 , \33203 , \33204 , \33205 , \33206 , \33207 , \33208 , \33209 , \33210 ,
         \33211 , \33212 , \33213 , \33214 , \33215 , \33216 , \33217 , \33218 , \33219 , \33220 ,
         \33221 , \33222 , \33223 , \33224 , \33225 , \33226 , \33227 , \33228 , \33229 , \33230 ,
         \33231 , \33232 , \33233 , \33234 , \33235 , \33236 , \33237 , \33238 , \33239 , \33240 ,
         \33241 , \33242 , \33243 , \33244 , \33245 , \33246 , \33247 , \33248 , \33249 , \33250 ,
         \33251 , \33252 , \33253 , \33254 , \33255 , \33256 , \33257 , \33258 , \33259 , \33260 ,
         \33261 , \33262 , \33263 , \33264 , \33265 , \33266 , \33267 , \33268 , \33269 , \33270 ,
         \33271 , \33272 , \33273 , \33274 , \33275 , \33276 , \33277 , \33278 , \33279 , \33280 ,
         \33281 , \33282 , \33283 , \33284 , \33285 , \33286 , \33287 , \33288 , \33289 , \33290 ,
         \33291 , \33292 , \33293 , \33294 , \33295 , \33296 , \33297 , \33298 , \33299 , \33300 ,
         \33301 , \33302 , \33303 , \33304 , \33305 , \33306 , \33307 , \33308 , \33309 , \33310 ,
         \33311 , \33312 , \33313 , \33314 , \33315 , \33316 , \33317 , \33318 , \33319 , \33320 ,
         \33321 , \33322 , \33323 , \33324 , \33325 , \33326 , \33327 , \33328 , \33329 , \33330 ,
         \33331 , \33332 , \33333 , \33334 , \33335 , \33336 , \33337 , \33338 , \33339 , \33340 ,
         \33341 , \33342 , \33343 , \33344 , \33345 , \33346 , \33347 , \33348 , \33349 , \33350 ,
         \33351 , \33352 , \33353 , \33354 , \33355 , \33356 , \33357 , \33358 , \33359 , \33360 ,
         \33361 , \33362 , \33363 , \33364 , \33365 , \33366 , \33367 , \33368 , \33369 , \33370 ,
         \33371 , \33372 , \33373 , \33374 , \33375 , \33376 , \33377 , \33378 , \33379 , \33380 ,
         \33381 , \33382 , \33383 , \33384 , \33385 , \33386 , \33387 , \33388 , \33389 , \33390 ,
         \33391 , \33392 , \33393 , \33394 , \33395 , \33396 , \33397 , \33398 , \33399 , \33400 ,
         \33401 , \33402 , \33403 , \33404 , \33405 , \33406 , \33407 , \33408 , \33409 , \33410 ,
         \33411 , \33412 , \33413 , \33414 , \33415 , \33416 , \33417 , \33418 , \33419 , \33420 ,
         \33421 , \33422 , \33423 , \33424 , \33425 , \33426 , \33427 , \33428 , \33429 , \33430 ,
         \33431 , \33432 , \33433 , \33434 , \33435 , \33436 , \33437 , \33438 , \33439 , \33440 ,
         \33441 , \33442 , \33443 , \33444 , \33445 , \33446 , \33447 , \33448 , \33449 , \33450 ,
         \33451 , \33452 , \33453 , \33454 , \33455 , \33456 , \33457 , \33458 , \33459 , \33460 ,
         \33461 , \33462 , \33463 , \33464 , \33465 , \33466 , \33467 , \33468 , \33469 , \33470 ,
         \33471 , \33472 , \33473 , \33474 , \33475 , \33476 , \33477 , \33478 , \33479 , \33480 ,
         \33481 , \33482 , \33483 , \33484 , \33485 , \33486 , \33487 , \33488 , \33489 , \33490 ,
         \33491 , \33492 , \33493 , \33494 , \33495 , \33496 , \33497 , \33498 , \33499 , \33500 ,
         \33501 , \33502 , \33503 , \33504 , \33505 , \33506 , \33507 , \33508 , \33509 , \33510 ,
         \33511 , \33512 , \33513 , \33514 , \33515 , \33516 , \33517 , \33518 , \33519 , \33520 ,
         \33521 , \33522 , \33523 , \33524 , \33525 , \33526 , \33527 , \33528 , \33529 , \33530 ,
         \33531 , \33532 , \33533 , \33534 , \33535 , \33536 , \33537 , \33538 , \33539 , \33540 ,
         \33541 , \33542 , \33543 , \33544 , \33545 , \33546 , \33547 , \33548 , \33549 , \33550 ,
         \33551 , \33552 , \33553 , \33554 , \33555 , \33556 , \33557 , \33558 , \33559 , \33560 ,
         \33561 , \33562 , \33563 , \33564 , \33565 , \33566 , \33567 , \33568 , \33569 , \33570 ,
         \33571 , \33572 , \33573 , \33574 , \33575 , \33576 , \33577 , \33578 , \33579 , \33580 ,
         \33581 , \33582 , \33583 , \33584 , \33585 , \33586 , \33587 , \33588 , \33589 , \33590 ,
         \33591 , \33592 , \33593 , \33594 , \33595 , \33596 , \33597 , \33598 , \33599 , \33600 ,
         \33601 , \33602 , \33603 , \33604 , \33605 , \33606 , \33607 , \33608 , \33609 , \33610 ,
         \33611 , \33612 , \33613 , \33614 , \33615 , \33616 , \33617 , \33618 , \33619 , \33620 ,
         \33621 , \33622 , \33623 , \33624 , \33625 , \33626 , \33627 , \33628 , \33629 , \33630 ,
         \33631 , \33632 , \33633 , \33634 , \33635 , \33636 , \33637 , \33638 , \33639 , \33640 ,
         \33641 , \33642 , \33643 , \33644 , \33645 , \33646 , \33647 , \33648 , \33649 , \33650 ,
         \33651 , \33652 , \33653 , \33654 , \33655 , \33656 , \33657 , \33658 , \33659 , \33660 ,
         \33661 , \33662 , \33663 , \33664 , \33665 , \33666 , \33667 , \33668 , \33669 , \33670 ,
         \33671 , \33672 , \33673 , \33674 , \33675 , \33676 , \33677 , \33678 , \33679 , \33680 ,
         \33681 , \33682 , \33683 , \33684 , \33685 , \33686 , \33687 , \33688 , \33689 , \33690 ,
         \33691 , \33692 , \33693 , \33694 , \33695 , \33696 , \33697 , \33698 , \33699 , \33700 ,
         \33701 , \33702 , \33703 , \33704 , \33705 , \33706 , \33707 , \33708 , \33709 , \33710 ,
         \33711 , \33712 , \33713 , \33714 , \33715 , \33716 , \33717 , \33718 , \33719 , \33720 ,
         \33721 , \33722 , \33723 , \33724 , \33725 , \33726 , \33727 , \33728 , \33729 , \33730 ,
         \33731 , \33732 , \33733 , \33734 , \33735 , \33736 , \33737 , \33738 , \33739 , \33740 ,
         \33741 , \33742 , \33743 , \33744 , \33745 , \33746 , \33747 , \33748 , \33749 , \33750 ,
         \33751 , \33752 , \33753 , \33754 , \33755 , \33756 , \33757 , \33758 , \33759 , \33760 ,
         \33761 , \33762 , \33763 , \33764 , \33765 , \33766 , \33767 , \33768 , \33769 , \33770 ,
         \33771 , \33772 , \33773 , \33774 , \33775 , \33776 , \33777 , \33778 , \33779 , \33780 ,
         \33781 , \33782 , \33783 , \33784 , \33785 , \33786 , \33787 , \33788 , \33789 , \33790 ,
         \33791 , \33792 , \33793 , \33794 , \33795 , \33796 , \33797 , \33798 , \33799 , \33800 ,
         \33801 , \33802 , \33803 , \33804 , \33805 , \33806 , \33807 , \33808 , \33809 , \33810 ,
         \33811 , \33812 , \33813 , \33814 , \33815 , \33816 , \33817 , \33818 , \33819 , \33820 ,
         \33821 , \33822 , \33823 , \33824 , \33825 , \33826 , \33827 , \33828 , \33829 , \33830 ,
         \33831 , \33832 , \33833 , \33834 , \33835 , \33836 , \33837 , \33838 , \33839 , \33840 ,
         \33841 , \33842 , \33843 , \33844 , \33845 , \33846 , \33847 , \33848 , \33849 , \33850 ,
         \33851 , \33852 , \33853 , \33854 , \33855 , \33856 , \33857 , \33858 , \33859 , \33860 ,
         \33861 , \33862 , \33863 , \33864 , \33865 , \33866 , \33867 , \33868 , \33869 , \33870 ,
         \33871 , \33872 , \33873 , \33874 , \33875 , \33876 , \33877 , \33878 , \33879 , \33880 ,
         \33881 , \33882 , \33883 , \33884 , \33885 , \33886 , \33887 , \33888 , \33889 , \33890 ,
         \33891 , \33892 , \33893 , \33894 , \33895 , \33896 , \33897 , \33898 , \33899 , \33900 ,
         \33901 , \33902 , \33903 , \33904 , \33905 , \33906 , \33907 , \33908 , \33909 , \33910 ,
         \33911 , \33912 , \33913 , \33914 , \33915 , \33916 , \33917 , \33918 , \33919 , \33920 ,
         \33921 , \33922 , \33923 , \33924 , \33925 , \33926 , \33927 , \33928 , \33929 , \33930 ,
         \33931 , \33932 , \33933 , \33934 , \33935 , \33936 , \33937 , \33938 , \33939 , \33940 ,
         \33941 , \33942 , \33943 , \33944 , \33945 , \33946 , \33947 , \33948 , \33949 , \33950 ,
         \33951 , \33952 , \33953 , \33954 , \33955 , \33956 , \33957 , \33958 , \33959 , \33960 ,
         \33961 , \33962 , \33963 , \33964 , \33965 , \33966 , \33967 , \33968 , \33969 , \33970 ,
         \33971 , \33972 , \33973 , \33974 , \33975 , \33976 , \33977 , \33978 , \33979 , \33980 ,
         \33981 , \33982 , \33983 , \33984 , \33985 , \33986 , \33987 , \33988 , \33989 , \33990 ,
         \33991 , \33992 , \33993 , \33994 , \33995 , \33996 , \33997 , \33998 , \33999 , \34000 ,
         \34001 , \34002 , \34003 , \34004 , \34005 , \34006 , \34007 , \34008 , \34009 , \34010 ,
         \34011 , \34012 , \34013 , \34014 , \34015 , \34016 , \34017 , \34018 , \34019 , \34020 ,
         \34021 , \34022 , \34023 , \34024 , \34025 , \34026 , \34027 , \34028 , \34029 , \34030 ,
         \34031 , \34032 , \34033 , \34034 , \34035 , \34036 , \34037 , \34038 , \34039 , \34040 ,
         \34041 , \34042 , \34043 , \34044 , \34045 , \34046 , \34047 , \34048 , \34049 , \34050 ,
         \34051 , \34052 , \34053 , \34054 , \34055 , \34056 , \34057 , \34058 , \34059 , \34060 ,
         \34061 , \34062 , \34063 , \34064 , \34065 , \34066 , \34067 , \34068 , \34069 , \34070 ,
         \34071 , \34072 , \34073 , \34074 , \34075 , \34076 , \34077 , \34078 , \34079 , \34080 ,
         \34081 , \34082 , \34083 , \34084 , \34085 , \34086 , \34087 , \34088 , \34089 , \34090 ,
         \34091 , \34092 , \34093 , \34094 , \34095 , \34096 , \34097 , \34098 , \34099 , \34100 ,
         \34101 , \34102 , \34103 , \34104 , \34105 , \34106 , \34107 , \34108 , \34109 , \34110 ,
         \34111 , \34112 , \34113 , \34114 , \34115 , \34116 , \34117 , \34118 , \34119 , \34120 ,
         \34121 , \34122 , \34123 , \34124 , \34125 , \34126 , \34127 , \34128 , \34129 , \34130 ,
         \34131 , \34132 , \34133 , \34134 , \34135 , \34136 , \34137 , \34138 , \34139 , \34140 ,
         \34141 , \34142 , \34143 , \34144 , \34145 , \34146 , \34147 , \34148 , \34149 , \34150 ,
         \34151 , \34152 , \34153 , \34154 , \34155 , \34156 , \34157 , \34158 , \34159 , \34160 ,
         \34161 , \34162 , \34163 , \34164 , \34165 , \34166 , \34167 , \34168 , \34169 , \34170 ,
         \34171 , \34172 , \34173 , \34174 , \34175 , \34176 , \34177 , \34178 , \34179 , \34180 ,
         \34181 , \34182 , \34183 , \34184 , \34185 , \34186 , \34187 , \34188 , \34189 , \34190 ,
         \34191 , \34192 , \34193 , \34194 , \34195 , \34196 , \34197 , \34198 , \34199 , \34200 ,
         \34201 , \34202 , \34203 , \34204 , \34205 , \34206 , \34207 , \34208 , \34209 , \34210 ,
         \34211 , \34212 , \34213 , \34214 , \34215 , \34216 , \34217 , \34218 , \34219 , \34220 ,
         \34221 , \34222 , \34223 , \34224 , \34225 , \34226 , \34227 , \34228 , \34229 , \34230 ,
         \34231 , \34232 , \34233 , \34234 , \34235 , \34236 , \34237 , \34238 , \34239 , \34240 ,
         \34241 , \34242 , \34243 , \34244 , \34245 , \34246 , \34247 , \34248 , \34249 , \34250 ,
         \34251 , \34252 , \34253 , \34254 , \34255 , \34256 , \34257 , \34258 , \34259 , \34260 ,
         \34261 , \34262 , \34263 , \34264 , \34265 , \34266 , \34267 , \34268 , \34269 , \34270 ,
         \34271 , \34272 , \34273 , \34274 , \34275 , \34276 , \34277 , \34278 , \34279 , \34280 ,
         \34281 , \34282 , \34283 , \34284 , \34285 , \34286 , \34287 , \34288 , \34289 , \34290 ,
         \34291 , \34292 , \34293 , \34294 , \34295 , \34296 , \34297 , \34298 , \34299 , \34300 ,
         \34301 , \34302 , \34303 , \34304 , \34305 , \34306 , \34307 , \34308 , \34309 , \34310 ,
         \34311 , \34312 , \34313 , \34314 , \34315 , \34316 , \34317 , \34318 , \34319 , \34320 ,
         \34321 , \34322 , \34323 , \34324 , \34325 , \34326 , \34327 , \34328 , \34329 , \34330 ,
         \34331 , \34332 , \34333 , \34334 , \34335 , \34336 , \34337 , \34338 , \34339 , \34340 ,
         \34341 , \34342 , \34343 , \34344 , \34345 , \34346 , \34347 , \34348 , \34349 , \34350 ,
         \34351 , \34352 , \34353 , \34354 , \34355 , \34356 , \34357 , \34358 , \34359 , \34360 ,
         \34361 , \34362 , \34363 , \34364 , \34365 , \34366 , \34367 , \34368 , \34369 , \34370 ,
         \34371 , \34372 , \34373 , \34374 , \34375 , \34376 , \34377 , \34378 , \34379 , \34380 ,
         \34381 , \34382 , \34383 , \34384 , \34385 , \34386 , \34387 , \34388 , \34389 , \34390 ,
         \34391 , \34392 , \34393 , \34394 , \34395 , \34396 , \34397 , \34398 , \34399 , \34400 ,
         \34401 , \34402 , \34403 , \34404 , \34405 , \34406 , \34407 , \34408 , \34409 , \34410 ,
         \34411 , \34412 , \34413 , \34414 , \34415 , \34416 , \34417 , \34418 , \34419 , \34420 ,
         \34421 , \34422 , \34423 , \34424 , \34425 , \34426 , \34427 , \34428 , \34429 , \34430 ,
         \34431 , \34432 , \34433 , \34434 , \34435 , \34436 , \34437 , \34438 , \34439 , \34440 ,
         \34441 , \34442 , \34443 , \34444 , \34445 , \34446 , \34447 , \34448 , \34449 , \34450 ,
         \34451 , \34452 , \34453 , \34454 , \34455 , \34456 , \34457 , \34458 , \34459 , \34460 ,
         \34461 , \34462 , \34463 , \34464 , \34465 , \34466 , \34467 , \34468 , \34469 , \34470 ,
         \34471 , \34472 , \34473 , \34474 , \34475 , \34476 , \34477 , \34478 , \34479 , \34480 ,
         \34481 , \34482 , \34483 , \34484 , \34485 , \34486 , \34487 , \34488 , \34489 , \34490 ,
         \34491 , \34492 , \34493 , \34494 , \34495 , \34496 , \34497 , \34498 , \34499 , \34500 ,
         \34501 , \34502 , \34503 , \34504 , \34505 , \34506 , \34507 , \34508 , \34509 , \34510 ,
         \34511 , \34512 , \34513 , \34514 , \34515 , \34516 , \34517 , \34518 , \34519 , \34520 ,
         \34521 , \34522 , \34523 , \34524 , \34525 , \34526 , \34527 , \34528 , \34529 , \34530 ,
         \34531 , \34532 , \34533 , \34534 , \34535 , \34536 , \34537 , \34538 , \34539 , \34540 ,
         \34541 , \34542 , \34543 , \34544 , \34545 , \34546 , \34547 , \34548 , \34549 , \34550 ,
         \34551 , \34552 , \34553 , \34554 , \34555 , \34556 , \34557 , \34558 , \34559 , \34560 ,
         \34561 , \34562 , \34563 , \34564 , \34565 , \34566 , \34567 , \34568 , \34569 , \34570 ,
         \34571 , \34572 , \34573 , \34574 , \34575 , \34576 , \34577 , \34578 , \34579 , \34580 ,
         \34581 , \34582 , \34583 , \34584 , \34585 , \34586 , \34587 , \34588 , \34589 , \34590 ,
         \34591 , \34592 , \34593 , \34594 , \34595 , \34596 , \34597 , \34598 , \34599 , \34600 ,
         \34601 , \34602 , \34603 , \34604 , \34605 , \34606 , \34607 , \34608 , \34609 , \34610 ,
         \34611 , \34612 , \34613 , \34614 , \34615 , \34616 , \34617 , \34618 , \34619 , \34620 ,
         \34621 , \34622 , \34623 , \34624 , \34625 , \34626 , \34627 , \34628 , \34629 , \34630 ,
         \34631 , \34632 , \34633 , \34634 , \34635 , \34636 , \34637 , \34638 , \34639 , \34640 ,
         \34641 , \34642 , \34643 , \34644 , \34645 , \34646 , \34647 , \34648 , \34649 , \34650 ,
         \34651 , \34652 , \34653 , \34654 , \34655 , \34656 , \34657 , \34658 , \34659 , \34660 ,
         \34661 , \34662 , \34663 , \34664 , \34665 , \34666 , \34667 , \34668 , \34669 , \34670 ,
         \34671 , \34672 , \34673 , \34674 , \34675 , \34676 , \34677 , \34678 , \34679 , \34680 ,
         \34681 , \34682 , \34683 , \34684 , \34685 , \34686 , \34687 , \34688 , \34689 , \34690 ,
         \34691 , \34692 , \34693 , \34694 , \34695 , \34696 , \34697 , \34698 , \34699 , \34700 ,
         \34701 , \34702 , \34703 , \34704 , \34705 , \34706 , \34707 , \34708 , \34709 , \34710 ,
         \34711 , \34712 , \34713 , \34714 , \34715 , \34716 , \34717 , \34718 , \34719 , \34720 ,
         \34721 , \34722 , \34723 , \34724 , \34725 , \34726 , \34727 , \34728 , \34729 , \34730 ,
         \34731 , \34732 , \34733 , \34734 , \34735 , \34736 , \34737 , \34738 , \34739 , \34740 ,
         \34741 , \34742 , \34743 , \34744 , \34745 , \34746 , \34747 , \34748 , \34749 , \34750 ,
         \34751 , \34752 , \34753 , \34754 , \34755 , \34756 , \34757 , \34758 , \34759 , \34760 ,
         \34761 , \34762 , \34763 , \34764 , \34765 , \34766 , \34767 , \34768 , \34769 , \34770 ,
         \34771 , \34772 , \34773 , \34774 , \34775 , \34776 , \34777 , \34778 , \34779 , \34780 ,
         \34781 , \34782 , \34783 , \34784 , \34785 , \34786 , \34787 , \34788 , \34789 , \34790 ,
         \34791 , \34792 , \34793 , \34794 , \34795 , \34796 , \34797 , \34798 , \34799 , \34800 ,
         \34801 , \34802 , \34803 , \34804 , \34805 , \34806 , \34807 , \34808 , \34809 , \34810 ,
         \34811 , \34812 , \34813 , \34814 , \34815 , \34816 , \34817 , \34818 , \34819 , \34820 ,
         \34821 , \34822 , \34823 , \34824 , \34825 , \34826 , \34827 , \34828 , \34829 , \34830 ,
         \34831 , \34832 , \34833 , \34834 , \34835 , \34836 , \34837 , \34838 , \34839 , \34840 ,
         \34841 , \34842 , \34843 , \34844 , \34845 , \34846 , \34847 , \34848 , \34849 , \34850 ,
         \34851 , \34852 , \34853 , \34854 , \34855 , \34856 , \34857 , \34858 , \34859 , \34860 ,
         \34861 , \34862 , \34863 , \34864 , \34865 , \34866 , \34867 , \34868 , \34869 , \34870 ,
         \34871 , \34872 , \34873 , \34874 , \34875 , \34876 , \34877 , \34878 , \34879 , \34880 ,
         \34881 , \34882 , \34883 , \34884 , \34885 , \34886 , \34887 , \34888 , \34889 , \34890 ,
         \34891 , \34892 , \34893 , \34894 , \34895 , \34896 , \34897 , \34898 , \34899 , \34900 ,
         \34901 , \34902 , \34903 , \34904 , \34905 , \34906 , \34907 , \34908 , \34909 , \34910 ,
         \34911 , \34912 , \34913 , \34914 , \34915 , \34916 , \34917 , \34918 , \34919 , \34920 ,
         \34921 , \34922 , \34923 , \34924 , \34925 , \34926 , \34927 , \34928 , \34929 , \34930 ,
         \34931 , \34932 , \34933 , \34934 , \34935 , \34936 , \34937 , \34938 , \34939 , \34940 ,
         \34941 , \34942 , \34943 , \34944 , \34945 , \34946 , \34947 , \34948 , \34949 , \34950 ,
         \34951 , \34952 , \34953 , \34954 , \34955 , \34956 , \34957 , \34958 , \34959 , \34960 ,
         \34961 , \34962 , \34963 , \34964 , \34965 , \34966 , \34967 , \34968 , \34969 , \34970 ,
         \34971 , \34972 , \34973 , \34974 , \34975 , \34976 , \34977 , \34978 , \34979 , \34980 ,
         \34981 , \34982 , \34983 , \34984 , \34985 , \34986 , \34987 , \34988 , \34989 , \34990 ,
         \34991 , \34992 , \34993 , \34994 , \34995 , \34996 , \34997 , \34998 , \34999 , \35000 ,
         \35001 , \35002 , \35003 , \35004 , \35005 , \35006 , \35007 , \35008 , \35009 , \35010 ,
         \35011 , \35012 , \35013 , \35014 , \35015 , \35016 , \35017 , \35018 , \35019 , \35020 ,
         \35021 , \35022 , \35023 , \35024 , \35025 , \35026 , \35027 , \35028 , \35029 , \35030 ,
         \35031 , \35032 , \35033 , \35034 , \35035 , \35036 , \35037 , \35038 , \35039 , \35040 ,
         \35041 , \35042 , \35043 , \35044 , \35045 , \35046 , \35047 , \35048 , \35049 , \35050 ,
         \35051 , \35052 , \35053 , \35054 , \35055 , \35056 , \35057 , \35058 , \35059 , \35060 ,
         \35061 , \35062 , \35063 , \35064 , \35065 , \35066 , \35067 , \35068 , \35069 , \35070 ,
         \35071 , \35072 , \35073 , \35074 , \35075 , \35076 , \35077 , \35078 , \35079 , \35080 ,
         \35081 , \35082 , \35083 , \35084 , \35085 , \35086 , \35087 , \35088 , \35089 , \35090 ,
         \35091 , \35092 , \35093 , \35094 , \35095 , \35096 , \35097 , \35098 , \35099 , \35100 ,
         \35101 , \35102 , \35103 , \35104 , \35105 , \35106 , \35107 , \35108 , \35109 , \35110 ,
         \35111 , \35112 , \35113 , \35114 , \35115 , \35116 , \35117 , \35118 , \35119 , \35120 ,
         \35121 , \35122 , \35123 , \35124 , \35125 , \35126 , \35127 , \35128 , \35129 , \35130 ,
         \35131 , \35132 , \35133 , \35134 , \35135 , \35136 , \35137 , \35138 , \35139 , \35140 ,
         \35141 , \35142 , \35143 , \35144 , \35145 , \35146 , \35147 , \35148 , \35149 , \35150 ,
         \35151 , \35152 , \35153 , \35154 , \35155 , \35156 , \35157 , \35158 , \35159 , \35160 ,
         \35161 , \35162 , \35163 , \35164 , \35165 , \35166 , \35167 , \35168 , \35169 , \35170 ,
         \35171 , \35172 , \35173 , \35174 , \35175 , \35176 , \35177 , \35178 , \35179 , \35180 ,
         \35181 , \35182 , \35183 , \35184 , \35185 , \35186 , \35187 , \35188 , \35189 , \35190 ,
         \35191 , \35192 , \35193 , \35194 , \35195 , \35196 , \35197 , \35198 , \35199 , \35200 ,
         \35201 , \35202 , \35203 , \35204 , \35205 , \35206 , \35207 , \35208 , \35209 , \35210 ,
         \35211 , \35212 , \35213 , \35214 , \35215 , \35216 , \35217 , \35218 , \35219 , \35220 ,
         \35221 , \35222 , \35223 , \35224 , \35225 , \35226 , \35227 , \35228 , \35229 , \35230 ,
         \35231 , \35232 , \35233 , \35234 , \35235 , \35236 , \35237 , \35238 , \35239 , \35240 ,
         \35241 , \35242 , \35243 , \35244 , \35245 , \35246 , \35247 , \35248 , \35249 , \35250 ,
         \35251 , \35252 , \35253 , \35254 , \35255 , \35256 , \35257 , \35258 , \35259 , \35260 ,
         \35261 , \35262 , \35263 , \35264 , \35265 , \35266 , \35267 , \35268 , \35269 , \35270 ,
         \35271 , \35272 , \35273 , \35274 , \35275 , \35276 , \35277 , \35278 , \35279 , \35280 ,
         \35281 , \35282 , \35283 , \35284 , \35285 , \35286 , \35287 , \35288 , \35289 , \35290 ,
         \35291 , \35292 , \35293 , \35294 , \35295 , \35296 , \35297 , \35298 , \35299 , \35300 ,
         \35301 , \35302 , \35303 , \35304 , \35305 , \35306 , \35307 , \35308 , \35309 , \35310 ,
         \35311 , \35312 , \35313 , \35314 , \35315 , \35316 , \35317 , \35318 , \35319 , \35320 ,
         \35321 , \35322 , \35323 , \35324 , \35325 , \35326 , \35327 , \35328 , \35329 , \35330 ,
         \35331 , \35332 , \35333 , \35334 , \35335 , \35336 , \35337 , \35338 , \35339 , \35340 ,
         \35341 , \35342 , \35343 , \35344 , \35345 , \35346 , \35347 , \35348 , \35349 , \35350 ,
         \35351 , \35352 , \35353 , \35354 , \35355 , \35356 , \35357 , \35358 , \35359 , \35360 ,
         \35361 , \35362 , \35363 , \35364 , \35365 , \35366 , \35367 , \35368 , \35369 , \35370 ,
         \35371 , \35372 , \35373 , \35374 , \35375 , \35376 , \35377 , \35378 , \35379 , \35380 ,
         \35381 , \35382 , \35383 , \35384 , \35385 , \35386 , \35387 , \35388 , \35389 , \35390 ,
         \35391 , \35392 , \35393 , \35394 , \35395 , \35396 , \35397 , \35398 , \35399 , \35400 ,
         \35401 , \35402 , \35403 , \35404 , \35405 , \35406 , \35407 , \35408 , \35409 , \35410 ,
         \35411 , \35412 , \35413 , \35414 , \35415 , \35416 , \35417 , \35418 , \35419 , \35420 ,
         \35421 , \35422 , \35423 , \35424 , \35425 , \35426 , \35427 , \35428 , \35429 , \35430 ,
         \35431 , \35432 , \35433 , \35434 , \35435 , \35436 , \35437 , \35438 , \35439 , \35440 ,
         \35441 , \35442 , \35443 , \35444 , \35445 , \35446 , \35447 , \35448 , \35449 , \35450 ,
         \35451 , \35452 , \35453 , \35454 , \35455 , \35456 , \35457 , \35458 , \35459 , \35460 ,
         \35461 , \35462 , \35463 , \35464 , \35465 , \35466 , \35467 , \35468 , \35469 , \35470 ,
         \35471 , \35472 , \35473 , \35474 , \35475 , \35476 , \35477 , \35478 , \35479 , \35480 ,
         \35481 , \35482 , \35483 , \35484 , \35485 , \35486 , \35487 , \35488 , \35489 , \35490 ,
         \35491 , \35492 , \35493 , \35494 , \35495 , \35496 , \35497 , \35498 , \35499 , \35500 ,
         \35501 , \35502 , \35503 , \35504 , \35505 , \35506 , \35507 , \35508 , \35509 , \35510 ,
         \35511 , \35512 , \35513 , \35514 , \35515 , \35516 , \35517 , \35518 , \35519 , \35520 ,
         \35521 , \35522 , \35523 , \35524 , \35525 , \35526 , \35527 , \35528 , \35529 , \35530 ,
         \35531 , \35532 , \35533 , \35534 , \35535 , \35536 , \35537 , \35538 , \35539 , \35540 ,
         \35541 , \35542 , \35543 , \35544 , \35545 , \35546 , \35547 , \35548 , \35549 , \35550 ,
         \35551 , \35552 , \35553 , \35554 , \35555 , \35556 , \35557 , \35558 , \35559 , \35560 ,
         \35561 , \35562 , \35563 , \35564 , \35565 , \35566 , \35567 , \35568 , \35569 , \35570 ,
         \35571 , \35572 , \35573 , \35574 , \35575 , \35576 , \35577 , \35578 , \35579 , \35580 ,
         \35581 , \35582 , \35583 , \35584 , \35585 , \35586 , \35587 , \35588 , \35589 , \35590 ,
         \35591 , \35592 , \35593 , \35594 , \35595 , \35596 , \35597 , \35598 , \35599 , \35600 ,
         \35601 , \35602 , \35603 , \35604 , \35605 , \35606 , \35607 , \35608 , \35609 , \35610 ,
         \35611 , \35612 , \35613 , \35614 , \35615 , \35616 , \35617 , \35618 , \35619 , \35620 ,
         \35621 , \35622 , \35623 , \35624 , \35625 , \35626 , \35627 , \35628 , \35629 , \35630 ,
         \35631 , \35632 , \35633 , \35634 , \35635 , \35636 , \35637 , \35638 , \35639 , \35640 ,
         \35641 , \35642 , \35643 , \35644 , \35645 , \35646 , \35647 , \35648 , \35649 , \35650 ,
         \35651 , \35652 , \35653 , \35654 , \35655 , \35656 , \35657 , \35658 , \35659 , \35660 ,
         \35661 , \35662 , \35663 , \35664 , \35665 , \35666 , \35667 , \35668 , \35669 , \35670 ,
         \35671 , \35672 , \35673 , \35674 , \35675 , \35676 , \35677 , \35678 , \35679 , \35680 ,
         \35681 , \35682 , \35683 , \35684 , \35685 , \35686 , \35687 , \35688 , \35689 , \35690 ,
         \35691 , \35692 , \35693 , \35694 , \35695 , \35696 , \35697 , \35698 , \35699 , \35700 ,
         \35701 , \35702 , \35703 , \35704 , \35705 , \35706 , \35707 , \35708 , \35709 , \35710 ,
         \35711 , \35712 , \35713 , \35714 , \35715 , \35716 , \35717 , \35718 , \35719 , \35720 ,
         \35721 , \35722 , \35723 , \35724 , \35725 , \35726 , \35727 , \35728 , \35729 , \35730 ,
         \35731 , \35732 , \35733 , \35734 , \35735 , \35736 , \35737 , \35738 , \35739 , \35740 ,
         \35741 , \35742 , \35743 , \35744 , \35745 , \35746 , \35747 , \35748 , \35749 , \35750 ,
         \35751 , \35752 , \35753 , \35754 , \35755 , \35756 , \35757 , \35758 , \35759 , \35760 ,
         \35761 , \35762 , \35763 , \35764 , \35765 , \35766 , \35767 , \35768 , \35769 , \35770 ,
         \35771 , \35772 , \35773 , \35774 , \35775 , \35776 , \35777 , \35778 , \35779 , \35780 ,
         \35781 , \35782 , \35783 , \35784 , \35785 , \35786 , \35787 , \35788 , \35789 , \35790 ,
         \35791 , \35792 , \35793 , \35794 , \35795 , \35796 , \35797 , \35798 , \35799 , \35800 ,
         \35801 , \35802 , \35803 , \35804 , \35805 , \35806 , \35807 , \35808 , \35809 , \35810 ,
         \35811 , \35812 , \35813 , \35814 , \35815 , \35816 , \35817 , \35818 , \35819 , \35820 ,
         \35821 , \35822 , \35823 , \35824 , \35825 , \35826 , \35827 , \35828 , \35829 , \35830 ,
         \35831 , \35832 , \35833 , \35834 , \35835 , \35836 , \35837 , \35838 , \35839 , \35840 ,
         \35841 , \35842 , \35843 , \35844 , \35845 , \35846 , \35847 , \35848 , \35849 , \35850 ,
         \35851 , \35852 , \35853 , \35854 , \35855 , \35856 , \35857 , \35858 , \35859 , \35860 ,
         \35861 , \35862 , \35863 , \35864 , \35865 , \35866 , \35867 , \35868 , \35869 , \35870 ,
         \35871 , \35872 , \35873 , \35874 , \35875 , \35876 , \35877 , \35878 , \35879 , \35880 ,
         \35881 , \35882 , \35883 , \35884 , \35885 , \35886 , \35887 , \35888 , \35889 , \35890 ,
         \35891 , \35892 , \35893 , \35894 , \35895 , \35896 , \35897 , \35898 , \35899 , \35900 ,
         \35901 , \35902 , \35903 , \35904 , \35905 , \35906 , \35907 , \35908 , \35909 , \35910 ,
         \35911 , \35912 , \35913 , \35914 , \35915 , \35916 , \35917 , \35918 , \35919 , \35920 ,
         \35921 , \35922 , \35923 , \35924 , \35925 , \35926 , \35927 , \35928 , \35929 , \35930 ,
         \35931 , \35932 , \35933 , \35934 , \35935 , \35936 , \35937 , \35938 , \35939 , \35940 ,
         \35941 , \35942 , \35943 , \35944 , \35945 , \35946 , \35947 , \35948 , \35949 , \35950 ,
         \35951 , \35952 , \35953 , \35954 , \35955 , \35956 , \35957 , \35958 , \35959 , \35960 ,
         \35961 , \35962 , \35963 , \35964 , \35965 , \35966 , \35967 , \35968 , \35969 , \35970 ,
         \35971 , \35972 , \35973 , \35974 , \35975 , \35976 , \35977 , \35978 , \35979 , \35980 ,
         \35981 , \35982 , \35983 , \35984 , \35985 , \35986 , \35987 , \35988 , \35989 , \35990 ,
         \35991 , \35992 , \35993 , \35994 , \35995 , \35996 , \35997 , \35998 , \35999 , \36000 ,
         \36001 , \36002 , \36003 , \36004 , \36005 , \36006 , \36007 , \36008 , \36009 , \36010 ,
         \36011 , \36012 , \36013 , \36014 , \36015 , \36016 , \36017 , \36018 , \36019 , \36020 ,
         \36021 , \36022 , \36023 , \36024 , \36025 , \36026 , \36027 , \36028 , \36029 , \36030 ,
         \36031 , \36032 , \36033 , \36034 , \36035 , \36036 , \36037 , \36038 , \36039 , \36040 ,
         \36041 , \36042 , \36043 , \36044 , \36045 , \36046 , \36047 , \36048 , \36049 , \36050 ,
         \36051 , \36052 , \36053 , \36054 , \36055 , \36056 , \36057 , \36058 , \36059 , \36060 ,
         \36061 , \36062 , \36063 , \36064 , \36065 , \36066 , \36067 , \36068 , \36069 , \36070 ,
         \36071 , \36072 , \36073 , \36074 , \36075 , \36076 , \36077 , \36078 , \36079 , \36080 ,
         \36081 , \36082 , \36083 , \36084 , \36085 , \36086 , \36087 , \36088 , \36089 , \36090 ,
         \36091 , \36092 , \36093 , \36094 , \36095 , \36096 , \36097 , \36098 , \36099 , \36100 ,
         \36101 , \36102 , \36103 , \36104 , \36105 , \36106 , \36107 , \36108 , \36109 , \36110 ,
         \36111 , \36112 , \36113 , \36114 , \36115 , \36116 , \36117 , \36118 , \36119 , \36120 ,
         \36121 , \36122 , \36123 , \36124 , \36125 , \36126 , \36127 , \36128 , \36129 , \36130 ,
         \36131 , \36132 , \36133 , \36134 , \36135 , \36136 , \36137 , \36138 , \36139 , \36140 ,
         \36141 , \36142 , \36143 , \36144 , \36145 , \36146 , \36147 , \36148 , \36149 , \36150 ,
         \36151 , \36152 , \36153 , \36154 , \36155 , \36156 , \36157 , \36158 , \36159 , \36160 ,
         \36161 , \36162 , \36163 , \36164 , \36165 , \36166 , \36167 , \36168 , \36169 , \36170 ,
         \36171 , \36172 , \36173 , \36174 , \36175 , \36176 , \36177 , \36178 , \36179 , \36180 ,
         \36181 , \36182 , \36183 , \36184 , \36185 , \36186 , \36187 , \36188 , \36189 , \36190 ,
         \36191 , \36192 , \36193 , \36194 , \36195 , \36196 , \36197 , \36198 , \36199 , \36200 ,
         \36201 , \36202 , \36203 , \36204 , \36205 , \36206 , \36207 , \36208 , \36209 , \36210 ,
         \36211 , \36212 , \36213 , \36214 , \36215 , \36216 , \36217 , \36218 , \36219 , \36220 ,
         \36221 , \36222 , \36223 , \36224 , \36225 , \36226 , \36227 , \36228 , \36229 , \36230 ,
         \36231 , \36232 , \36233 , \36234 , \36235 , \36236 , \36237 , \36238 , \36239 , \36240 ,
         \36241 , \36242 , \36243 , \36244 , \36245 , \36246 , \36247 , \36248 , \36249 , \36250 ,
         \36251 , \36252 , \36253 , \36254 , \36255 , \36256 , \36257 , \36258 , \36259 , \36260 ,
         \36261 , \36262 , \36263 , \36264 , \36265 , \36266 , \36267 , \36268 , \36269 , \36270 ,
         \36271 , \36272 , \36273 , \36274 , \36275 , \36276 , \36277 , \36278 , \36279 , \36280 ,
         \36281 , \36282 , \36283 , \36284 , \36285 , \36286 , \36287 , \36288 , \36289 , \36290 ,
         \36291 , \36292 , \36293 , \36294 , \36295 , \36296 , \36297 , \36298 , \36299 , \36300 ,
         \36301 , \36302 , \36303 , \36304 , \36305 , \36306 , \36307 , \36308 , \36309 , \36310 ,
         \36311 , \36312 , \36313 , \36314 , \36315 , \36316 , \36317 , \36318 , \36319 , \36320 ,
         \36321 , \36322 , \36323 , \36324 , \36325 , \36326 , \36327 , \36328 , \36329 , \36330 ,
         \36331 , \36332 , \36333 , \36334 , \36335 , \36336 , \36337 , \36338 , \36339 , \36340 ,
         \36341 , \36342 , \36343 , \36344 , \36345 , \36346 , \36347 , \36348 , \36349 , \36350 ,
         \36351 , \36352 , \36353 , \36354 , \36355 , \36356 , \36357 , \36358 , \36359 , \36360 ,
         \36361 , \36362 , \36363 , \36364 , \36365 , \36366 , \36367 , \36368 , \36369 , \36370 ,
         \36371 , \36372 , \36373 , \36374 , \36375 , \36376 , \36377 , \36378 , \36379 , \36380 ,
         \36381 , \36382 , \36383 , \36384 , \36385 , \36386 , \36387 , \36388 , \36389 , \36390 ,
         \36391 , \36392 , \36393 , \36394 , \36395 , \36396 , \36397 , \36398 , \36399 , \36400 ,
         \36401 , \36402 , \36403 , \36404 , \36405 , \36406 , \36407 , \36408 , \36409 , \36410 ,
         \36411 , \36412 , \36413 , \36414 , \36415 , \36416 , \36417 , \36418 , \36419 , \36420 ,
         \36421 , \36422 , \36423 , \36424 , \36425 , \36426 , \36427 , \36428 , \36429 , \36430 ,
         \36431 , \36432 , \36433 , \36434 , \36435 , \36436 , \36437 , \36438 , \36439 , \36440 ,
         \36441 , \36442 , \36443 , \36444 , \36445 , \36446 , \36447 , \36448 , \36449 , \36450 ,
         \36451 , \36452 , \36453 , \36454 , \36455 , \36456 , \36457 , \36458 , \36459 , \36460 ,
         \36461 , \36462 , \36463 , \36464 , \36465 , \36466 , \36467 , \36468 , \36469 , \36470 ,
         \36471 , \36472 , \36473 , \36474 , \36475 , \36476 , \36477 , \36478 , \36479 , \36480 ,
         \36481 , \36482 , \36483 , \36484 , \36485 , \36486 , \36487 , \36488 , \36489 , \36490 ,
         \36491 , \36492 , \36493 , \36494 , \36495 , \36496 , \36497 , \36498 , \36499 , \36500 ,
         \36501 , \36502 , \36503 , \36504 , \36505 , \36506 , \36507 , \36508 , \36509 , \36510 ,
         \36511 , \36512 , \36513 , \36514 , \36515 , \36516 , \36517 , \36518 , \36519 , \36520 ,
         \36521 , \36522 , \36523 , \36524 , \36525 , \36526 , \36527 , \36528 , \36529 , \36530 ,
         \36531 , \36532 , \36533 , \36534 , \36535 , \36536 , \36537 , \36538 , \36539 , \36540 ,
         \36541 , \36542 , \36543 , \36544 , \36545 , \36546 , \36547 , \36548 , \36549 , \36550 ,
         \36551 , \36552 , \36553 , \36554 , \36555 , \36556 , \36557 , \36558 , \36559 , \36560 ,
         \36561 , \36562 , \36563 , \36564 , \36565 , \36566 , \36567 , \36568 , \36569 , \36570 ,
         \36571 , \36572 , \36573 , \36574 , \36575 , \36576 , \36577 , \36578 , \36579 , \36580 ,
         \36581 , \36582 , \36583 , \36584 , \36585 , \36586 , \36587 , \36588 , \36589 , \36590 ,
         \36591 , \36592 , \36593 , \36594 , \36595 , \36596 , \36597 , \36598 , \36599 , \36600 ,
         \36601 , \36602 , \36603 , \36604 , \36605 , \36606 , \36607 , \36608 , \36609 , \36610 ,
         \36611 , \36612 , \36613 , \36614 , \36615 , \36616 , \36617 , \36618 , \36619 , \36620 ,
         \36621 , \36622 , \36623 , \36624 , \36625 , \36626 , \36627 , \36628 , \36629 , \36630 ,
         \36631 , \36632 , \36633 , \36634 , \36635 , \36636 , \36637 , \36638 , \36639 , \36640 ,
         \36641 , \36642 , \36643 , \36644 , \36645 , \36646 , \36647 , \36648 , \36649 , \36650 ,
         \36651 , \36652 , \36653 , \36654 , \36655 , \36656 , \36657 , \36658 , \36659 , \36660 ,
         \36661 , \36662 , \36663 , \36664 , \36665 , \36666 , \36667 , \36668 , \36669 , \36670 ,
         \36671 , \36672 , \36673 , \36674 , \36675 , \36676 , \36677 , \36678 , \36679 , \36680 ,
         \36681 , \36682 , \36683 , \36684 , \36685 , \36686 , \36687 , \36688 , \36689 , \36690 ,
         \36691 , \36692 , \36693 , \36694 , \36695 , \36696 , \36697 , \36698 , \36699 , \36700 ,
         \36701 , \36702 , \36703 , \36704 , \36705 , \36706 , \36707 , \36708 , \36709 , \36710 ,
         \36711 , \36712 , \36713 , \36714 , \36715 , \36716 , \36717 , \36718 , \36719 , \36720 ,
         \36721 , \36722 , \36723 , \36724 , \36725 , \36726 , \36727 , \36728 , \36729 , \36730 ,
         \36731 , \36732 , \36733 , \36734 , \36735 , \36736 , \36737 , \36738 , \36739 , \36740 ,
         \36741 , \36742 , \36743 , \36744 , \36745 , \36746 , \36747 , \36748 , \36749 , \36750 ,
         \36751 , \36752 , \36753 , \36754 , \36755 , \36756 , \36757 , \36758 , \36759 , \36760 ,
         \36761 , \36762 , \36763 , \36764 , \36765 , \36766 , \36767 , \36768 , \36769 , \36770 ,
         \36771 , \36772 , \36773 , \36774 , \36775 , \36776 , \36777 , \36778 , \36779 , \36780 ,
         \36781 , \36782 , \36783 , \36784 , \36785 , \36786 , \36787 , \36788 , \36789 , \36790 ,
         \36791 , \36792 , \36793 , \36794 , \36795 , \36796 , \36797 , \36798 , \36799 , \36800 ,
         \36801 , \36802 , \36803 , \36804 , \36805 , \36806 , \36807 , \36808 , \36809 , \36810 ,
         \36811 , \36812 , \36813 , \36814 , \36815 , \36816 , \36817 , \36818 , \36819 , \36820 ,
         \36821 , \36822 , \36823 , \36824 , \36825 , \36826 , \36827 , \36828 , \36829 , \36830 ,
         \36831 , \36832 , \36833 , \36834 , \36835 , \36836 , \36837 , \36838 , \36839 , \36840 ,
         \36841 , \36842 , \36843 , \36844 , \36845 , \36846 , \36847 , \36848 , \36849 , \36850 ,
         \36851 , \36852 , \36853 , \36854 , \36855 , \36856 , \36857 , \36858 , \36859 , \36860 ,
         \36861 , \36862 , \36863 , \36864 , \36865 , \36866 , \36867 , \36868 , \36869 , \36870 ,
         \36871 , \36872 , \36873 , \36874 , \36875 , \36876 , \36877 , \36878 , \36879 , \36880 ,
         \36881 , \36882 , \36883 , \36884 , \36885 , \36886 , \36887 , \36888 , \36889 , \36890 ,
         \36891 , \36892 , \36893 , \36894 , \36895 , \36896 , \36897 , \36898 , \36899 , \36900 ,
         \36901 , \36902 , \36903 , \36904 , \36905 , \36906 , \36907 , \36908 , \36909 , \36910 ,
         \36911 , \36912 , \36913 , \36914 , \36915 , \36916 , \36917 , \36918 , \36919 , \36920 ,
         \36921 , \36922 , \36923 , \36924 , \36925 , \36926 , \36927 , \36928 , \36929 , \36930 ,
         \36931 , \36932 , \36933 , \36934 , \36935 , \36936 , \36937 , \36938 , \36939 , \36940 ,
         \36941 , \36942 , \36943 , \36944 , \36945 , \36946 , \36947 , \36948 , \36949 , \36950 ,
         \36951 , \36952 , \36953 , \36954 , \36955 , \36956 , \36957 , \36958 , \36959 , \36960 ,
         \36961 , \36962 , \36963 , \36964 , \36965 , \36966 , \36967 , \36968 , \36969 , \36970 ,
         \36971 , \36972 , \36973 , \36974 , \36975 , \36976 , \36977 , \36978 , \36979 , \36980 ,
         \36981 , \36982 , \36983 , \36984 , \36985 , \36986 , \36987 , \36988 , \36989 , \36990 ,
         \36991 , \36992 , \36993 , \36994 , \36995 , \36996 , \36997 , \36998 , \36999 , \37000 ,
         \37001 , \37002 , \37003 , \37004 , \37005 , \37006 , \37007 , \37008 , \37009 , \37010 ,
         \37011 , \37012 , \37013 , \37014 , \37015 , \37016 , \37017 , \37018 , \37019 , \37020 ,
         \37021 , \37022 , \37023 , \37024 , \37025 , \37026 , \37027 , \37028 , \37029 , \37030 ,
         \37031 , \37032 , \37033 , \37034 , \37035 , \37036 , \37037 , \37038 , \37039 , \37040 ,
         \37041 , \37042 , \37043 , \37044 , \37045 , \37046 , \37047 , \37048 , \37049 , \37050 ,
         \37051 , \37052 , \37053 , \37054 , \37055 , \37056 , \37057 , \37058 , \37059 , \37060 ,
         \37061 , \37062 , \37063 , \37064 , \37065 , \37066 , \37067 , \37068 , \37069 , \37070 ,
         \37071 , \37072 , \37073 , \37074 , \37075 , \37076 , \37077 , \37078 , \37079 , \37080 ,
         \37081 , \37082 , \37083 , \37084 , \37085 , \37086 , \37087 , \37088 , \37089 , \37090 ,
         \37091 , \37092 , \37093 , \37094 , \37095 , \37096 , \37097 , \37098 , \37099 , \37100 ,
         \37101 , \37102 , \37103 , \37104 , \37105 , \37106 , \37107 , \37108 , \37109 , \37110 ,
         \37111 , \37112 , \37113 , \37114 , \37115 , \37116 , \37117 , \37118 , \37119 , \37120 ,
         \37121 , \37122 , \37123 , \37124 , \37125 , \37126 , \37127 , \37128 , \37129 , \37130 ,
         \37131 , \37132 , \37133 , \37134 , \37135 , \37136 , \37137 , \37138 , \37139 , \37140 ,
         \37141 , \37142 , \37143 , \37144 , \37145 , \37146 , \37147 , \37148 , \37149 , \37150 ,
         \37151 , \37152 , \37153 , \37154 , \37155 , \37156 , \37157 , \37158 , \37159 , \37160 ,
         \37161 , \37162 , \37163 , \37164 , \37165 , \37166 , \37167 , \37168 , \37169 , \37170 ,
         \37171 , \37172 , \37173 , \37174 , \37175 , \37176 , \37177 , \37178 , \37179 , \37180 ,
         \37181 , \37182 , \37183 , \37184 , \37185 , \37186 , \37187 , \37188 , \37189 , \37190 ,
         \37191 , \37192 , \37193 , \37194 , \37195 , \37196 , \37197 , \37198 , \37199 , \37200 ,
         \37201 , \37202 , \37203 , \37204 , \37205 , \37206 , \37207 , \37208 , \37209 , \37210 ,
         \37211 , \37212 , \37213 , \37214 , \37215 , \37216 , \37217 , \37218 , \37219 , \37220 ,
         \37221 , \37222 , \37223 , \37224 , \37225 , \37226 , \37227 , \37228 , \37229 , \37230 ,
         \37231 , \37232 , \37233 , \37234 , \37235 , \37236 , \37237 , \37238 , \37239 , \37240 ,
         \37241 , \37242 , \37243 , \37244 , \37245 , \37246 , \37247 , \37248 , \37249 , \37250 ,
         \37251 , \37252 , \37253 , \37254 , \37255 , \37256 , \37257 , \37258 , \37259 , \37260 ,
         \37261 , \37262 , \37263 , \37264 , \37265 , \37266 , \37267 , \37268 , \37269 , \37270 ,
         \37271 , \37272 , \37273 , \37274 , \37275 , \37276 , \37277 , \37278 , \37279 , \37280 ,
         \37281 , \37282 , \37283 , \37284 , \37285 , \37286 , \37287 , \37288 , \37289 , \37290 ,
         \37291 , \37292 , \37293 , \37294 , \37295 , \37296 , \37297 , \37298 , \37299 , \37300 ,
         \37301 , \37302 , \37303 , \37304 , \37305 , \37306 , \37307 , \37308 , \37309 , \37310 ,
         \37311 , \37312 , \37313 , \37314 , \37315 , \37316 , \37317 , \37318 , \37319 , \37320 ,
         \37321 , \37322 , \37323 , \37324 , \37325 , \37326 , \37327 , \37328 , \37329 , \37330 ,
         \37331 , \37332 , \37333 , \37334 , \37335 , \37336 , \37337 , \37338 , \37339 , \37340 ,
         \37341 , \37342 , \37343 , \37344 , \37345 , \37346 , \37347 , \37348 , \37349 , \37350 ,
         \37351 , \37352 , \37353 , \37354 , \37355 , \37356 , \37357 , \37358 , \37359 , \37360 ,
         \37361 , \37362 , \37363 , \37364 , \37365 , \37366 , \37367 , \37368 , \37369 , \37370 ,
         \37371 , \37372 , \37373 , \37374 , \37375 , \37376 , \37377 , \37378 , \37379 , \37380 ,
         \37381 , \37382 , \37383 , \37384 , \37385 , \37386 , \37387 , \37388 , \37389 , \37390 ,
         \37391 , \37392 , \37393 , \37394 , \37395 , \37396 , \37397 , \37398 , \37399 , \37400 ,
         \37401 , \37402 , \37403 , \37404 , \37405 , \37406 , \37407 , \37408 , \37409 , \37410 ,
         \37411 , \37412 , \37413 , \37414 , \37415 , \37416 , \37417 , \37418 , \37419 , \37420 ,
         \37421 , \37422 , \37423 , \37424 , \37425 , \37426 , \37427 , \37428 , \37429 , \37430 ,
         \37431 , \37432 , \37433 , \37434 , \37435 , \37436 , \37437 , \37438 , \37439 , \37440 ,
         \37441 , \37442 , \37443 , \37444 , \37445 , \37446 , \37447 , \37448 , \37449 , \37450 ,
         \37451 , \37452 , \37453 , \37454 , \37455 , \37456 , \37457 , \37458 , \37459 , \37460 ,
         \37461 , \37462 , \37463 , \37464 , \37465 , \37466 , \37467 , \37468 , \37469 , \37470 ,
         \37471 , \37472 , \37473 , \37474 , \37475 , \37476 , \37477 , \37478 , \37479 , \37480 ,
         \37481 , \37482 , \37483 , \37484 , \37485 , \37486 , \37487 , \37488 , \37489 , \37490 ,
         \37491 , \37492 , \37493 , \37494 , \37495 , \37496 , \37497 , \37498 , \37499 , \37500 ,
         \37501 , \37502 , \37503 , \37504 , \37505 , \37506 , \37507 , \37508 , \37509 , \37510 ,
         \37511 , \37512 , \37513 , \37514 , \37515 , \37516 , \37517 , \37518 , \37519 , \37520 ,
         \37521 , \37522 , \37523 , \37524 , \37525 , \37526 , \37527 , \37528 , \37529 , \37530 ,
         \37531 , \37532 , \37533 , \37534 , \37535 , \37536 , \37537 , \37538 , \37539 , \37540 ,
         \37541 , \37542 , \37543 , \37544 , \37545 , \37546 , \37547 , \37548 , \37549 , \37550 ,
         \37551 , \37552 , \37553 , \37554 , \37555 , \37556 , \37557 , \37558 , \37559 , \37560 ,
         \37561 , \37562 , \37563 , \37564 , \37565 , \37566 , \37567 , \37568 , \37569 , \37570 ,
         \37571 , \37572 , \37573 , \37574 , \37575 , \37576 , \37577 , \37578 , \37579 , \37580 ,
         \37581 , \37582 , \37583 , \37584 , \37585 , \37586 , \37587 , \37588 , \37589 , \37590 ,
         \37591 , \37592 , \37593 , \37594 , \37595 , \37596 , \37597 , \37598 , \37599 , \37600 ,
         \37601 , \37602 , \37603 , \37604 , \37605 , \37606 , \37607 , \37608 , \37609 , \37610 ,
         \37611 , \37612 , \37613 , \37614 , \37615 , \37616 , \37617 , \37618 , \37619 , \37620 ,
         \37621 , \37622 , \37623 , \37624 , \37625 , \37626 , \37627 , \37628 , \37629 , \37630 ,
         \37631 , \37632 , \37633 , \37634 , \37635 , \37636 , \37637 , \37638 , \37639 , \37640 ,
         \37641 , \37642 , \37643 , \37644 , \37645 , \37646 , \37647 , \37648 , \37649 , \37650 ,
         \37651 , \37652 , \37653 , \37654 , \37655 , \37656 , \37657 , \37658 , \37659 , \37660 ,
         \37661 , \37662 , \37663 , \37664 , \37665 , \37666 , \37667 , \37668 , \37669 , \37670 ,
         \37671 , \37672 , \37673 , \37674 , \37675 , \37676 , \37677 , \37678 , \37679 , \37680 ,
         \37681 , \37682 , \37683 , \37684 , \37685 , \37686 , \37687 , \37688 , \37689 , \37690 ,
         \37691 , \37692 , \37693 , \37694 , \37695 , \37696 , \37697 , \37698 , \37699 , \37700 ,
         \37701 , \37702 , \37703 , \37704 , \37705 , \37706 , \37707 , \37708 , \37709 , \37710 ,
         \37711 , \37712 , \37713 , \37714 , \37715 , \37716 , \37717 , \37718 , \37719 , \37720 ,
         \37721 , \37722 , \37723 , \37724 , \37725 , \37726 , \37727 , \37728 , \37729 , \37730 ,
         \37731 , \37732 , \37733 , \37734 , \37735 , \37736 , \37737 , \37738 , \37739 , \37740 ,
         \37741 , \37742 , \37743 , \37744 , \37745 , \37746 , \37747 , \37748 , \37749 , \37750 ,
         \37751 , \37752 , \37753 , \37754 , \37755 , \37756 , \37757 , \37758 , \37759 , \37760 ,
         \37761 , \37762 , \37763 , \37764 , \37765 , \37766 , \37767 , \37768 , \37769 , \37770 ,
         \37771 , \37772 , \37773 , \37774 , \37775 , \37776 , \37777 , \37778 , \37779 , \37780 ,
         \37781 , \37782 , \37783 , \37784 , \37785 , \37786 , \37787 , \37788 , \37789 , \37790 ,
         \37791 , \37792 , \37793 , \37794 , \37795 , \37796 , \37797 , \37798 , \37799 , \37800 ,
         \37801 , \37802 , \37803 , \37804 , \37805 , \37806 , \37807 , \37808 , \37809 , \37810 ,
         \37811 , \37812 , \37813 , \37814 , \37815 , \37816 , \37817 , \37818 , \37819 , \37820 ,
         \37821 , \37822 , \37823 , \37824 , \37825 , \37826 , \37827 , \37828 , \37829 , \37830 ,
         \37831 , \37832 , \37833 , \37834 , \37835 , \37836 , \37837 , \37838 , \37839 , \37840 ,
         \37841 , \37842 , \37843 , \37844 , \37845 , \37846 , \37847 , \37848 , \37849 , \37850 ,
         \37851 , \37852 , \37853 , \37854 , \37855 , \37856 , \37857 , \37858 , \37859 , \37860 ,
         \37861 , \37862 , \37863 , \37864 , \37865 , \37866 , \37867 , \37868 , \37869 , \37870 ,
         \37871 , \37872 , \37873 , \37874 , \37875 , \37876 , \37877 , \37878 , \37879 , \37880 ,
         \37881 , \37882 , \37883 , \37884 , \37885 , \37886 , \37887 , \37888 , \37889 , \37890 ,
         \37891 , \37892 , \37893 , \37894 , \37895 , \37896 , \37897 , \37898 , \37899 , \37900 ,
         \37901 , \37902 , \37903 , \37904 , \37905 , \37906 , \37907 , \37908 , \37909 , \37910 ,
         \37911 , \37912 , \37913 , \37914 , \37915 , \37916 , \37917 , \37918 , \37919 , \37920 ,
         \37921 , \37922 , \37923 , \37924 , \37925 , \37926 , \37927 , \37928 , \37929 , \37930 ,
         \37931 , \37932 , \37933 , \37934 , \37935 , \37936 , \37937 , \37938 , \37939 , \37940 ,
         \37941 , \37942 , \37943 , \37944 , \37945 , \37946 , \37947 , \37948 , \37949 , \37950 ,
         \37951 , \37952 , \37953 , \37954 , \37955 , \37956 , \37957 , \37958 , \37959 , \37960 ,
         \37961 , \37962 , \37963 , \37964 , \37965 , \37966 , \37967 , \37968 , \37969 , \37970 ,
         \37971 , \37972 , \37973 , \37974 , \37975 , \37976 , \37977 , \37978 , \37979 , \37980 ,
         \37981 , \37982 , \37983 , \37984 , \37985 , \37986 , \37987 , \37988 , \37989 , \37990 ,
         \37991 , \37992 , \37993 , \37994 , \37995 , \37996 , \37997 , \37998 , \37999 , \38000 ,
         \38001 , \38002 , \38003 , \38004 , \38005 , \38006 , \38007 , \38008 , \38009 , \38010 ,
         \38011 , \38012 , \38013 , \38014 , \38015 , \38016 , \38017 , \38018 , \38019 , \38020 ,
         \38021 , \38022 , \38023 , \38024 , \38025 , \38026 , \38027 , \38028 , \38029 , \38030 ,
         \38031 , \38032 , \38033 , \38034 , \38035 , \38036 , \38037 , \38038 , \38039 , \38040 ,
         \38041 , \38042 , \38043 , \38044 , \38045 , \38046 , \38047 , \38048 , \38049 , \38050 ,
         \38051 , \38052 , \38053 , \38054 , \38055 , \38056 , \38057 , \38058 , \38059 , \38060 ,
         \38061 , \38062 , \38063 , \38064 , \38065 , \38066 , \38067 , \38068 , \38069 , \38070 ,
         \38071 , \38072 , \38073 , \38074 , \38075 , \38076 , \38077 , \38078 , \38079 , \38080 ,
         \38081 , \38082 , \38083 , \38084 , \38085 , \38086 , \38087 , \38088 , \38089 , \38090 ,
         \38091 , \38092 , \38093 , \38094 , \38095 , \38096 , \38097 , \38098 , \38099 , \38100 ,
         \38101 , \38102 , \38103 , \38104 , \38105 , \38106 , \38107 , \38108 , \38109 , \38110 ,
         \38111 , \38112 , \38113 , \38114 , \38115 , \38116 , \38117 , \38118 , \38119 , \38120 ,
         \38121 , \38122 , \38123 , \38124 , \38125 , \38126 , \38127 , \38128 , \38129 , \38130 ,
         \38131 , \38132 , \38133 , \38134 , \38135 , \38136 , \38137 , \38138 , \38139 , \38140 ,
         \38141 , \38142 , \38143 , \38144 , \38145 , \38146 , \38147 , \38148 , \38149 , \38150 ,
         \38151 , \38152 , \38153 , \38154 , \38155 , \38156 , \38157 , \38158 , \38159 , \38160 ,
         \38161 , \38162 , \38163 , \38164 , \38165 , \38166 , \38167 , \38168 , \38169 , \38170 ,
         \38171 , \38172 , \38173 , \38174 , \38175 , \38176 , \38177 , \38178 , \38179 , \38180 ,
         \38181 , \38182 , \38183 , \38184 , \38185 , \38186 , \38187 , \38188 , \38189 , \38190 ,
         \38191 , \38192 , \38193 , \38194 , \38195 , \38196 , \38197 , \38198 , \38199 , \38200 ,
         \38201 , \38202 , \38203 , \38204 , \38205 , \38206 , \38207 , \38208 , \38209 , \38210 ,
         \38211 , \38212 , \38213 , \38214 , \38215 , \38216 , \38217 , \38218 , \38219 , \38220 ,
         \38221 , \38222 , \38223 , \38224 , \38225 , \38226 , \38227 , \38228 , \38229 , \38230 ,
         \38231 , \38232 , \38233 , \38234 , \38235 , \38236 , \38237 , \38238 , \38239 , \38240 ,
         \38241 , \38242 , \38243 , \38244 , \38245 , \38246 , \38247 , \38248 , \38249 , \38250 ,
         \38251 , \38252 , \38253 , \38254 , \38255 , \38256 , \38257 , \38258 , \38259 , \38260 ,
         \38261 , \38262 , \38263 , \38264 , \38265 , \38266 , \38267 , \38268 , \38269 , \38270 ,
         \38271 , \38272 , \38273 , \38274 , \38275 , \38276 , \38277 , \38278 , \38279 , \38280 ,
         \38281 , \38282 , \38283 , \38284 , \38285 , \38286 , \38287 , \38288 , \38289 , \38290 ,
         \38291 , \38292 , \38293 , \38294 , \38295 , \38296 , \38297 , \38298 , \38299 , \38300 ,
         \38301 , \38302 , \38303 , \38304 , \38305 , \38306 , \38307 , \38308 , \38309 , \38310 ,
         \38311 , \38312 , \38313 , \38314 , \38315 , \38316 , \38317 , \38318 , \38319 , \38320 ,
         \38321 , \38322 , \38323 , \38324 , \38325 , \38326 , \38327 , \38328 , \38329 , \38330 ,
         \38331 , \38332 , \38333 , \38334 , \38335 , \38336 , \38337 , \38338 , \38339 , \38340 ,
         \38341 , \38342 , \38343 , \38344 , \38345 , \38346 , \38347 , \38348 , \38349 , \38350 ,
         \38351 , \38352 , \38353 , \38354 , \38355 , \38356 , \38357 , \38358 , \38359 , \38360 ,
         \38361 , \38362 , \38363 , \38364 , \38365 , \38366 , \38367 , \38368 , \38369 , \38370 ,
         \38371 , \38372 , \38373 , \38374 , \38375 , \38376 , \38377 , \38378 , \38379 , \38380 ,
         \38381 , \38382 , \38383 , \38384 , \38385 , \38386 , \38387 , \38388 , \38389 , \38390 ,
         \38391 , \38392 , \38393 , \38394 , \38395 , \38396 , \38397 , \38398 , \38399 , \38400 ,
         \38401 , \38402 , \38403 , \38404 , \38405 , \38406 , \38407 , \38408 , \38409 , \38410 ,
         \38411 , \38412 , \38413 , \38414 , \38415 , \38416 , \38417 , \38418 , \38419 , \38420 ,
         \38421 , \38422 , \38423 , \38424 , \38425 , \38426 , \38427 , \38428 , \38429 , \38430 ,
         \38431 , \38432 , \38433 , \38434 , \38435 , \38436 , \38437 , \38438 , \38439 , \38440 ,
         \38441 , \38442 , \38443 , \38444 , \38445 , \38446 , \38447 , \38448 , \38449 , \38450 ,
         \38451 , \38452 , \38453 , \38454 , \38455 , \38456 , \38457 , \38458 , \38459 , \38460 ,
         \38461 , \38462 , \38463 , \38464 , \38465 , \38466 , \38467 , \38468 , \38469 , \38470 ,
         \38471 , \38472 , \38473 , \38474 , \38475 , \38476 , \38477 , \38478 , \38479 , \38480 ,
         \38481 , \38482 , \38483 , \38484 , \38485 , \38486 , \38487 , \38488 , \38489 , \38490 ,
         \38491 , \38492 , \38493 , \38494 , \38495 , \38496 , \38497 , \38498 , \38499 , \38500 ,
         \38501 , \38502 , \38503 , \38504 , \38505 , \38506 , \38507 , \38508 , \38509 , \38510 ,
         \38511 , \38512 , \38513 , \38514 , \38515 , \38516 , \38517 , \38518 , \38519 , \38520 ,
         \38521 , \38522 , \38523 , \38524 , \38525 , \38526 , \38527 , \38528 , \38529 , \38530 ,
         \38531 , \38532 , \38533 , \38534 , \38535 , \38536 , \38537 , \38538 , \38539 , \38540 ,
         \38541 , \38542 , \38543 , \38544 , \38545 , \38546 , \38547 , \38548 , \38549 , \38550 ,
         \38551 , \38552 , \38553 , \38554 , \38555 , \38556 , \38557 , \38558 , \38559 , \38560 ,
         \38561 , \38562 , \38563 , \38564 , \38565 , \38566 , \38567 , \38568 , \38569 , \38570 ,
         \38571 , \38572 , \38573 , \38574 , \38575 , \38576 , \38577 , \38578 , \38579 , \38580 ,
         \38581 , \38582 , \38583 , \38584 , \38585 , \38586 , \38587 , \38588 , \38589 , \38590 ,
         \38591 , \38592 , \38593 , \38594 , \38595 , \38596 , \38597 , \38598 , \38599 , \38600 ,
         \38601 , \38602 , \38603 , \38604 , \38605 , \38606 , \38607 , \38608 , \38609 , \38610 ,
         \38611 , \38612 , \38613 , \38614 , \38615 , \38616 , \38617 , \38618 , \38619 , \38620 ,
         \38621 , \38622 , \38623 , \38624 , \38625 , \38626 , \38627 , \38628 , \38629 , \38630 ,
         \38631 , \38632 , \38633 , \38634 , \38635 , \38636 , \38637 , \38638 , \38639 , \38640 ,
         \38641 , \38642 , \38643 , \38644 , \38645 , \38646 , \38647 , \38648 , \38649 , \38650 ,
         \38651 , \38652 , \38653 , \38654 , \38655 , \38656 , \38657 , \38658 , \38659 , \38660 ,
         \38661 , \38662 , \38663 , \38664 , \38665 , \38666 , \38667 , \38668 , \38669 , \38670 ,
         \38671 , \38672 , \38673 , \38674 , \38675 , \38676 , \38677 , \38678 , \38679 , \38680 ,
         \38681 , \38682 , \38683 , \38684 , \38685 , \38686 , \38687 , \38688 , \38689 , \38690 ,
         \38691 , \38692 , \38693 , \38694 , \38695 , \38696 , \38697 , \38698 , \38699 , \38700 ,
         \38701 , \38702 , \38703 , \38704 , \38705 , \38706 , \38707 , \38708 , \38709 , \38710 ,
         \38711 , \38712 , \38713 , \38714 , \38715 , \38716 , \38717 , \38718 , \38719 , \38720 ,
         \38721 , \38722 , \38723 , \38724 , \38725 , \38726 , \38727 , \38728 , \38729 , \38730 ,
         \38731 , \38732 , \38733 , \38734 , \38735 , \38736 , \38737 , \38738 , \38739 , \38740 ,
         \38741 , \38742 , \38743 , \38744 , \38745 , \38746 , \38747 , \38748 , \38749 , \38750 ,
         \38751 , \38752 , \38753 , \38754 , \38755 , \38756 , \38757 , \38758 , \38759 , \38760 ,
         \38761 , \38762 , \38763 , \38764 , \38765 , \38766 , \38767 , \38768 , \38769 , \38770 ,
         \38771 , \38772 , \38773 , \38774 , \38775 , \38776 , \38777 , \38778 , \38779 , \38780 ,
         \38781 , \38782 , \38783 , \38784 , \38785 , \38786 , \38787 , \38788 , \38789 , \38790 ,
         \38791 , \38792 , \38793 , \38794 , \38795 , \38796 , \38797 , \38798 , \38799 , \38800 ,
         \38801 , \38802 , \38803 , \38804 , \38805 , \38806 , \38807 , \38808 , \38809 , \38810 ,
         \38811 , \38812 , \38813 , \38814 , \38815 , \38816 , \38817 , \38818 , \38819 , \38820 ,
         \38821 , \38822 , \38823 , \38824 , \38825 , \38826 , \38827 , \38828 , \38829 , \38830 ,
         \38831 , \38832 , \38833 , \38834 , \38835 , \38836 , \38837 , \38838 , \38839 , \38840 ,
         \38841 , \38842 , \38843 , \38844 , \38845 , \38846 , \38847 , \38848 , \38849 , \38850 ,
         \38851 , \38852 , \38853 , \38854 , \38855 , \38856 , \38857 , \38858 , \38859 , \38860 ,
         \38861 , \38862 , \38863 , \38864 , \38865 , \38866 , \38867 , \38868 , \38869 , \38870 ,
         \38871 , \38872 , \38873 , \38874 , \38875 , \38876 , \38877 , \38878 , \38879 , \38880 ,
         \38881 , \38882 , \38883 , \38884 , \38885 , \38886 , \38887 , \38888 , \38889 , \38890 ,
         \38891 , \38892 , \38893 , \38894 , \38895 , \38896 , \38897 , \38898 , \38899 , \38900 ,
         \38901 , \38902 , \38903 , \38904 , \38905 , \38906 , \38907 , \38908 , \38909 , \38910 ,
         \38911 , \38912 , \38913 , \38914 , \38915 , \38916 , \38917 , \38918 , \38919 , \38920 ,
         \38921 , \38922 , \38923 , \38924 , \38925 , \38926 , \38927 , \38928 , \38929 , \38930 ,
         \38931 , \38932 , \38933 , \38934 , \38935 , \38936 , \38937 , \38938 , \38939 , \38940 ,
         \38941 , \38942 , \38943 , \38944 , \38945 , \38946 , \38947 , \38948 , \38949 , \38950 ,
         \38951 , \38952 , \38953 , \38954 , \38955 , \38956 , \38957 , \38958 , \38959 , \38960 ,
         \38961 , \38962 , \38963 , \38964 , \38965 , \38966 , \38967 , \38968 , \38969 , \38970 ,
         \38971 , \38972 , \38973 , \38974 , \38975 , \38976 , \38977 , \38978 , \38979 , \38980 ,
         \38981 , \38982 , \38983 , \38984 , \38985 , \38986 , \38987 , \38988 , \38989 , \38990 ,
         \38991 , \38992 , \38993 , \38994 , \38995 , \38996 , \38997 , \38998 , \38999 , \39000 ,
         \39001 , \39002 , \39003 , \39004 , \39005 , \39006 , \39007 , \39008 , \39009 , \39010 ,
         \39011 , \39012 , \39013 , \39014 , \39015 , \39016 , \39017 , \39018 , \39019 , \39020 ,
         \39021 , \39022 , \39023 , \39024 , \39025 , \39026 , \39027 , \39028 , \39029 , \39030 ,
         \39031 , \39032 , \39033 , \39034 , \39035 , \39036 , \39037 , \39038 , \39039 , \39040 ,
         \39041 , \39042 , \39043 , \39044 , \39045 , \39046 , \39047 , \39048 , \39049 , \39050 ,
         \39051 , \39052 , \39053 , \39054 , \39055 , \39056 , \39057 , \39058 , \39059 , \39060 ,
         \39061 , \39062 , \39063 , \39064 , \39065 , \39066 , \39067 , \39068 , \39069 , \39070 ,
         \39071 , \39072 , \39073 , \39074 , \39075 , \39076 , \39077 , \39078 , \39079 , \39080 ,
         \39081 , \39082 , \39083 , \39084 , \39085 , \39086 , \39087 , \39088 , \39089 , \39090 ,
         \39091 , \39092 , \39093 , \39094 , \39095 , \39096 , \39097 , \39098 , \39099 , \39100 ,
         \39101 , \39102 , \39103 , \39104 , \39105 , \39106 , \39107 , \39108 , \39109 , \39110 ,
         \39111 , \39112 , \39113 , \39114 , \39115 , \39116 , \39117 , \39118 , \39119 , \39120 ,
         \39121 , \39122 , \39123 , \39124 , \39125 , \39126 , \39127 , \39128 , \39129 , \39130 ,
         \39131 , \39132 , \39133 , \39134 , \39135 , \39136 , \39137 , \39138 , \39139 , \39140 ,
         \39141 , \39142 , \39143 , \39144 , \39145 , \39146 , \39147 , \39148 , \39149 , \39150 ,
         \39151 , \39152 , \39153 , \39154 , \39155 , \39156 , \39157 , \39158 , \39159 , \39160 ,
         \39161 , \39162 , \39163 , \39164 , \39165 , \39166 , \39167 , \39168 , \39169 , \39170 ,
         \39171 , \39172 , \39173 , \39174 , \39175 , \39176 , \39177 , \39178 , \39179 , \39180 ,
         \39181 , \39182 , \39183 , \39184 , \39185 , \39186 , \39187 , \39188 , \39189 , \39190 ,
         \39191 , \39192 , \39193 , \39194 , \39195 , \39196 , \39197 , \39198 , \39199 , \39200 ,
         \39201 , \39202 , \39203 , \39204 , \39205 , \39206 , \39207 , \39208 , \39209 , \39210 ,
         \39211 , \39212 , \39213 , \39214 , \39215 , \39216 , \39217 , \39218 , \39219 , \39220 ,
         \39221 , \39222 , \39223 , \39224 , \39225 , \39226 , \39227 , \39228 , \39229 , \39230 ,
         \39231 , \39232 , \39233 , \39234 , \39235 , \39236 , \39237 , \39238 , \39239 , \39240 ,
         \39241 , \39242 , \39243 , \39244 , \39245 , \39246 , \39247 , \39248 , \39249 , \39250 ,
         \39251 , \39252 , \39253 , \39254 , \39255 , \39256 , \39257 , \39258 , \39259 , \39260 ,
         \39261 , \39262 , \39263 , \39264 , \39265 , \39266 , \39267 , \39268 , \39269 , \39270 ,
         \39271 , \39272 , \39273 , \39274 , \39275 , \39276 , \39277 , \39278 , \39279 , \39280 ,
         \39281 , \39282 , \39283 , \39284 , \39285 , \39286 , \39287 , \39288 , \39289 , \39290 ,
         \39291 , \39292 , \39293 , \39294 , \39295 , \39296 , \39297 , \39298 , \39299 , \39300 ,
         \39301 , \39302 , \39303 , \39304 , \39305 , \39306 , \39307 , \39308 , \39309 , \39310 ,
         \39311 , \39312 , \39313 , \39314 , \39315 , \39316 , \39317 , \39318 , \39319 , \39320 ,
         \39321 , \39322 , \39323 , \39324 , \39325 , \39326 , \39327 , \39328 , \39329 , \39330 ,
         \39331 , \39332 , \39333 , \39334 , \39335 , \39336 , \39337 , \39338 , \39339 , \39340 ,
         \39341 , \39342 , \39343 , \39344 , \39345 , \39346 , \39347 , \39348 , \39349 , \39350 ,
         \39351 , \39352 , \39353 , \39354 , \39355 , \39356 , \39357 , \39358 , \39359 , \39360 ,
         \39361 , \39362 , \39363 , \39364 , \39365 , \39366 , \39367 , \39368 , \39369 , \39370 ,
         \39371 , \39372 , \39373 , \39374 , \39375 , \39376 , \39377 , \39378 , \39379 , \39380 ,
         \39381 , \39382 , \39383 , \39384 , \39385 , \39386 , \39387 , \39388 , \39389 , \39390 ,
         \39391 , \39392 , \39393 , \39394 , \39395 , \39396 , \39397 , \39398 , \39399 , \39400 ,
         \39401 , \39402 , \39403 , \39404 , \39405 , \39406 , \39407 , \39408 , \39409 , \39410 ,
         \39411 , \39412 , \39413 , \39414 , \39415 , \39416 , \39417 , \39418 , \39419 , \39420 ,
         \39421 , \39422 , \39423 , \39424 , \39425 , \39426 , \39427 , \39428 , \39429 , \39430 ,
         \39431 , \39432 , \39433 , \39434 , \39435 , \39436 , \39437 , \39438 , \39439 , \39440 ,
         \39441 , \39442 , \39443 , \39444 , \39445 , \39446 , \39447 , \39448 , \39449 , \39450 ,
         \39451 , \39452 , \39453 , \39454 , \39455 , \39456 , \39457 , \39458 , \39459 , \39460 ,
         \39461 , \39462 , \39463 , \39464 , \39465 , \39466 , \39467 , \39468 , \39469 , \39470 ,
         \39471 , \39472 , \39473 , \39474 , \39475 , \39476 , \39477 , \39478 , \39479 , \39480 ,
         \39481 , \39482 , \39483 , \39484 , \39485 , \39486 , \39487 , \39488 , \39489 , \39490 ,
         \39491 , \39492 , \39493 , \39494 , \39495 , \39496 , \39497 , \39498 , \39499 , \39500 ,
         \39501 , \39502 , \39503 , \39504 , \39505 , \39506 , \39507 , \39508 , \39509 , \39510 ,
         \39511 , \39512 , \39513 , \39514 , \39515 , \39516 , \39517 , \39518 , \39519 , \39520 ,
         \39521 , \39522 , \39523 , \39524 , \39525 , \39526 , \39527 , \39528 , \39529 , \39530 ,
         \39531 , \39532 , \39533 , \39534 , \39535 , \39536 , \39537 , \39538 , \39539 , \39540 ,
         \39541 , \39542 , \39543 , \39544 , \39545 , \39546 , \39547 , \39548 , \39549 , \39550 ,
         \39551 , \39552 , \39553 , \39554 , \39555 , \39556 , \39557 , \39558 , \39559 , \39560 ,
         \39561 , \39562 , \39563 , \39564 , \39565 , \39566 , \39567 , \39568 , \39569 , \39570 ,
         \39571 , \39572 , \39573 , \39574 , \39575 , \39576 , \39577 , \39578 , \39579 , \39580 ,
         \39581 , \39582 , \39583 , \39584 , \39585 , \39586 , \39587 , \39588 , \39589 , \39590 ,
         \39591 , \39592 , \39593 , \39594 , \39595 , \39596 , \39597 , \39598 , \39599 , \39600 ,
         \39601 , \39602 , \39603 , \39604 , \39605 , \39606 , \39607 , \39608 , \39609 , \39610 ,
         \39611 , \39612 , \39613 , \39614 , \39615 , \39616 , \39617 , \39618 , \39619 , \39620 ,
         \39621 , \39622 , \39623 , \39624 , \39625 , \39626 , \39627 , \39628 , \39629 , \39630 ,
         \39631 , \39632 , \39633 , \39634 , \39635 , \39636 , \39637 , \39638 , \39639 , \39640 ,
         \39641 , \39642 , \39643 , \39644 , \39645 , \39646 , \39647 , \39648 , \39649 , \39650 ,
         \39651 , \39652 , \39653 , \39654 , \39655 , \39656 , \39657 , \39658 , \39659 , \39660 ,
         \39661 , \39662 , \39663 , \39664 , \39665 , \39666 , \39667 , \39668 , \39669 , \39670 ,
         \39671 , \39672 , \39673 , \39674 , \39675 , \39676 , \39677 , \39678 , \39679 , \39680 ,
         \39681 , \39682 , \39683 , \39684 , \39685 , \39686 , \39687 , \39688 , \39689 , \39690 ,
         \39691 , \39692 , \39693 , \39694 , \39695 , \39696 , \39697 , \39698 , \39699 , \39700 ,
         \39701 , \39702 , \39703 , \39704 , \39705 , \39706 , \39707 , \39708 , \39709 , \39710 ,
         \39711 , \39712 , \39713 , \39714 , \39715 , \39716 , \39717 , \39718 , \39719 , \39720 ,
         \39721 , \39722 , \39723 , \39724 , \39725 , \39726 , \39727 , \39728 , \39729 , \39730 ,
         \39731 , \39732 , \39733 , \39734 , \39735 , \39736 , \39737 , \39738 , \39739 , \39740 ,
         \39741 , \39742 , \39743 , \39744 , \39745 , \39746 , \39747 , \39748 , \39749 , \39750 ,
         \39751 , \39752 , \39753 , \39754 , \39755 , \39756 , \39757 , \39758 , \39759 , \39760 ,
         \39761 , \39762 , \39763 , \39764 , \39765 , \39766 , \39767 , \39768 , \39769 , \39770 ,
         \39771 , \39772 , \39773 , \39774 , \39775 , \39776 , \39777 , \39778 , \39779 , \39780 ,
         \39781 , \39782 , \39783 , \39784 , \39785 , \39786 , \39787 , \39788 , \39789 , \39790 ,
         \39791 , \39792 , \39793 , \39794 , \39795 , \39796 , \39797 , \39798 , \39799 , \39800 ,
         \39801 , \39802 , \39803 , \39804 , \39805 , \39806 , \39807 , \39808 , \39809 , \39810 ,
         \39811 , \39812 , \39813 , \39814 , \39815 , \39816 , \39817 , \39818 , \39819 , \39820 ,
         \39821 , \39822 , \39823 , \39824 , \39825 , \39826 , \39827 , \39828 , \39829 , \39830 ,
         \39831 , \39832 , \39833 , \39834 , \39835 , \39836 , \39837 , \39838 , \39839 , \39840 ,
         \39841 , \39842 , \39843 , \39844 , \39845 , \39846 , \39847 , \39848 , \39849 , \39850 ,
         \39851 , \39852 , \39853 , \39854 , \39855 , \39856 , \39857 , \39858 , \39859 , \39860 ,
         \39861 , \39862 , \39863 , \39864 , \39865 , \39866 , \39867 , \39868 , \39869 , \39870 ,
         \39871 , \39872 , \39873 , \39874 , \39875 , \39876 , \39877 , \39878 , \39879 , \39880 ,
         \39881 , \39882 , \39883 , \39884 , \39885 , \39886 , \39887 , \39888 , \39889 , \39890 ,
         \39891 , \39892 , \39893 , \39894 , \39895 , \39896 , \39897 , \39898 , \39899 , \39900 ,
         \39901 , \39902 , \39903 , \39904 , \39905 , \39906 , \39907 , \39908 , \39909 , \39910 ,
         \39911 , \39912 , \39913 , \39914 , \39915 , \39916 , \39917 , \39918 , \39919 , \39920 ,
         \39921 , \39922 , \39923 , \39924 , \39925 , \39926 , \39927 , \39928 , \39929 , \39930 ,
         \39931 , \39932 , \39933 , \39934 , \39935 , \39936 , \39937 , \39938 , \39939 , \39940 ,
         \39941 , \39942 , \39943 , \39944 , \39945 , \39946 , \39947 , \39948 , \39949 , \39950 ,
         \39951 , \39952 , \39953 , \39954 , \39955 , \39956 , \39957 , \39958 , \39959 , \39960 ,
         \39961 , \39962 , \39963 , \39964 , \39965 , \39966 , \39967 , \39968 , \39969 , \39970 ,
         \39971 , \39972 , \39973 , \39974 , \39975 , \39976 , \39977 , \39978 , \39979 , \39980 ,
         \39981 , \39982 , \39983 , \39984 , \39985 , \39986 , \39987 , \39988 , \39989 , \39990 ,
         \39991 , \39992 , \39993 , \39994 , \39995 , \39996 , \39997 , \39998 , \39999 , \40000 ,
         \40001 , \40002 , \40003 , \40004 , \40005 , \40006 , \40007 , \40008 , \40009 , \40010 ,
         \40011 , \40012 , \40013 , \40014 , \40015 , \40016 , \40017 , \40018 , \40019 , \40020 ,
         \40021 , \40022 , \40023 , \40024 , \40025 , \40026 , \40027 , \40028 , \40029 , \40030 ,
         \40031 , \40032 , \40033 , \40034 , \40035 , \40036 , \40037 , \40038 , \40039 , \40040 ,
         \40041 , \40042 , \40043 , \40044 , \40045 , \40046 , \40047 , \40048 , \40049 , \40050 ,
         \40051 , \40052 , \40053 , \40054 , \40055 , \40056 , \40057 , \40058 , \40059 , \40060 ,
         \40061 , \40062 , \40063 , \40064 , \40065 , \40066 , \40067 , \40068 , \40069 , \40070 ,
         \40071 , \40072 , \40073 , \40074 , \40075 , \40076 , \40077 , \40078 , \40079 , \40080 ,
         \40081 , \40082 , \40083 , \40084 , \40085 , \40086 , \40087 , \40088 , \40089 , \40090 ,
         \40091 , \40092 , \40093 , \40094 , \40095 , \40096 , \40097 , \40098 , \40099 , \40100 ,
         \40101 , \40102 , \40103 , \40104 , \40105 , \40106 , \40107 , \40108 , \40109 , \40110 ,
         \40111 , \40112 , \40113 , \40114 , \40115 , \40116 , \40117 , \40118 , \40119 , \40120 ,
         \40121 , \40122 , \40123 , \40124 , \40125 , \40126 , \40127 , \40128 , \40129 , \40130 ,
         \40131 , \40132 , \40133 , \40134 , \40135 , \40136 , \40137 , \40138 , \40139 , \40140 ,
         \40141 , \40142 , \40143 , \40144 , \40145 , \40146 , \40147 , \40148 , \40149 , \40150 ,
         \40151 , \40152 , \40153 , \40154 , \40155 , \40156 , \40157 , \40158 , \40159 , \40160 ,
         \40161 , \40162 , \40163 , \40164 , \40165 , \40166 , \40167 , \40168 , \40169 , \40170 ,
         \40171 , \40172 , \40173 , \40174 , \40175 , \40176 , \40177 , \40178 , \40179 , \40180 ,
         \40181 , \40182 , \40183 , \40184 , \40185 , \40186 , \40187 , \40188 , \40189 , \40190 ,
         \40191 , \40192 , \40193 , \40194 , \40195 , \40196 , \40197 , \40198 , \40199 , \40200 ,
         \40201 , \40202 , \40203 , \40204 , \40205 , \40206 , \40207 , \40208 , \40209 , \40210 ,
         \40211 , \40212 , \40213 , \40214 , \40215 , \40216 , \40217 , \40218 , \40219 , \40220 ,
         \40221 , \40222 , \40223 , \40224 , \40225 , \40226 , \40227 , \40228 , \40229 , \40230 ,
         \40231 , \40232 , \40233 , \40234 , \40235 , \40236 , \40237 , \40238 , \40239 , \40240 ,
         \40241 , \40242 , \40243 , \40244 , \40245 , \40246 , \40247 , \40248 , \40249 , \40250 ,
         \40251 , \40252 , \40253 , \40254 , \40255 , \40256 , \40257 , \40258 , \40259 , \40260 ,
         \40261 , \40262 , \40263 , \40264 , \40265 , \40266 , \40267 , \40268 , \40269 , \40270 ,
         \40271 , \40272 , \40273 , \40274 , \40275 , \40276 , \40277 , \40278 , \40279 , \40280 ,
         \40281 , \40282 , \40283 , \40284 , \40285 , \40286 , \40287 , \40288 , \40289 , \40290 ,
         \40291 , \40292 , \40293 , \40294 , \40295 , \40296 , \40297 , \40298 , \40299 , \40300 ,
         \40301 , \40302 , \40303 , \40304 , \40305 , \40306 , \40307 , \40308 , \40309 , \40310 ,
         \40311 , \40312 , \40313 , \40314 , \40315 , \40316 , \40317 , \40318 , \40319 , \40320 ,
         \40321 , \40322 , \40323 , \40324 , \40325 , \40326 , \40327 , \40328 , \40329 , \40330 ,
         \40331 , \40332 , \40333 , \40334 , \40335 , \40336 , \40337 , \40338 , \40339 , \40340 ,
         \40341 , \40342 , \40343 , \40344 , \40345 , \40346 , \40347 , \40348 , \40349 , \40350 ,
         \40351 , \40352 , \40353 , \40354 , \40355 , \40356 , \40357 , \40358 , \40359 , \40360 ,
         \40361 , \40362 , \40363 , \40364 , \40365 , \40366 , \40367 , \40368 , \40369 , \40370 ,
         \40371 , \40372 , \40373 , \40374 , \40375 , \40376 , \40377 , \40378 , \40379 , \40380 ,
         \40381 , \40382 , \40383 , \40384 , \40385 , \40386 , \40387 , \40388 , \40389 , \40390 ,
         \40391 , \40392 , \40393 , \40394 , \40395 , \40396 , \40397 , \40398 , \40399 , \40400 ,
         \40401 , \40402 , \40403 , \40404 , \40405 , \40406 , \40407 , \40408 , \40409 , \40410 ,
         \40411 , \40412 , \40413 , \40414 , \40415 , \40416 , \40417 , \40418 , \40419 , \40420 ,
         \40421 , \40422 , \40423 , \40424 , \40425 , \40426 , \40427 , \40428 , \40429 , \40430 ,
         \40431 , \40432 , \40433 , \40434 , \40435 , \40436 , \40437 , \40438 , \40439 , \40440 ,
         \40441 , \40442 , \40443 , \40444 , \40445 , \40446 , \40447 , \40448 , \40449 , \40450 ,
         \40451 , \40452 , \40453 , \40454 , \40455 , \40456 , \40457 , \40458 , \40459 , \40460 ,
         \40461 , \40462 , \40463 , \40464 , \40465 , \40466 , \40467 , \40468 , \40469 , \40470 ,
         \40471 , \40472 , \40473 , \40474 , \40475 , \40476 , \40477 , \40478 , \40479 , \40480 ,
         \40481 , \40482 , \40483 , \40484 , \40485 , \40486 , \40487 , \40488 , \40489 , \40490 ,
         \40491 , \40492 , \40493 , \40494 , \40495 , \40496 , \40497 , \40498 , \40499 , \40500 ,
         \40501 , \40502 , \40503 , \40504 , \40505 , \40506 , \40507 , \40508 , \40509 , \40510 ,
         \40511 , \40512 , \40513 , \40514 , \40515 , \40516 , \40517 , \40518 , \40519 , \40520 ,
         \40521 , \40522 , \40523 , \40524 , \40525 , \40526 , \40527 , \40528 , \40529 , \40530 ,
         \40531 , \40532 , \40533 , \40534 , \40535 , \40536 , \40537 , \40538 , \40539 , \40540 ,
         \40541 , \40542 , \40543 , \40544 , \40545 , \40546 , \40547 , \40548 , \40549 , \40550 ,
         \40551 , \40552 , \40553 , \40554 , \40555 , \40556 , \40557 , \40558 , \40559 , \40560 ,
         \40561 , \40562 , \40563 , \40564 , \40565 , \40566 , \40567 , \40568 , \40569 , \40570 ,
         \40571 , \40572 , \40573 , \40574 , \40575 , \40576 , \40577 , \40578 , \40579 , \40580 ,
         \40581 , \40582 , \40583 , \40584 , \40585 , \40586 , \40587 , \40588 , \40589 , \40590 ,
         \40591 , \40592 , \40593 , \40594 , \40595 , \40596 , \40597 , \40598 , \40599 , \40600 ,
         \40601 , \40602 , \40603 , \40604 , \40605 , \40606 , \40607 , \40608 , \40609 , \40610 ,
         \40611 , \40612 , \40613 , \40614 , \40615 , \40616 , \40617 , \40618 , \40619 , \40620 ,
         \40621 , \40622 , \40623 , \40624 , \40625 , \40626 , \40627 , \40628 , \40629 , \40630 ,
         \40631 , \40632 , \40633 , \40634 , \40635 , \40636 , \40637 , \40638 , \40639 , \40640 ,
         \40641 , \40642 , \40643 , \40644 , \40645 , \40646 , \40647 , \40648 , \40649 , \40650 ,
         \40651 , \40652 , \40653 , \40654 , \40655 , \40656 , \40657 , \40658 , \40659 , \40660 ,
         \40661 , \40662 , \40663 , \40664 , \40665 , \40666 , \40667 , \40668 , \40669 , \40670 ,
         \40671 , \40672 , \40673 , \40674 , \40675 , \40676 , \40677 , \40678 , \40679 , \40680 ,
         \40681 , \40682 , \40683 , \40684 , \40685 , \40686 , \40687 , \40688 , \40689 , \40690 ,
         \40691 , \40692 , \40693 , \40694 , \40695 , \40696 , \40697 , \40698 , \40699 , \40700 ,
         \40701 , \40702 , \40703 , \40704 , \40705 , \40706 , \40707 , \40708 , \40709 , \40710 ,
         \40711 , \40712 , \40713 , \40714 , \40715 , \40716 , \40717 , \40718 , \40719 , \40720 ,
         \40721 , \40722 , \40723 , \40724 , \40725 , \40726 , \40727 , \40728 , \40729 , \40730 ,
         \40731 , \40732 , \40733 , \40734 , \40735 , \40736 , \40737 , \40738 , \40739 , \40740 ,
         \40741 , \40742 , \40743 , \40744 , \40745 , \40746 , \40747 , \40748 , \40749 , \40750 ,
         \40751 , \40752 , \40753 , \40754 , \40755 , \40756 , \40757 , \40758 , \40759 , \40760 ,
         \40761 , \40762 , \40763 , \40764 , \40765 , \40766 , \40767 , \40768 , \40769 , \40770 ,
         \40771 , \40772 , \40773 , \40774 , \40775 , \40776 , \40777 , \40778 , \40779 , \40780 ,
         \40781 , \40782 , \40783 , \40784 , \40785 , \40786 , \40787 , \40788 , \40789 , \40790 ,
         \40791 , \40792 , \40793 , \40794 , \40795 , \40796 , \40797 , \40798 , \40799 , \40800 ,
         \40801 , \40802 , \40803 , \40804 , \40805 , \40806 , \40807 , \40808 , \40809 , \40810 ,
         \40811 , \40812 , \40813 , \40814 , \40815 , \40816 , \40817 , \40818 , \40819 , \40820 ,
         \40821 , \40822 , \40823 , \40824 , \40825 , \40826 , \40827 , \40828 , \40829 , \40830 ,
         \40831 , \40832 , \40833 , \40834 , \40835 , \40836 , \40837 , \40838 , \40839 , \40840 ,
         \40841 , \40842 , \40843 , \40844 , \40845 , \40846 , \40847 , \40848 , \40849 , \40850 ,
         \40851 , \40852 , \40853 , \40854 , \40855 , \40856 , \40857 , \40858 , \40859 , \40860 ,
         \40861 , \40862 , \40863 , \40864 , \40865 , \40866 , \40867 , \40868 , \40869 , \40870 ,
         \40871 , \40872 , \40873 , \40874 , \40875 , \40876 , \40877 , \40878 , \40879 , \40880 ,
         \40881 , \40882 , \40883 , \40884 , \40885 , \40886 , \40887 , \40888 , \40889 , \40890 ,
         \40891 , \40892 , \40893 , \40894 , \40895 , \40896 , \40897 , \40898 , \40899 , \40900 ,
         \40901 , \40902 , \40903 , \40904 , \40905 , \40906 , \40907 , \40908 , \40909 , \40910 ,
         \40911 , \40912 , \40913 , \40914 , \40915 , \40916 , \40917 , \40918 , \40919 , \40920 ,
         \40921 , \40922 , \40923 , \40924 , \40925 , \40926 , \40927 , \40928 , \40929 , \40930 ,
         \40931 , \40932 , \40933 , \40934 , \40935 , \40936 , \40937 , \40938 , \40939 , \40940 ,
         \40941 , \40942 , \40943 , \40944 , \40945 , \40946 , \40947 , \40948 , \40949 , \40950 ,
         \40951 , \40952 , \40953 , \40954 , \40955 , \40956 , \40957 , \40958 , \40959 , \40960 ,
         \40961 , \40962 , \40963 , \40964 , \40965 , \40966 , \40967 , \40968 , \40969 , \40970 ,
         \40971 , \40972 , \40973 , \40974 , \40975 , \40976 , \40977 , \40978 , \40979 , \40980 ,
         \40981 , \40982 , \40983 , \40984 , \40985 , \40986 , \40987 , \40988 , \40989 , \40990 ,
         \40991 , \40992 , \40993 , \40994 , \40995 , \40996 , \40997 , \40998 , \40999 , \41000 ,
         \41001 , \41002 , \41003 , \41004 , \41005 , \41006 , \41007 , \41008 , \41009 , \41010 ,
         \41011 , \41012 , \41013 , \41014 , \41015 , \41016 , \41017 , \41018 , \41019 , \41020 ,
         \41021 , \41022 , \41023 , \41024 , \41025 , \41026 , \41027 , \41028 , \41029 , \41030 ,
         \41031 , \41032 , \41033 , \41034 , \41035 , \41036 , \41037 , \41038 , \41039 , \41040 ,
         \41041 , \41042 , \41043 , \41044 , \41045 , \41046 , \41047 , \41048 , \41049 , \41050 ,
         \41051 , \41052 , \41053 , \41054 , \41055 , \41056 , \41057 , \41058 , \41059 , \41060 ,
         \41061 , \41062 , \41063 , \41064 , \41065 , \41066 , \41067 , \41068 , \41069 , \41070 ,
         \41071 , \41072 , \41073 , \41074 , \41075 , \41076 , \41077 , \41078 , \41079 , \41080 ,
         \41081 , \41082 , \41083 , \41084 , \41085 , \41086 , \41087 , \41088 , \41089 , \41090 ,
         \41091 , \41092 , \41093 , \41094 , \41095 , \41096 , \41097 , \41098 , \41099 , \41100 ,
         \41101 , \41102 , \41103 , \41104 , \41105 , \41106 , \41107 , \41108 , \41109 , \41110 ,
         \41111 , \41112 , \41113 , \41114 , \41115 , \41116 , \41117 , \41118 , \41119 , \41120 ,
         \41121 , \41122 , \41123 , \41124 , \41125 , \41126 , \41127 , \41128 , \41129 , \41130 ,
         \41131 , \41132 , \41133 , \41134 , \41135 , \41136 , \41137 , \41138 , \41139 , \41140 ,
         \41141 , \41142 , \41143 , \41144 , \41145 , \41146 , \41147 , \41148 , \41149 , \41150 ,
         \41151 , \41152 , \41153 , \41154 , \41155 , \41156 , \41157 , \41158 , \41159 , \41160 ,
         \41161 , \41162 , \41163 , \41164 , \41165 , \41166 , \41167 , \41168 , \41169 , \41170 ,
         \41171 , \41172 , \41173 , \41174 , \41175 , \41176 , \41177 , \41178 , \41179 , \41180 ,
         \41181 , \41182 , \41183 , \41184 , \41185 , \41186 , \41187 , \41188 , \41189 , \41190 ,
         \41191 , \41192 , \41193 , \41194 , \41195 , \41196 , \41197 , \41198 , \41199 , \41200 ,
         \41201 , \41202 , \41203 , \41204 , \41205 , \41206 , \41207 , \41208 , \41209 , \41210 ,
         \41211 , \41212 , \41213 , \41214 , \41215 , \41216 , \41217 , \41218 , \41219 , \41220 ,
         \41221 , \41222 , \41223 , \41224 , \41225 , \41226 , \41227 , \41228 , \41229 , \41230 ,
         \41231 , \41232 , \41233 , \41234 , \41235 , \41236 , \41237 , \41238 , \41239 , \41240 ,
         \41241 , \41242 , \41243 , \41244 , \41245 , \41246 , \41247 , \41248 , \41249 , \41250 ,
         \41251 , \41252 , \41253 , \41254 , \41255 , \41256 , \41257 , \41258 , \41259 , \41260 ,
         \41261 , \41262 , \41263 , \41264 , \41265 , \41266 , \41267 , \41268 , \41269 , \41270 ,
         \41271 , \41272 , \41273 , \41274 , \41275 , \41276 , \41277 , \41278 , \41279 , \41280 ,
         \41281 , \41282 , \41283 , \41284 , \41285 , \41286 , \41287 , \41288 , \41289 , \41290 ,
         \41291 , \41292 , \41293 , \41294 , \41295 , \41296 , \41297 , \41298 , \41299 , \41300 ,
         \41301 , \41302 , \41303 , \41304 , \41305 , \41306 , \41307 , \41308 , \41309 , \41310 ,
         \41311 , \41312 , \41313 , \41314 , \41315 , \41316 , \41317 , \41318 , \41319 , \41320 ,
         \41321 , \41322 , \41323 , \41324 , \41325 , \41326 , \41327 , \41328 , \41329 , \41330 ,
         \41331 , \41332 , \41333 , \41334 , \41335 , \41336 , \41337 , \41338 , \41339 , \41340 ,
         \41341 , \41342 , \41343 , \41344 , \41345 , \41346 , \41347 , \41348 , \41349 , \41350 ,
         \41351 , \41352 , \41353 , \41354 , \41355 , \41356 , \41357 , \41358 , \41359 , \41360 ,
         \41361 , \41362 , \41363 , \41364 , \41365 , \41366 , \41367 , \41368 , \41369 , \41370 ,
         \41371 , \41372 , \41373 , \41374 , \41375 , \41376 , \41377 , \41378 , \41379 , \41380 ,
         \41381 , \41382 , \41383 , \41384 , \41385 , \41386 , \41387 , \41388 , \41389 , \41390 ,
         \41391 , \41392 , \41393 , \41394 , \41395 , \41396 , \41397 , \41398 , \41399 , \41400 ,
         \41401 , \41402 , \41403 , \41404 , \41405 , \41406 , \41407 , \41408 , \41409 , \41410 ,
         \41411 , \41412 , \41413 , \41414 , \41415 , \41416 , \41417 , \41418 , \41419 , \41420 ,
         \41421 , \41422 , \41423 , \41424 , \41425 , \41426 , \41427 , \41428 , \41429 , \41430 ,
         \41431 , \41432 , \41433 , \41434 , \41435 , \41436 , \41437 , \41438 , \41439 , \41440 ,
         \41441 , \41442 , \41443 , \41444 , \41445 , \41446 , \41447 , \41448 , \41449 , \41450 ,
         \41451 , \41452 , \41453 , \41454 , \41455 , \41456 , \41457 , \41458 , \41459 , \41460 ,
         \41461 , \41462 , \41463 , \41464 , \41465 , \41466 , \41467 , \41468 , \41469 , \41470 ,
         \41471 , \41472 , \41473 , \41474 , \41475 , \41476 , \41477 , \41478 , \41479 , \41480 ,
         \41481 , \41482 , \41483 , \41484 , \41485 , \41486 , \41487 , \41488 , \41489 , \41490 ,
         \41491 , \41492 , \41493 , \41494 , \41495 , \41496 , \41497 , \41498 , \41499 , \41500 ,
         \41501 , \41502 , \41503 , \41504 , \41505 , \41506 , \41507 , \41508 , \41509 , \41510 ,
         \41511 , \41512 , \41513 , \41514 , \41515 , \41516 , \41517 , \41518 , \41519 , \41520 ,
         \41521 , \41522 , \41523 , \41524 , \41525 , \41526 , \41527 , \41528 , \41529 , \41530 ,
         \41531 , \41532 , \41533 , \41534 , \41535 , \41536 , \41537 , \41538 , \41539 , \41540 ,
         \41541 , \41542 , \41543 , \41544 , \41545 , \41546 , \41547 , \41548 , \41549 , \41550 ,
         \41551 , \41552 , \41553 , \41554 , \41555 , \41556 , \41557 , \41558 , \41559 , \41560 ,
         \41561 , \41562 , \41563 , \41564 , \41565 , \41566 , \41567 , \41568 , \41569 , \41570 ,
         \41571 , \41572 , \41573 , \41574 , \41575 , \41576 , \41577 , \41578 , \41579 , \41580 ,
         \41581 , \41582 , \41583 , \41584 , \41585 , \41586 , \41587 , \41588 , \41589 , \41590 ,
         \41591 , \41592 , \41593 , \41594 , \41595 , \41596 , \41597 , \41598 , \41599 , \41600 ,
         \41601 , \41602 , \41603 , \41604 , \41605 , \41606 , \41607 , \41608 , \41609 , \41610 ,
         \41611 , \41612 , \41613 , \41614 , \41615 , \41616 , \41617 , \41618 , \41619 , \41620 ,
         \41621 , \41622 , \41623 , \41624 , \41625 , \41626 , \41627 , \41628 , \41629 , \41630 ,
         \41631 , \41632 , \41633 , \41634 , \41635 , \41636 , \41637 , \41638 , \41639 , \41640 ,
         \41641 , \41642 , \41643 , \41644 , \41645 , \41646 , \41647 , \41648 , \41649 , \41650 ,
         \41651 , \41652 , \41653 , \41654 , \41655 , \41656 , \41657 , \41658 , \41659 , \41660 ,
         \41661 , \41662 , \41663 , \41664 , \41665 , \41666 , \41667 , \41668 , \41669 , \41670 ,
         \41671 , \41672 , \41673 , \41674 , \41675 , \41676 , \41677 , \41678 , \41679 , \41680 ,
         \41681 , \41682 , \41683 , \41684 , \41685 , \41686 , \41687 , \41688 , \41689 , \41690 ,
         \41691 , \41692 , \41693 , \41694 , \41695 , \41696 , \41697 , \41698 , \41699 , \41700 ,
         \41701 , \41702 , \41703 , \41704 , \41705 , \41706 , \41707 , \41708 , \41709 , \41710 ,
         \41711 , \41712 , \41713 , \41714 , \41715 , \41716 , \41717 , \41718 , \41719 , \41720 ,
         \41721 , \41722 , \41723 , \41724 , \41725 , \41726 , \41727 , \41728 , \41729 , \41730 ,
         \41731 , \41732 , \41733 , \41734 , \41735 , \41736 , \41737 , \41738 , \41739 , \41740 ,
         \41741 , \41742 , \41743 , \41744 , \41745 , \41746 , \41747 , \41748 , \41749 , \41750 ,
         \41751 , \41752 , \41753 , \41754 , \41755 , \41756 , \41757 , \41758 , \41759 , \41760 ,
         \41761 , \41762 , \41763 , \41764 , \41765 , \41766 , \41767 , \41768 , \41769 , \41770 ,
         \41771 , \41772 , \41773 , \41774 , \41775 , \41776 , \41777 , \41778 , \41779 , \41780 ,
         \41781 , \41782 , \41783 , \41784 , \41785 , \41786 , \41787 , \41788 , \41789 , \41790 ,
         \41791 , \41792 , \41793 , \41794 , \41795 , \41796 , \41797 , \41798 , \41799 , \41800 ,
         \41801 , \41802 , \41803 , \41804 , \41805 , \41806 , \41807 , \41808 , \41809 , \41810 ,
         \41811 , \41812 , \41813 , \41814 , \41815 , \41816 , \41817 , \41818 , \41819 , \41820 ,
         \41821 , \41822 , \41823 , \41824 , \41825 , \41826 , \41827 , \41828 , \41829 , \41830 ,
         \41831 , \41832 , \41833 , \41834 , \41835 , \41836 , \41837 , \41838 , \41839 , \41840 ,
         \41841 , \41842 , \41843 , \41844 , \41845 , \41846 , \41847 , \41848 , \41849 , \41850 ,
         \41851 , \41852 , \41853 , \41854 , \41855 , \41856 , \41857 , \41858 , \41859 , \41860 ,
         \41861 , \41862 , \41863 , \41864 , \41865 , \41866 , \41867 , \41868 , \41869 , \41870 ,
         \41871 , \41872 , \41873 , \41874 , \41875 , \41876 , \41877 , \41878 , \41879 , \41880 ,
         \41881 , \41882 , \41883 , \41884 , \41885 , \41886 , \41887 , \41888 , \41889 , \41890 ,
         \41891 , \41892 , \41893 , \41894 , \41895 , \41896 , \41897 , \41898 , \41899 , \41900 ,
         \41901 , \41902 , \41903 , \41904 , \41905 , \41906 , \41907 , \41908 , \41909 , \41910 ,
         \41911 , \41912 , \41913 , \41914 , \41915 , \41916 , \41917 , \41918 , \41919 , \41920 ,
         \41921 , \41922 , \41923 , \41924 , \41925 , \41926 , \41927 , \41928 , \41929 , \41930 ,
         \41931 , \41932 , \41933 , \41934 , \41935 , \41936 , \41937 , \41938 , \41939 , \41940 ,
         \41941 , \41942 , \41943 , \41944 , \41945 , \41946 , \41947 , \41948 , \41949 , \41950 ,
         \41951 , \41952 , \41953 , \41954 , \41955 , \41956 , \41957 , \41958 , \41959 , \41960 ,
         \41961 , \41962 , \41963 , \41964 , \41965 , \41966 , \41967 , \41968 , \41969 , \41970 ,
         \41971 , \41972 , \41973 , \41974 , \41975 , \41976 , \41977 , \41978 , \41979 , \41980 ,
         \41981 , \41982 , \41983 , \41984 , \41985 , \41986 , \41987 , \41988 , \41989 , \41990 ,
         \41991 , \41992 , \41993 , \41994 , \41995 , \41996 , \41997 , \41998 , \41999 , \42000 ,
         \42001 , \42002 , \42003 , \42004 , \42005 , \42006 , \42007 , \42008 , \42009 , \42010 ,
         \42011 , \42012 , \42013 , \42014 , \42015 , \42016 , \42017 , \42018 , \42019 , \42020 ,
         \42021 , \42022 , \42023 , \42024 , \42025 , \42026 , \42027 , \42028 , \42029 , \42030 ,
         \42031 , \42032 , \42033 , \42034 , \42035 , \42036 , \42037 , \42038 , \42039 , \42040 ,
         \42041 , \42042 , \42043 , \42044 , \42045 , \42046 , \42047 , \42048 , \42049 , \42050 ,
         \42051 , \42052 , \42053 , \42054 , \42055 , \42056 , \42057 , \42058 , \42059 , \42060 ,
         \42061 , \42062 , \42063 , \42064 , \42065 , \42066 , \42067 , \42068 , \42069 , \42070 ,
         \42071 , \42072 , \42073 , \42074 , \42075 , \42076 , \42077 , \42078 , \42079 , \42080 ,
         \42081 , \42082 , \42083 , \42084 , \42085 , \42086 , \42087 , \42088 , \42089 , \42090 ,
         \42091 , \42092 , \42093 , \42094 , \42095 , \42096 , \42097 , \42098 , \42099 , \42100 ,
         \42101 , \42102 , \42103 , \42104 , \42105 , \42106 , \42107 , \42108 , \42109 , \42110 ,
         \42111 , \42112 , \42113 , \42114 , \42115 , \42116 , \42117 , \42118 , \42119 , \42120 ,
         \42121 , \42122 , \42123 , \42124 , \42125 , \42126 , \42127 , \42128 , \42129 , \42130 ,
         \42131 , \42132 , \42133 , \42134 , \42135 , \42136 , \42137 , \42138 , \42139 , \42140 ,
         \42141 , \42142 , \42143 , \42144 , \42145 , \42146 , \42147 , \42148 , \42149 , \42150 ,
         \42151 , \42152 , \42153 , \42154 , \42155 , \42156 , \42157 , \42158 , \42159 , \42160 ,
         \42161 , \42162 , \42163 , \42164 , \42165 , \42166 , \42167 , \42168 , \42169 , \42170 ,
         \42171 , \42172 , \42173 , \42174 , \42175 , \42176 , \42177 , \42178 , \42179 , \42180 ,
         \42181 , \42182 , \42183 , \42184 , \42185 , \42186 , \42187 , \42188 , \42189 , \42190 ,
         \42191 , \42192 , \42193 , \42194 , \42195 , \42196 , \42197 , \42198 , \42199 , \42200 ,
         \42201 , \42202 , \42203 , \42204 , \42205 , \42206 , \42207 , \42208 , \42209 , \42210 ,
         \42211 , \42212 , \42213 , \42214 , \42215 , \42216 , \42217 , \42218 , \42219 , \42220 ,
         \42221 , \42222 , \42223 , \42224 , \42225 , \42226 , \42227 , \42228 , \42229 , \42230 ,
         \42231 , \42232 , \42233 , \42234 , \42235 , \42236 , \42237 , \42238 , \42239 , \42240 ,
         \42241 , \42242 , \42243 , \42244 , \42245 , \42246 , \42247 , \42248 , \42249 , \42250 ,
         \42251 , \42252 , \42253 , \42254 , \42255 , \42256 , \42257 , \42258 , \42259 , \42260 ,
         \42261 , \42262 , \42263 , \42264 , \42265 , \42266 , \42267 , \42268 , \42269 , \42270 ,
         \42271 , \42272 , \42273 , \42274 , \42275 , \42276 , \42277 , \42278 , \42279 , \42280 ,
         \42281 , \42282 , \42283 , \42284 , \42285 , \42286 , \42287 , \42288 , \42289 , \42290 ,
         \42291 , \42292 , \42293 , \42294 , \42295 , \42296 , \42297 , \42298 , \42299 , \42300 ,
         \42301 , \42302 , \42303 , \42304 , \42305 , \42306 , \42307 , \42308 , \42309 , \42310 ,
         \42311 , \42312 , \42313 , \42314 , \42315 , \42316 , \42317 , \42318 , \42319 , \42320 ,
         \42321 , \42322 , \42323 , \42324 , \42325 , \42326 , \42327 , \42328 , \42329 , \42330 ,
         \42331 , \42332 , \42333 , \42334 , \42335 , \42336 , \42337 , \42338 , \42339 , \42340 ,
         \42341 , \42342 , \42343 , \42344 , \42345 , \42346 , \42347 , \42348 , \42349 , \42350 ,
         \42351 , \42352 , \42353 , \42354 , \42355 , \42356 , \42357 , \42358 , \42359 , \42360 ,
         \42361 , \42362 , \42363 , \42364 , \42365 , \42366 , \42367 , \42368 , \42369 , \42370 ,
         \42371 , \42372 , \42373 , \42374 , \42375 , \42376 , \42377 , \42378 , \42379 , \42380 ,
         \42381 , \42382 , \42383 , \42384 , \42385 , \42386 , \42387 , \42388 , \42389 , \42390 ,
         \42391 , \42392 , \42393 , \42394 , \42395 , \42396 , \42397 , \42398 , \42399 , \42400 ,
         \42401 , \42402 , \42403 , \42404 , \42405 , \42406 , \42407 , \42408 , \42409 , \42410 ,
         \42411 , \42412 , \42413 , \42414 , \42415 , \42416 , \42417 , \42418 , \42419 , \42420 ,
         \42421 , \42422 , \42423 , \42424 , \42425 , \42426 , \42427 , \42428 , \42429 , \42430 ,
         \42431 , \42432 , \42433 , \42434 , \42435 , \42436 , \42437 , \42438 , \42439 , \42440 ,
         \42441 , \42442 , \42443 , \42444 , \42445 , \42446 , \42447 , \42448 , \42449 , \42450 ,
         \42451 , \42452 , \42453 , \42454 , \42455 , \42456 , \42457 , \42458 , \42459 , \42460 ,
         \42461 , \42462 , \42463 , \42464 , \42465 , \42466 , \42467 , \42468 , \42469 , \42470 ,
         \42471 , \42472 , \42473 , \42474 , \42475 , \42476 , \42477 , \42478 , \42479 , \42480 ,
         \42481 , \42482 , \42483 , \42484 , \42485 , \42486 , \42487 , \42488 , \42489 , \42490 ,
         \42491 , \42492 , \42493 , \42494 , \42495 , \42496 , \42497 , \42498 , \42499 , \42500 ,
         \42501 , \42502 , \42503 , \42504 , \42505 , \42506 , \42507 , \42508 , \42509 , \42510 ,
         \42511 , \42512 , \42513 , \42514 , \42515 , \42516 , \42517 , \42518 , \42519 , \42520 ,
         \42521 , \42522 , \42523 , \42524 , \42525 , \42526 , \42527 , \42528 , \42529 , \42530 ,
         \42531 , \42532 , \42533 , \42534 , \42535 , \42536 , \42537 , \42538 , \42539 , \42540 ,
         \42541 , \42542 , \42543 , \42544 , \42545 , \42546 , \42547 , \42548 , \42549 , \42550 ,
         \42551 , \42552 , \42553 , \42554 , \42555 , \42556 , \42557 , \42558 , \42559 , \42560 ,
         \42561 , \42562 , \42563 , \42564 , \42565 , \42566 , \42567 , \42568 , \42569 , \42570 ,
         \42571 , \42572 , \42573 , \42574 , \42575 , \42576 , \42577 , \42578 , \42579 , \42580 ,
         \42581 , \42582 , \42583 , \42584 , \42585 , \42586 , \42587 , \42588 , \42589 , \42590 ,
         \42591 , \42592 , \42593 , \42594 , \42595 , \42596 , \42597 , \42598 , \42599 , \42600 ,
         \42601 , \42602 , \42603 , \42604 , \42605 , \42606 , \42607 , \42608 , \42609 , \42610 ,
         \42611 , \42612 , \42613 , \42614 , \42615 , \42616 , \42617 , \42618 , \42619 , \42620 ,
         \42621 , \42622 , \42623 , \42624 , \42625 , \42626 , \42627 , \42628 , \42629 , \42630 ,
         \42631 , \42632 , \42633 , \42634 , \42635 , \42636 , \42637 , \42638 , \42639 , \42640 ,
         \42641 , \42642 , \42643 , \42644 , \42645 , \42646 , \42647 , \42648 , \42649 , \42650 ,
         \42651 , \42652 , \42653 , \42654 , \42655 , \42656 , \42657 , \42658 , \42659 , \42660 ,
         \42661 , \42662 , \42663 , \42664 , \42665 , \42666 , \42667 , \42668 , \42669 , \42670 ,
         \42671 , \42672 , \42673 , \42674 , \42675 , \42676 , \42677 , \42678 , \42679 , \42680 ,
         \42681 , \42682 , \42683 , \42684 , \42685 , \42686 , \42687 , \42688 , \42689 , \42690 ,
         \42691 , \42692 , \42693 , \42694 , \42695 , \42696 , \42697 , \42698 , \42699 , \42700 ,
         \42701 , \42702 , \42703 , \42704 , \42705 , \42706 , \42707 , \42708 , \42709 , \42710 ,
         \42711 , \42712 , \42713 , \42714 , \42715 , \42716 , \42717 , \42718 , \42719 , \42720 ,
         \42721 , \42722 , \42723 , \42724 , \42725 , \42726 , \42727 , \42728 , \42729 , \42730 ,
         \42731 , \42732 , \42733 , \42734 , \42735 , \42736 , \42737 , \42738 , \42739 , \42740 ,
         \42741 , \42742 , \42743 , \42744 , \42745 , \42746 , \42747 , \42748 , \42749 , \42750 ,
         \42751 , \42752 , \42753 , \42754 , \42755 , \42756 , \42757 , \42758 , \42759 , \42760 ,
         \42761 , \42762 , \42763 , \42764 , \42765 , \42766 , \42767 , \42768 , \42769 , \42770 ,
         \42771 , \42772 , \42773 , \42774 , \42775 , \42776 , \42777 , \42778 , \42779 , \42780 ,
         \42781 , \42782 , \42783 , \42784 , \42785 , \42786 , \42787 , \42788 , \42789 , \42790 ,
         \42791 , \42792 , \42793 , \42794 , \42795 , \42796 , \42797 , \42798 , \42799 , \42800 ,
         \42801 , \42802 , \42803 , \42804 , \42805 , \42806 , \42807 , \42808 , \42809 , \42810 ,
         \42811 , \42812 , \42813 , \42814 , \42815 , \42816 , \42817 , \42818 , \42819 , \42820 ,
         \42821 , \42822 , \42823 , \42824 , \42825 , \42826 , \42827 , \42828 , \42829 , \42830 ,
         \42831 , \42832 , \42833 , \42834 , \42835 , \42836 , \42837 , \42838 , \42839 , \42840 ,
         \42841 , \42842 , \42843 , \42844 , \42845 , \42846 , \42847 , \42848 , \42849 , \42850 ,
         \42851 , \42852 , \42853 , \42854 , \42855 , \42856 , \42857 , \42858 , \42859 , \42860 ,
         \42861 , \42862 , \42863 , \42864 , \42865 , \42866 , \42867 , \42868 , \42869 , \42870 ,
         \42871 , \42872 , \42873 , \42874 , \42875 , \42876 , \42877 , \42878 , \42879 , \42880 ,
         \42881 , \42882 , \42883 , \42884 , \42885 , \42886 , \42887 , \42888 , \42889 , \42890 ,
         \42891 , \42892 , \42893 , \42894 , \42895 , \42896 , \42897 , \42898 , \42899 , \42900 ,
         \42901 , \42902 , \42903 , \42904 , \42905 , \42906 , \42907 , \42908 , \42909 , \42910 ,
         \42911 , \42912 , \42913 , \42914 , \42915 , \42916 , \42917 , \42918 , \42919 , \42920 ,
         \42921 , \42922 , \42923 , \42924 , \42925 , \42926 , \42927 , \42928 , \42929 , \42930 ,
         \42931 , \42932 , \42933 , \42934 , \42935 , \42936 , \42937 , \42938 , \42939 , \42940 ,
         \42941 , \42942 , \42943 , \42944 , \42945 , \42946 , \42947 , \42948 , \42949 , \42950 ,
         \42951 , \42952 , \42953 , \42954 , \42955 , \42956 , \42957 , \42958 , \42959 , \42960 ,
         \42961 , \42962 , \42963 , \42964 , \42965 , \42966 , \42967 , \42968 , \42969 , \42970 ,
         \42971 , \42972 , \42973 , \42974 , \42975 , \42976 , \42977 , \42978 , \42979 , \42980 ,
         \42981 , \42982 , \42983 , \42984 , \42985 , \42986 , \42987 , \42988 , \42989 , \42990 ,
         \42991 , \42992 , \42993 , \42994 , \42995 , \42996 , \42997 , \42998 , \42999 , \43000 ,
         \43001 , \43002 , \43003 , \43004 , \43005 , \43006 , \43007 , \43008 , \43009 , \43010 ,
         \43011 , \43012 , \43013 , \43014 , \43015 , \43016 , \43017 , \43018 , \43019 , \43020 ,
         \43021 , \43022 , \43023 , \43024 , \43025 , \43026 , \43027 , \43028 , \43029 , \43030 ,
         \43031 , \43032 , \43033 , \43034 , \43035 , \43036 , \43037 , \43038 , \43039 , \43040 ,
         \43041 , \43042 , \43043 , \43044 , \43045 , \43046 , \43047 , \43048 , \43049 , \43050 ,
         \43051 , \43052 , \43053 , \43054 , \43055 , \43056 , \43057 , \43058 , \43059 , \43060 ,
         \43061 , \43062 , \43063 , \43064 , \43065 , \43066 , \43067 , \43068 , \43069 , \43070 ,
         \43071 , \43072 , \43073 , \43074 , \43075 , \43076 , \43077 , \43078 , \43079 , \43080 ,
         \43081 , \43082 , \43083 , \43084 , \43085 , \43086 , \43087 , \43088 , \43089 , \43090 ,
         \43091 , \43092 , \43093 , \43094 , \43095 , \43096 , \43097 , \43098 , \43099 , \43100 ,
         \43101 , \43102 , \43103 , \43104 , \43105 , \43106 , \43107 , \43108 , \43109 , \43110 ,
         \43111 , \43112 , \43113 , \43114 , \43115 , \43116 , \43117 , \43118 , \43119 , \43120 ,
         \43121 , \43122 , \43123 , \43124 , \43125 , \43126 , \43127 , \43128 , \43129 , \43130 ,
         \43131 , \43132 , \43133 , \43134 , \43135 , \43136 , \43137 , \43138 , \43139 , \43140 ,
         \43141 , \43142 , \43143 , \43144 , \43145 , \43146 , \43147 , \43148 , \43149 , \43150 ,
         \43151 , \43152 , \43153 , \43154 , \43155 , \43156 , \43157 , \43158 , \43159 , \43160 ,
         \43161 , \43162 , \43163 , \43164 , \43165 , \43166 , \43167 , \43168 , \43169 , \43170 ,
         \43171 , \43172 , \43173 , \43174 , \43175 , \43176 , \43177 , \43178 , \43179 , \43180 ,
         \43181 , \43182 , \43183 , \43184 , \43185 , \43186 , \43187 , \43188 , \43189 , \43190 ,
         \43191 , \43192 , \43193 , \43194 , \43195 , \43196 , \43197 , \43198 , \43199 , \43200 ,
         \43201 , \43202 , \43203 , \43204 , \43205 , \43206 , \43207 , \43208 , \43209 , \43210 ,
         \43211 , \43212 , \43213 , \43214 , \43215 , \43216 , \43217 , \43218 , \43219 , \43220 ,
         \43221 , \43222 , \43223 , \43224 , \43225 , \43226 , \43227 , \43228 , \43229 , \43230 ,
         \43231 , \43232 , \43233 , \43234 , \43235 , \43236 , \43237 , \43238 , \43239 , \43240 ,
         \43241 , \43242 , \43243 , \43244 , \43245 , \43246 , \43247 , \43248 , \43249 , \43250 ,
         \43251 , \43252 , \43253 , \43254 , \43255 , \43256 , \43257 , \43258 , \43259 , \43260 ,
         \43261 , \43262 , \43263 , \43264 , \43265 , \43266 , \43267 , \43268 , \43269 , \43270 ,
         \43271 , \43272 , \43273 , \43274 , \43275 , \43276 , \43277 , \43278 , \43279 , \43280 ,
         \43281 , \43282 , \43283 , \43284 , \43285 , \43286 , \43287 , \43288 , \43289 , \43290 ,
         \43291 , \43292 , \43293 , \43294 , \43295 , \43296 , \43297 , \43298 , \43299 , \43300 ,
         \43301 , \43302 , \43303 , \43304 , \43305 , \43306 , \43307 , \43308 , \43309 , \43310 ,
         \43311 , \43312 , \43313 , \43314 , \43315 , \43316 , \43317 , \43318 , \43319 , \43320 ,
         \43321 , \43322 , \43323 , \43324 , \43325 , \43326 , \43327 , \43328 , \43329 , \43330 ,
         \43331 , \43332 , \43333 , \43334 , \43335 , \43336 , \43337 , \43338 , \43339 , \43340 ,
         \43341 , \43342 , \43343 , \43344 , \43345 , \43346 , \43347 , \43348 , \43349 , \43350 ,
         \43351 , \43352 , \43353 , \43354 , \43355 , \43356 , \43357 , \43358 , \43359 , \43360 ,
         \43361 , \43362 , \43363 , \43364 , \43365 , \43366 , \43367 , \43368 , \43369 , \43370 ,
         \43371 , \43372 , \43373 , \43374 , \43375 , \43376 , \43377 , \43378 , \43379 , \43380 ,
         \43381 , \43382 , \43383 , \43384 , \43385 , \43386 , \43387 , \43388 , \43389 , \43390 ,
         \43391 , \43392 , \43393 , \43394 , \43395 , \43396 , \43397 , \43398 , \43399 , \43400 ,
         \43401 , \43402 , \43403 , \43404 , \43405 , \43406 , \43407 , \43408 , \43409 , \43410 ,
         \43411 , \43412 , \43413 , \43414 , \43415 , \43416 , \43417 , \43418 , \43419 , \43420 ,
         \43421 , \43422 , \43423 , \43424 , \43425 , \43426 , \43427 , \43428 , \43429 , \43430 ,
         \43431 , \43432 , \43433 , \43434 , \43435 , \43436 , \43437 , \43438 , \43439 , \43440 ,
         \43441 , \43442 , \43443 , \43444 , \43445 , \43446 , \43447 , \43448 , \43449 , \43450 ,
         \43451 , \43452 , \43453 , \43454 , \43455 , \43456 , \43457 , \43458 , \43459 , \43460 ,
         \43461 , \43462 , \43463 , \43464 , \43465 , \43466 , \43467 , \43468 , \43469 , \43470 ,
         \43471 , \43472 , \43473 , \43474 , \43475 , \43476 , \43477 , \43478 , \43479 , \43480 ,
         \43481 , \43482 , \43483 , \43484 , \43485 , \43486 , \43487 , \43488 , \43489 , \43490 ,
         \43491 , \43492 , \43493 , \43494 , \43495 , \43496 , \43497 , \43498 , \43499 , \43500 ,
         \43501 , \43502 , \43503 , \43504 , \43505 , \43506 , \43507 , \43508 , \43509 , \43510 ,
         \43511 , \43512 , \43513 , \43514 , \43515 , \43516 , \43517 , \43518 , \43519 , \43520 ,
         \43521 , \43522 , \43523 , \43524 , \43525 , \43526 , \43527 , \43528 , \43529 , \43530 ,
         \43531 , \43532 , \43533 , \43534 , \43535 , \43536 , \43537 , \43538 , \43539 , \43540 ,
         \43541 , \43542 , \43543 , \43544 , \43545 , \43546 , \43547 , \43548 , \43549 , \43550 ,
         \43551 , \43552 , \43553 , \43554 , \43555 , \43556 , \43557 , \43558 , \43559 , \43560 ,
         \43561 , \43562 , \43563 , \43564 , \43565 , \43566 , \43567 , \43568 , \43569 , \43570 ,
         \43571 , \43572 , \43573 , \43574 , \43575 , \43576 , \43577 , \43578 , \43579 , \43580 ,
         \43581 , \43582 , \43583 , \43584 , \43585 , \43586 , \43587 , \43588 , \43589 , \43590 ,
         \43591 , \43592 , \43593 , \43594 , \43595 , \43596 , \43597 , \43598 , \43599 , \43600 ,
         \43601 , \43602 , \43603 , \43604 , \43605 , \43606 , \43607 , \43608 , \43609 , \43610 ,
         \43611 , \43612 , \43613 , \43614 , \43615 , \43616 , \43617 , \43618 , \43619 , \43620 ,
         \43621 , \43622 , \43623 , \43624 , \43625 , \43626 , \43627 , \43628 , \43629 , \43630 ,
         \43631 , \43632 , \43633 , \43634 , \43635 , \43636 , \43637 , \43638 , \43639 , \43640 ,
         \43641 , \43642 , \43643 , \43644 , \43645 , \43646 , \43647 , \43648 , \43649 , \43650 ,
         \43651 , \43652 , \43653 , \43654 , \43655 , \43656 , \43657 , \43658 , \43659 , \43660 ,
         \43661 , \43662 , \43663 , \43664 , \43665 , \43666 , \43667 , \43668 , \43669 , \43670 ,
         \43671 , \43672 , \43673 , \43674 , \43675 , \43676 , \43677 , \43678 , \43679 , \43680 ,
         \43681 , \43682 , \43683 , \43684 , \43685 , \43686 , \43687 , \43688 , \43689 , \43690 ,
         \43691 , \43692 , \43693 , \43694 , \43695 , \43696 , \43697 , \43698 , \43699 , \43700 ,
         \43701 , \43702 , \43703 , \43704 , \43705 , \43706 , \43707 , \43708 , \43709 , \43710 ,
         \43711 , \43712 , \43713 , \43714 , \43715 , \43716 , \43717 , \43718 , \43719 , \43720 ,
         \43721 , \43722 , \43723 , \43724 , \43725 , \43726 , \43727 , \43728 , \43729 , \43730 ,
         \43731 , \43732 , \43733 , \43734 , \43735 , \43736 , \43737 , \43738 , \43739 , \43740 ,
         \43741 , \43742 , \43743 , \43744 , \43745 , \43746 , \43747 , \43748 , \43749 , \43750 ,
         \43751 , \43752 , \43753 , \43754 , \43755 , \43756 , \43757 , \43758 , \43759 , \43760 ,
         \43761 , \43762 , \43763 , \43764 , \43765 , \43766 , \43767 , \43768 , \43769 , \43770 ,
         \43771 , \43772 , \43773 , \43774 , \43775 , \43776 , \43777 , \43778 , \43779 , \43780 ,
         \43781 , \43782 , \43783 , \43784 , \43785 , \43786 , \43787 , \43788 , \43789 , \43790 ,
         \43791 , \43792 , \43793 , \43794 , \43795 , \43796 , \43797 , \43798 , \43799 , \43800 ,
         \43801 , \43802 , \43803 , \43804 , \43805 , \43806 , \43807 , \43808 , \43809 , \43810 ,
         \43811 , \43812 , \43813 , \43814 , \43815 , \43816 , \43817 , \43818 , \43819 , \43820 ,
         \43821 , \43822 , \43823 , \43824 , \43825 , \43826 , \43827 , \43828 , \43829 , \43830 ,
         \43831 , \43832 , \43833 , \43834 , \43835 , \43836 , \43837 , \43838 , \43839 , \43840 ,
         \43841 , \43842 , \43843 , \43844 , \43845 , \43846 , \43847 , \43848 , \43849 , \43850 ,
         \43851 , \43852 , \43853 , \43854 , \43855 , \43856 , \43857 , \43858 , \43859 , \43860 ,
         \43861 , \43862 , \43863 , \43864 , \43865 , \43866 , \43867 , \43868 , \43869 , \43870 ,
         \43871 , \43872 , \43873 , \43874 , \43875 , \43876 , \43877 , \43878 , \43879 , \43880 ,
         \43881 , \43882 , \43883 , \43884 , \43885 , \43886 , \43887 , \43888 , \43889 , \43890 ,
         \43891 , \43892 , \43893 , \43894 , \43895 , \43896 , \43897 , \43898 , \43899 , \43900 ,
         \43901 , \43902 , \43903 , \43904 , \43905 , \43906 , \43907 , \43908 , \43909 , \43910 ,
         \43911 , \43912 , \43913 , \43914 , \43915 , \43916 , \43917 , \43918 , \43919 , \43920 ,
         \43921 , \43922 , \43923 , \43924 , \43925 , \43926 , \43927 , \43928 , \43929 , \43930 ,
         \43931 , \43932 , \43933 , \43934 , \43935 , \43936 , \43937 , \43938 , \43939 , \43940 ,
         \43941 , \43942 , \43943 , \43944 , \43945 , \43946 , \43947 , \43948 , \43949 , \43950 ,
         \43951 , \43952 , \43953 , \43954 , \43955 , \43956 , \43957 , \43958 , \43959 , \43960 ,
         \43961 , \43962 , \43963 , \43964 , \43965 , \43966 , \43967 , \43968 , \43969 , \43970 ,
         \43971 , \43972 , \43973 , \43974 , \43975 , \43976 , \43977 , \43978 , \43979 , \43980 ,
         \43981 , \43982 , \43983 , \43984 , \43985 , \43986 , \43987 , \43988 , \43989 , \43990 ,
         \43991 , \43992 , \43993 , \43994 , \43995 , \43996 , \43997 , \43998 , \43999 , \44000 ,
         \44001 , \44002 , \44003 , \44004 , \44005 , \44006 , \44007 , \44008 , \44009 , \44010 ,
         \44011 , \44012 , \44013 , \44014 , \44015 , \44016 , \44017 , \44018 , \44019 , \44020 ,
         \44021 , \44022 , \44023 , \44024 , \44025 , \44026 , \44027 , \44028 , \44029 , \44030 ,
         \44031 , \44032 , \44033 , \44034 , \44035 , \44036 , \44037 , \44038 , \44039 , \44040 ,
         \44041 , \44042 , \44043 , \44044 , \44045 , \44046 , \44047 , \44048 , \44049 , \44050 ,
         \44051 , \44052 , \44053 , \44054 , \44055 , \44056 , \44057 , \44058 , \44059 , \44060 ,
         \44061 , \44062 , \44063 , \44064 , \44065 , \44066 , \44067 , \44068 , \44069 , \44070 ,
         \44071 , \44072 , \44073 , \44074 , \44075 , \44076 , \44077 , \44078 , \44079 , \44080 ,
         \44081 , \44082 , \44083 , \44084 , \44085 , \44086 , \44087 , \44088 , \44089 , \44090 ,
         \44091 , \44092 , \44093 , \44094 , \44095 , \44096 , \44097 , \44098 , \44099 , \44100 ,
         \44101 , \44102 , \44103 , \44104 , \44105 , \44106 , \44107 , \44108 , \44109 , \44110 ,
         \44111 , \44112 , \44113 , \44114 , \44115 , \44116 , \44117 , \44118 , \44119 , \44120 ,
         \44121 , \44122 , \44123 , \44124 , \44125 , \44126 , \44127 , \44128 , \44129 , \44130 ,
         \44131 , \44132 , \44133 , \44134 , \44135 , \44136 , \44137 , \44138 , \44139 , \44140 ,
         \44141 , \44142 , \44143 , \44144 , \44145 , \44146 , \44147 , \44148 , \44149 , \44150 ,
         \44151 , \44152 , \44153 , \44154 , \44155 , \44156 , \44157 , \44158 , \44159 , \44160 ,
         \44161 , \44162 , \44163 , \44164 , \44165 , \44166 , \44167 , \44168 , \44169 , \44170 ,
         \44171 , \44172 , \44173 , \44174 , \44175 , \44176 , \44177 , \44178 , \44179 , \44180 ,
         \44181 , \44182 , \44183 , \44184 , \44185 , \44186 , \44187 , \44188 , \44189 , \44190 ,
         \44191 , \44192 , \44193 , \44194 , \44195 , \44196 , \44197 , \44198 , \44199 , \44200 ,
         \44201 , \44202 , \44203 , \44204 , \44205 , \44206 , \44207 , \44208 , \44209 , \44210 ,
         \44211 , \44212 , \44213 , \44214 , \44215 , \44216 , \44217 , \44218 , \44219 , \44220 ,
         \44221 , \44222 , \44223 , \44224 , \44225 , \44226 , \44227 , \44228 , \44229 , \44230 ,
         \44231 , \44232 , \44233 , \44234 , \44235 , \44236 , \44237 , \44238 , \44239 , \44240 ,
         \44241 , \44242 , \44243 , \44244 , \44245 , \44246 , \44247 , \44248 , \44249 , \44250 ,
         \44251 , \44252 , \44253 , \44254 , \44255 , \44256 , \44257 , \44258 , \44259 , \44260 ,
         \44261 , \44262 , \44263 , \44264 , \44265 , \44266 , \44267 , \44268 , \44269 , \44270 ,
         \44271 , \44272 , \44273 , \44274 , \44275 , \44276 , \44277 , \44278 , \44279 , \44280 ,
         \44281 , \44282 , \44283 , \44284 , \44285 , \44286 , \44287 , \44288 , \44289 , \44290 ,
         \44291 , \44292 , \44293 , \44294 , \44295 , \44296 , \44297 , \44298 , \44299 , \44300 ,
         \44301 , \44302 , \44303 , \44304 , \44305 , \44306 , \44307 , \44308 , \44309 , \44310 ,
         \44311 , \44312 , \44313 , \44314 , \44315 , \44316 , \44317 , \44318 , \44319 , \44320 ,
         \44321 , \44322 , \44323 , \44324 , \44325 , \44326 , \44327 , \44328 , \44329 , \44330 ,
         \44331 , \44332 , \44333 , \44334 , \44335 , \44336 , \44337 , \44338 , \44339 , \44340 ,
         \44341 , \44342 , \44343 , \44344 , \44345 , \44346 , \44347 , \44348 , \44349 , \44350 ,
         \44351 , \44352 , \44353 , \44354 , \44355 , \44356 , \44357 , \44358 , \44359 , \44360 ,
         \44361 , \44362 , \44363 , \44364 , \44365 , \44366 , \44367 , \44368 , \44369 , \44370 ,
         \44371 , \44372 , \44373 , \44374 , \44375 , \44376 , \44377 , \44378 , \44379 , \44380 ,
         \44381 , \44382 , \44383 , \44384 , \44385 , \44386 , \44387 , \44388 , \44389 , \44390 ,
         \44391 , \44392 , \44393 , \44394 , \44395 , \44396 , \44397 , \44398 , \44399 , \44400 ,
         \44401 , \44402 , \44403 , \44404 , \44405 , \44406 , \44407 , \44408 , \44409 , \44410 ,
         \44411 , \44412 , \44413 , \44414 , \44415 , \44416 , \44417 , \44418 , \44419 , \44420 ,
         \44421 , \44422 , \44423 , \44424 , \44425 , \44426 , \44427 , \44428 , \44429 , \44430 ,
         \44431 , \44432 , \44433 , \44434 , \44435 , \44436 , \44437 , \44438 , \44439 , \44440 ,
         \44441 , \44442 , \44443 , \44444 , \44445 , \44446 , \44447 , \44448 , \44449 , \44450 ,
         \44451 , \44452 , \44453 , \44454 , \44455 , \44456 , \44457 , \44458 , \44459 , \44460 ,
         \44461 , \44462 , \44463 , \44464 , \44465 , \44466 , \44467 , \44468 , \44469 , \44470 ,
         \44471 , \44472 , \44473 , \44474 , \44475 , \44476 , \44477 , \44478 , \44479 , \44480 ,
         \44481 , \44482 , \44483 , \44484 , \44485 , \44486 , \44487 , \44488 , \44489 , \44490 ,
         \44491 , \44492 , \44493 , \44494 , \44495 , \44496 , \44497 , \44498 , \44499 , \44500 ,
         \44501 , \44502 , \44503 , \44504 , \44505 , \44506 , \44507 , \44508 , \44509 , \44510 ,
         \44511 , \44512 , \44513 , \44514 , \44515 , \44516 , \44517 , \44518 , \44519 , \44520 ,
         \44521 , \44522 , \44523 , \44524 , \44525 , \44526 , \44527 , \44528 , \44529 , \44530 ,
         \44531 , \44532 , \44533 , \44534 , \44535 , \44536 , \44537 , \44538 , \44539 , \44540 ,
         \44541 , \44542 , \44543 , \44544 , \44545 , \44546 , \44547 , \44548 , \44549 , \44550 ,
         \44551 , \44552 , \44553 , \44554 , \44555 , \44556 , \44557 , \44558 , \44559 , \44560 ,
         \44561 , \44562 , \44563 , \44564 , \44565 , \44566 , \44567 , \44568 , \44569 , \44570 ,
         \44571 , \44572 , \44573 , \44574 , \44575 , \44576 , \44577 , \44578 , \44579 , \44580 ,
         \44581 , \44582 , \44583 , \44584 , \44585 , \44586 , \44587 , \44588 , \44589 , \44590 ,
         \44591 , \44592 , \44593 , \44594 , \44595 , \44596 , \44597 , \44598 , \44599 , \44600 ,
         \44601 , \44602 , \44603 , \44604 , \44605 , \44606 , \44607 , \44608 , \44609 , \44610 ,
         \44611 , \44612 , \44613 , \44614 , \44615 , \44616 , \44617 , \44618 , \44619 , \44620 ,
         \44621 , \44622 , \44623 , \44624 , \44625 , \44626 , \44627 , \44628 , \44629 , \44630 ,
         \44631 , \44632 , \44633 , \44634 , \44635 , \44636 , \44637 , \44638 , \44639 , \44640 ,
         \44641 , \44642 , \44643 , \44644 , \44645 , \44646 , \44647 , \44648 , \44649 , \44650 ,
         \44651 , \44652 , \44653 , \44654 , \44655 , \44656 , \44657 , \44658 , \44659 , \44660 ,
         \44661 , \44662 , \44663 , \44664 , \44665 , \44666 , \44667 , \44668 , \44669 , \44670 ,
         \44671 , \44672 , \44673 , \44674 , \44675 , \44676 , \44677 , \44678 , \44679 , \44680 ,
         \44681 , \44682 , \44683 , \44684 , \44685 , \44686 , \44687 , \44688 , \44689 , \44690 ,
         \44691 , \44692 , \44693 , \44694 , \44695 , \44696 , \44697 , \44698 , \44699 , \44700 ,
         \44701 , \44702 , \44703 , \44704 , \44705 , \44706 , \44707 , \44708 , \44709 , \44710 ,
         \44711 , \44712 , \44713 , \44714 , \44715 , \44716 , \44717 , \44718 , \44719 , \44720 ,
         \44721 , \44722 , \44723 , \44724 , \44725 , \44726 , \44727 , \44728 , \44729 , \44730 ,
         \44731 , \44732 , \44733 , \44734 , \44735 , \44736 , \44737 , \44738 , \44739 , \44740 ,
         \44741 , \44742 , \44743 , \44744 , \44745 , \44746 , \44747 , \44748 , \44749 , \44750 ,
         \44751 , \44752 , \44753 , \44754 , \44755 , \44756 , \44757 , \44758 , \44759 , \44760 ,
         \44761 , \44762 , \44763 , \44764 , \44765 , \44766 , \44767 , \44768 , \44769 , \44770 ,
         \44771 , \44772 , \44773 , \44774 , \44775 , \44776 , \44777 , \44778 , \44779 , \44780 ,
         \44781 , \44782 , \44783 , \44784 , \44785 , \44786 , \44787 , \44788 , \44789 , \44790 ,
         \44791 , \44792 , \44793 , \44794 , \44795 , \44796 , \44797 , \44798 , \44799 , \44800 ,
         \44801 , \44802 , \44803 , \44804 , \44805 , \44806 , \44807 , \44808 , \44809 , \44810 ,
         \44811 , \44812 , \44813 , \44814 , \44815 , \44816 , \44817 , \44818 , \44819 , \44820 ,
         \44821 , \44822 , \44823 , \44824 , \44825 , \44826 , \44827 , \44828 , \44829 , \44830 ,
         \44831 , \44832 , \44833 , \44834 , \44835 , \44836 , \44837 , \44838 , \44839 , \44840 ,
         \44841 , \44842 , \44843 , \44844 , \44845 , \44846 , \44847 , \44848 , \44849 , \44850 ,
         \44851 , \44852 , \44853 , \44854 , \44855 , \44856 , \44857 , \44858 , \44859 , \44860 ,
         \44861 , \44862 , \44863 , \44864 , \44865 , \44866 , \44867 , \44868 , \44869 , \44870 ,
         \44871 , \44872 , \44873 , \44874 , \44875 , \44876 , \44877 , \44878 , \44879 , \44880 ,
         \44881 , \44882 , \44883 , \44884 , \44885 , \44886 , \44887 , \44888 , \44889 , \44890 ,
         \44891 , \44892 , \44893 , \44894 , \44895 , \44896 , \44897 , \44898 , \44899 , \44900 ,
         \44901 , \44902 , \44903 , \44904 , \44905 , \44906 , \44907 , \44908 , \44909 , \44910 ,
         \44911 , \44912 , \44913 , \44914 , \44915 , \44916 , \44917 , \44918 , \44919 , \44920 ,
         \44921 , \44922 , \44923 , \44924 , \44925 , \44926 , \44927 , \44928 , \44929 , \44930 ,
         \44931 , \44932 , \44933 , \44934 , \44935 , \44936 , \44937 , \44938 , \44939 , \44940 ,
         \44941 , \44942 , \44943 , \44944 , \44945 , \44946 , \44947 , \44948 , \44949 , \44950 ,
         \44951 , \44952 , \44953 , \44954 , \44955 , \44956 , \44957 , \44958 , \44959 , \44960 ,
         \44961 , \44962 , \44963 , \44964 , \44965 , \44966 , \44967 , \44968 , \44969 , \44970 ,
         \44971 , \44972 , \44973 , \44974 , \44975 , \44976 , \44977 , \44978 , \44979 , \44980 ,
         \44981 , \44982 , \44983 , \44984 , \44985 , \44986 , \44987 , \44988 , \44989 , \44990 ,
         \44991 , \44992 , \44993 , \44994 , \44995 , \44996 , \44997 , \44998 , \44999 , \45000 ,
         \45001 , \45002 , \45003 , \45004 , \45005 , \45006 , \45007 , \45008 , \45009 , \45010 ,
         \45011 , \45012 , \45013 , \45014 , \45015 , \45016 , \45017 , \45018 , \45019 , \45020 ,
         \45021 , \45022 , \45023 , \45024 , \45025 , \45026 , \45027 , \45028 , \45029 , \45030 ,
         \45031 , \45032 , \45033 , \45034 , \45035 , \45036 , \45037 , \45038 , \45039 , \45040 ,
         \45041 , \45042 , \45043 , \45044 , \45045 , \45046 , \45047 , \45048 , \45049 , \45050 ,
         \45051 , \45052 , \45053 , \45054 , \45055 , \45056 , \45057 , \45058 , \45059 , \45060 ,
         \45061 , \45062 , \45063 , \45064 , \45065 , \45066 , \45067 , \45068 , \45069 , \45070 ,
         \45071 , \45072 , \45073 , \45074 , \45075 , \45076 , \45077 , \45078 , \45079 , \45080 ,
         \45081 , \45082 , \45083 , \45084 , \45085 , \45086 , \45087 , \45088 , \45089 , \45090 ,
         \45091 , \45092 , \45093 , \45094 , \45095 , \45096 , \45097 , \45098 , \45099 , \45100 ,
         \45101 , \45102 , \45103 , \45104 , \45105 , \45106 , \45107 , \45108 , \45109 , \45110 ,
         \45111 , \45112 , \45113 , \45114 , \45115 , \45116 , \45117 , \45118 , \45119 , \45120 ,
         \45121 , \45122 , \45123 , \45124 , \45125 , \45126 , \45127 , \45128 , \45129 , \45130 ,
         \45131 , \45132 , \45133 , \45134 , \45135 , \45136 , \45137 , \45138 , \45139 , \45140 ,
         \45141 , \45142 , \45143 , \45144 , \45145 , \45146 , \45147 , \45148 , \45149 , \45150 ,
         \45151 , \45152 , \45153 , \45154 , \45155 , \45156 , \45157 , \45158 , \45159 , \45160 ,
         \45161 , \45162 , \45163 , \45164 , \45165 , \45166 , \45167 , \45168 , \45169 , \45170 ,
         \45171 , \45172 , \45173 , \45174 , \45175 , \45176 , \45177 , \45178 , \45179 , \45180 ,
         \45181 , \45182 , \45183 , \45184 , \45185 , \45186 , \45187 , \45188 , \45189 , \45190 ,
         \45191 , \45192 , \45193 , \45194 , \45195 , \45196 , \45197 , \45198 , \45199 , \45200 ,
         \45201 , \45202 , \45203 , \45204 , \45205 , \45206 , \45207 , \45208 , \45209 , \45210 ,
         \45211 , \45212 , \45213 , \45214 , \45215 , \45216 , \45217 , \45218 , \45219 , \45220 ,
         \45221 , \45222 , \45223 , \45224 , \45225 , \45226 , \45227 , \45228 , \45229 , \45230 ,
         \45231 , \45232 , \45233 , \45234 , \45235 , \45236 , \45237 , \45238 , \45239 , \45240 ,
         \45241 , \45242 , \45243 , \45244 , \45245 , \45246 , \45247 , \45248 , \45249 , \45250 ,
         \45251 , \45252 , \45253 , \45254 , \45255 , \45256 , \45257 , \45258 , \45259 , \45260 ,
         \45261 , \45262 , \45263 , \45264 , \45265 , \45266 , \45267 , \45268 , \45269 , \45270 ,
         \45271 , \45272 , \45273 , \45274 , \45275 , \45276 , \45277 , \45278 , \45279 , \45280 ,
         \45281 , \45282 , \45283 , \45284 , \45285 , \45286 , \45287 , \45288 , \45289 , \45290 ,
         \45291 , \45292 , \45293 , \45294 , \45295 , \45296 , \45297 , \45298 , \45299 , \45300 ,
         \45301 , \45302 , \45303 , \45304 , \45305 , \45306 , \45307 , \45308 , \45309 , \45310 ,
         \45311 , \45312 , \45313 , \45314 , \45315 , \45316 , \45317 , \45318 , \45319 , \45320 ,
         \45321 , \45322 , \45323 , \45324 , \45325 , \45326 , \45327 , \45328 , \45329 , \45330 ,
         \45331 , \45332 , \45333 , \45334 , \45335 , \45336 , \45337 , \45338 , \45339 , \45340 ,
         \45341 , \45342 , \45343 , \45344 , \45345 , \45346 , \45347 , \45348 , \45349 , \45350 ,
         \45351 , \45352 , \45353 , \45354 , \45355 , \45356 , \45357 , \45358 , \45359 , \45360 ,
         \45361 , \45362 , \45363 , \45364 , \45365 , \45366 , \45367 , \45368 , \45369 , \45370 ,
         \45371 , \45372 , \45373 , \45374 , \45375 , \45376 , \45377 , \45378 , \45379 , \45380 ,
         \45381 , \45382 , \45383 , \45384 , \45385 , \45386 , \45387 , \45388 , \45389 , \45390 ,
         \45391 , \45392 , \45393 , \45394 , \45395 , \45396 , \45397 , \45398 , \45399 , \45400 ,
         \45401 , \45402 , \45403 , \45404 , \45405 , \45406 , \45407 , \45408 , \45409 , \45410 ,
         \45411 , \45412 , \45413 , \45414 , \45415 , \45416 , \45417 , \45418 , \45419 , \45420 ,
         \45421 , \45422 , \45423 , \45424 , \45425 , \45426 , \45427 , \45428 , \45429 , \45430 ,
         \45431 , \45432 , \45433 , \45434 , \45435 , \45436 , \45437 , \45438 , \45439 , \45440 ,
         \45441 , \45442 , \45443 , \45444 , \45445 , \45446 , \45447 , \45448 , \45449 , \45450 ,
         \45451 , \45452 , \45453 , \45454 , \45455 , \45456 , \45457 , \45458 , \45459 , \45460 ,
         \45461 , \45462 , \45463 , \45464 , \45465 , \45466 , \45467 , \45468 , \45469 , \45470 ,
         \45471 , \45472 , \45473 , \45474 , \45475 , \45476 , \45477 , \45478 , \45479 , \45480 ,
         \45481 , \45482 , \45483 , \45484 , \45485 , \45486 , \45487 , \45488 , \45489 , \45490 ,
         \45491 , \45492 ;
buf \U$labajz4591 ( R_101_8a8e950, \44291 );
buf \U$labajz4592 ( R_102_8a8f868, \44319 );
buf \U$labajz4593 ( R_103_8a8f910, \44329 );
buf \U$labajz4594 ( R_104_8a8f9b8, \44342 );
buf \U$labajz4595 ( R_105_8a8fa60, \44356 );
buf \U$labajz4596 ( R_106_8a8fb08, \44378 );
buf \U$labajz4597 ( R_107_8a8fbb0, \44386 );
buf \U$labajz4598 ( R_108_8a8fc58, \44400 );
buf \U$labajz4599 ( R_109_8a8fd00, \44413 );
buf \U$labajz4600 ( R_10a_8a8fda8, \44443 );
buf \U$labajz4601 ( R_10b_8a8fe50, \44457 );
buf \U$labajz4602 ( R_10c_8a8fef8, \44466 );
buf \U$labajz4603 ( R_10d_8a8ffa0, \44487 );
buf \U$labajz4604 ( R_10e_8a90048, \44502 );
buf \U$labajz4605 ( R_10f_8a900f0, \44508 );
buf \U$labajz4606 ( R_110_8a90198, \44528 );
buf \U$labajz4607 ( R_111_8a90240, \44548 );
buf \U$labajz4608 ( R_112_8a902e8, \44553 );
buf \U$labajz4609 ( R_113_8a90390, \44567 );
buf \U$labajz4610 ( R_114_8a90438, \44582 );
buf \U$labajz4611 ( R_115_8a904e0, \44587 );
buf \U$labajz4612 ( R_116_8a90588, \44621 );
buf \U$labajz4613 ( R_117_8a90630, \44629 );
buf \U$labajz4614 ( R_118_8a906d8, \44645 );
buf \U$labajz4615 ( R_119_8a90780, \44658 );
buf \U$labajz4616 ( R_11a_8a90828, \44666 );
buf \U$labajz4617 ( R_11b_8a908d0, \44687 );
buf \U$labajz4618 ( R_11c_8a90978, \44705 );
buf \U$labajz4619 ( R_11d_8a90a20, \44727 );
buf \U$labajz4620 ( R_11e_8a90ac8, \44731 );
buf \U$labajz4621 ( R_11f_8a90b70, \44741 );
buf \U$labajz4622 ( R_120_8a90c18, \44749 );
buf \U$labajz4623 ( R_121_8a90cc0, \44790 );
buf \U$labajz4624 ( R_122_8a90d68, \44806 );
buf \U$labajz4625 ( R_123_8a90e10, \44817 );
buf \U$labajz4626 ( R_124_8a90eb8, \44837 );
buf \U$labajz4627 ( R_125_8a90f60, \44847 );
buf \U$labajz4628 ( R_126_8a91008, \44862 );
buf \U$labajz4629 ( R_127_8a910b0, \44872 );
buf \U$labajz4630 ( R_128_8a91158, \44898 );
buf \U$labajz4631 ( R_129_8a91200, \44910 );
buf \U$labajz4632 ( R_12a_8a912a8, \44924 );
buf \U$labajz4633 ( R_12b_8a91350, \44936 );
buf \U$labajz4634 ( R_12c_8a913f8, \44958 );
buf \U$labajz4635 ( R_12d_8a914a0, \44968 );
buf \U$labajz4636 ( R_12e_8a91548, \44980 );
buf \U$labajz4637 ( R_12f_8a915f0, \44993 );
buf \U$labajz4638 ( R_130_8a91698, \45022 );
buf \U$labajz4639 ( R_131_8a91740, \45032 );
buf \U$labajz4640 ( R_132_8a917e8, \45047 );
buf \U$labajz4641 ( R_133_8a91890, \45057 );
buf \U$labajz4642 ( R_134_8a91938, \45080 );
buf \U$labajz4643 ( R_135_8a919e0, \45090 );
buf \U$labajz4644 ( R_136_8a91a88, \45105 );
buf \U$labajz4645 ( R_137_8a91b30, \45115 );
buf \U$labajz4646 ( R_138_8a91bd8, \45141 );
buf \U$labajz4647 ( R_139_8a91c80, \45151 );
buf \U$labajz4648 ( R_13a_8a91d28, \45164 );
buf \U$labajz4649 ( R_13b_8a91dd0, \45174 );
buf \U$labajz4650 ( R_13c_8a91e78, \45195 );
buf \U$labajz4651 ( R_13d_8a91f20, \45205 );
buf \U$labajz4652 ( R_13e_8a91fc8, \45219 );
buf \U$labajz4653 ( R_13f_8a92070, \45226 );
buf \U$labajz4654 ( R_140_8a92118, \45247 );
buf \U$labajz4655 ( R_141_8a921c0, \45258 );
buf \U$labajz4656 ( R_142_8a92268, \45274 );
buf \U$labajz4657 ( R_143_8a92310, \45285 );
buf \U$labajz4658 ( R_144_8a923b8, \45304 );
buf \U$labajz4659 ( R_145_8a92460, \45314 );
buf \U$labajz4660 ( R_146_8a92508, \45325 );
buf \U$labajz4661 ( R_147_8a925b0, \45333 );
buf \U$labajz4662 ( R_148_8a92658, \45353 );
buf \U$labajz4663 ( R_149_8a92700, \45365 );
buf \U$labajz4664 ( R_14a_8a927a8, \45382 );
buf \U$labajz4665 ( R_14b_8a92850, \45389 );
buf \U$labajz4666 ( R_14c_8a928f8, \45411 );
buf \U$labajz4667 ( R_14d_8a929a0, \45422 );
buf \U$labajz4668 ( R_14e_8a92a48, \45437 );
buf \U$labajz4669 ( R_14f_8a92af0, \45444 );
buf \U$labajz4670 ( R_150_8a92b98, \45456 );
buf \U$labajz4671 ( R_151_8a92c40, \45462 );
buf \U$labajz4672 ( R_152_8a92ce8, \45468 );
buf \U$labajz4673 ( R_153_8a92d90, \45474 );
buf \U$labajz4674 ( R_154_8a92e38, \45480 );
buf \U$labajz4675 ( R_155_8a92ee0, \45492 );
or \U$1 ( \344 , RI986e350_15, RI986e3c8_16);
not \U$2 ( \345 , \344 );
or \U$3 ( \346 , RI986e260_13, RI986e2d8_14);
not \U$4 ( \347 , \346 );
or \U$5 ( \348 , RI986e080_9, RI986e0f8_10);
not \U$6 ( \349 , \348 );
or \U$7 ( \350 , RI986e170_11, RI986e1e8_12);
not \U$8 ( \351 , \350 );
or \U$9 ( \352 , RI986dcc0_1, RI986dd38_2);
not \U$10 ( \353 , \352 );
not \U$11 ( \354 , RI986dea0_5);
not \U$12 ( \355 , RI986df18_6);
or \U$13 ( \356 , \354 , \355 );
nor \U$14 ( \357 , RI986dea0_5, RI986df18_6);
nand \U$15 ( \358 , RI986df90_7, RI986e008_8);
or \U$16 ( \359 , \357 , \358 );
nand \U$17 ( \360 , \356 , \359 );
not \U$18 ( \361 , \360 );
or \U$19 ( \362 , RI986de28_4, RI986ddb0_3);
not \U$20 ( \363 , \362 );
or \U$21 ( \364 , \361 , \363 );
nand \U$22 ( \365 , RI986ddb0_3, RI986de28_4);
nand \U$23 ( \366 , \364 , \365 );
not \U$24 ( \367 , \366 );
or \U$25 ( \368 , \353 , \367 );
nand \U$26 ( \369 , RI986dcc0_1, RI986dd38_2);
nand \U$27 ( \370 , \368 , \369 );
not \U$28 ( \371 , \370 );
or \U$29 ( \372 , \351 , \371 );
nand \U$30 ( \373 , RI986e170_11, RI986e1e8_12);
nand \U$31 ( \374 , \372 , \373 );
not \U$32 ( \375 , \374 );
or \U$33 ( \376 , \349 , \375 );
nand \U$34 ( \377 , RI986e080_9, RI986e0f8_10);
nand \U$35 ( \378 , \376 , \377 );
not \U$36 ( \379 , \378 );
or \U$37 ( \380 , \347 , \379 );
nand \U$38 ( \381 , RI986e260_13, RI986e2d8_14);
nand \U$39 ( \382 , \380 , \381 );
not \U$40 ( \383 , \382 );
nor \U$41 ( \384 , RI986ef80_41, RI986eff8_42);
nor \U$42 ( \385 , RI986f070_43, RI986f0e8_44);
nor \U$43 ( \386 , \384 , \385 );
or \U$44 ( \387 , RI986f250_47, RI986f2c8_48);
or \U$45 ( \388 , RI986f160_45, RI986f1d8_46);
and \U$46 ( \389 , \386 , \387 , \388 );
not \U$47 ( \390 , \389 );
not \U$48 ( \391 , RI986e878_26);
not \U$49 ( \392 , RI986e800_25);
or \U$50 ( \393 , \391 , \392 );
nor \U$51 ( \394 , RI986e9e0_29, RI986ea58_30);
nand \U$52 ( \395 , RI986ead0_31, RI986eb48_32);
or \U$53 ( \396 , \394 , \395 );
nand \U$54 ( \397 , RI986e9e0_29, RI986ea58_30);
nand \U$55 ( \398 , \396 , \397 );
nand \U$56 ( \399 , RI986e8f0_27, RI986e968_28);
not \U$57 ( \400 , \399 );
or \U$58 ( \401 , \398 , \400 );
not \U$59 ( \402 , RI986e800_25);
not \U$60 ( \403 , RI986e878_26);
and \U$61 ( \404 , \402 , \403 );
nor \U$62 ( \405 , RI986e8f0_27, RI986e968_28);
nor \U$63 ( \406 , \404 , \405 );
nand \U$64 ( \407 , \401 , \406 );
nand \U$65 ( \408 , \393 , \407 );
or \U$66 ( \409 , RI986ebc0_33, RI986ec38_34);
or \U$67 ( \410 , RI986ecb0_35, RI986ed28_36);
or \U$68 ( \411 , RI986eda0_37, RI986ee18_38);
not \U$69 ( \412 , RI986ee90_39);
not \U$70 ( \413 , RI986ef08_40);
nand \U$71 ( \414 , \412 , \413 );
and \U$72 ( \415 , \409 , \410 , \411 , \414 );
nand \U$73 ( \416 , \408 , \415 );
not \U$74 ( \417 , \409 );
nor \U$75 ( \418 , RI986eda0_37, RI986ee18_38);
nand \U$76 ( \419 , RI986ee90_39, RI986ef08_40);
or \U$77 ( \420 , \418 , \419 );
nand \U$78 ( \421 , RI986eda0_37, RI986ee18_38);
nand \U$79 ( \422 , \420 , \421 );
not \U$80 ( \423 , \422 );
or \U$81 ( \424 , \417 , \423 );
nand \U$82 ( \425 , RI986ebc0_33, RI986ec38_34);
nand \U$83 ( \426 , \424 , \425 );
nand \U$84 ( \427 , \426 , \410 );
nand \U$85 ( \428 , RI986ecb0_35, RI986ed28_36);
nand \U$86 ( \429 , \416 , \427 , \428 );
not \U$87 ( \430 , \429 );
or \U$88 ( \431 , \390 , \430 );
not \U$89 ( \432 , \388 );
not \U$90 ( \433 , \387 );
nand \U$91 ( \434 , RI986f070_43, RI986f0e8_44);
or \U$92 ( \435 , \384 , \434 );
nand \U$93 ( \436 , RI986ef80_41, RI986eff8_42);
nand \U$94 ( \437 , \435 , \436 );
not \U$95 ( \438 , \437 );
or \U$96 ( \439 , \433 , \438 );
nand \U$97 ( \440 , RI986f250_47, RI986f2c8_48);
nand \U$98 ( \441 , \439 , \440 );
not \U$99 ( \442 , \441 );
or \U$100 ( \443 , \432 , \442 );
nand \U$101 ( \444 , RI986f160_45, RI986f1d8_46);
nand \U$102 ( \445 , \443 , \444 );
not \U$103 ( \446 , \445 );
nand \U$104 ( \447 , \431 , \446 );
or \U$105 ( \448 , RI986e710_23, RI986e788_24);
or \U$106 ( \449 , RI986e620_21, RI986e698_22);
nand \U$107 ( \450 , \448 , \449 );
or \U$108 ( \451 , RI986e530_19, RI986e5a8_20);
or \U$109 ( \452 , RI986e440_17, RI986e4b8_18);
nand \U$110 ( \453 , \451 , \452 );
nor \U$111 ( \454 , \450 , \453 );
buf \U$112 ( \455 , \454 );
nand \U$113 ( \456 , \447 , \455 );
not \U$114 ( \457 , \456 );
not \U$115 ( \458 , RI986ffe8_76);
not \U$116 ( \459 , RI986ff70_75);
nand \U$117 ( \460 , \458 , \459 );
not \U$118 ( \461 , RI9870060_77);
not \U$119 ( \462 , RI98700d8_78);
nand \U$120 ( \463 , \461 , \462 );
not \U$121 ( \464 , RI986fe80_73);
not \U$122 ( \465 , RI986fef8_74);
nand \U$123 ( \466 , \464 , \465 );
not \U$124 ( \467 , RI9870150_79);
not \U$125 ( \468 , RI98701c8_80);
nand \U$126 ( \469 , \467 , \468 );
nand \U$127 ( \470 , \460 , \463 , \466 , \469 );
not \U$128 ( \471 , \470 );
not \U$129 ( \472 , \471 );
not \U$130 ( \473 , RI986fca0_69);
not \U$131 ( \474 , RI986fd18_70);
nand \U$132 ( \475 , \473 , \474 );
not \U$133 ( \476 , \475 );
nor \U$134 ( \477 , RI986fd90_71, RI986fe08_72);
not \U$135 ( \478 , \477 );
not \U$136 ( \479 , \478 );
nor \U$137 ( \480 , \476 , \479 );
not \U$138 ( \481 , \480 );
or \U$139 ( \482 , RI986fbb0_67, RI986fc28_68);
nand \U$140 ( \483 , \482 , RI986fac0_65, RI986fb38_66);
nand \U$141 ( \484 , RI986fbb0_67, RI986fc28_68);
nand \U$142 ( \485 , \483 , \484 );
not \U$143 ( \486 , \485 );
or \U$144 ( \487 , \481 , \486 );
nand \U$145 ( \488 , RI986fd90_71, RI986fe08_72);
not \U$146 ( \489 , \488 );
and \U$147 ( \490 , \475 , \489 );
and \U$148 ( \491 , RI986fca0_69, RI986fd18_70);
nor \U$149 ( \492 , \490 , \491 );
nand \U$150 ( \493 , \487 , \492 );
not \U$151 ( \494 , \493 );
or \U$152 ( \495 , \472 , \494 );
nor \U$153 ( \496 , RI9870240_81, RI98702b8_82);
nor \U$154 ( \497 , RI9870330_83, RI98703a8_84);
nor \U$155 ( \498 , \496 , \497 );
not \U$156 ( \499 , \498 );
nand \U$157 ( \500 , RI9870420_85, RI9870498_86);
nor \U$158 ( \501 , RI9870510_87, RI9870588_88);
or \U$159 ( \502 , \500 , \501 );
nand \U$160 ( \503 , RI9870510_87, RI9870588_88);
nand \U$161 ( \504 , \502 , \503 );
not \U$162 ( \505 , \504 );
or \U$163 ( \506 , \499 , \505 );
not \U$164 ( \507 , RI9870240_81);
not \U$165 ( \508 , RI98702b8_82);
nand \U$166 ( \509 , \507 , \508 );
nand \U$167 ( \510 , RI9870330_83, RI98703a8_84);
not \U$168 ( \511 , \510 );
and \U$169 ( \512 , \509 , \511 );
nor \U$170 ( \513 , \507 , \508 );
nor \U$171 ( \514 , \512 , \513 );
nand \U$172 ( \515 , \506 , \514 );
nor \U$173 ( \516 , RI986fbb0_67, RI986fc28_68);
not \U$174 ( \517 , \516 );
nor \U$175 ( \518 , RI986fac0_65, RI986fb38_66);
not \U$176 ( \519 , \518 );
not \U$177 ( \520 , RI986fca0_69);
nand \U$178 ( \521 , \520 , \474 );
nand \U$179 ( \522 , \517 , \519 , \478 , \521 );
not \U$180 ( \523 , \522 );
not \U$181 ( \524 , RI98707e0_93);
not \U$182 ( \525 , RI9870858_94);
nand \U$183 ( \526 , \524 , \525 );
nor \U$184 ( \527 , RI9870600_89, RI9870678_90);
not \U$185 ( \528 , \527 );
nor \U$186 ( \529 , RI98708d0_95, RI9870948_96);
not \U$187 ( \530 , \529 );
not \U$188 ( \531 , RI9870768_92);
not \U$189 ( \532 , RI98706f0_91);
nand \U$190 ( \533 , \531 , \532 );
and \U$191 ( \534 , \526 , \528 , \530 , \533 );
nand \U$192 ( \535 , \515 , \523 , \534 , \471 );
nand \U$193 ( \536 , \495 , \535 );
nor \U$194 ( \537 , RI9871050_111, RI98710c8_112);
nor \U$195 ( \538 , RI9870e70_107, RI9870ee8_108);
nor \U$196 ( \539 , RI9870ba0_101, RI9870c18_102);
nor \U$197 ( \540 , \537 , \538 , \539 );
nor \U$198 ( \541 , RI9870f60_109, RI9870fd8_110);
nor \U$199 ( \542 , RI9870ab0_99, RI9870b28_100);
nor \U$200 ( \543 , \541 , \542 );
nor \U$201 ( \544 , RI98709c0_97, RI9870a38_98);
nor \U$202 ( \545 , RI9870d80_105, RI9870df8_106);
nor \U$203 ( \546 , \544 , \545 );
or \U$204 ( \547 , RI9870c90_103, RI9870d08_104);
and \U$205 ( \548 , \540 , \543 , \546 , \547 );
not \U$206 ( \549 , RI9871398_118);
not \U$207 ( \550 , RI9871320_117);
nand \U$208 ( \551 , \549 , \550 );
not \U$209 ( \552 , RI9871230_115);
not \U$210 ( \553 , RI98712a8_116);
nand \U$211 ( \554 , \552 , \553 );
not \U$212 ( \555 , RI9871140_113);
not \U$213 ( \556 , RI98711b8_114);
nand \U$214 ( \557 , \555 , \556 );
not \U$215 ( \558 , RI9871410_119);
not \U$216 ( \559 , RI9871488_120);
nand \U$217 ( \560 , \558 , \559 );
nand \U$218 ( \561 , \551 , \554 , \557 , \560 );
nor \U$219 ( \562 , RI98716e0_125, RI9871758_126);
nor \U$220 ( \563 , RI98717d0_127, RI9871848_128);
nor \U$221 ( \564 , \562 , \563 );
nor \U$222 ( \565 , RI98715f0_123, RI9871668_124);
nor \U$223 ( \566 , RI9871500_121, RI9871578_122);
nor \U$224 ( \567 , \565 , \566 );
nand \U$225 ( \568 , \564 , \567 );
nor \U$226 ( \569 , \561 , \568 );
and \U$227 ( \570 , \548 , \569 );
nand \U$228 ( \571 , \536 , \570 );
not \U$229 ( \572 , \548 );
nor \U$230 ( \573 , RI98707e0_93, RI9870858_94);
nor \U$231 ( \574 , \573 , \529 );
not \U$232 ( \575 , \574 );
nand \U$233 ( \576 , RI98706f0_91, RI9870768_92);
or \U$234 ( \577 , \527 , \576 );
nand \U$235 ( \578 , RI9870600_89, RI9870678_90);
nand \U$236 ( \579 , \577 , \578 );
not \U$237 ( \580 , \579 );
or \U$238 ( \581 , \575 , \580 );
nand \U$239 ( \582 , RI98708d0_95, RI9870948_96);
not \U$240 ( \583 , \582 );
and \U$241 ( \584 , \526 , \583 );
and \U$242 ( \585 , RI98707e0_93, RI9870858_94);
nor \U$243 ( \586 , \584 , \585 );
nand \U$244 ( \587 , \581 , \586 );
not \U$245 ( \588 , \587 );
nor \U$246 ( \589 , \522 , \470 );
not \U$247 ( \590 , \589 );
or \U$248 ( \591 , \588 , \590 );
nor \U$249 ( \592 , RI9870150_79, RI98701c8_80);
nor \U$250 ( \593 , RI9870060_77, RI98700d8_78);
nor \U$251 ( \594 , \592 , \593 );
not \U$252 ( \595 , \594 );
nand \U$253 ( \596 , RI986ff70_75, RI986ffe8_76);
not \U$254 ( \597 , \596 );
not \U$255 ( \598 , \597 );
not \U$256 ( \599 , RI986fef8_74);
nand \U$257 ( \600 , \464 , \599 );
not \U$258 ( \601 , \600 );
or \U$259 ( \602 , \598 , \601 );
nand \U$260 ( \603 , RI986fe80_73, RI986fef8_74);
nand \U$261 ( \604 , \602 , \603 );
not \U$262 ( \605 , \604 );
or \U$263 ( \606 , \595 , \605 );
nand \U$264 ( \607 , RI9870060_77, RI98700d8_78);
or \U$265 ( \608 , \592 , \607 );
nand \U$266 ( \609 , RI9870150_79, RI98701c8_80);
nand \U$267 ( \610 , \608 , \609 );
not \U$268 ( \611 , \610 );
nand \U$269 ( \612 , \606 , \611 );
not \U$270 ( \613 , \612 );
nand \U$271 ( \614 , \591 , \613 );
not \U$272 ( \615 , \614 );
or \U$273 ( \616 , \572 , \615 );
nand \U$274 ( \617 , RI98709c0_97, RI9870a38_98);
not \U$275 ( \618 , \617 );
nand \U$276 ( \619 , RI9870f60_109, RI9870fd8_110);
or \U$277 ( \620 , \542 , \619 );
nand \U$278 ( \621 , RI9870ab0_99, RI9870b28_100);
nand \U$279 ( \622 , \620 , \621 );
nand \U$280 ( \623 , RI9870d80_105, RI9870df8_106);
not \U$281 ( \624 , \623 );
or \U$282 ( \625 , \622 , \624 );
nand \U$283 ( \626 , \625 , \546 );
not \U$284 ( \627 , \626 );
or \U$285 ( \628 , \618 , \627 );
nor \U$286 ( \629 , RI9870ba0_101, RI9870c18_102);
nor \U$287 ( \630 , \538 , \537 , \629 );
not \U$288 ( \631 , \630 );
not \U$289 ( \632 , \547 );
nor \U$290 ( \633 , \631 , \632 );
nand \U$291 ( \634 , \628 , \633 );
nand \U$292 ( \635 , \616 , \634 );
buf \U$293 ( \636 , \569 );
nand \U$294 ( \637 , \635 , \636 );
not \U$295 ( \638 , \561 );
nor \U$296 ( \639 , \568 , \632 );
or \U$297 ( \640 , RI9871050_111, RI98710c8_112);
not \U$298 ( \641 , \640 );
nand \U$299 ( \642 , RI9870e70_107, RI9870ee8_108);
or \U$300 ( \643 , \539 , \642 );
nand \U$301 ( \644 , RI9870ba0_101, RI9870c18_102);
nand \U$302 ( \645 , \643 , \644 );
not \U$303 ( \646 , \645 );
or \U$304 ( \647 , \641 , \646 );
nand \U$305 ( \648 , RI9871050_111, RI98710c8_112);
nand \U$306 ( \649 , \647 , \648 );
nand \U$307 ( \650 , \638 , \639 , \649 );
nand \U$308 ( \651 , RI9870c90_103, RI9870d08_104);
nor \U$309 ( \652 , \568 , \651 );
nand \U$310 ( \653 , \638 , \652 );
not \U$311 ( \654 , \566 );
not \U$312 ( \655 , \654 );
nor \U$313 ( \656 , RI98717d0_127, RI9871848_128);
nand \U$314 ( \657 , RI98716e0_125, RI9871758_126);
or \U$315 ( \658 , \656 , \657 );
nand \U$316 ( \659 , RI98717d0_127, RI9871848_128);
nand \U$317 ( \660 , \658 , \659 );
not \U$318 ( \661 , \660 );
or \U$319 ( \662 , \655 , \661 );
nand \U$320 ( \663 , RI9871500_121, RI9871578_122);
nand \U$321 ( \664 , \662 , \663 );
not \U$322 ( \665 , \565 );
nand \U$323 ( \666 , \664 , \665 );
and \U$324 ( \667 , \650 , \653 , \666 );
not \U$325 ( \668 , \568 );
not \U$326 ( \669 , \551 );
nor \U$327 ( \670 , RI9871140_113, RI98711b8_114);
nand \U$328 ( \671 , RI9871230_115, RI98712a8_116);
or \U$329 ( \672 , \670 , \671 );
nand \U$330 ( \673 , RI9871140_113, RI98711b8_114);
nand \U$331 ( \674 , \672 , \673 );
not \U$332 ( \675 , \674 );
or \U$333 ( \676 , \669 , \675 );
nand \U$334 ( \677 , RI9871320_117, RI9871398_118);
nand \U$335 ( \678 , \676 , \677 );
nand \U$336 ( \679 , \668 , \678 , \560 );
not \U$337 ( \680 , \679 );
not \U$338 ( \681 , \668 );
nand \U$339 ( \682 , RI9871410_119, RI9871488_120);
or \U$340 ( \683 , \681 , \682 );
nand \U$341 ( \684 , RI98715f0_123, RI9871668_124);
nand \U$342 ( \685 , \683 , \684 );
nor \U$343 ( \686 , \680 , \685 );
nand \U$344 ( \687 , \571 , \637 , \667 , \686 );
nor \U$345 ( \688 , RI986ead0_31, RI986eb48_32);
nor \U$346 ( \689 , \688 , \394 );
and \U$347 ( \690 , \689 , \406 );
nand \U$348 ( \691 , \415 , \690 );
nand \U$349 ( \692 , \389 , \454 );
nor \U$350 ( \693 , \691 , \692 );
nand \U$351 ( \694 , \687 , \693 );
not \U$352 ( \695 , \694 );
or \U$353 ( \696 , \457 , \695 );
nor \U$354 ( \697 , RI986df90_7, RI986e008_8);
nor \U$355 ( \698 , \697 , \357 );
and \U$356 ( \699 , \698 , \352 , \362 );
and \U$357 ( \700 , \699 , \350 );
nor \U$358 ( \701 , RI986f700_57, RI986f778_58);
not \U$359 ( \702 , \701 );
or \U$360 ( \703 , RI986f868_60, RI986f7f0_59);
or \U$361 ( \704 , RI986f9d0_63, RI986fa48_64);
and \U$362 ( \705 , \702 , \703 , \704 );
nor \U$363 ( \706 , RI986f340_49, RI986f3b8_50);
nor \U$364 ( \707 , RI986f430_51, RI986f4a8_52);
nor \U$365 ( \708 , \706 , \707 );
or \U$366 ( \709 , RI986f598_54, RI986f520_53);
or \U$367 ( \710 , RI986f688_56, RI986f610_55);
and \U$368 ( \711 , \708 , \709 , \710 );
or \U$369 ( \712 , RI986f8e0_61, RI986f958_62);
nand \U$370 ( \713 , \705 , \711 , \712 );
not \U$371 ( \714 , \713 );
and \U$372 ( \715 , \700 , \714 , \348 , \346 );
nand \U$373 ( \716 , \696 , \715 );
or \U$374 ( \717 , RI986e620_21, RI986e698_22);
not \U$375 ( \718 , \717 );
or \U$376 ( \719 , RI986e788_24, RI986e710_23);
not \U$377 ( \720 , \719 );
nor \U$378 ( \721 , RI986e440_17, RI986e4b8_18);
nand \U$379 ( \722 , RI986e530_19, RI986e5a8_20);
or \U$380 ( \723 , \721 , \722 );
nand \U$381 ( \724 , RI986e440_17, RI986e4b8_18);
nand \U$382 ( \725 , \723 , \724 );
not \U$383 ( \726 , \725 );
or \U$384 ( \727 , \720 , \726 );
nand \U$385 ( \728 , RI986e710_23, RI986e788_24);
nand \U$386 ( \729 , \727 , \728 );
not \U$387 ( \730 , \729 );
or \U$388 ( \731 , \718 , \730 );
nand \U$389 ( \732 , RI986e620_21, RI986e698_22);
nand \U$390 ( \733 , \731 , \732 );
not \U$391 ( \734 , \733 );
nor \U$392 ( \735 , \734 , \713 );
not \U$393 ( \736 , \711 );
not \U$394 ( \737 , \712 );
not \U$395 ( \738 , \704 );
not \U$396 ( \739 , RI986f700_57);
not \U$397 ( \740 , RI986f778_58);
or \U$398 ( \741 , \739 , \740 );
nand \U$399 ( \742 , RI986f7f0_59, RI986f868_60);
or \U$400 ( \743 , \701 , \742 );
nand \U$401 ( \744 , \741 , \743 );
not \U$402 ( \745 , \744 );
or \U$403 ( \746 , \738 , \745 );
nand \U$404 ( \747 , RI986f9d0_63, RI986fa48_64);
nand \U$405 ( \748 , \746 , \747 );
not \U$406 ( \749 , \748 );
or \U$407 ( \750 , \737 , \749 );
nand \U$408 ( \751 , RI986f8e0_61, RI986f958_62);
nand \U$409 ( \752 , \750 , \751 );
not \U$410 ( \753 , \752 );
or \U$411 ( \754 , \736 , \753 );
not \U$412 ( \755 , \710 );
not \U$413 ( \756 , \709 );
nand \U$414 ( \757 , RI986f430_51, RI986f4a8_52);
or \U$415 ( \758 , \706 , \757 );
nand \U$416 ( \759 , RI986f340_49, RI986f3b8_50);
nand \U$417 ( \760 , \758 , \759 );
not \U$418 ( \761 , \760 );
or \U$419 ( \762 , \756 , \761 );
nand \U$420 ( \763 , RI986f520_53, RI986f598_54);
nand \U$421 ( \764 , \762 , \763 );
not \U$422 ( \765 , \764 );
or \U$423 ( \766 , \755 , \765 );
nand \U$424 ( \767 , RI986f610_55, RI986f688_56);
nand \U$425 ( \768 , \766 , \767 );
not \U$426 ( \769 , \768 );
nand \U$427 ( \770 , \754 , \769 );
or \U$428 ( \771 , \735 , \770 );
and \U$429 ( \772 , \699 , \350 , \348 , \346 );
nand \U$430 ( \773 , \771 , \772 );
nand \U$431 ( \774 , \383 , \716 , \773 );
not \U$432 ( \775 , \774 );
or \U$433 ( \776 , \345 , \775 );
nand \U$434 ( \777 , RI986e350_15, RI986e3c8_16);
nand \U$435 ( \778 , \776 , \777 );
not \U$436 ( \779 , \778 );
not \U$437 ( \780 , \779 );
xor \U$438 ( \781 , \780 , RI98719b0_131);
and \U$439 ( \782 , RI9871aa0_133, RI9871a28_132);
not \U$440 ( \783 , RI9871aa0_133);
not \U$441 ( \784 , RI9871a28_132);
and \U$442 ( \785 , \783 , \784 );
or \U$443 ( \786 , \782 , \785 );
and \U$444 ( \787 , RI98719b0_131, RI9871a28_132);
not \U$445 ( \788 , RI98719b0_131);
and \U$446 ( \789 , \788 , \784 );
nor \U$447 ( \790 , \787 , \789 );
and \U$448 ( \791 , \786 , \790 );
not \U$449 ( \792 , \791 );
not \U$450 ( \793 , \792 );
buf \U$451 ( \794 , \793 );
and \U$452 ( \795 , \781 , \794 );
not \U$453 ( \796 , \786 );
buf \U$454 ( \797 , \796 );
and \U$455 ( \798 , \797 , RI98719b0_131);
nor \U$456 ( \799 , \795 , \798 );
not \U$457 ( \800 , \708 );
and \U$458 ( \801 , \705 , \712 );
not \U$459 ( \802 , \801 );
not \U$460 ( \803 , \456 );
nor \U$461 ( \804 , \803 , \733 );
nand \U$462 ( \805 , \694 , \804 );
not \U$463 ( \806 , \805 );
or \U$464 ( \807 , \802 , \806 );
not \U$465 ( \808 , \752 );
nand \U$466 ( \809 , \807 , \808 );
not \U$467 ( \810 , \809 );
or \U$468 ( \811 , \800 , \810 );
not \U$469 ( \812 , \760 );
nand \U$470 ( \813 , \811 , \812 );
nand \U$471 ( \814 , \709 , \763 );
and \U$472 ( \815 , \813 , \814 );
not \U$473 ( \816 , \813 );
not \U$474 ( \817 , \814 );
and \U$475 ( \818 , \816 , \817 );
nor \U$476 ( \819 , \815 , \818 );
buf \U$477 ( \820 , \819 );
not \U$478 ( \821 , \820 );
and \U$479 ( \822 , RI9871d70_139, \821 );
not \U$480 ( \823 , RI9871d70_139);
not \U$481 ( \824 , \821 );
and \U$482 ( \825 , \823 , \824 );
nor \U$483 ( \826 , \822 , \825 );
and \U$484 ( \827 , RI9872130_147, RI9872220_149);
not \U$485 ( \828 , RI9872130_147);
not \U$486 ( \829 , RI9872220_149);
and \U$487 ( \830 , \828 , \829 );
nor \U$488 ( \831 , \827 , \830 );
buf \U$489 ( \832 , \831 );
and \U$490 ( \833 , \826 , \832 );
not \U$491 ( \834 , \707 );
not \U$492 ( \835 , \834 );
not \U$493 ( \836 , \809 );
or \U$494 ( \837 , \835 , \836 );
nand \U$495 ( \838 , \837 , \757 );
not \U$496 ( \839 , \759 );
nor \U$497 ( \840 , \839 , \706 );
and \U$498 ( \841 , \838 , \840 );
not \U$499 ( \842 , \838 );
not \U$500 ( \843 , \840 );
and \U$501 ( \844 , \842 , \843 );
nor \U$502 ( \845 , \841 , \844 );
buf \U$503 ( \846 , \845 );
buf \U$504 ( \847 , \846 );
not \U$505 ( \848 , \847 );
and \U$506 ( \849 , RI9871d70_139, \848 );
not \U$507 ( \850 , RI9871d70_139);
and \U$508 ( \851 , \850 , \847 );
nor \U$509 ( \852 , \849 , \851 );
not \U$510 ( \853 , \831 );
and \U$511 ( \854 , RI9871d70_139, RI9872220_149);
not \U$512 ( \855 , RI9871d70_139);
and \U$513 ( \856 , \855 , \829 );
nor \U$514 ( \857 , \854 , \856 );
and \U$515 ( \858 , \853 , \857 );
buf \U$516 ( \859 , \858 );
not \U$517 ( \860 , \859 );
nor \U$518 ( \861 , \852 , \860 );
nor \U$519 ( \862 , \833 , \861 );
xor \U$520 ( \863 , \799 , \862 );
and \U$521 ( \864 , RI9871c80_137, RI98721a8_148);
not \U$522 ( \865 , RI9871c80_137);
not \U$523 ( \866 , RI98721a8_148);
and \U$524 ( \867 , \865 , \866 );
nor \U$525 ( \868 , \864 , \867 );
not \U$526 ( \869 , \868 );
and \U$527 ( \870 , RI9872130_147, RI98721a8_148);
not \U$528 ( \871 , RI9872130_147);
and \U$529 ( \872 , \871 , \866 );
nor \U$530 ( \873 , \870 , \872 );
nand \U$531 ( \874 , \869 , \873 );
not \U$532 ( \875 , \874 );
buf \U$533 ( \876 , \875 );
not \U$534 ( \877 , \876 );
nand \U$535 ( \878 , \710 , \767 );
not \U$536 ( \879 , \878 );
not \U$537 ( \880 , \879 );
not \U$538 ( \881 , \709 );
and \U$539 ( \882 , \809 , \708 );
not \U$540 ( \883 , \882 );
or \U$541 ( \884 , \881 , \883 );
not \U$542 ( \885 , \764 );
nand \U$543 ( \886 , \884 , \885 );
not \U$544 ( \887 , \886 );
not \U$545 ( \888 , \887 );
or \U$546 ( \889 , \880 , \888 );
nand \U$547 ( \890 , \886 , \878 );
nand \U$548 ( \891 , \889 , \890 );
not \U$549 ( \892 , \891 );
buf \U$550 ( \893 , \892 );
buf \U$551 ( \894 , \893 );
not \U$552 ( \895 , \894 );
and \U$553 ( \896 , RI9872130_147, \895 );
not \U$554 ( \897 , RI9872130_147);
and \U$555 ( \898 , \897 , \894 );
nor \U$556 ( \899 , \896 , \898 );
not \U$557 ( \900 , \899 );
or \U$558 ( \901 , \877 , \900 );
not \U$559 ( \902 , \697 );
and \U$560 ( \903 , \902 , \358 );
not \U$561 ( \904 , \714 );
nand \U$562 ( \905 , \694 , \456 );
not \U$563 ( \906 , \905 );
or \U$564 ( \907 , \904 , \906 );
nor \U$565 ( \908 , \735 , \770 );
nand \U$566 ( \909 , \907 , \908 );
and \U$567 ( \910 , \903 , \909 );
not \U$568 ( \911 , \903 );
not \U$569 ( \912 , \909 );
and \U$570 ( \913 , \911 , \912 );
or \U$571 ( \914 , \910 , \913 );
buf \U$572 ( \915 , \914 );
buf \U$573 ( \916 , \915 );
not \U$574 ( \917 , \916 );
not \U$575 ( \918 , \917 );
not \U$576 ( \919 , RI9872130_147);
and \U$577 ( \920 , \918 , \919 );
not \U$578 ( \921 , \918 );
and \U$579 ( \922 , \921 , RI9872130_147);
nor \U$580 ( \923 , \920 , \922 );
buf \U$581 ( \924 , \868 );
nand \U$582 ( \925 , \923 , \924 );
nand \U$583 ( \926 , \901 , \925 );
not \U$584 ( \927 , \926 );
xor \U$585 ( \928 , \863 , \927 );
not \U$586 ( \929 , \928 );
not \U$587 ( \930 , \929 );
not \U$588 ( \931 , \799 );
not \U$589 ( \932 , \832 );
or \U$590 ( \933 , \852 , \932 );
not \U$591 ( \934 , RI9871d70_139);
buf \U$592 ( \935 , \809 );
not \U$593 ( \936 , \935 );
nand \U$594 ( \937 , \834 , \757 );
not \U$595 ( \938 , \937 );
and \U$596 ( \939 , \936 , \938 );
and \U$597 ( \940 , \935 , \937 );
nor \U$598 ( \941 , \939 , \940 );
not \U$599 ( \942 , \941 );
buf \U$600 ( \943 , \942 );
buf \U$601 ( \944 , \943 );
not \U$602 ( \945 , \944 );
not \U$603 ( \946 , \945 );
not \U$604 ( \947 , \946 );
or \U$605 ( \948 , \934 , \947 );
or \U$606 ( \949 , \946 , RI9871d70_139);
nand \U$607 ( \950 , \948 , \949 );
or \U$608 ( \951 , \950 , \860 );
nand \U$609 ( \952 , \933 , \951 );
not \U$610 ( \953 , \952 );
or \U$611 ( \954 , \931 , \953 );
not \U$612 ( \955 , RI986fb38_66);
not \U$613 ( \956 , RI9870420_85);
not \U$614 ( \957 , RI9870510_87);
nand \U$615 ( \958 , \956 , \957 , RI98708d0_95, RI9870600_89);
nand \U$616 ( \959 , \507 , \532 , RI9870330_83, RI98707e0_93);
nor \U$617 ( \960 , \958 , \959 );
nor \U$618 ( \961 , RI986fe80_73, RI986ff70_75);
nor \U$619 ( \962 , RI9870060_77, RI9870150_79);
nand \U$620 ( \963 , \961 , \962 );
nand \U$621 ( \964 , \473 , RI986fac0_65, RI986fbb0_67, RI986fd90_71);
nor \U$622 ( \965 , \963 , \964 );
and \U$623 ( \966 , \960 , \965 );
nor \U$624 ( \967 , RI9871410_119, RI9871500_121);
nor \U$625 ( \968 , RI98715f0_123, RI98716e0_125);
nor \U$626 ( \969 , RI9871230_115, RI9871320_117);
nor \U$627 ( \970 , RI9871140_113, RI98717d0_127);
nand \U$628 ( \971 , \967 , \968 , \969 , \970 );
nor \U$629 ( \972 , RI98709c0_97, RI9870ab0_99);
nor \U$630 ( \973 , RI9870ba0_101, RI9870c90_103);
nor \U$631 ( \974 , RI9870d80_105, RI9870e70_107);
nor \U$632 ( \975 , RI9870f60_109, RI9871050_111);
nand \U$633 ( \976 , \972 , \973 , \974 , \975 );
nor \U$634 ( \977 , \971 , \976 );
nor \U$635 ( \978 , RI986e800_25, RI986e8f0_27);
nor \U$636 ( \979 , RI986e9e0_29, RI986ead0_31);
nor \U$637 ( \980 , RI986ebc0_33, RI986ecb0_35);
nor \U$638 ( \981 , RI986eda0_37, RI986ee90_39);
nand \U$639 ( \982 , \978 , \979 , \980 , \981 );
nor \U$640 ( \983 , RI986dcc0_1, RI986ddb0_3);
nor \U$641 ( \984 , RI986dea0_5, RI986e080_9);
nor \U$642 ( \985 , RI986df90_7, RI986e170_11);
nor \U$643 ( \986 , RI986e260_13, RI986e350_15);
nand \U$644 ( \987 , \983 , \984 , \985 , \986 );
nor \U$645 ( \988 , \982 , \987 );
nor \U$646 ( \989 , RI986f340_49, RI986f520_53);
nor \U$647 ( \990 , RI986f610_55, RI986f700_57);
nor \U$648 ( \991 , RI986f430_51, RI986f7f0_59);
nor \U$649 ( \992 , RI986f8e0_61, RI986f9d0_63);
nand \U$650 ( \993 , \989 , \990 , \991 , \992 );
nor \U$651 ( \994 , RI986e440_17, RI986e710_23);
nor \U$652 ( \995 , RI986e530_19, RI986ef80_41);
nor \U$653 ( \996 , RI986e620_21, RI986f070_43);
nor \U$654 ( \997 , RI986f160_45, RI986f250_47);
nand \U$655 ( \998 , \994 , \995 , \996 , \997 );
nor \U$656 ( \999 , \993 , \998 );
nand \U$657 ( \1000 , \966 , \977 , \988 , \999 );
not \U$658 ( \1001 , \1000 );
not \U$659 ( \1002 , \1001 );
or \U$660 ( \1003 , \955 , \1002 );
nand \U$661 ( \1004 , \1000 , RI9871ed8_142);
nand \U$662 ( \1005 , \1003 , \1004 );
nor \U$663 ( \1006 , \1005 , RI9871f50_143);
not \U$664 ( \1007 , \1006 );
nand \U$665 ( \1008 , \1005 , RI9871f50_143);
not \U$666 ( \1009 , RI9871f50_143);
and \U$667 ( \1010 , RI9871e60_141, \1009 );
not \U$668 ( \1011 , RI9871e60_141);
and \U$669 ( \1012 , \1011 , RI9871f50_143);
or \U$670 ( \1013 , \1010 , \1012 );
not \U$671 ( \1014 , \1013 );
nand \U$672 ( \1015 , \1007 , \1008 , \1014 );
not \U$673 ( \1016 , \1015 );
buf \U$674 ( \1017 , \1016 );
buf \U$675 ( \1018 , \1017 );
not \U$676 ( \1019 , \1018 );
buf \U$677 ( \1020 , \687 );
not \U$678 ( \1021 , \691 );
and \U$679 ( \1022 , \1020 , \1021 , \389 );
buf \U$680 ( \1023 , \447 );
or \U$681 ( \1024 , \1022 , \1023 );
not \U$682 ( \1025 , \453 );
nand \U$683 ( \1026 , \1024 , \1025 );
not \U$684 ( \1027 , \719 );
or \U$685 ( \1028 , \1026 , \1027 );
not \U$686 ( \1029 , \729 );
nand \U$687 ( \1030 , \1028 , \1029 );
not \U$688 ( \1031 , \1030 );
and \U$689 ( \1032 , \717 , \732 );
not \U$690 ( \1033 , \1032 );
and \U$691 ( \1034 , \1031 , \1033 );
not \U$692 ( \1035 , \1031 );
and \U$693 ( \1036 , \1035 , \1032 );
nor \U$694 ( \1037 , \1034 , \1036 );
buf \U$695 ( \1038 , \1037 );
buf \U$696 ( \1039 , \1038 );
not \U$697 ( \1040 , \1039 );
buf \U$698 ( \1041 , \1040 );
buf \U$699 ( \1042 , \1005 );
not \U$700 ( \1043 , \1042 );
not \U$701 ( \1044 , \1043 );
not \U$702 ( \1045 , \1044 );
and \U$703 ( \1046 , \1041 , \1045 );
buf \U$704 ( \1047 , \1039 );
and \U$705 ( \1048 , \1047 , \1044 );
nor \U$706 ( \1049 , \1046 , \1048 );
not \U$707 ( \1050 , \1049 );
or \U$708 ( \1051 , \1019 , \1050 );
nand \U$709 ( \1052 , \703 , \742 );
not \U$710 ( \1053 , \1052 );
not \U$711 ( \1054 , \1053 );
buf \U$712 ( \1055 , \805 );
not \U$713 ( \1056 , \1055 );
not \U$714 ( \1057 , \1056 );
or \U$715 ( \1058 , \1054 , \1057 );
nand \U$716 ( \1059 , \1055 , \1052 );
nand \U$717 ( \1060 , \1058 , \1059 );
buf \U$718 ( \1061 , \1060 );
buf \U$719 ( \1062 , \1061 );
and \U$720 ( \1063 , \1062 , \1045 );
not \U$721 ( \1064 , \1062 );
and \U$722 ( \1065 , \1064 , \1044 );
nor \U$723 ( \1066 , \1063 , \1065 );
buf \U$724 ( \1067 , \1013 );
not \U$725 ( \1068 , \1067 );
or \U$726 ( \1069 , \1066 , \1068 );
nand \U$727 ( \1070 , \1051 , \1069 );
not \U$728 ( \1071 , \1070 );
and \U$729 ( \1072 , RI98718c0_129, RI9871938_130);
not \U$730 ( \1073 , RI98718c0_129);
not \U$731 ( \1074 , RI9871938_130);
and \U$732 ( \1075 , \1073 , \1074 );
nor \U$733 ( \1076 , \1072 , \1075 );
not \U$734 ( \1077 , \1076 );
not \U$735 ( \1078 , RI98719b0_131);
nand \U$736 ( \1079 , \1074 , \1078 );
nand \U$737 ( \1080 , RI9871938_130, RI98719b0_131);
and \U$738 ( \1081 , \1079 , \1080 );
nor \U$739 ( \1082 , \1077 , \1081 );
buf \U$740 ( \1083 , \1082 );
not \U$741 ( \1084 , \1083 );
not \U$742 ( \1085 , \700 );
not \U$743 ( \1086 , \909 );
or \U$744 ( \1087 , \1085 , \1086 );
not \U$745 ( \1088 , \374 );
nand \U$746 ( \1089 , \1087 , \1088 );
not \U$747 ( \1090 , \1089 );
nand \U$748 ( \1091 , \348 , \377 );
not \U$749 ( \1092 , \1091 );
and \U$750 ( \1093 , \1090 , \1092 );
not \U$751 ( \1094 , \1090 );
and \U$752 ( \1095 , \1094 , \1091 );
nor \U$753 ( \1096 , \1093 , \1095 );
buf \U$754 ( \1097 , \1096 );
buf \U$755 ( \1098 , \1097 );
and \U$756 ( \1099 , RI98718c0_129, \1098 );
not \U$757 ( \1100 , RI98718c0_129);
not \U$758 ( \1101 , \1092 );
not \U$759 ( \1102 , \1090 );
or \U$760 ( \1103 , \1101 , \1102 );
nand \U$761 ( \1104 , \1089 , \1091 );
nand \U$762 ( \1105 , \1103 , \1104 );
buf \U$763 ( \1106 , \1105 );
and \U$764 ( \1107 , \1100 , \1106 );
or \U$765 ( \1108 , \1099 , \1107 );
not \U$766 ( \1109 , \1108 );
or \U$767 ( \1110 , \1084 , \1109 );
not \U$768 ( \1111 , RI98718c0_129);
nand \U$769 ( \1112 , \346 , \381 );
not \U$770 ( \1113 , \1112 );
not \U$771 ( \1114 , \1113 );
and \U$772 ( \1115 , \700 , \348 );
not \U$773 ( \1116 , \1115 );
not \U$774 ( \1117 , \909 );
or \U$775 ( \1118 , \1116 , \1117 );
not \U$776 ( \1119 , \378 );
nand \U$777 ( \1120 , \1118 , \1119 );
not \U$778 ( \1121 , \1120 );
not \U$779 ( \1122 , \1121 );
or \U$780 ( \1123 , \1114 , \1122 );
nand \U$781 ( \1124 , \1120 , \1112 );
nand \U$782 ( \1125 , \1123 , \1124 );
buf \U$783 ( \1126 , \1125 );
not \U$784 ( \1127 , \1126 );
buf \U$785 ( \1128 , \1127 );
not \U$786 ( \1129 , \1128 );
and \U$787 ( \1130 , \1111 , \1129 );
not \U$788 ( \1131 , \1111 );
and \U$789 ( \1132 , \1131 , \1128 );
nor \U$790 ( \1133 , \1130 , \1132 );
buf \U$791 ( \1134 , \1081 );
buf \U$792 ( \1135 , \1134 );
buf \U$793 ( \1136 , \1135 );
not \U$794 ( \1137 , \1136 );
or \U$795 ( \1138 , \1133 , \1137 );
nand \U$796 ( \1139 , \1110 , \1138 );
not \U$797 ( \1140 , RI9872040_145);
not \U$798 ( \1141 , \1000 );
or \U$799 ( \1142 , \1140 , \1141 );
nand \U$800 ( \1143 , \1141 , RI9871ed8_142);
nand \U$801 ( \1144 , \1142 , \1143 );
not \U$802 ( \1145 , \1144 );
not \U$803 ( \1146 , \1005 );
nand \U$804 ( \1147 , \1145 , \1146 );
not \U$805 ( \1148 , RI9872040_145);
not \U$806 ( \1149 , \1141 );
or \U$807 ( \1150 , \1148 , \1149 );
not \U$808 ( \1151 , \1141 );
nand \U$809 ( \1152 , \1151 , RI9871fc8_144);
nand \U$810 ( \1153 , \1150 , \1152 );
not \U$811 ( \1154 , \1153 );
or \U$812 ( \1155 , \1147 , \1154 );
not \U$813 ( \1156 , \1153 );
not \U$814 ( \1157 , \1146 );
buf \U$815 ( \1158 , \1144 );
nand \U$816 ( \1159 , \1156 , \1157 , \1158 );
nand \U$817 ( \1160 , \1155 , \1159 );
buf \U$818 ( \1161 , \1160 );
buf \U$819 ( \1162 , \1161 );
not \U$820 ( \1163 , \1162 );
not \U$821 ( \1164 , \1153 );
not \U$822 ( \1165 , \1164 );
not \U$823 ( \1166 , \1165 );
not \U$824 ( \1167 , \724 );
nor \U$825 ( \1168 , \1167 , \721 );
not \U$826 ( \1169 , \1168 );
or \U$827 ( \1170 , RI986e530_19, RI986e5a8_20);
not \U$828 ( \1171 , \1170 );
not \U$829 ( \1172 , \389 );
not \U$830 ( \1173 , \1021 );
not \U$831 ( \1174 , \687 );
or \U$832 ( \1175 , \1173 , \1174 );
not \U$833 ( \1176 , \429 );
nand \U$834 ( \1177 , \1175 , \1176 );
not \U$835 ( \1178 , \1177 );
or \U$836 ( \1179 , \1172 , \1178 );
nand \U$837 ( \1180 , \1179 , \446 );
not \U$838 ( \1181 , \1180 );
or \U$839 ( \1182 , \1171 , \1181 );
nand \U$840 ( \1183 , \1182 , \722 );
not \U$841 ( \1184 , \1183 );
not \U$842 ( \1185 , \1184 );
or \U$843 ( \1186 , \1169 , \1185 );
not \U$844 ( \1187 , \1168 );
nand \U$845 ( \1188 , \1187 , \1183 );
nand \U$846 ( \1189 , \1186 , \1188 );
not \U$847 ( \1190 , \1189 );
buf \U$848 ( \1191 , \1190 );
and \U$849 ( \1192 , \1166 , \1191 );
not \U$850 ( \1193 , \1166 );
not \U$851 ( \1194 , \1191 );
and \U$852 ( \1195 , \1193 , \1194 );
nor \U$853 ( \1196 , \1192 , \1195 );
not \U$854 ( \1197 , \1196 );
or \U$855 ( \1198 , \1163 , \1197 );
not \U$856 ( \1199 , \1165 );
not \U$857 ( \1200 , \1199 );
not \U$858 ( \1201 , \725 );
nand \U$859 ( \1202 , \1201 , \1026 );
not \U$860 ( \1203 , \1202 );
nand \U$861 ( \1204 , \719 , \728 );
not \U$862 ( \1205 , \1204 );
and \U$863 ( \1206 , \1203 , \1205 );
and \U$864 ( \1207 , \1202 , \1204 );
nor \U$865 ( \1208 , \1206 , \1207 );
buf \U$866 ( \1209 , \1208 );
buf \U$867 ( \1210 , \1209 );
not \U$868 ( \1211 , \1210 );
buf \U$869 ( \1212 , \1211 );
xor \U$870 ( \1213 , \1200 , \1212 );
not \U$871 ( \1214 , \1144 );
not \U$872 ( \1215 , \1042 );
or \U$873 ( \1216 , \1214 , \1215 );
or \U$874 ( \1217 , \1042 , \1158 );
nand \U$875 ( \1218 , \1216 , \1217 );
buf \U$876 ( \1219 , \1218 );
not \U$877 ( \1220 , \1219 );
nand \U$878 ( \1221 , \1213 , \1220 );
nand \U$879 ( \1222 , \1198 , \1221 );
xor \U$880 ( \1223 , \1139 , \1222 );
not \U$881 ( \1224 , \1223 );
or \U$882 ( \1225 , \1071 , \1224 );
nand \U$883 ( \1226 , \1222 , \1139 );
nand \U$884 ( \1227 , \1225 , \1226 );
xor \U$885 ( \1228 , \952 , \799 );
nand \U$886 ( \1229 , \1227 , \1228 );
nand \U$887 ( \1230 , \954 , \1229 );
not \U$888 ( \1231 , \1230 );
or \U$889 ( \1232 , \930 , \1231 );
not \U$890 ( \1233 , \928 );
not \U$891 ( \1234 , \1230 );
and \U$892 ( \1235 , \1233 , \1234 );
and \U$893 ( \1236 , \928 , \1230 );
nor \U$894 ( \1237 , \1235 , \1236 );
not \U$895 ( \1238 , \1237 );
not \U$896 ( \1239 , \950 );
not \U$897 ( \1240 , \932 );
and \U$898 ( \1241 , \1239 , \1240 );
not \U$899 ( \1242 , \705 );
not \U$900 ( \1243 , \805 );
or \U$901 ( \1244 , \1242 , \1243 );
not \U$902 ( \1245 , \748 );
nand \U$903 ( \1246 , \1244 , \1245 );
nand \U$904 ( \1247 , \712 , \751 );
and \U$905 ( \1248 , \1246 , \1247 );
not \U$906 ( \1249 , \1246 );
not \U$907 ( \1250 , \1247 );
and \U$908 ( \1251 , \1249 , \1250 );
nor \U$909 ( \1252 , \1248 , \1251 );
buf \U$910 ( \1253 , \1252 );
not \U$911 ( \1254 , \1253 );
and \U$912 ( \1255 , RI9871d70_139, \1254 );
not \U$913 ( \1256 , RI9871d70_139);
not \U$914 ( \1257 , \1254 );
and \U$915 ( \1258 , \1256 , \1257 );
nor \U$916 ( \1259 , \1255 , \1258 );
and \U$917 ( \1260 , \1259 , \859 );
nor \U$918 ( \1261 , \1241 , \1260 );
xor \U$919 ( \1262 , RI986dea0_5, RI986df18_6);
not \U$920 ( \1263 , \1262 );
not \U$921 ( \1264 , \902 );
not \U$922 ( \1265 , \909 );
or \U$923 ( \1266 , \1264 , \1265 );
nand \U$924 ( \1267 , \1266 , \358 );
not \U$925 ( \1268 , \1267 );
not \U$926 ( \1269 , \1268 );
or \U$927 ( \1270 , \1263 , \1269 );
not \U$928 ( \1271 , \1262 );
nand \U$929 ( \1272 , \1267 , \1271 );
nand \U$930 ( \1273 , \1270 , \1272 );
buf \U$931 ( \1274 , \1273 );
buf \U$932 ( \1275 , \1274 );
not \U$933 ( \1276 , \1275 );
not \U$934 ( \1277 , RI9871b18_134);
and \U$935 ( \1278 , \1276 , \1277 );
and \U$936 ( \1279 , \1275 , RI9871b18_134);
nor \U$937 ( \1280 , \1278 , \1279 );
not \U$938 ( \1281 , \1280 );
not \U$939 ( \1282 , \1281 );
not \U$940 ( \1283 , RI9871b18_134);
not \U$941 ( \1284 , RI9871b90_135);
and \U$942 ( \1285 , \1283 , \1284 );
and \U$943 ( \1286 , RI9871b18_134, RI9871b90_135);
nand \U$944 ( \1287 , RI9871b90_135, RI9871c08_136);
not \U$945 ( \1288 , \1287 );
nor \U$946 ( \1289 , RI9871b90_135, RI9871c08_136);
nor \U$947 ( \1290 , \1288 , \1289 );
nor \U$948 ( \1291 , \1285 , \1286 , \1290 );
buf \U$949 ( \1292 , \1291 );
not \U$950 ( \1293 , \1292 );
not \U$951 ( \1294 , \1293 );
and \U$952 ( \1295 , \1282 , \1294 );
not \U$953 ( \1296 , \698 );
not \U$954 ( \1297 , \909 );
or \U$955 ( \1298 , \1296 , \1297 );
not \U$956 ( \1299 , \360 );
nand \U$957 ( \1300 , \1298 , \1299 );
nand \U$958 ( \1301 , \362 , \365 );
not \U$959 ( \1302 , \1301 );
and \U$960 ( \1303 , \1300 , \1302 );
not \U$961 ( \1304 , \1300 );
and \U$962 ( \1305 , \1304 , \1301 );
nor \U$963 ( \1306 , \1303 , \1305 );
not \U$964 ( \1307 , \1306 );
buf \U$965 ( \1308 , \1307 );
not \U$966 ( \1309 , \1308 );
not \U$967 ( \1310 , \1309 );
not \U$968 ( \1311 , \1310 );
and \U$969 ( \1312 , RI9871b18_134, \1311 );
not \U$970 ( \1313 , RI9871b18_134);
not \U$971 ( \1314 , \1300 );
not \U$972 ( \1315 , \1301 );
and \U$973 ( \1316 , \1314 , \1315 );
and \U$974 ( \1317 , \1300 , \1301 );
nor \U$975 ( \1318 , \1316 , \1317 );
buf \U$976 ( \1319 , \1318 );
buf \U$977 ( \1320 , \1319 );
and \U$978 ( \1321 , \1313 , \1320 );
nor \U$979 ( \1322 , \1312 , \1321 );
buf \U$980 ( \1323 , \1290 );
and \U$981 ( \1324 , \1322 , \1323 );
nor \U$982 ( \1325 , \1295 , \1324 );
xor \U$983 ( \1326 , \1261 , \1325 );
not \U$984 ( \1327 , \703 );
nor \U$985 ( \1328 , \1327 , \701 );
not \U$986 ( \1329 , \1328 );
not \U$987 ( \1330 , \805 );
or \U$988 ( \1331 , \1329 , \1330 );
not \U$989 ( \1332 , \744 );
nand \U$990 ( \1333 , \1331 , \1332 );
not \U$991 ( \1334 , \1333 );
nand \U$992 ( \1335 , \704 , \747 );
not \U$993 ( \1336 , \1335 );
and \U$994 ( \1337 , \1334 , \1336 );
and \U$995 ( \1338 , \1333 , \1335 );
nor \U$996 ( \1339 , \1337 , \1338 );
buf \U$997 ( \1340 , \1339 );
not \U$998 ( \1341 , \1340 );
and \U$999 ( \1342 , RI9871e60_141, \1341 );
not \U$1000 ( \1343 , RI9871e60_141);
buf \U$1001 ( \1344 , \1340 );
and \U$1002 ( \1345 , \1343 , \1344 );
nor \U$1003 ( \1346 , \1342 , \1345 );
not \U$1004 ( \1347 , RI9871d70_139);
not \U$1005 ( \1348 , RI9871de8_140);
nand \U$1006 ( \1349 , \1347 , \1348 );
nand \U$1007 ( \1350 , RI9871d70_139, RI9871de8_140);
and \U$1008 ( \1351 , \1349 , \1350 );
buf \U$1009 ( \1352 , \1351 );
buf \U$1010 ( \1353 , \1352 );
and \U$1011 ( \1354 , \1346 , \1353 );
not \U$1012 ( \1355 , \703 );
not \U$1013 ( \1356 , \805 );
or \U$1014 ( \1357 , \1355 , \1356 );
nand \U$1015 ( \1358 , \1357 , \742 );
xor \U$1016 ( \1359 , RI986f700_57, RI986f778_58);
and \U$1017 ( \1360 , \1358 , \1359 );
not \U$1018 ( \1361 , \1358 );
not \U$1019 ( \1362 , \1359 );
and \U$1020 ( \1363 , \1361 , \1362 );
nor \U$1021 ( \1364 , \1360 , \1363 );
buf \U$1022 ( \1365 , \1364 );
not \U$1023 ( \1366 , \1365 );
not \U$1024 ( \1367 , RI9871e60_141);
and \U$1025 ( \1368 , \1366 , \1367 );
not \U$1026 ( \1369 , \1365 );
not \U$1027 ( \1370 , \1369 );
buf \U$1028 ( \1371 , \1370 );
and \U$1029 ( \1372 , \1371 , RI9871e60_141);
nor \U$1030 ( \1373 , \1368 , \1372 );
not \U$1031 ( \1374 , \1351 );
and \U$1032 ( \1375 , RI9871e60_141, RI9871de8_140);
not \U$1033 ( \1376 , RI9871e60_141);
and \U$1034 ( \1377 , \1376 , \1348 );
nor \U$1035 ( \1378 , \1375 , \1377 );
and \U$1036 ( \1379 , \1374 , \1378 );
buf \U$1037 ( \1380 , \1379 );
buf \U$1038 ( \1381 , \1380 );
buf \U$1039 ( \1382 , \1381 );
and \U$1040 ( \1383 , \1373 , \1382 );
nor \U$1041 ( \1384 , \1354 , \1383 );
and \U$1042 ( \1385 , \1326 , \1384 );
and \U$1043 ( \1386 , \1261 , \1325 );
nor \U$1044 ( \1387 , \1385 , \1386 );
not \U$1045 ( \1388 , \1387 );
nand \U$1046 ( \1389 , RI9872298_150, RI9872310_151);
and \U$1047 ( \1390 , \1389 , RI9871aa0_133);
and \U$1048 ( \1391 , \344 , \777 );
xor \U$1049 ( \1392 , \1391 , \774 );
buf \U$1050 ( \1393 , \1392 );
buf \U$1051 ( \1394 , \1393 );
xor \U$1052 ( \1395 , \1394 , RI98719b0_131);
not \U$1053 ( \1396 , \1395 );
not \U$1054 ( \1397 , \1396 );
not \U$1055 ( \1398 , \794 );
not \U$1056 ( \1399 , \1398 );
and \U$1057 ( \1400 , \1397 , \1399 );
and \U$1058 ( \1401 , \781 , \797 );
nor \U$1059 ( \1402 , \1400 , \1401 );
xnor \U$1060 ( \1403 , \1390 , \1402 );
not \U$1061 ( \1404 , \699 );
not \U$1062 ( \1405 , \909 );
or \U$1063 ( \1406 , \1404 , \1405 );
not \U$1064 ( \1407 , \370 );
nand \U$1065 ( \1408 , \1406 , \1407 );
nand \U$1066 ( \1409 , \350 , \373 );
not \U$1067 ( \1410 , \1409 );
and \U$1068 ( \1411 , \1408 , \1410 );
not \U$1069 ( \1412 , \1408 );
and \U$1070 ( \1413 , \1412 , \1409 );
nor \U$1071 ( \1414 , \1411 , \1413 );
buf \U$1072 ( \1415 , \1414 );
not \U$1073 ( \1416 , \1415 );
not \U$1074 ( \1417 , \1416 );
not \U$1075 ( \1418 , \1417 );
and \U$1076 ( \1419 , RI9871c08_136, \1418 );
not \U$1077 ( \1420 , RI9871c08_136);
and \U$1078 ( \1421 , \1420 , \1417 );
nor \U$1079 ( \1422 , \1419 , \1421 );
and \U$1080 ( \1423 , RI98718c0_129, RI98720b8_146);
not \U$1081 ( \1424 , RI98718c0_129);
not \U$1082 ( \1425 , RI98720b8_146);
and \U$1083 ( \1426 , \1424 , \1425 );
nor \U$1084 ( \1427 , \1423 , \1426 );
buf \U$1085 ( \1428 , \1427 );
buf \U$1086 ( \1429 , \1428 );
buf \U$1087 ( \1430 , \1429 );
buf \U$1088 ( \1431 , \1430 );
not \U$1089 ( \1432 , \1431 );
or \U$1090 ( \1433 , \1422 , \1432 );
and \U$1091 ( \1434 , \698 , \362 );
not \U$1092 ( \1435 , \1434 );
not \U$1093 ( \1436 , \909 );
or \U$1094 ( \1437 , \1435 , \1436 );
not \U$1095 ( \1438 , \366 );
nand \U$1096 ( \1439 , \1437 , \1438 );
not \U$1097 ( \1440 , \1439 );
nand \U$1098 ( \1441 , \352 , \369 );
not \U$1099 ( \1442 , \1441 );
and \U$1100 ( \1443 , \1440 , \1442 );
and \U$1101 ( \1444 , \1439 , \1441 );
nor \U$1102 ( \1445 , \1443 , \1444 );
buf \U$1103 ( \1446 , \1445 );
buf \U$1104 ( \1447 , \1446 );
xor \U$1105 ( \1448 , \1447 , RI9871c08_136);
and \U$1106 ( \1449 , RI9871c08_136, RI98720b8_146);
not \U$1107 ( \1450 , RI9871c08_136);
and \U$1108 ( \1451 , \1450 , \1425 );
nor \U$1109 ( \1452 , \1449 , \1451 );
not \U$1110 ( \1453 , \1452 );
nor \U$1111 ( \1454 , \1453 , \1427 );
buf \U$1112 ( \1455 , \1454 );
buf \U$1113 ( \1456 , \1455 );
not \U$1114 ( \1457 , \1456 );
or \U$1115 ( \1458 , \1448 , \1457 );
nand \U$1116 ( \1459 , \1433 , \1458 );
not \U$1117 ( \1460 , \1459 );
or \U$1118 ( \1461 , \1403 , \1460 );
or \U$1119 ( \1462 , \1402 , \1390 );
nand \U$1120 ( \1463 , \1461 , \1462 );
not \U$1121 ( \1464 , \1463 );
and \U$1122 ( \1465 , RI9872130_147, \824 );
not \U$1123 ( \1466 , RI9872130_147);
and \U$1124 ( \1467 , \1466 , \821 );
nor \U$1125 ( \1468 , \1465 , \1467 );
not \U$1126 ( \1469 , \1468 );
not \U$1127 ( \1470 , \924 );
not \U$1128 ( \1471 , \1470 );
and \U$1129 ( \1472 , \1469 , \1471 );
xnor \U$1130 ( \1473 , \848 , RI9872130_147);
and \U$1131 ( \1474 , \1473 , \876 );
nor \U$1132 ( \1475 , \1472 , \1474 );
not \U$1133 ( \1476 , \1475 );
not \U$1134 ( \1477 , \1476 );
buf \U$1135 ( \1478 , \1180 );
not \U$1136 ( \1479 , \1478 );
nand \U$1137 ( \1480 , \1170 , \722 );
not \U$1138 ( \1481 , \1480 );
and \U$1139 ( \1482 , \1479 , \1481 );
and \U$1140 ( \1483 , \1478 , \1480 );
nor \U$1141 ( \1484 , \1482 , \1483 );
buf \U$1142 ( \1485 , \1484 );
not \U$1143 ( \1486 , \1485 );
not \U$1144 ( \1487 , \1486 );
nor \U$1145 ( \1488 , \1487 , \1166 );
and \U$1146 ( \1489 , RI9871b18_134, RI9871cf8_138);
not \U$1147 ( \1490 , RI9871b18_134);
not \U$1148 ( \1491 , RI9871cf8_138);
and \U$1149 ( \1492 , \1490 , \1491 );
nor \U$1150 ( \1493 , \1489 , \1492 );
not \U$1151 ( \1494 , \1493 );
and \U$1152 ( \1495 , RI9871c80_137, RI9871cf8_138);
not \U$1153 ( \1496 , RI9871c80_137);
and \U$1154 ( \1497 , \1496 , \1491 );
nor \U$1155 ( \1498 , \1495 , \1497 );
nand \U$1156 ( \1499 , \1494 , \1498 );
not \U$1157 ( \1500 , \1499 );
buf \U$1158 ( \1501 , \1500 );
not \U$1159 ( \1502 , \1501 );
and \U$1160 ( \1503 , RI9871c80_137, \895 );
not \U$1161 ( \1504 , RI9871c80_137);
not \U$1162 ( \1505 , \891 );
buf \U$1163 ( \1506 , \1505 );
and \U$1164 ( \1507 , \1504 , \1506 );
nor \U$1165 ( \1508 , \1503 , \1507 );
not \U$1166 ( \1509 , \1508 );
or \U$1167 ( \1510 , \1502 , \1509 );
and \U$1168 ( \1511 , RI9871c80_137, \918 );
not \U$1169 ( \1512 , RI9871c80_137);
not \U$1170 ( \1513 , \916 );
and \U$1171 ( \1514 , \1512 , \1513 );
nor \U$1172 ( \1515 , \1511 , \1514 );
not \U$1173 ( \1516 , \1515 );
not \U$1174 ( \1517 , \1494 );
buf \U$1175 ( \1518 , \1517 );
nand \U$1176 ( \1519 , \1516 , \1518 );
nand \U$1177 ( \1520 , \1510 , \1519 );
xor \U$1178 ( \1521 , \1488 , \1520 );
not \U$1179 ( \1522 , \1521 );
or \U$1180 ( \1523 , \1477 , \1522 );
nand \U$1181 ( \1524 , \1520 , \1488 );
nand \U$1182 ( \1525 , \1523 , \1524 );
not \U$1183 ( \1526 , \1525 );
not \U$1184 ( \1527 , \1526 );
or \U$1185 ( \1528 , \1464 , \1527 );
not \U$1186 ( \1529 , \1463 );
nand \U$1187 ( \1530 , \1529 , \1525 );
nand \U$1188 ( \1531 , \1528 , \1530 );
not \U$1189 ( \1532 , \1531 );
or \U$1190 ( \1533 , \1388 , \1532 );
nand \U$1191 ( \1534 , \1525 , \1463 );
nand \U$1192 ( \1535 , \1533 , \1534 );
nand \U$1193 ( \1536 , \1238 , \1535 );
nand \U$1194 ( \1537 , \1232 , \1536 );
and \U$1195 ( \1538 , RI9871b18_134, \1106 );
not \U$1196 ( \1539 , RI9871b18_134);
and \U$1197 ( \1540 , \1539 , \1097 );
or \U$1198 ( \1541 , \1538 , \1540 );
not \U$1199 ( \1542 , \1541 );
not \U$1200 ( \1543 , \1323 );
not \U$1201 ( \1544 , \1543 );
and \U$1202 ( \1545 , \1542 , \1544 );
xor \U$1203 ( \1546 , \1417 , RI9871b18_134);
and \U$1204 ( \1547 , \1546 , \1292 );
nor \U$1205 ( \1548 , \1545 , \1547 );
not \U$1206 ( \1549 , \943 );
not \U$1207 ( \1550 , \1549 );
not \U$1208 ( \1551 , \1550 );
not \U$1209 ( \1552 , RI9871e60_141);
and \U$1210 ( \1553 , \1551 , \1552 );
and \U$1211 ( \1554 , \1550 , RI9871e60_141);
nor \U$1212 ( \1555 , \1553 , \1554 );
not \U$1213 ( \1556 , \1555 );
not \U$1214 ( \1557 , \1556 );
not \U$1215 ( \1558 , \1382 );
not \U$1216 ( \1559 , \1558 );
and \U$1217 ( \1560 , \1557 , \1559 );
xor \U$1218 ( \1561 , RI9871e60_141, \847 );
and \U$1219 ( \1562 , \1561 , \1353 );
nor \U$1220 ( \1563 , \1560 , \1562 );
xnor \U$1221 ( \1564 , \1548 , \1563 );
xnor \U$1222 ( \1565 , \894 , RI9871d70_139);
and \U$1223 ( \1566 , \1565 , \832 );
and \U$1224 ( \1567 , \826 , \859 );
nor \U$1225 ( \1568 , \1566 , \1567 );
xor \U$1226 ( \1569 , \1564 , \1568 );
xor \U$1227 ( \1570 , \799 , \862 );
not \U$1228 ( \1571 , \926 );
and \U$1229 ( \1572 , \1570 , \1571 );
and \U$1230 ( \1573 , \799 , \862 );
or \U$1231 ( \1574 , \1572 , \1573 );
not \U$1232 ( \1575 , \1574 );
xor \U$1233 ( \1576 , \1569 , \1575 );
not \U$1234 ( \1577 , \1518 );
not \U$1235 ( \1578 , \1272 );
nor \U$1236 ( \1579 , \1267 , \1271 );
nor \U$1237 ( \1580 , \1578 , \1579 );
buf \U$1238 ( \1581 , \1580 );
not \U$1239 ( \1582 , \1581 );
not \U$1240 ( \1583 , \1582 );
not \U$1241 ( \1584 , RI9871c80_137);
and \U$1242 ( \1585 , \1583 , \1584 );
not \U$1243 ( \1586 , \1583 );
and \U$1244 ( \1587 , \1586 , RI9871c80_137);
nor \U$1245 ( \1588 , \1585 , \1587 );
not \U$1246 ( \1589 , \1588 );
or \U$1247 ( \1590 , \1577 , \1589 );
not \U$1248 ( \1591 , \1501 );
or \U$1249 ( \1592 , \1515 , \1591 );
nand \U$1250 ( \1593 , \1590 , \1592 );
not \U$1251 ( \1594 , \1220 );
not \U$1252 ( \1595 , \1041 );
xor \U$1253 ( \1596 , \1200 , \1595 );
not \U$1254 ( \1597 , \1596 );
or \U$1255 ( \1598 , \1594 , \1597 );
nand \U$1256 ( \1599 , \1213 , \1162 );
nand \U$1257 ( \1600 , \1598 , \1599 );
xor \U$1258 ( \1601 , \1593 , \1600 );
not \U$1259 ( \1602 , \1067 );
not \U$1260 ( \1603 , \1365 );
not \U$1261 ( \1604 , \1603 );
buf \U$1262 ( \1605 , \1604 );
not \U$1263 ( \1606 , \1605 );
and \U$1264 ( \1607 , \1606 , \1045 );
and \U$1265 ( \1608 , \1605 , \1044 );
nor \U$1266 ( \1609 , \1607 , \1608 );
not \U$1267 ( \1610 , \1609 );
or \U$1268 ( \1611 , \1602 , \1610 );
not \U$1269 ( \1612 , \1018 );
or \U$1270 ( \1613 , \1066 , \1612 );
nand \U$1271 ( \1614 , \1611 , \1613 );
and \U$1272 ( \1615 , \1601 , \1614 );
and \U$1273 ( \1616 , \1593 , \1600 );
nor \U$1274 ( \1617 , \1615 , \1616 );
and \U$1275 ( \1618 , \1098 , RI9871c08_136);
not \U$1276 ( \1619 , RI9871c08_136);
and \U$1277 ( \1620 , \1106 , \1619 );
nor \U$1278 ( \1621 , \1618 , \1620 );
or \U$1279 ( \1622 , \1621 , \1432 );
or \U$1280 ( \1623 , \1422 , \1457 );
nand \U$1281 ( \1624 , \1622 , \1623 );
not \U$1282 ( \1625 , \1624 );
nand \U$1283 ( \1626 , \924 , \899 );
not \U$1284 ( \1627 , \1468 );
nand \U$1285 ( \1628 , \1627 , \876 );
and \U$1286 ( \1629 , \1626 , \1628 );
nand \U$1287 ( \1630 , \1194 , \1165 );
and \U$1288 ( \1631 , \1629 , \1630 );
not \U$1289 ( \1632 , \1629 );
not \U$1290 ( \1633 , \1630 );
and \U$1291 ( \1634 , \1632 , \1633 );
nor \U$1292 ( \1635 , \1631 , \1634 );
not \U$1293 ( \1636 , \1635 );
or \U$1294 ( \1637 , \1625 , \1636 );
not \U$1295 ( \1638 , \1629 );
nand \U$1296 ( \1639 , \1638 , \1633 );
nand \U$1297 ( \1640 , \1637 , \1639 );
and \U$1298 ( \1641 , \1617 , \1640 );
not \U$1299 ( \1642 , \1617 );
not \U$1300 ( \1643 , \1640 );
and \U$1301 ( \1644 , \1642 , \1643 );
or \U$1302 ( \1645 , \1641 , \1644 );
not \U$1303 ( \1646 , \1645 );
and \U$1304 ( \1647 , RI9871b18_134, \1447 );
not \U$1305 ( \1648 , RI9871b18_134);
not \U$1306 ( \1649 , \1447 );
and \U$1307 ( \1650 , \1648 , \1649 );
nor \U$1308 ( \1651 , \1647 , \1650 );
not \U$1309 ( \1652 , \1651 );
not \U$1310 ( \1653 , \1543 );
and \U$1311 ( \1654 , \1652 , \1653 );
and \U$1312 ( \1655 , \1322 , \1292 );
nor \U$1313 ( \1656 , \1654 , \1655 );
not \U$1314 ( \1657 , \1656 );
buf \U$1315 ( \1658 , \1253 );
not \U$1316 ( \1659 , \1658 );
and \U$1317 ( \1660 , RI9871e60_141, \1659 );
not \U$1318 ( \1661 , RI9871e60_141);
and \U$1319 ( \1662 , \1661 , \1257 );
nor \U$1320 ( \1663 , \1660 , \1662 );
and \U$1321 ( \1664 , \1663 , \1353 );
and \U$1322 ( \1665 , \1346 , \1381 );
nor \U$1323 ( \1666 , \1664 , \1665 );
not \U$1324 ( \1667 , \1666 );
and \U$1325 ( \1668 , \1657 , \1667 );
xor \U$1326 ( \1669 , \1656 , \1666 );
and \U$1327 ( \1670 , \1111 , \1394 );
not \U$1328 ( \1671 , \1111 );
not \U$1329 ( \1672 , \1394 );
and \U$1330 ( \1673 , \1671 , \1672 );
nor \U$1331 ( \1674 , \1670 , \1673 );
or \U$1332 ( \1675 , \1674 , \1137 );
not \U$1333 ( \1676 , \1083 );
or \U$1334 ( \1677 , \1133 , \1676 );
nand \U$1335 ( \1678 , \1675 , \1677 );
and \U$1336 ( \1679 , \1669 , \1678 );
nor \U$1337 ( \1680 , \1668 , \1679 );
or \U$1338 ( \1681 , \1646 , \1680 );
or \U$1339 ( \1682 , \1643 , \1617 );
nand \U$1340 ( \1683 , \1681 , \1682 );
xor \U$1341 ( \1684 , \1576 , \1683 );
xor \U$1342 ( \1685 , \1537 , \1684 );
and \U$1343 ( \1686 , RI9871a28_132, RI9871aa0_133);
nor \U$1344 ( \1687 , \1686 , \1078 );
not \U$1345 ( \1688 , \1083 );
or \U$1346 ( \1689 , \1674 , \1688 );
buf \U$1347 ( \1690 , \778 );
not \U$1348 ( \1691 , \1690 );
not \U$1349 ( \1692 , \1691 );
not \U$1350 ( \1693 , \1692 );
and \U$1351 ( \1694 , \1693 , RI98718c0_129);
and \U$1352 ( \1695 , \1692 , \1111 );
nor \U$1353 ( \1696 , \1694 , \1695 );
or \U$1354 ( \1697 , \1696 , \1137 );
nand \U$1355 ( \1698 , \1689 , \1697 );
not \U$1356 ( \1699 , \1698 );
and \U$1357 ( \1700 , \1687 , \1699 );
not \U$1358 ( \1701 , \1687 );
and \U$1359 ( \1702 , \1701 , \1698 );
nor \U$1360 ( \1703 , \1700 , \1702 );
not \U$1361 ( \1704 , \1323 );
not \U$1362 ( \1705 , \1546 );
or \U$1363 ( \1706 , \1704 , \1705 );
or \U$1364 ( \1707 , \1651 , \1293 );
nand \U$1365 ( \1708 , \1706 , \1707 );
xnor \U$1366 ( \1709 , \1703 , \1708 );
not \U$1367 ( \1710 , \1596 );
not \U$1368 ( \1711 , \1162 );
or \U$1369 ( \1712 , \1710 , \1711 );
buf \U$1370 ( \1713 , \1061 );
not \U$1371 ( \1714 , \1713 );
and \U$1372 ( \1715 , \1714 , \1200 );
not \U$1373 ( \1716 , \1165 );
and \U$1374 ( \1717 , \1062 , \1716 );
nor \U$1375 ( \1718 , \1715 , \1717 );
not \U$1376 ( \1719 , \1220 );
or \U$1377 ( \1720 , \1718 , \1719 );
nand \U$1378 ( \1721 , \1712 , \1720 );
and \U$1379 ( \1722 , \1200 , \1212 );
xor \U$1380 ( \1723 , \1721 , \1722 );
not \U$1381 ( \1724 , \1125 );
buf \U$1382 ( \1725 , \1724 );
not \U$1383 ( \1726 , \1725 );
xnor \U$1384 ( \1727 , \1726 , RI9871c08_136);
or \U$1385 ( \1728 , \1727 , \1432 );
or \U$1386 ( \1729 , \1621 , \1457 );
nand \U$1387 ( \1730 , \1728 , \1729 );
not \U$1388 ( \1731 , \1730 );
and \U$1389 ( \1732 , \1723 , \1731 );
not \U$1390 ( \1733 , \1723 );
and \U$1391 ( \1734 , \1733 , \1730 );
nor \U$1392 ( \1735 , \1732 , \1734 );
xor \U$1393 ( \1736 , \1709 , \1735 );
not \U$1394 ( \1737 , \1501 );
not \U$1395 ( \1738 , \1588 );
or \U$1396 ( \1739 , \1737 , \1738 );
not \U$1397 ( \1740 , \1308 );
buf \U$1398 ( \1741 , \1740 );
and \U$1399 ( \1742 , \1584 , \1741 );
not \U$1400 ( \1743 , \1584 );
and \U$1401 ( \1744 , \1743 , \1320 );
nor \U$1402 ( \1745 , \1742 , \1744 );
not \U$1403 ( \1746 , \1518 );
or \U$1404 ( \1747 , \1745 , \1746 );
nand \U$1405 ( \1748 , \1739 , \1747 );
not \U$1406 ( \1749 , \1748 );
and \U$1407 ( \1750 , \1555 , \1353 );
and \U$1408 ( \1751 , \1663 , \1382 );
nor \U$1409 ( \1752 , \1750 , \1751 );
not \U$1410 ( \1753 , \1752 );
and \U$1411 ( \1754 , \1749 , \1753 );
and \U$1412 ( \1755 , \1748 , \1752 );
nor \U$1413 ( \1756 , \1754 , \1755 );
and \U$1414 ( \1757 , \1609 , \1018 );
not \U$1415 ( \1758 , \1044 );
and \U$1416 ( \1759 , \1340 , \1758 );
and \U$1417 ( \1760 , \1341 , \1044 );
nor \U$1418 ( \1761 , \1759 , \1760 );
and \U$1419 ( \1762 , \1761 , \1067 );
nor \U$1420 ( \1763 , \1757 , \1762 );
xor \U$1421 ( \1764 , \1756 , \1763 );
xor \U$1422 ( \1765 , \1736 , \1764 );
not \U$1423 ( \1766 , \1765 );
xnor \U$1424 ( \1767 , \1669 , \1678 );
not \U$1425 ( \1768 , \1767 );
not \U$1426 ( \1769 , \1768 );
xor \U$1427 ( \1770 , \1593 , \1600 );
xor \U$1428 ( \1771 , \1770 , \1614 );
xor \U$1429 ( \1772 , \1624 , \1635 );
xor \U$1430 ( \1773 , \1771 , \1772 );
not \U$1431 ( \1774 , \1773 );
or \U$1432 ( \1775 , \1769 , \1774 );
nand \U$1433 ( \1776 , \1772 , \1771 );
nand \U$1434 ( \1777 , \1775 , \1776 );
not \U$1435 ( \1778 , \1777 );
not \U$1436 ( \1779 , \1680 );
not \U$1437 ( \1780 , \1645 );
or \U$1438 ( \1781 , \1779 , \1780 );
or \U$1439 ( \1782 , \1645 , \1680 );
nand \U$1440 ( \1783 , \1781 , \1782 );
not \U$1441 ( \1784 , \1783 );
not \U$1442 ( \1785 , \1784 );
or \U$1443 ( \1786 , \1778 , \1785 );
not \U$1444 ( \1787 , \1777 );
nand \U$1445 ( \1788 , \1783 , \1787 );
nand \U$1446 ( \1789 , \1786 , \1788 );
not \U$1447 ( \1790 , \1789 );
or \U$1448 ( \1791 , \1766 , \1790 );
or \U$1449 ( \1792 , \1784 , \1787 );
nand \U$1450 ( \1793 , \1791 , \1792 );
and \U$1451 ( \1794 , \1685 , \1793 );
and \U$1452 ( \1795 , \1537 , \1684 );
nor \U$1453 ( \1796 , \1794 , \1795 );
not \U$1454 ( \1797 , \1796 );
not \U$1455 ( \1798 , \1518 );
buf \U$1456 ( \1799 , \1447 );
not \U$1457 ( \1800 , RI9871c80_137);
and \U$1458 ( \1801 , \1799 , \1800 );
not \U$1459 ( \1802 , \1799 );
and \U$1460 ( \1803 , \1802 , RI9871c80_137);
nor \U$1461 ( \1804 , \1801 , \1803 );
not \U$1462 ( \1805 , \1804 );
or \U$1463 ( \1806 , \1798 , \1805 );
or \U$1464 ( \1807 , \1745 , \1591 );
nand \U$1465 ( \1808 , \1806 , \1807 );
not \U$1466 ( \1809 , \1162 );
or \U$1467 ( \1810 , \1718 , \1809 );
and \U$1468 ( \1811 , \1371 , \1199 );
not \U$1469 ( \1812 , \1371 );
and \U$1470 ( \1813 , \1812 , \1165 );
nor \U$1471 ( \1814 , \1811 , \1813 );
or \U$1472 ( \1815 , \1814 , \1719 );
nand \U$1473 ( \1816 , \1810 , \1815 );
xor \U$1474 ( \1817 , \1808 , \1816 );
and \U$1475 ( \1818 , \1761 , \1018 );
and \U$1476 ( \1819 , \1257 , \1758 );
not \U$1477 ( \1820 , \1257 );
and \U$1478 ( \1821 , \1820 , \1044 );
nor \U$1479 ( \1822 , \1819 , \1821 );
and \U$1480 ( \1823 , \1822 , \1067 );
nor \U$1481 ( \1824 , \1818 , \1823 );
not \U$1482 ( \1825 , \1824 );
xor \U$1483 ( \1826 , \1817 , \1825 );
not \U$1484 ( \1827 , \1826 );
and \U$1485 ( \1828 , \1723 , \1730 );
and \U$1486 ( \1829 , \1721 , \1722 );
nor \U$1487 ( \1830 , \1828 , \1829 );
not \U$1488 ( \1831 , \876 );
not \U$1489 ( \1832 , \923 );
or \U$1490 ( \1833 , \1831 , \1832 );
not \U$1491 ( \1834 , \1582 );
not \U$1492 ( \1835 , \1834 );
not \U$1493 ( \1836 , RI9872130_147);
and \U$1494 ( \1837 , \1835 , \1836 );
not \U$1495 ( \1838 , \1582 );
and \U$1496 ( \1839 , \1838 , RI9872130_147);
nor \U$1497 ( \1840 , \1837 , \1839 );
not \U$1498 ( \1841 , \1840 );
nand \U$1499 ( \1842 , \1841 , \924 );
nand \U$1500 ( \1843 , \1833 , \1842 );
and \U$1501 ( \1844 , \1200 , \1595 );
xor \U$1502 ( \1845 , \1843 , \1844 );
not \U$1503 ( \1846 , \1845 );
not \U$1504 ( \1847 , \1727 );
not \U$1505 ( \1848 , \1457 );
and \U$1506 ( \1849 , \1847 , \1848 );
not \U$1507 ( \1850 , RI9871c08_136);
and \U$1508 ( \1851 , \1850 , \1672 );
not \U$1509 ( \1852 , \1850 );
and \U$1510 ( \1853 , \1852 , \1394 );
nor \U$1511 ( \1854 , \1851 , \1853 );
and \U$1512 ( \1855 , \1854 , \1431 );
nor \U$1513 ( \1856 , \1849 , \1855 );
not \U$1514 ( \1857 , \1856 );
and \U$1515 ( \1858 , \1846 , \1857 );
and \U$1516 ( \1859 , \1845 , \1856 );
nor \U$1517 ( \1860 , \1858 , \1859 );
and \U$1518 ( \1861 , \1830 , \1860 );
not \U$1519 ( \1862 , \1830 );
not \U$1520 ( \1863 , \1860 );
and \U$1521 ( \1864 , \1862 , \1863 );
nor \U$1522 ( \1865 , \1861 , \1864 );
not \U$1523 ( \1866 , \1865 );
or \U$1524 ( \1867 , \1827 , \1866 );
or \U$1525 ( \1868 , \1830 , \1860 );
nand \U$1526 ( \1869 , \1867 , \1868 );
not \U$1527 ( \1870 , \1699 );
not \U$1528 ( \1871 , \1687 );
and \U$1529 ( \1872 , \1870 , \1871 );
and \U$1530 ( \1873 , \1703 , \1708 );
nor \U$1531 ( \1874 , \1872 , \1873 );
or \U$1532 ( \1875 , \1696 , \1676 );
or \U$1533 ( \1876 , \1137 , \1111 );
nand \U$1534 ( \1877 , \1875 , \1876 );
not \U$1535 ( \1878 , \1877 );
and \U$1536 ( \1879 , \1874 , \1878 );
not \U$1537 ( \1880 , \1874 );
and \U$1538 ( \1881 , \1880 , \1877 );
nor \U$1539 ( \1882 , \1879 , \1881 );
or \U$1540 ( \1883 , \1756 , \1763 );
not \U$1541 ( \1884 , \1748 );
or \U$1542 ( \1885 , \1884 , \1752 );
nand \U$1543 ( \1886 , \1883 , \1885 );
not \U$1544 ( \1887 , \1886 );
or \U$1545 ( \1888 , \1882 , \1887 );
or \U$1546 ( \1889 , \1874 , \1877 );
nand \U$1547 ( \1890 , \1888 , \1889 );
xor \U$1548 ( \1891 , \1869 , \1890 );
or \U$1549 ( \1892 , \1564 , \1568 );
or \U$1550 ( \1893 , \1563 , \1548 );
nand \U$1551 ( \1894 , \1892 , \1893 );
not \U$1552 ( \1895 , \1844 );
not \U$1553 ( \1896 , \1843 );
or \U$1554 ( \1897 , \1895 , \1896 );
not \U$1555 ( \1898 , \1856 );
nand \U$1556 ( \1899 , \1898 , \1845 );
nand \U$1557 ( \1900 , \1897 , \1899 );
xor \U$1558 ( \1901 , \1894 , \1900 );
not \U$1559 ( \1902 , \1541 );
not \U$1560 ( \1903 , \1293 );
and \U$1561 ( \1904 , \1902 , \1903 );
and \U$1562 ( \1905 , RI9871b18_134, \1726 );
not \U$1563 ( \1906 , RI9871b18_134);
and \U$1564 ( \1907 , \1906 , \1128 );
nor \U$1565 ( \1908 , \1905 , \1907 );
and \U$1566 ( \1909 , \1908 , \1323 );
nor \U$1567 ( \1910 , \1904 , \1909 );
nand \U$1568 ( \1911 , \1062 , \1200 );
xor \U$1569 ( \1912 , \1910 , \1911 );
and \U$1570 ( \1913 , \916 , \1347 );
and \U$1571 ( \1914 , \1513 , RI9871d70_139);
nor \U$1572 ( \1915 , \1913 , \1914 );
and \U$1573 ( \1916 , \1915 , \832 );
and \U$1574 ( \1917 , \1565 , \859 );
nor \U$1575 ( \1918 , \1916 , \1917 );
xor \U$1576 ( \1919 , \1912 , \1918 );
not \U$1577 ( \1920 , \1919 );
xor \U$1578 ( \1921 , \1901 , \1920 );
xor \U$1579 ( \1922 , \1891 , \1921 );
not \U$1580 ( \1923 , \1735 );
not \U$1581 ( \1924 , \1709 );
and \U$1582 ( \1925 , \1923 , \1924 );
and \U$1583 ( \1926 , \1736 , \1764 );
nor \U$1584 ( \1927 , \1925 , \1926 );
and \U$1585 ( \1928 , \1882 , \1886 );
not \U$1586 ( \1929 , \1882 );
and \U$1587 ( \1930 , \1929 , \1887 );
nor \U$1588 ( \1931 , \1928 , \1930 );
xnor \U$1589 ( \1932 , \1927 , \1931 );
xnor \U$1590 ( \1933 , \1865 , \1826 );
or \U$1591 ( \1934 , \1932 , \1933 );
or \U$1592 ( \1935 , \1927 , \1931 );
nand \U$1593 ( \1936 , \1934 , \1935 );
and \U$1594 ( \1937 , RI9872130_147, \1320 );
not \U$1595 ( \1938 , RI9872130_147);
and \U$1596 ( \1939 , \1938 , \1311 );
nor \U$1597 ( \1940 , \1937 , \1939 );
or \U$1598 ( \1941 , \1940 , \1470 );
not \U$1599 ( \1942 , \876 );
or \U$1600 ( \1943 , \1840 , \1942 );
nand \U$1601 ( \1944 , \1941 , \1943 );
not \U$1602 ( \1945 , \1944 );
not \U$1603 ( \1946 , \1814 );
not \U$1604 ( \1947 , \1809 );
and \U$1605 ( \1948 , \1946 , \1947 );
not \U$1606 ( \1949 , \1344 );
nand \U$1607 ( \1950 , \1949 , \1165 );
nand \U$1608 ( \1951 , \1344 , \1199 );
and \U$1609 ( \1952 , \1950 , \1951 );
and \U$1610 ( \1953 , \1952 , \1220 );
nor \U$1611 ( \1954 , \1948 , \1953 );
not \U$1612 ( \1955 , \1954 );
and \U$1613 ( \1956 , \1945 , \1955 );
and \U$1614 ( \1957 , \1944 , \1954 );
nor \U$1615 ( \1958 , \1956 , \1957 );
and \U$1616 ( \1959 , \1822 , \1018 );
not \U$1617 ( \1960 , \944 );
xor \U$1618 ( \1961 , \1045 , \1960 );
and \U$1619 ( \1962 , \1961 , \1067 );
nor \U$1620 ( \1963 , \1959 , \1962 );
xor \U$1621 ( \1964 , \1958 , \1963 );
and \U$1622 ( \1965 , \1854 , \1456 );
xor \U$1623 ( \1966 , \780 , RI9871c08_136);
and \U$1624 ( \1967 , \1966 , \1431 );
nor \U$1625 ( \1968 , \1965 , \1967 );
and \U$1626 ( \1969 , \1688 , \1137 );
nor \U$1627 ( \1970 , \1969 , \1111 );
xnor \U$1628 ( \1971 , \1968 , \1970 );
and \U$1629 ( \1972 , \1800 , \1418 );
not \U$1630 ( \1973 , \1800 );
and \U$1631 ( \1974 , \1973 , \1417 );
nor \U$1632 ( \1975 , \1972 , \1974 );
and \U$1633 ( \1976 , \1975 , \1518 );
and \U$1634 ( \1977 , \1804 , \1501 );
nor \U$1635 ( \1978 , \1976 , \1977 );
xor \U$1636 ( \1979 , \1971 , \1978 );
xnor \U$1637 ( \1980 , \1964 , \1979 );
xor \U$1638 ( \1981 , \1808 , \1816 );
not \U$1639 ( \1982 , \1824 );
and \U$1640 ( \1983 , \1981 , \1982 );
and \U$1641 ( \1984 , \1808 , \1816 );
or \U$1642 ( \1985 , \1983 , \1984 );
not \U$1643 ( \1986 , \1985 );
xnor \U$1644 ( \1987 , \821 , RI9871e60_141);
not \U$1645 ( \1988 , \1987 );
not \U$1646 ( \1989 , \1353 );
not \U$1647 ( \1990 , \1989 );
and \U$1648 ( \1991 , \1988 , \1990 );
and \U$1649 ( \1992 , \1561 , \1382 );
nor \U$1650 ( \1993 , \1991 , \1992 );
and \U$1651 ( \1994 , \1993 , \1877 );
not \U$1652 ( \1995 , \1993 );
and \U$1653 ( \1996 , \1995 , \1878 );
nor \U$1654 ( \1997 , \1994 , \1996 );
xnor \U$1655 ( \1998 , \1986 , \1997 );
not \U$1656 ( \1999 , \1998 );
xor \U$1657 ( \2000 , \1980 , \1999 );
not \U$1658 ( \2001 , \2000 );
xor \U$1659 ( \2002 , \1569 , \1575 );
and \U$1660 ( \2003 , \2002 , \1683 );
and \U$1661 ( \2004 , \1569 , \1575 );
or \U$1662 ( \2005 , \2003 , \2004 );
not \U$1663 ( \2006 , \2005 );
or \U$1664 ( \2007 , \2001 , \2006 );
or \U$1665 ( \2008 , \2005 , \2000 );
nand \U$1666 ( \2009 , \2007 , \2008 );
xor \U$1667 ( \2010 , \1936 , \2009 );
xor \U$1668 ( \2011 , \1922 , \2010 );
not \U$1669 ( \2012 , \2011 );
or \U$1670 ( \2013 , \1797 , \2012 );
or \U$1671 ( \2014 , \2011 , \1796 );
nand \U$1672 ( \2015 , \2013 , \2014 );
not \U$1673 ( \2016 , \2015 );
and \U$1674 ( \2017 , \1403 , \1460 );
not \U$1675 ( \2018 , \1403 );
and \U$1676 ( \2019 , \2018 , \1459 );
nor \U$1677 ( \2020 , \2017 , \2019 );
xor \U$1678 ( \2021 , \1261 , \1325 );
xor \U$1679 ( \2022 , \2021 , \1384 );
not \U$1680 ( \2023 , \2022 );
xor \U$1681 ( \2024 , \2020 , \2023 );
xor \U$1682 ( \2025 , \1223 , \1070 );
and \U$1683 ( \2026 , \2024 , \2025 );
and \U$1684 ( \2027 , \2020 , \2023 );
nor \U$1685 ( \2028 , \2026 , \2027 );
not \U$1686 ( \2029 , \2028 );
not \U$1687 ( \2030 , \2029 );
xnor \U$1688 ( \2031 , \1227 , \1228 );
not \U$1689 ( \2032 , \2031 );
not \U$1690 ( \2033 , \1448 );
not \U$1691 ( \2034 , \1432 );
and \U$1692 ( \2035 , \2033 , \2034 );
and \U$1693 ( \2036 , RI9871c08_136, \1741 );
not \U$1694 ( \2037 , RI9871c08_136);
buf \U$1695 ( \2038 , \1320 );
and \U$1696 ( \2039 , \2037 , \2038 );
nor \U$1697 ( \2040 , \2036 , \2039 );
and \U$1698 ( \2041 , \2040 , \1456 );
nor \U$1699 ( \2042 , \2035 , \2041 );
and \U$1700 ( \2043 , RI98719b0_131, \1128 );
not \U$1701 ( \2044 , RI98719b0_131);
and \U$1702 ( \2045 , \2044 , \1726 );
nor \U$1703 ( \2046 , \2043 , \2045 );
not \U$1704 ( \2047 , \2046 );
not \U$1705 ( \2048 , \1398 );
and \U$1706 ( \2049 , \2047 , \2048 );
and \U$1707 ( \2050 , \1395 , \797 );
nor \U$1708 ( \2051 , \2049 , \2050 );
xor \U$1709 ( \2052 , \2042 , \2051 );
xnor \U$1710 ( \2053 , \1341 , RI9871d70_139);
not \U$1711 ( \2054 , \2053 );
not \U$1712 ( \2055 , \860 );
and \U$1713 ( \2056 , \2054 , \2055 );
and \U$1714 ( \2057 , \1259 , \832 );
nor \U$1715 ( \2058 , \2056 , \2057 );
and \U$1716 ( \2059 , \2052 , \2058 );
and \U$1717 ( \2060 , \2042 , \2051 );
nor \U$1718 ( \2061 , \2059 , \2060 );
not \U$1719 ( \2062 , \2061 );
xor \U$1720 ( \2063 , RI9872298_150, RI9872310_151);
not \U$1721 ( \2064 , \2063 );
and \U$1722 ( \2065 , RI9871aa0_133, RI9872298_150);
not \U$1723 ( \2066 , RI9871aa0_133);
not \U$1724 ( \2067 , RI9872298_150);
and \U$1725 ( \2068 , \2066 , \2067 );
nor \U$1726 ( \2069 , \2065 , \2068 );
and \U$1727 ( \2070 , \2064 , \2069 );
buf \U$1728 ( \2071 , \2070 );
buf \U$1729 ( \2072 , \2071 );
not \U$1730 ( \2073 , \2072 );
not \U$1731 ( \2074 , \2073 );
not \U$1732 ( \2075 , \2074 );
not \U$1733 ( \2076 , RI9871aa0_133);
not \U$1734 ( \2077 , \2076 );
not \U$1735 ( \2078 , \780 );
or \U$1736 ( \2079 , \2077 , \2078 );
not \U$1737 ( \2080 , RI9871aa0_133);
or \U$1738 ( \2081 , \1692 , \2080 );
nand \U$1739 ( \2082 , \2079 , \2081 );
not \U$1740 ( \2083 , \2082 );
or \U$1741 ( \2084 , \2075 , \2083 );
buf \U$1742 ( \2085 , \2063 );
not \U$1743 ( \2086 , \2085 );
not \U$1744 ( \2087 , \2086 );
nand \U$1745 ( \2088 , \2087 , RI9871aa0_133);
nand \U$1746 ( \2089 , \2084 , \2088 );
xnor \U$1747 ( \2090 , \1417 , RI98718c0_129);
not \U$1748 ( \2091 , \2090 );
not \U$1749 ( \2092 , \1688 );
and \U$1750 ( \2093 , \2091 , \2092 );
and \U$1751 ( \2094 , \1108 , \1136 );
nor \U$1752 ( \2095 , \2093 , \2094 );
not \U$1753 ( \2096 , \2095 );
not \U$1754 ( \2097 , \2096 );
nand \U$1755 ( \2098 , \388 , \444 );
not \U$1756 ( \2099 , \2098 );
and \U$1757 ( \2100 , \386 , \387 );
not \U$1758 ( \2101 , \2100 );
not \U$1759 ( \2102 , \1177 );
or \U$1760 ( \2103 , \2101 , \2102 );
not \U$1761 ( \2104 , \441 );
nand \U$1762 ( \2105 , \2103 , \2104 );
not \U$1763 ( \2106 , \2105 );
or \U$1764 ( \2107 , \2099 , \2106 );
or \U$1765 ( \2108 , \2098 , \2105 );
nand \U$1766 ( \2109 , \2107 , \2108 );
buf \U$1767 ( \2110 , \2109 );
buf \U$1768 ( \2111 , \2110 );
and \U$1769 ( \2112 , \2111 , \1200 );
not \U$1770 ( \2113 , \1220 );
not \U$1771 ( \2114 , \1196 );
or \U$1772 ( \2115 , \2113 , \2114 );
buf \U$1773 ( \2116 , \1485 );
and \U$1774 ( \2117 , \2116 , \1165 );
not \U$1775 ( \2118 , \2116 );
and \U$1776 ( \2119 , \2118 , \1199 );
nor \U$1777 ( \2120 , \2117 , \2119 );
or \U$1778 ( \2121 , \2120 , \1809 );
nand \U$1779 ( \2122 , \2115 , \2121 );
xor \U$1780 ( \2123 , \2112 , \2122 );
not \U$1781 ( \2124 , \2123 );
or \U$1782 ( \2125 , \2097 , \2124 );
nand \U$1783 ( \2126 , \2122 , \2112 );
nand \U$1784 ( \2127 , \2125 , \2126 );
xor \U$1785 ( \2128 , \2089 , \2127 );
not \U$1786 ( \2129 , \2128 );
or \U$1787 ( \2130 , \2062 , \2129 );
nand \U$1788 ( \2131 , \2127 , \2089 );
nand \U$1789 ( \2132 , \2130 , \2131 );
not \U$1790 ( \2133 , \2132 );
or \U$1791 ( \2134 , \2032 , \2133 );
or \U$1792 ( \2135 , \2132 , \2031 );
nand \U$1793 ( \2136 , \2134 , \2135 );
not \U$1794 ( \2137 , \2136 );
or \U$1795 ( \2138 , \2030 , \2137 );
not \U$1796 ( \2139 , \2031 );
nand \U$1797 ( \2140 , \2139 , \2132 );
nand \U$1798 ( \2141 , \2138 , \2140 );
not \U$1799 ( \2142 , \1535 );
not \U$1800 ( \2143 , \1237 );
and \U$1801 ( \2144 , \2142 , \2143 );
and \U$1802 ( \2145 , \1535 , \1237 );
nor \U$1803 ( \2146 , \2144 , \2145 );
xor \U$1804 ( \2147 , \2141 , \2146 );
not \U$1805 ( \2148 , \2147 );
xor \U$1806 ( \2149 , \1789 , \1765 );
not \U$1807 ( \2150 , \2149 );
not \U$1808 ( \2151 , \2150 );
and \U$1809 ( \2152 , \2148 , \2151 );
not \U$1810 ( \2153 , \2146 );
and \U$1811 ( \2154 , \2141 , \2153 );
nor \U$1812 ( \2155 , \2152 , \2154 );
not \U$1813 ( \2156 , \2155 );
not \U$1814 ( \2157 , \2156 );
xor \U$1815 ( \2158 , \1932 , \1933 );
not \U$1816 ( \2159 , \1793 );
and \U$1817 ( \2160 , \1685 , \2159 );
not \U$1818 ( \2161 , \1685 );
and \U$1819 ( \2162 , \2161 , \1793 );
nor \U$1820 ( \2163 , \2160 , \2162 );
and \U$1821 ( \2164 , \2158 , \2163 );
not \U$1822 ( \2165 , \2158 );
not \U$1823 ( \2166 , \2163 );
and \U$1824 ( \2167 , \2165 , \2166 );
or \U$1825 ( \2168 , \2164 , \2167 );
not \U$1826 ( \2169 , \2168 );
or \U$1827 ( \2170 , \2157 , \2169 );
nand \U$1828 ( \2171 , \2166 , \2158 );
nand \U$1829 ( \2172 , \2170 , \2171 );
not \U$1830 ( \2173 , \2172 );
nand \U$1831 ( \2174 , \2016 , \2173 );
or \U$1832 ( \2175 , \1986 , \1997 );
or \U$1833 ( \2176 , \1993 , \1878 );
nand \U$1834 ( \2177 , \2175 , \2176 );
and \U$1835 ( \2178 , \1901 , \1920 );
and \U$1836 ( \2179 , \1894 , \1900 );
nor \U$1837 ( \2180 , \2178 , \2179 );
not \U$1838 ( \2181 , \2180 );
and \U$1839 ( \2182 , \2177 , \2181 );
not \U$1840 ( \2183 , \2177 );
and \U$1841 ( \2184 , \2183 , \2180 );
nor \U$1842 ( \2185 , \2182 , \2184 );
or \U$1843 ( \2186 , \1971 , \1978 );
or \U$1844 ( \2187 , \1968 , \1970 );
nand \U$1845 ( \2188 , \2186 , \2187 );
xor \U$1846 ( \2189 , \1910 , \1911 );
and \U$1847 ( \2190 , \2189 , \1918 );
and \U$1848 ( \2191 , \1910 , \1911 );
nor \U$1849 ( \2192 , \2190 , \2191 );
xor \U$1850 ( \2193 , \2188 , \2192 );
or \U$1851 ( \2194 , \1958 , \1963 );
not \U$1852 ( \2195 , \1944 );
or \U$1853 ( \2196 , \2195 , \1954 );
nand \U$1854 ( \2197 , \2194 , \2196 );
xor \U$1855 ( \2198 , \2193 , \2197 );
xor \U$1856 ( \2199 , \2185 , \2198 );
not \U$1857 ( \2200 , \2199 );
not \U$1858 ( \2201 , \1936 );
not \U$1859 ( \2202 , \2009 );
or \U$1860 ( \2203 , \2201 , \2202 );
not \U$1861 ( \2204 , \2000 );
nand \U$1862 ( \2205 , \2204 , \2005 );
nand \U$1863 ( \2206 , \2203 , \2205 );
not \U$1864 ( \2207 , \2206 );
or \U$1865 ( \2208 , \2200 , \2207 );
xor \U$1866 ( \2209 , \2206 , \2199 );
not \U$1867 ( \2210 , \2209 );
not \U$1868 ( \2211 , \847 );
not \U$1869 ( \2212 , \2211 );
not \U$1870 ( \2213 , \1045 );
and \U$1871 ( \2214 , \2212 , \2213 );
not \U$1872 ( \2215 , \846 );
buf \U$1873 ( \2216 , \2215 );
and \U$1874 ( \2217 , \2216 , \1045 );
nor \U$1875 ( \2218 , \2214 , \2217 );
not \U$1876 ( \2219 , \2218 );
not \U$1877 ( \2220 , \2219 );
not \U$1878 ( \2221 , \1068 );
and \U$1879 ( \2222 , \2220 , \2221 );
and \U$1880 ( \2223 , \1961 , \1018 );
nor \U$1881 ( \2224 , \2222 , \2223 );
not \U$1882 ( \2225 , \2224 );
and \U$1883 ( \2226 , \1966 , \1456 );
and \U$1884 ( \2227 , \1431 , RI9871c08_136);
nor \U$1885 ( \2228 , \2226 , \2227 );
not \U$1886 ( \2229 , \2228 );
and \U$1887 ( \2230 , \2225 , \2229 );
and \U$1888 ( \2231 , \2224 , \2228 );
nor \U$1889 ( \2232 , \2230 , \2231 );
not \U$1890 ( \2233 , \1987 );
not \U$1891 ( \2234 , \1558 );
and \U$1892 ( \2235 , \2233 , \2234 );
and \U$1893 ( \2236 , RI9871e60_141, \895 );
not \U$1894 ( \2237 , RI9871e60_141);
and \U$1895 ( \2238 , \2237 , \894 );
nor \U$1896 ( \2239 , \2236 , \2238 );
and \U$1897 ( \2240 , \2239 , \1353 );
nor \U$1898 ( \2241 , \2235 , \2240 );
xor \U$1899 ( \2242 , \2232 , \2241 );
not \U$1900 ( \2243 , RI9871d70_139);
and \U$1901 ( \2244 , \2243 , \1583 );
not \U$1902 ( \2245 , \2243 );
and \U$1903 ( \2246 , \2245 , \1275 );
nor \U$1904 ( \2247 , \2244 , \2246 );
and \U$1905 ( \2248 , \2247 , \832 );
and \U$1906 ( \2249 , \1915 , \859 );
nor \U$1907 ( \2250 , \2248 , \2249 );
not \U$1908 ( \2251 , \2250 );
and \U$1909 ( \2252 , \1106 , \1584 );
not \U$1910 ( \2253 , \1106 );
and \U$1911 ( \2254 , \2253 , RI9871c80_137);
nor \U$1912 ( \2255 , \2252 , \2254 );
not \U$1913 ( \2256 , \2255 );
not \U$1914 ( \2257 , \1746 );
and \U$1915 ( \2258 , \2256 , \2257 );
and \U$1916 ( \2259 , \1975 , \1501 );
nor \U$1917 ( \2260 , \2258 , \2259 );
xor \U$1918 ( \2261 , \1394 , RI9871b18_134);
not \U$1919 ( \2262 , \2261 );
not \U$1920 ( \2263 , \2262 );
not \U$1921 ( \2264 , \1543 );
and \U$1922 ( \2265 , \2263 , \2264 );
and \U$1923 ( \2266 , \1908 , \1292 );
nor \U$1924 ( \2267 , \2265 , \2266 );
xor \U$1925 ( \2268 , \2260 , \2267 );
not \U$1926 ( \2269 , \2268 );
or \U$1927 ( \2270 , \2251 , \2269 );
or \U$1928 ( \2271 , \2268 , \2250 );
nand \U$1929 ( \2272 , \2270 , \2271 );
xor \U$1930 ( \2273 , \2242 , \2272 );
not \U$1931 ( \2274 , \924 );
xnor \U$1932 ( \2275 , \1447 , RI9872130_147);
not \U$1933 ( \2276 , \2275 );
or \U$1934 ( \2277 , \2274 , \2276 );
not \U$1935 ( \2278 , \1940 );
nand \U$1936 ( \2279 , \2278 , \876 );
nand \U$1937 ( \2280 , \2277 , \2279 );
and \U$1938 ( \2281 , \1605 , \1165 );
xnor \U$1939 ( \2282 , \2280 , \2281 );
and \U$1940 ( \2283 , \1952 , \1162 );
and \U$1941 ( \2284 , \1257 , \1716 );
nand \U$1942 ( \2285 , \1659 , \1200 );
not \U$1943 ( \2286 , \2285 );
nor \U$1944 ( \2287 , \2284 , \2286 );
and \U$1945 ( \2288 , \2287 , \1220 );
nor \U$1946 ( \2289 , \2283 , \2288 );
xor \U$1947 ( \2290 , \2282 , \2289 );
xnor \U$1948 ( \2291 , \2273 , \2290 );
not \U$1949 ( \2292 , \1980 );
not \U$1950 ( \2293 , \1998 );
and \U$1951 ( \2294 , \2292 , \2293 );
and \U$1952 ( \2295 , \1964 , \1979 );
nor \U$1953 ( \2296 , \2294 , \2295 );
xor \U$1954 ( \2297 , \2291 , \2296 );
and \U$1955 ( \2298 , \1869 , \1890 );
and \U$1956 ( \2299 , \1891 , \1921 );
nor \U$1957 ( \2300 , \2298 , \2299 );
xor \U$1958 ( \2301 , \2297 , \2300 );
or \U$1959 ( \2302 , \2210 , \2301 );
nand \U$1960 ( \2303 , \2208 , \2302 );
xor \U$1961 ( \2304 , \2291 , \2296 );
and \U$1962 ( \2305 , \2304 , \2300 );
and \U$1963 ( \2306 , \2291 , \2296 );
or \U$1964 ( \2307 , \2305 , \2306 );
xor \U$1965 ( \2308 , \2188 , \2192 );
and \U$1966 ( \2309 , \2308 , \2197 );
and \U$1967 ( \2310 , \2188 , \2192 );
nor \U$1968 ( \2311 , \2309 , \2310 );
not \U$1969 ( \2312 , RI9871d70_139);
and \U$1970 ( \2313 , \2312 , \1320 );
not \U$1971 ( \2314 , \2312 );
and \U$1972 ( \2315 , \2314 , \1741 );
nor \U$1973 ( \2316 , \2313 , \2315 );
and \U$1974 ( \2317 , \2316 , \832 );
and \U$1975 ( \2318 , \2247 , \859 );
nor \U$1976 ( \2319 , \2317 , \2318 );
xor \U$1977 ( \2320 , \2319 , \1950 );
or \U$1978 ( \2321 , \944 , \1200 );
nand \U$1979 ( \2322 , \944 , \1200 );
nand \U$1980 ( \2323 , \2321 , \2322 );
not \U$1981 ( \2324 , \2323 );
not \U$1982 ( \2325 , \1719 );
and \U$1983 ( \2326 , \2324 , \2325 );
and \U$1984 ( \2327 , \2287 , \1162 );
nor \U$1985 ( \2328 , \2326 , \2327 );
xor \U$1986 ( \2329 , \2320 , \2328 );
xor \U$1987 ( \2330 , \2311 , \2329 );
not \U$1988 ( \2331 , \2282 );
not \U$1989 ( \2332 , \2289 );
and \U$1990 ( \2333 , \2331 , \2332 );
and \U$1991 ( \2334 , \2280 , \2281 );
nor \U$1992 ( \2335 , \2333 , \2334 );
and \U$1993 ( \2336 , \2335 , \2228 );
not \U$1994 ( \2337 , \2335 );
not \U$1995 ( \2338 , \2228 );
and \U$1996 ( \2339 , \2337 , \2338 );
nor \U$1997 ( \2340 , \2336 , \2339 );
not \U$1998 ( \2341 , \2268 );
or \U$1999 ( \2342 , \2341 , \2250 );
or \U$2000 ( \2343 , \2260 , \2267 );
nand \U$2001 ( \2344 , \2342 , \2343 );
xnor \U$2002 ( \2345 , \2340 , \2344 );
xor \U$2003 ( \2346 , \2330 , \2345 );
xor \U$2004 ( \2347 , \2307 , \2346 );
and \U$2005 ( \2348 , \2185 , \2198 );
and \U$2006 ( \2349 , \2181 , \2177 );
nor \U$2007 ( \2350 , \2348 , \2349 );
and \U$2008 ( \2351 , \2273 , \2290 );
and \U$2009 ( \2352 , \2272 , \2242 );
nor \U$2010 ( \2353 , \2351 , \2352 );
or \U$2011 ( \2354 , \2232 , \2241 );
or \U$2012 ( \2355 , \2224 , \2338 );
nand \U$2013 ( \2356 , \2354 , \2355 );
nand \U$2014 ( \2357 , RI98718c0_129, RI98720b8_146);
and \U$2015 ( \2358 , \2357 , RI9871c08_136);
not \U$2016 ( \2359 , RI9871b18_134);
not \U$2017 ( \2360 , \1690 );
not \U$2018 ( \2361 , \2360 );
not \U$2019 ( \2362 , \2361 );
or \U$2020 ( \2363 , \2359 , \2362 );
or \U$2021 ( \2364 , \1692 , RI9871b18_134);
nand \U$2022 ( \2365 , \2363 , \2364 );
not \U$2023 ( \2366 , \2365 );
not \U$2024 ( \2367 , \1543 );
and \U$2025 ( \2368 , \2366 , \2367 );
and \U$2026 ( \2369 , \2261 , \1292 );
nor \U$2027 ( \2370 , \2368 , \2369 );
xor \U$2028 ( \2371 , \2358 , \2370 );
and \U$2029 ( \2372 , \1418 , \919 );
and \U$2030 ( \2373 , \1417 , RI9872130_147);
nor \U$2031 ( \2374 , \2372 , \2373 );
and \U$2032 ( \2375 , \2374 , \924 );
and \U$2033 ( \2376 , \2275 , \876 );
nor \U$2034 ( \2377 , \2375 , \2376 );
not \U$2035 ( \2378 , \2377 );
and \U$2036 ( \2379 , \2371 , \2378 );
not \U$2037 ( \2380 , \2371 );
and \U$2038 ( \2381 , \2380 , \2377 );
nor \U$2039 ( \2382 , \2379 , \2381 );
xor \U$2040 ( \2383 , \2356 , \2382 );
and \U$2041 ( \2384 , RI9871e60_141, \916 );
not \U$2042 ( \2385 , RI9871e60_141);
and \U$2043 ( \2386 , \2385 , \1513 );
nor \U$2044 ( \2387 , \2384 , \2386 );
not \U$2045 ( \2388 , \2387 );
not \U$2046 ( \2389 , \1989 );
and \U$2047 ( \2390 , \2388 , \2389 );
and \U$2048 ( \2391 , \2239 , \1382 );
nor \U$2049 ( \2392 , \2390 , \2391 );
not \U$2050 ( \2393 , \2255 );
not \U$2051 ( \2394 , \1591 );
and \U$2052 ( \2395 , \2393 , \2394 );
and \U$2053 ( \2396 , RI9871c80_137, \1129 );
not \U$2054 ( \2397 , RI9871c80_137);
not \U$2055 ( \2398 , \1125 );
buf \U$2056 ( \2399 , \2398 );
and \U$2057 ( \2400 , \2397 , \2399 );
nor \U$2058 ( \2401 , \2396 , \2400 );
and \U$2059 ( \2402 , \2401 , \1518 );
nor \U$2060 ( \2403 , \2395 , \2402 );
xor \U$2061 ( \2404 , \2392 , \2403 );
and \U$2062 ( \2405 , \2218 , \1018 );
xor \U$2063 ( \2406 , \1758 , \824 );
and \U$2064 ( \2407 , \2406 , \1067 );
nor \U$2065 ( \2408 , \2405 , \2407 );
xor \U$2066 ( \2409 , \2404 , \2408 );
not \U$2067 ( \2410 , \2409 );
xnor \U$2068 ( \2411 , \2383 , \2410 );
xnor \U$2069 ( \2412 , \2353 , \2411 );
xnor \U$2070 ( \2413 , \2350 , \2412 );
xor \U$2071 ( \2414 , \2347 , \2413 );
not \U$2072 ( \2415 , \2414 );
or \U$2073 ( \2416 , \2303 , \2415 );
xor \U$2074 ( \2417 , \2311 , \2329 );
and \U$2075 ( \2418 , \2417 , \2345 );
and \U$2076 ( \2419 , \2311 , \2329 );
nor \U$2077 ( \2420 , \2418 , \2419 );
xor \U$2078 ( \2421 , \2392 , \2403 );
and \U$2079 ( \2422 , \2421 , \2408 );
and \U$2080 ( \2423 , \2392 , \2403 );
nor \U$2081 ( \2424 , \2422 , \2423 );
xor \U$2082 ( \2425 , \2319 , \1950 );
and \U$2083 ( \2426 , \2425 , \2328 );
and \U$2084 ( \2427 , \2319 , \1950 );
nor \U$2085 ( \2428 , \2426 , \2427 );
xor \U$2086 ( \2429 , \2424 , \2428 );
and \U$2087 ( \2430 , RI9872130_147, \1106 );
not \U$2088 ( \2431 , RI9872130_147);
and \U$2089 ( \2432 , \2431 , \1098 );
nor \U$2090 ( \2433 , \2430 , \2432 );
and \U$2091 ( \2434 , \2433 , \924 );
and \U$2092 ( \2435 , \2374 , \876 );
nor \U$2093 ( \2436 , \2434 , \2435 );
and \U$2094 ( \2437 , \1367 , \1275 );
not \U$2095 ( \2438 , \1367 );
and \U$2096 ( \2439 , \2438 , \1834 );
nor \U$2097 ( \2440 , \2437 , \2439 );
or \U$2098 ( \2441 , \2440 , \1989 );
or \U$2099 ( \2442 , \2387 , \1558 );
nand \U$2100 ( \2443 , \2441 , \2442 );
and \U$2101 ( \2444 , \2436 , \2443 );
not \U$2102 ( \2445 , \2436 );
not \U$2103 ( \2446 , \2443 );
and \U$2104 ( \2447 , \2445 , \2446 );
nor \U$2105 ( \2448 , \2444 , \2447 );
and \U$2106 ( \2449 , \2406 , \1018 );
and \U$2107 ( \2450 , \894 , \1758 );
and \U$2108 ( \2451 , \895 , \1044 );
nor \U$2109 ( \2452 , \2450 , \2451 );
and \U$2110 ( \2453 , \2452 , \1067 );
nor \U$2111 ( \2454 , \2449 , \2453 );
xor \U$2112 ( \2455 , \2448 , \2454 );
xor \U$2113 ( \2456 , \2429 , \2455 );
and \U$2114 ( \2457 , \2383 , \2410 );
and \U$2115 ( \2458 , \2356 , \2382 );
nor \U$2116 ( \2459 , \2457 , \2458 );
not \U$2117 ( \2460 , \2459 );
and \U$2118 ( \2461 , \2456 , \2460 );
not \U$2119 ( \2462 , \2456 );
and \U$2120 ( \2463 , \2462 , \2459 );
nor \U$2121 ( \2464 , \2461 , \2463 );
not \U$2122 ( \2465 , \2378 );
not \U$2123 ( \2466 , \2371 );
or \U$2124 ( \2467 , \2465 , \2466 );
or \U$2125 ( \2468 , \2370 , \2358 );
nand \U$2126 ( \2469 , \2467 , \2468 );
or \U$2127 ( \2470 , \2323 , \1809 );
not \U$2128 ( \2471 , \1199 );
not \U$2129 ( \2472 , \848 );
or \U$2130 ( \2473 , \2471 , \2472 );
nand \U$2131 ( \2474 , \847 , \1200 );
nand \U$2132 ( \2475 , \2473 , \2474 );
or \U$2133 ( \2476 , \2475 , \1719 );
nand \U$2134 ( \2477 , \2470 , \2476 );
or \U$2135 ( \2478 , \2365 , \1293 );
not \U$2136 ( \2479 , RI9871b18_134);
or \U$2137 ( \2480 , \1543 , \2479 );
nand \U$2138 ( \2481 , \2478 , \2480 );
and \U$2139 ( \2482 , \2477 , \2481 );
not \U$2140 ( \2483 , \2477 );
not \U$2141 ( \2484 , \2481 );
and \U$2142 ( \2485 , \2483 , \2484 );
nor \U$2143 ( \2486 , \2482 , \2485 );
not \U$2144 ( \2487 , \2486 );
and \U$2145 ( \2488 , \2469 , \2487 );
not \U$2146 ( \2489 , \2469 );
and \U$2147 ( \2490 , \2489 , \2486 );
nor \U$2148 ( \2491 , \2488 , \2490 );
buf \U$2149 ( \2492 , \1446 );
and \U$2150 ( \2493 , \2492 , \1347 );
and \U$2151 ( \2494 , \1649 , RI9871d70_139);
nor \U$2152 ( \2495 , \2493 , \2494 );
and \U$2153 ( \2496 , \2495 , \832 );
and \U$2154 ( \2497 , \2316 , \859 );
nor \U$2155 ( \2498 , \2496 , \2497 );
xor \U$2156 ( \2499 , \2498 , \2285 );
not \U$2157 ( \2500 , \1501 );
not \U$2158 ( \2501 , \2401 );
or \U$2159 ( \2502 , \2500 , \2501 );
and \U$2160 ( \2503 , RI9871c80_137, \1672 );
not \U$2161 ( \2504 , RI9871c80_137);
and \U$2162 ( \2505 , \2504 , \1394 );
nor \U$2163 ( \2506 , \2503 , \2505 );
or \U$2164 ( \2507 , \2506 , \1746 );
nand \U$2165 ( \2508 , \2502 , \2507 );
xor \U$2166 ( \2509 , \2499 , \2508 );
xor \U$2167 ( \2510 , \2491 , \2509 );
not \U$2168 ( \2511 , \2344 );
not \U$2169 ( \2512 , \2340 );
or \U$2170 ( \2513 , \2511 , \2512 );
or \U$2171 ( \2514 , \2335 , \2228 );
nand \U$2172 ( \2515 , \2513 , \2514 );
xor \U$2173 ( \2516 , \2510 , \2515 );
xor \U$2174 ( \2517 , \2464 , \2516 );
xor \U$2175 ( \2518 , \2420 , \2517 );
or \U$2176 ( \2519 , \2350 , \2412 );
or \U$2177 ( \2520 , \2353 , \2411 );
nand \U$2178 ( \2521 , \2519 , \2520 );
xor \U$2179 ( \2522 , \2518 , \2521 );
xor \U$2180 ( \2523 , \2307 , \2346 );
and \U$2181 ( \2524 , \2523 , \2413 );
and \U$2182 ( \2525 , \2307 , \2346 );
nor \U$2183 ( \2526 , \2524 , \2525 );
nor \U$2184 ( \2527 , \2522 , \2526 );
not \U$2185 ( \2528 , \2527 );
nand \U$2186 ( \2529 , \2416 , \2528 );
and \U$2187 ( \2530 , \2301 , \2209 );
not \U$2188 ( \2531 , \2301 );
and \U$2189 ( \2532 , \2531 , \2210 );
or \U$2190 ( \2533 , \2530 , \2532 );
not \U$2191 ( \2534 , \1922 );
not \U$2192 ( \2535 , \2010 );
or \U$2193 ( \2536 , \2534 , \2535 );
not \U$2194 ( \2537 , \1796 );
nand \U$2195 ( \2538 , \2537 , \2011 );
nand \U$2196 ( \2539 , \2536 , \2538 );
nor \U$2197 ( \2540 , \2533 , \2539 );
nor \U$2198 ( \2541 , \2529 , \2540 );
and \U$2199 ( \2542 , \2174 , \2541 );
xor \U$2200 ( \2543 , \2420 , \2517 );
and \U$2201 ( \2544 , \2543 , \2521 );
and \U$2202 ( \2545 , \2420 , \2517 );
nor \U$2203 ( \2546 , \2544 , \2545 );
xor \U$2204 ( \2547 , \2424 , \2428 );
and \U$2205 ( \2548 , \2547 , \2455 );
and \U$2206 ( \2549 , \2424 , \2428 );
nor \U$2207 ( \2550 , \2548 , \2549 );
or \U$2208 ( \2551 , \2448 , \2454 );
or \U$2209 ( \2552 , \2436 , \2446 );
nand \U$2210 ( \2553 , \2551 , \2552 );
not \U$2211 ( \2554 , \2506 );
not \U$2212 ( \2555 , \1591 );
and \U$2213 ( \2556 , \2554 , \2555 );
and \U$2214 ( \2557 , \1693 , \1584 );
and \U$2215 ( \2558 , \1692 , RI9871c80_137);
nor \U$2216 ( \2559 , \2557 , \2558 );
and \U$2217 ( \2560 , \2559 , \1518 );
nor \U$2218 ( \2561 , \2556 , \2560 );
and \U$2219 ( \2562 , \1293 , \1543 );
nor \U$2220 ( \2563 , \2562 , \2479 );
xnor \U$2221 ( \2564 , \2561 , \2563 );
and \U$2222 ( \2565 , RI9871d70_139, \1418 );
not \U$2223 ( \2566 , RI9871d70_139);
and \U$2224 ( \2567 , \2566 , \1417 );
nor \U$2225 ( \2568 , \2565 , \2567 );
not \U$2226 ( \2569 , \2568 );
not \U$2227 ( \2570 , \932 );
and \U$2228 ( \2571 , \2569 , \2570 );
and \U$2229 ( \2572 , \2495 , \859 );
nor \U$2230 ( \2573 , \2571 , \2572 );
xor \U$2231 ( \2574 , \2564 , \2573 );
xor \U$2232 ( \2575 , \2553 , \2574 );
not \U$2233 ( \2576 , \2508 );
not \U$2234 ( \2577 , \2499 );
or \U$2235 ( \2578 , \2576 , \2577 );
or \U$2236 ( \2579 , \2498 , \2285 );
nand \U$2237 ( \2580 , \2578 , \2579 );
xor \U$2238 ( \2581 , \2575 , \2580 );
and \U$2239 ( \2582 , \2550 , \2581 );
not \U$2240 ( \2583 , \2550 );
not \U$2241 ( \2584 , \2581 );
and \U$2242 ( \2585 , \2583 , \2584 );
nor \U$2243 ( \2586 , \2582 , \2585 );
and \U$2244 ( \2587 , \2510 , \2515 );
and \U$2245 ( \2588 , \2491 , \2509 );
nor \U$2246 ( \2589 , \2587 , \2588 );
xnor \U$2247 ( \2590 , \2586 , \2589 );
and \U$2248 ( \2591 , \1367 , \1311 );
not \U$2249 ( \2592 , \1367 );
and \U$2250 ( \2593 , \2592 , \1320 );
nor \U$2251 ( \2594 , \2591 , \2593 );
not \U$2252 ( \2595 , \1353 );
or \U$2253 ( \2596 , \2594 , \2595 );
or \U$2254 ( \2597 , \2440 , \1558 );
nand \U$2255 ( \2598 , \2596 , \2597 );
not \U$2256 ( \2599 , \2322 );
and \U$2257 ( \2600 , \2598 , \2599 );
not \U$2258 ( \2601 , \2598 );
and \U$2259 ( \2602 , \2601 , \2322 );
nor \U$2260 ( \2603 , \2600 , \2602 );
not \U$2261 ( \2604 , \2603 );
not \U$2262 ( \2605 , \2399 );
and \U$2263 ( \2606 , RI9872130_147, \2605 );
not \U$2264 ( \2607 , RI9872130_147);
and \U$2265 ( \2608 , \2607 , \1128 );
nor \U$2266 ( \2609 , \2606 , \2608 );
and \U$2267 ( \2610 , \2609 , \924 );
and \U$2268 ( \2611 , \2433 , \876 );
nor \U$2269 ( \2612 , \2610 , \2611 );
not \U$2270 ( \2613 , \2612 );
and \U$2271 ( \2614 , \2604 , \2613 );
and \U$2272 ( \2615 , \2603 , \2612 );
nor \U$2273 ( \2616 , \2614 , \2615 );
xor \U$2274 ( \2617 , \1165 , \821 );
not \U$2275 ( \2618 , \2617 );
not \U$2276 ( \2619 , \1220 );
or \U$2277 ( \2620 , \2618 , \2619 );
or \U$2278 ( \2621 , \2475 , \1809 );
nand \U$2279 ( \2622 , \2620 , \2621 );
not \U$2280 ( \2623 , \2622 );
and \U$2281 ( \2624 , \2623 , \2481 );
and \U$2282 ( \2625 , \2622 , \2484 );
nor \U$2283 ( \2626 , \2624 , \2625 );
and \U$2284 ( \2627 , \2452 , \1018 );
and \U$2285 ( \2628 , \916 , \1045 );
and \U$2286 ( \2629 , \1513 , \1044 );
nor \U$2287 ( \2630 , \2628 , \2629 );
and \U$2288 ( \2631 , \2630 , \1067 );
nor \U$2289 ( \2632 , \2627 , \2631 );
xnor \U$2290 ( \2633 , \2626 , \2632 );
xor \U$2291 ( \2634 , \2616 , \2633 );
and \U$2292 ( \2635 , \2469 , \2487 );
and \U$2293 ( \2636 , \2477 , \2484 );
nor \U$2294 ( \2637 , \2635 , \2636 );
xor \U$2295 ( \2638 , \2634 , \2637 );
xor \U$2296 ( \2639 , \2590 , \2638 );
and \U$2297 ( \2640 , \2464 , \2516 );
and \U$2298 ( \2641 , \2456 , \2460 );
nor \U$2299 ( \2642 , \2640 , \2641 );
xor \U$2300 ( \2643 , \2639 , \2642 );
nand \U$2301 ( \2644 , \2546 , \2643 );
xor \U$2302 ( \2645 , \2590 , \2638 );
and \U$2303 ( \2646 , \2645 , \2642 );
and \U$2304 ( \2647 , \2590 , \2638 );
nor \U$2305 ( \2648 , \2646 , \2647 );
xor \U$2306 ( \2649 , \2616 , \2633 );
and \U$2307 ( \2650 , \2649 , \2637 );
and \U$2308 ( \2651 , \2616 , \2633 );
nor \U$2309 ( \2652 , \2650 , \2651 );
not \U$2310 ( \2653 , \2599 );
not \U$2311 ( \2654 , \2598 );
or \U$2312 ( \2655 , \2653 , \2654 );
not \U$2313 ( \2656 , \2612 );
nand \U$2314 ( \2657 , \2656 , \2603 );
nand \U$2315 ( \2658 , \2655 , \2657 );
and \U$2316 ( \2659 , \2559 , \1501 );
and \U$2317 ( \2660 , \1518 , RI9871c80_137);
nor \U$2318 ( \2661 , \2659 , \2660 );
and \U$2319 ( \2662 , \2658 , \2661 );
not \U$2320 ( \2663 , \2658 );
not \U$2321 ( \2664 , \2661 );
and \U$2322 ( \2665 , \2663 , \2664 );
nor \U$2323 ( \2666 , \2662 , \2665 );
or \U$2324 ( \2667 , \2564 , \2573 );
or \U$2325 ( \2668 , \2561 , \2563 );
nand \U$2326 ( \2669 , \2667 , \2668 );
xor \U$2327 ( \2670 , \2666 , \2669 );
xor \U$2328 ( \2671 , \2553 , \2574 );
and \U$2329 ( \2672 , \2671 , \2580 );
and \U$2330 ( \2673 , \2553 , \2574 );
or \U$2331 ( \2674 , \2672 , \2673 );
xor \U$2332 ( \2675 , \2670 , \2674 );
not \U$2333 ( \2676 , \2594 );
not \U$2334 ( \2677 , \1558 );
and \U$2335 ( \2678 , \2676 , \2677 );
and \U$2336 ( \2679 , \1447 , \1367 );
not \U$2337 ( \2680 , \2492 );
and \U$2338 ( \2681 , \2680 , RI9871e60_141);
nor \U$2339 ( \2682 , \2679 , \2681 );
and \U$2340 ( \2683 , \2682 , \1353 );
nor \U$2341 ( \2684 , \2678 , \2683 );
and \U$2342 ( \2685 , \2630 , \1018 );
and \U$2343 ( \2686 , \1834 , \1045 );
and \U$2344 ( \2687 , \1275 , \1044 );
nor \U$2345 ( \2688 , \2686 , \2687 );
and \U$2346 ( \2689 , \2688 , \1067 );
nor \U$2347 ( \2690 , \2685 , \2689 );
xnor \U$2348 ( \2691 , \2684 , \2690 );
xnor \U$2349 ( \2692 , \1672 , RI9872130_147);
and \U$2350 ( \2693 , \2692 , \924 );
and \U$2351 ( \2694 , \2609 , \876 );
nor \U$2352 ( \2695 , \2693 , \2694 );
xor \U$2353 ( \2696 , \2691 , \2695 );
or \U$2354 ( \2697 , \2626 , \2632 );
or \U$2355 ( \2698 , \2623 , \2484 );
nand \U$2356 ( \2699 , \2697 , \2698 );
xor \U$2357 ( \2700 , \2696 , \2699 );
and \U$2358 ( \2701 , \1098 , RI9871d70_139);
and \U$2359 ( \2702 , \1106 , \1347 );
nor \U$2360 ( \2703 , \2701 , \2702 );
or \U$2361 ( \2704 , \2703 , \932 );
or \U$2362 ( \2705 , \2568 , \860 );
nand \U$2363 ( \2706 , \2704 , \2705 );
not \U$2364 ( \2707 , \2474 );
xor \U$2365 ( \2708 , \2706 , \2707 );
and \U$2366 ( \2709 , \2617 , \1162 );
and \U$2367 ( \2710 , \894 , \1166 );
and \U$2368 ( \2711 , \895 , \1165 );
nor \U$2369 ( \2712 , \2710 , \2711 );
and \U$2370 ( \2713 , \2712 , \1220 );
nor \U$2371 ( \2714 , \2709 , \2713 );
not \U$2372 ( \2715 , \2714 );
and \U$2373 ( \2716 , \2708 , \2715 );
not \U$2374 ( \2717 , \2708 );
and \U$2375 ( \2718 , \2717 , \2714 );
nor \U$2376 ( \2719 , \2716 , \2718 );
xor \U$2377 ( \2720 , \2700 , \2719 );
xor \U$2378 ( \2721 , \2675 , \2720 );
xor \U$2379 ( \2722 , \2652 , \2721 );
or \U$2380 ( \2723 , \2586 , \2589 );
or \U$2381 ( \2724 , \2550 , \2584 );
nand \U$2382 ( \2725 , \2723 , \2724 );
xor \U$2383 ( \2726 , \2722 , \2725 );
or \U$2384 ( \2727 , \2648 , \2726 );
and \U$2385 ( \2728 , \2644 , \2727 );
xor \U$2386 ( \2729 , \2652 , \2721 );
and \U$2387 ( \2730 , \2729 , \2725 );
and \U$2388 ( \2731 , \2652 , \2721 );
nor \U$2389 ( \2732 , \2730 , \2731 );
and \U$2390 ( \2733 , \2675 , \2720 );
and \U$2391 ( \2734 , \2670 , \2674 );
nor \U$2392 ( \2735 , \2733 , \2734 );
and \U$2393 ( \2736 , \2708 , \2715 );
and \U$2394 ( \2737 , \2706 , \2707 );
nor \U$2395 ( \2738 , \2736 , \2737 );
and \U$2396 ( \2739 , \2692 , \876 );
xnor \U$2397 ( \2740 , \1693 , RI9872130_147);
and \U$2398 ( \2741 , \2740 , \924 );
nor \U$2399 ( \2742 , \2739 , \2741 );
and \U$2400 ( \2743 , \1591 , \1746 );
nor \U$2401 ( \2744 , \2743 , \1584 );
xor \U$2402 ( \2745 , \2742 , \2744 );
xnor \U$2403 ( \2746 , \1418 , RI9871e60_141);
and \U$2404 ( \2747 , \2746 , \1353 );
and \U$2405 ( \2748 , \2682 , \1382 );
nor \U$2406 ( \2749 , \2747 , \2748 );
xor \U$2407 ( \2750 , \2745 , \2749 );
xor \U$2408 ( \2751 , \2738 , \2750 );
and \U$2409 ( \2752 , \2712 , \1162 );
or \U$2410 ( \2753 , \1513 , \1166 );
or \U$2411 ( \2754 , \916 , \1165 );
nand \U$2412 ( \2755 , \2753 , \2754 );
and \U$2413 ( \2756 , \2755 , \1220 );
nor \U$2414 ( \2757 , \2752 , \2756 );
not \U$2415 ( \2758 , \2703 );
not \U$2416 ( \2759 , \860 );
and \U$2417 ( \2760 , \2758 , \2759 );
xnor \U$2418 ( \2761 , \2399 , RI9871d70_139);
and \U$2419 ( \2762 , \2761 , \832 );
nor \U$2420 ( \2763 , \2760 , \2762 );
xor \U$2421 ( \2764 , \2757 , \2763 );
and \U$2422 ( \2765 , \1758 , \1311 );
not \U$2423 ( \2766 , \1758 );
and \U$2424 ( \2767 , \2766 , \1320 );
nor \U$2425 ( \2768 , \2765 , \2767 );
not \U$2426 ( \2769 , \2768 );
not \U$2427 ( \2770 , \1068 );
and \U$2428 ( \2771 , \2769 , \2770 );
and \U$2429 ( \2772 , \2688 , \1018 );
nor \U$2430 ( \2773 , \2771 , \2772 );
xor \U$2431 ( \2774 , \2764 , \2773 );
xor \U$2432 ( \2775 , \2751 , \2774 );
xor \U$2433 ( \2776 , \2735 , \2775 );
and \U$2434 ( \2777 , \2666 , \2669 );
and \U$2435 ( \2778 , \2658 , \2661 );
nor \U$2436 ( \2779 , \2777 , \2778 );
or \U$2437 ( \2780 , \2691 , \2695 );
or \U$2438 ( \2781 , \2684 , \2690 );
nand \U$2439 ( \2782 , \2780 , \2781 );
and \U$2440 ( \2783 , \1165 , \821 );
and \U$2441 ( \2784 , \2783 , \2664 );
not \U$2442 ( \2785 , \2783 );
and \U$2443 ( \2786 , \2785 , \2661 );
nor \U$2444 ( \2787 , \2784 , \2786 );
xnor \U$2445 ( \2788 , \2782 , \2787 );
xor \U$2446 ( \2789 , \2779 , \2788 );
and \U$2447 ( \2790 , \2700 , \2719 );
and \U$2448 ( \2791 , \2699 , \2696 );
nor \U$2449 ( \2792 , \2790 , \2791 );
xor \U$2450 ( \2793 , \2789 , \2792 );
xor \U$2451 ( \2794 , \2776 , \2793 );
nand \U$2452 ( \2795 , \2732 , \2794 );
and \U$2453 ( \2796 , \2542 , \2728 , \2795 );
not \U$2454 ( \2797 , \2796 );
and \U$2455 ( \2798 , \2147 , \2149 );
not \U$2456 ( \2799 , \2147 );
and \U$2457 ( \2800 , \2799 , \2150 );
or \U$2458 ( \2801 , \2798 , \2800 );
not \U$2459 ( \2802 , \2801 );
not \U$2460 ( \2803 , \2802 );
not \U$2461 ( \2804 , \1767 );
not \U$2462 ( \2805 , \1773 );
or \U$2463 ( \2806 , \2804 , \2805 );
or \U$2464 ( \2807 , \1773 , \1767 );
nand \U$2465 ( \2808 , \2806 , \2807 );
not \U$2466 ( \2809 , \2808 );
xor \U$2467 ( \2810 , \1387 , \1531 );
and \U$2468 ( \2811 , \1473 , \924 );
xnor \U$2469 ( \2812 , \1550 , RI9872130_147);
not \U$2470 ( \2813 , \2812 );
and \U$2471 ( \2814 , \2813 , \876 );
nor \U$2472 ( \2815 , \2811 , \2814 );
xor \U$2473 ( \2816 , \2089 , \2815 );
not \U$2474 ( \2817 , \1518 );
not \U$2475 ( \2818 , \1508 );
or \U$2476 ( \2819 , \2817 , \2818 );
and \U$2477 ( \2820 , RI9871c80_137, \821 );
not \U$2478 ( \2821 , RI9871c80_137);
and \U$2479 ( \2822 , \2821 , \824 );
nor \U$2480 ( \2823 , \2820 , \2822 );
nand \U$2481 ( \2824 , \2823 , \1501 );
nand \U$2482 ( \2825 , \2819 , \2824 );
not \U$2483 ( \2826 , \2825 );
and \U$2484 ( \2827 , \2816 , \2826 );
and \U$2485 ( \2828 , \2089 , \2815 );
or \U$2486 ( \2829 , \2827 , \2828 );
not \U$2487 ( \2830 , \2829 );
not \U$2488 ( \2831 , \2830 );
not \U$2489 ( \2832 , \1292 );
and \U$2490 ( \2833 , \918 , \2479 );
not \U$2491 ( \2834 , \918 );
and \U$2492 ( \2835 , \2834 , RI9871b18_134);
nor \U$2493 ( \2836 , \2833 , \2835 );
not \U$2494 ( \2837 , \2836 );
or \U$2495 ( \2838 , \2832 , \2837 );
nand \U$2496 ( \2839 , \1280 , \1323 );
nand \U$2497 ( \2840 , \2838 , \2839 );
not \U$2498 ( \2841 , \2840 );
not \U$2499 ( \2842 , \1062 );
and \U$2500 ( \2843 , RI9871e60_141, \2842 );
not \U$2501 ( \2844 , RI9871e60_141);
and \U$2502 ( \2845 , \2844 , \1062 );
nor \U$2503 ( \2846 , \2843 , \2845 );
not \U$2504 ( \2847 , \2846 );
not \U$2505 ( \2848 , \1558 );
and \U$2506 ( \2849 , \2847 , \2848 );
and \U$2507 ( \2850 , \1373 , \1353 );
nor \U$2508 ( \2851 , \2849 , \2850 );
not \U$2509 ( \2852 , \2851 );
and \U$2510 ( \2853 , \2841 , \2852 );
and \U$2511 ( \2854 , \2840 , \2851 );
nor \U$2512 ( \2855 , \2853 , \2854 );
and \U$2513 ( \2856 , \1212 , \1044 );
not \U$2514 ( \2857 , \1212 );
and \U$2515 ( \2858 , \2857 , \1045 );
nor \U$2516 ( \2859 , \2856 , \2858 );
and \U$2517 ( \2860 , \2859 , \1018 );
and \U$2518 ( \2861 , \1049 , \1067 );
nor \U$2519 ( \2862 , \2860 , \2861 );
or \U$2520 ( \2863 , \2855 , \2862 );
not \U$2521 ( \2864 , \2840 );
or \U$2522 ( \2865 , \2864 , \2851 );
nand \U$2523 ( \2866 , \2863 , \2865 );
not \U$2524 ( \2867 , \2866 );
not \U$2525 ( \2868 , \1475 );
not \U$2526 ( \2869 , \1521 );
or \U$2527 ( \2870 , \2868 , \2869 );
or \U$2528 ( \2871 , \1521 , \1475 );
nand \U$2529 ( \2872 , \2870 , \2871 );
not \U$2530 ( \2873 , \2872 );
not \U$2531 ( \2874 , \2873 );
or \U$2532 ( \2875 , \2867 , \2874 );
not \U$2533 ( \2876 , \2866 );
nand \U$2534 ( \2877 , \2876 , \2872 );
nand \U$2535 ( \2878 , \2875 , \2877 );
not \U$2536 ( \2879 , \2878 );
or \U$2537 ( \2880 , \2831 , \2879 );
nand \U$2538 ( \2881 , \2872 , \2866 );
nand \U$2539 ( \2882 , \2880 , \2881 );
xor \U$2540 ( \2883 , \2810 , \2882 );
not \U$2541 ( \2884 , \2883 );
or \U$2542 ( \2885 , \2809 , \2884 );
nand \U$2543 ( \2886 , \2810 , \2882 );
nand \U$2544 ( \2887 , \2885 , \2886 );
not \U$2545 ( \2888 , \2887 );
not \U$2546 ( \2889 , \2888 );
and \U$2547 ( \2890 , \2803 , \2889 );
xnor \U$2548 ( \2891 , \2801 , \2888 );
not \U$2549 ( \2892 , \2808 );
and \U$2550 ( \2893 , \2883 , \2892 );
not \U$2551 ( \2894 , \2883 );
and \U$2552 ( \2895 , \2894 , \2808 );
nor \U$2553 ( \2896 , \2893 , \2895 );
not \U$2554 ( \2897 , \2896 );
not \U$2555 ( \2898 , \2897 );
not \U$2556 ( \2899 , \2136 );
not \U$2557 ( \2900 , \2028 );
and \U$2558 ( \2901 , \2899 , \2900 );
and \U$2559 ( \2902 , \2028 , \2136 );
nor \U$2560 ( \2903 , \2901 , \2902 );
not \U$2561 ( \2904 , \2903 );
xor \U$2562 ( \2905 , \2128 , \2061 );
not \U$2563 ( \2906 , \2905 );
not \U$2564 ( \2907 , \797 );
not \U$2565 ( \2908 , \2046 );
not \U$2566 ( \2909 , \2908 );
or \U$2567 ( \2910 , \2907 , \2909 );
xnor \U$2568 ( \2911 , \1097 , RI98719b0_131);
nand \U$2569 ( \2912 , \2911 , \793 );
nand \U$2570 ( \2913 , \2910 , \2912 );
and \U$2571 ( \2914 , RI9871e60_141, \1047 );
not \U$2572 ( \2915 , RI9871e60_141);
and \U$2573 ( \2916 , \2915 , \1041 );
nor \U$2574 ( \2917 , \2914 , \2916 );
not \U$2575 ( \2918 , \2917 );
not \U$2576 ( \2919 , \1382 );
or \U$2577 ( \2920 , \2918 , \2919 );
or \U$2578 ( \2921 , \2846 , \1989 );
nand \U$2579 ( \2922 , \2920 , \2921 );
xor \U$2580 ( \2923 , \2913 , \2922 );
and \U$2581 ( \2924 , \1191 , \1044 );
not \U$2582 ( \2925 , \1191 );
and \U$2583 ( \2926 , \2925 , \1045 );
or \U$2584 ( \2927 , \2924 , \2926 );
and \U$2585 ( \2928 , \2927 , \1018 );
and \U$2586 ( \2929 , \2859 , \1067 );
nor \U$2587 ( \2930 , \2928 , \2929 );
not \U$2588 ( \2931 , \2930 );
and \U$2589 ( \2932 , \2923 , \2931 );
and \U$2590 ( \2933 , \2913 , \2922 );
or \U$2591 ( \2934 , \2932 , \2933 );
not \U$2592 ( \2935 , \2934 );
not \U$2593 ( \2936 , \386 );
not \U$2594 ( \2937 , \1177 );
or \U$2595 ( \2938 , \2936 , \2937 );
not \U$2596 ( \2939 , \437 );
nand \U$2597 ( \2940 , \2938 , \2939 );
nand \U$2598 ( \2941 , \387 , \440 );
and \U$2599 ( \2942 , \2940 , \2941 );
not \U$2600 ( \2943 , \2940 );
not \U$2601 ( \2944 , \2941 );
and \U$2602 ( \2945 , \2943 , \2944 );
nor \U$2603 ( \2946 , \2942 , \2945 );
buf \U$2604 ( \2947 , \2946 );
not \U$2605 ( \2948 , \2947 );
and \U$2606 ( \2949 , \1200 , \2948 );
not \U$2607 ( \2950 , \1323 );
not \U$2608 ( \2951 , \2836 );
or \U$2609 ( \2952 , \2950 , \2951 );
and \U$2610 ( \2953 , RI9871b18_134, \894 );
not \U$2611 ( \2954 , RI9871b18_134);
not \U$2612 ( \2955 , \1506 );
and \U$2613 ( \2956 , \2954 , \2955 );
nor \U$2614 ( \2957 , \2953 , \2956 );
not \U$2615 ( \2958 , \2957 );
nand \U$2616 ( \2959 , \2958 , \1292 );
nand \U$2617 ( \2960 , \2952 , \2959 );
xor \U$2618 ( \2961 , \2949 , \2960 );
not \U$2619 ( \2962 , \2111 );
and \U$2620 ( \2963 , \2962 , \1165 );
not \U$2621 ( \2964 , \2962 );
and \U$2622 ( \2965 , \2964 , \1199 );
nor \U$2623 ( \2966 , \2963 , \2965 );
or \U$2624 ( \2967 , \2966 , \1809 );
or \U$2625 ( \2968 , \1719 , \2120 );
nand \U$2626 ( \2969 , \2967 , \2968 );
and \U$2627 ( \2970 , \2961 , \2969 );
and \U$2628 ( \2971 , \2949 , \2960 );
nor \U$2629 ( \2972 , \2970 , \2971 );
not \U$2630 ( \2973 , \2972 );
nand \U$2631 ( \2974 , RI98726d0_159, RI9872748_160);
and \U$2632 ( \2975 , \2974 , RI9872310_151);
not \U$2633 ( \2976 , \2975 );
not \U$2634 ( \2977 , \2976 );
not \U$2635 ( \2978 , \2087 );
not \U$2636 ( \2979 , \2082 );
or \U$2637 ( \2980 , \2978 , \2979 );
not \U$2638 ( \2981 , \2076 );
buf \U$2639 ( \2982 , \1393 );
not \U$2640 ( \2983 , \2982 );
or \U$2641 ( \2984 , \2981 , \2983 );
or \U$2642 ( \2985 , \1394 , \2080 );
nand \U$2643 ( \2986 , \2984 , \2985 );
nand \U$2644 ( \2987 , \2986 , \2074 );
nand \U$2645 ( \2988 , \2980 , \2987 );
not \U$2646 ( \2989 , \2988 );
or \U$2647 ( \2990 , \2977 , \2989 );
not \U$2648 ( \2991 , \2988 );
not \U$2649 ( \2992 , \2975 );
and \U$2650 ( \2993 , \2991 , \2992 );
and \U$2651 ( \2994 , \2988 , \2975 );
nor \U$2652 ( \2995 , \2993 , \2994 );
not \U$2653 ( \2996 , \2995 );
or \U$2654 ( \2997 , \2090 , \1137 );
and \U$2655 ( \2998 , RI98718c0_129, \1799 );
not \U$2656 ( \2999 , RI98718c0_129);
and \U$2657 ( \3000 , \2999 , \2680 );
nor \U$2658 ( \3001 , \2998 , \3000 );
or \U$2659 ( \3002 , \3001 , \1688 );
nand \U$2660 ( \3003 , \2997 , \3002 );
nand \U$2661 ( \3004 , \2996 , \3003 );
nand \U$2662 ( \3005 , \2990 , \3004 );
not \U$2663 ( \3006 , \3005 );
or \U$2664 ( \3007 , \2973 , \3006 );
or \U$2665 ( \3008 , \2972 , \3005 );
nand \U$2666 ( \3009 , \3007 , \3008 );
not \U$2667 ( \3010 , \3009 );
or \U$2668 ( \3011 , \2935 , \3010 );
not \U$2669 ( \3012 , \2972 );
nand \U$2670 ( \3013 , \3012 , \3005 );
nand \U$2671 ( \3014 , \3011 , \3013 );
xor \U$2672 ( \3015 , \2089 , \2815 );
not \U$2673 ( \3016 , \2825 );
xor \U$2674 ( \3017 , \3015 , \3016 );
not \U$2675 ( \3018 , \3017 );
not \U$2676 ( \3019 , \3018 );
not \U$2677 ( \3020 , \2095 );
not \U$2678 ( \3021 , \2123 );
or \U$2679 ( \3022 , \3020 , \3021 );
or \U$2680 ( \3023 , \2123 , \2095 );
nand \U$2681 ( \3024 , \3022 , \3023 );
and \U$2682 ( \3025 , \2040 , \1431 );
and \U$2683 ( \3026 , RI9871c08_136, \1275 );
not \U$2684 ( \3027 , RI9871c08_136);
and \U$2685 ( \3028 , \3027 , \1838 );
nor \U$2686 ( \3029 , \3026 , \3028 );
and \U$2687 ( \3030 , \3029 , \1456 );
nor \U$2688 ( \3031 , \3025 , \3030 );
not \U$2689 ( \3032 , \3031 );
or \U$2690 ( \3033 , \2812 , \1470 );
and \U$2691 ( \3034 , \919 , \1659 );
not \U$2692 ( \3035 , \919 );
and \U$2693 ( \3036 , \3035 , \1253 );
nor \U$2694 ( \3037 , \3034 , \3036 );
or \U$2695 ( \3038 , \3037 , \1942 );
nand \U$2696 ( \3039 , \3033 , \3038 );
not \U$2697 ( \3040 , \3039 );
not \U$2698 ( \3041 , \3040 );
and \U$2699 ( \3042 , \3032 , \3041 );
not \U$2700 ( \3043 , \3039 );
not \U$2701 ( \3044 , \3031 );
or \U$2702 ( \3045 , \3043 , \3044 );
or \U$2703 ( \3046 , \3031 , \3039 );
nand \U$2704 ( \3047 , \3045 , \3046 );
not \U$2705 ( \3048 , \859 );
and \U$2706 ( \3049 , RI9871d70_139, \1605 );
not \U$2707 ( \3050 , RI9871d70_139);
and \U$2708 ( \3051 , \3050 , \1606 );
nor \U$2709 ( \3052 , \3049 , \3051 );
not \U$2710 ( \3053 , \3052 );
or \U$2711 ( \3054 , \3048 , \3053 );
or \U$2712 ( \3055 , \2053 , \932 );
nand \U$2713 ( \3056 , \3054 , \3055 );
and \U$2714 ( \3057 , \3047 , \3056 );
nor \U$2715 ( \3058 , \3042 , \3057 );
and \U$2716 ( \3059 , \3024 , \3058 );
not \U$2717 ( \3060 , \3024 );
not \U$2718 ( \3061 , \3058 );
and \U$2719 ( \3062 , \3060 , \3061 );
or \U$2720 ( \3063 , \3059 , \3062 );
not \U$2721 ( \3064 , \3063 );
or \U$2722 ( \3065 , \3019 , \3064 );
nand \U$2723 ( \3066 , \3024 , \3061 );
nand \U$2724 ( \3067 , \3065 , \3066 );
xor \U$2725 ( \3068 , \3014 , \3067 );
not \U$2726 ( \3069 , \3068 );
or \U$2727 ( \3070 , \2906 , \3069 );
nand \U$2728 ( \3071 , \3014 , \3067 );
nand \U$2729 ( \3072 , \3070 , \3071 );
not \U$2730 ( \3073 , \3072 );
or \U$2731 ( \3074 , \2904 , \3073 );
or \U$2732 ( \3075 , \3072 , \2903 );
nand \U$2733 ( \3076 , \3074 , \3075 );
not \U$2734 ( \3077 , \3076 );
or \U$2735 ( \3078 , \2898 , \3077 );
not \U$2736 ( \3079 , \2903 );
nand \U$2737 ( \3080 , \3079 , \3072 );
nand \U$2738 ( \3081 , \3078 , \3080 );
and \U$2739 ( \3082 , \2891 , \3081 );
nor \U$2740 ( \3083 , \2890 , \3082 );
and \U$2741 ( \3084 , \2168 , \2155 );
not \U$2742 ( \3085 , \2168 );
and \U$2743 ( \3086 , \3085 , \2156 );
nor \U$2744 ( \3087 , \3084 , \3086 );
nand \U$2745 ( \3088 , \3083 , \3087 );
not \U$2746 ( \3089 , \3088 );
xor \U$2747 ( \3090 , \2020 , \2023 );
xor \U$2748 ( \3091 , \3090 , \2025 );
not \U$2749 ( \3092 , \3091 );
xor \U$2750 ( \3093 , \2042 , \2051 );
xor \U$2751 ( \3094 , \3093 , \2058 );
not \U$2752 ( \3095 , \3094 );
not \U$2753 ( \3096 , \2862 );
and \U$2754 ( \3097 , \2855 , \3096 );
not \U$2755 ( \3098 , \2855 );
and \U$2756 ( \3099 , \3098 , \2862 );
nor \U$2757 ( \3100 , \3097 , \3099 );
not \U$2758 ( \3101 , \3100 );
or \U$2759 ( \3102 , \3095 , \3101 );
and \U$2760 ( \3103 , \3029 , \1431 );
and \U$2761 ( \3104 , RI9871c08_136, \1513 );
not \U$2762 ( \3105 , RI9871c08_136);
and \U$2763 ( \3106 , \3105 , \916 );
nor \U$2764 ( \3107 , \3104 , \3106 );
and \U$2765 ( \3108 , \3107 , \1456 );
nor \U$2766 ( \3109 , \3103 , \3108 );
not \U$2767 ( \3110 , \3109 );
not \U$2768 ( \3111 , \3110 );
and \U$2769 ( \3112 , \3052 , \832 );
and \U$2770 ( \3113 , RI9871d70_139, \1713 );
not \U$2771 ( \3114 , RI9871d70_139);
and \U$2772 ( \3115 , \3114 , \1714 );
nor \U$2773 ( \3116 , \3113 , \3115 );
and \U$2774 ( \3117 , \3116 , \859 );
nor \U$2775 ( \3118 , \3112 , \3117 );
not \U$2776 ( \3119 , \3118 );
not \U$2777 ( \3120 , \1353 );
not \U$2778 ( \3121 , \2917 );
or \U$2779 ( \3122 , \3120 , \3121 );
not \U$2780 ( \3123 , RI9871e60_141);
and \U$2781 ( \3124 , \3123 , \1212 );
not \U$2782 ( \3125 , \3123 );
not \U$2783 ( \3126 , \1209 );
not \U$2784 ( \3127 , \3126 );
not \U$2785 ( \3128 , \3127 );
not \U$2786 ( \3129 , \3128 );
buf \U$2787 ( \3130 , \3129 );
and \U$2788 ( \3131 , \3125 , \3130 );
nor \U$2789 ( \3132 , \3124 , \3131 );
or \U$2790 ( \3133 , \3132 , \1558 );
nand \U$2791 ( \3134 , \3122 , \3133 );
not \U$2792 ( \3135 , \3134 );
or \U$2793 ( \3136 , \3119 , \3135 );
or \U$2794 ( \3137 , \3134 , \3118 );
nand \U$2795 ( \3138 , \3136 , \3137 );
not \U$2796 ( \3139 , \3138 );
or \U$2797 ( \3140 , \3111 , \3139 );
not \U$2798 ( \3141 , \3118 );
nand \U$2799 ( \3142 , \3141 , \3134 );
nand \U$2800 ( \3143 , \3140 , \3142 );
not \U$2801 ( \3144 , \3143 );
and \U$2802 ( \3145 , \1800 , \847 );
not \U$2803 ( \3146 , \1800 );
and \U$2804 ( \3147 , \3146 , \848 );
nor \U$2805 ( \3148 , \3145 , \3147 );
not \U$2806 ( \3149 , \3148 );
not \U$2807 ( \3150 , \1591 );
and \U$2808 ( \3151 , \3149 , \3150 );
and \U$2809 ( \3152 , \2823 , \1518 );
nor \U$2810 ( \3153 , \3151 , \3152 );
not \U$2811 ( \3154 , RI9872310_151);
not \U$2812 ( \3155 , RI9872748_160);
and \U$2813 ( \3156 , \3154 , \3155 );
and \U$2814 ( \3157 , RI9872310_151, RI9872748_160);
and \U$2815 ( \3158 , RI98726d0_159, RI9872748_160);
not \U$2816 ( \3159 , RI98726d0_159);
and \U$2817 ( \3160 , \3159 , \3155 );
nor \U$2818 ( \3161 , \3158 , \3160 );
nor \U$2819 ( \3162 , \3156 , \3157 , \3161 );
buf \U$2820 ( \3163 , \3162 );
buf \U$2821 ( \3164 , \3163 );
not \U$2822 ( \3165 , \3164 );
xor \U$2823 ( \3166 , RI9872310_151, \1692 );
not \U$2824 ( \3167 , \3166 );
or \U$2825 ( \3168 , \3165 , \3167 );
buf \U$2826 ( \3169 , \3161 );
buf \U$2827 ( \3170 , \3169 );
nand \U$2828 ( \3171 , \3170 , RI9872310_151);
nand \U$2829 ( \3172 , \3168 , \3171 );
not \U$2830 ( \3173 , \3172 );
and \U$2831 ( \3174 , \3153 , \3173 );
not \U$2832 ( \3175 , \3153 );
and \U$2833 ( \3176 , \3175 , \3172 );
nor \U$2834 ( \3177 , \3174 , \3176 );
not \U$2835 ( \3178 , \3177 );
or \U$2836 ( \3179 , \3144 , \3178 );
not \U$2837 ( \3180 , \3153 );
nand \U$2838 ( \3181 , \3180 , \3172 );
nand \U$2839 ( \3182 , \3179 , \3181 );
nand \U$2840 ( \3183 , \3102 , \3182 );
or \U$2841 ( \3184 , \3100 , \3094 );
and \U$2842 ( \3185 , \3183 , \3184 );
not \U$2843 ( \3186 , \3185 );
xor \U$2844 ( \3187 , \2830 , \2878 );
not \U$2845 ( \3188 , \3187 );
or \U$2846 ( \3189 , \3186 , \3188 );
or \U$2847 ( \3190 , \3187 , \3185 );
nand \U$2848 ( \3191 , \3189 , \3190 );
not \U$2849 ( \3192 , \3191 );
or \U$2850 ( \3193 , \3092 , \3192 );
not \U$2851 ( \3194 , \3185 );
nand \U$2852 ( \3195 , \3194 , \3187 );
nand \U$2853 ( \3196 , \3193 , \3195 );
and \U$2854 ( \3197 , \3076 , \2897 );
not \U$2855 ( \3198 , \3076 );
and \U$2856 ( \3199 , \3198 , \2896 );
nor \U$2857 ( \3200 , \3197 , \3199 );
xor \U$2858 ( \3201 , \3196 , \3200 );
xor \U$2859 ( \3202 , \3185 , \3091 );
xnor \U$2860 ( \3203 , \3202 , \3187 );
not \U$2861 ( \3204 , \3203 );
xor \U$2862 ( \3205 , \3047 , \3056 );
not \U$2863 ( \3206 , \3205 );
xor \U$2864 ( \3207 , \2995 , \3003 );
not \U$2865 ( \3208 , \3207 );
xor \U$2866 ( \3209 , \2913 , \2922 );
not \U$2867 ( \3210 , \2930 );
xor \U$2868 ( \3211 , \3209 , \3210 );
not \U$2869 ( \3212 , \3211 );
or \U$2870 ( \3213 , \3208 , \3212 );
or \U$2871 ( \3214 , \3211 , \3207 );
nand \U$2872 ( \3215 , \3213 , \3214 );
not \U$2873 ( \3216 , \3215 );
or \U$2874 ( \3217 , \3206 , \3216 );
not \U$2875 ( \3218 , \3207 );
nand \U$2876 ( \3219 , \3218 , \3211 );
nand \U$2877 ( \3220 , \3217 , \3219 );
or \U$2878 ( \3221 , \3148 , \1746 );
and \U$2879 ( \3222 , \945 , RI9871c80_137);
and \U$2880 ( \3223 , \944 , \1800 );
nor \U$2881 ( \3224 , \3222 , \3223 );
or \U$2882 ( \3225 , \3224 , \1591 );
nand \U$2883 ( \3226 , \3221 , \3225 );
xor \U$2884 ( \3227 , RI986ef80_41, RI986eff8_42);
not \U$2885 ( \3228 , \3227 );
not \U$2886 ( \3229 , \385 );
not \U$2887 ( \3230 , \3229 );
not \U$2888 ( \3231 , \1177 );
or \U$2889 ( \3232 , \3230 , \3231 );
nand \U$2890 ( \3233 , \3232 , \434 );
not \U$2891 ( \3234 , \3233 );
not \U$2892 ( \3235 , \3234 );
or \U$2893 ( \3236 , \3228 , \3235 );
not \U$2894 ( \3237 , \3227 );
nand \U$2895 ( \3238 , \3233 , \3237 );
nand \U$2896 ( \3239 , \3236 , \3238 );
buf \U$2897 ( \3240 , \3239 );
and \U$2898 ( \3241 , \1200 , \3240 );
xor \U$2899 ( \3242 , \3226 , \3241 );
not \U$2900 ( \3243 , \2911 );
not \U$2901 ( \3244 , \797 );
or \U$2902 ( \3245 , \3243 , \3244 );
and \U$2903 ( \3246 , \1418 , RI98719b0_131);
and \U$2904 ( \3247 , \1417 , \1078 );
nor \U$2905 ( \3248 , \3246 , \3247 );
or \U$2906 ( \3249 , \3248 , \792 );
nand \U$2907 ( \3250 , \3245 , \3249 );
and \U$2908 ( \3251 , \3242 , \3250 );
and \U$2909 ( \3252 , \3226 , \3241 );
nor \U$2910 ( \3253 , \3251 , \3252 );
not \U$2911 ( \3254 , \3253 );
xor \U$2912 ( \3255 , \1200 , \2948 );
not \U$2913 ( \3256 , \3255 );
or \U$2914 ( \3257 , \3256 , \1809 );
or \U$2915 ( \3258 , \2966 , \1719 );
nand \U$2916 ( \3259 , \3257 , \3258 );
or \U$2917 ( \3260 , \2957 , \1543 );
and \U$2918 ( \3261 , RI9871b18_134, \824 );
not \U$2919 ( \3262 , RI9871b18_134);
and \U$2920 ( \3263 , \3262 , \821 );
nor \U$2921 ( \3264 , \3261 , \3263 );
or \U$2922 ( \3265 , \3264 , \1293 );
nand \U$2923 ( \3266 , \3260 , \3265 );
xor \U$2924 ( \3267 , \3259 , \3266 );
not \U$2925 ( \3268 , \1067 );
not \U$2926 ( \3269 , \2927 );
or \U$2927 ( \3270 , \3268 , \3269 );
buf \U$2928 ( \3271 , \1146 );
not \U$2929 ( \3272 , \3271 );
and \U$2930 ( \3273 , \3272 , \2116 );
not \U$2931 ( \3274 , \3272 );
not \U$2932 ( \3275 , \1485 );
and \U$2933 ( \3276 , \3274 , \3275 );
nor \U$2934 ( \3277 , \3273 , \3276 );
or \U$2935 ( \3278 , \3277 , \1612 );
nand \U$2936 ( \3279 , \3270 , \3278 );
and \U$2937 ( \3280 , \3267 , \3279 );
and \U$2938 ( \3281 , \3259 , \3266 );
nor \U$2939 ( \3282 , \3280 , \3281 );
nor \U$2940 ( \3283 , \3001 , \1137 );
and \U$2941 ( \3284 , RI98718c0_129, \2038 );
not \U$2942 ( \3285 , RI98718c0_129);
and \U$2943 ( \3286 , \3285 , \1311 );
nor \U$2944 ( \3287 , \3284 , \3286 );
nor \U$2945 ( \3288 , \3287 , \1688 );
or \U$2946 ( \3289 , \3283 , \3288 );
or \U$2947 ( \3290 , \3037 , \1470 );
and \U$2948 ( \3291 , \1344 , RI9872130_147);
not \U$2949 ( \3292 , \1344 );
and \U$2950 ( \3293 , \3292 , \919 );
nor \U$2951 ( \3294 , \3291 , \3293 );
or \U$2952 ( \3295 , \3294 , \1942 );
nand \U$2953 ( \3296 , \3290 , \3295 );
xnor \U$2954 ( \3297 , \3289 , \3296 );
not \U$2955 ( \3298 , \3297 );
and \U$2956 ( \3299 , \2986 , \2087 );
and \U$2957 ( \3300 , RI9871aa0_133, \1129 );
not \U$2958 ( \3301 , RI9871aa0_133);
and \U$2959 ( \3302 , \3301 , \2399 );
nor \U$2960 ( \3303 , \3300 , \3302 );
and \U$2961 ( \3304 , \3303 , \2074 );
nor \U$2962 ( \3305 , \3299 , \3304 );
not \U$2963 ( \3306 , \3305 );
and \U$2964 ( \3307 , \3298 , \3306 );
and \U$2965 ( \3308 , \3289 , \3296 );
nor \U$2966 ( \3309 , \3307 , \3308 );
and \U$2967 ( \3310 , \3282 , \3309 );
not \U$2968 ( \3311 , \3282 );
not \U$2969 ( \3312 , \3309 );
and \U$2970 ( \3313 , \3311 , \3312 );
nor \U$2971 ( \3314 , \3310 , \3313 );
nand \U$2972 ( \3315 , \3254 , \3314 );
not \U$2973 ( \3316 , \3282 );
nand \U$2974 ( \3317 , \3316 , \3312 );
nand \U$2975 ( \3318 , \3315 , \3317 );
xor \U$2976 ( \3319 , \3220 , \3318 );
xor \U$2977 ( \3320 , \3009 , \2934 );
and \U$2978 ( \3321 , \3319 , \3320 );
and \U$2979 ( \3322 , \3220 , \3318 );
nor \U$2980 ( \3323 , \3321 , \3322 );
not \U$2981 ( \3324 , \3323 );
xor \U$2982 ( \3325 , \3068 , \2905 );
not \U$2983 ( \3326 , \3325 );
and \U$2984 ( \3327 , \3324 , \3326 );
and \U$2985 ( \3328 , \3325 , \3323 );
nor \U$2986 ( \3329 , \3327 , \3328 );
not \U$2987 ( \3330 , \3329 );
not \U$2988 ( \3331 , \3330 );
or \U$2989 ( \3332 , \3204 , \3331 );
not \U$2990 ( \3333 , \3323 );
nand \U$2991 ( \3334 , \3333 , \3325 );
nand \U$2992 ( \3335 , \3332 , \3334 );
and \U$2993 ( \3336 , \3201 , \3335 );
and \U$2994 ( \3337 , \3196 , \3200 );
nor \U$2995 ( \3338 , \3336 , \3337 );
not \U$2996 ( \3339 , \2891 );
not \U$2997 ( \3340 , \3081 );
not \U$2998 ( \3341 , \3340 );
and \U$2999 ( \3342 , \3339 , \3341 );
and \U$3000 ( \3343 , \2891 , \3340 );
nor \U$3001 ( \3344 , \3342 , \3343 );
nand \U$3002 ( \3345 , \3338 , \3344 );
xor \U$3003 ( \3346 , \2949 , \2960 );
xor \U$3004 ( \3347 , \3346 , \2969 );
not \U$3005 ( \3348 , \3347 );
not \U$3006 ( \3349 , \3348 );
xor \U$3007 ( \3350 , \3143 , \3177 );
not \U$3008 ( \3351 , \3350 );
or \U$3009 ( \3352 , \3349 , \3351 );
or \U$3010 ( \3353 , \3350 , \3348 );
nand \U$3011 ( \3354 , \3352 , \3353 );
not \U$3012 ( \3355 , \3354 );
not \U$3013 ( \3356 , \3173 );
or \U$3014 ( \3357 , \3224 , \1746 );
and \U$3015 ( \3358 , \1257 , RI9871c80_137);
and \U$3016 ( \3359 , \1659 , \1584 );
nor \U$3017 ( \3360 , \3358 , \3359 );
or \U$3018 ( \3361 , \1591 , \3360 );
nand \U$3019 ( \3362 , \3357 , \3361 );
not \U$3020 ( \3363 , \3362 );
or \U$3021 ( \3364 , \3294 , \1470 );
not \U$3022 ( \3365 , \1366 );
and \U$3023 ( \3366 , \919 , \3365 );
not \U$3024 ( \3367 , \919 );
and \U$3025 ( \3368 , \3367 , \1606 );
nor \U$3026 ( \3369 , \3366 , \3368 );
not \U$3027 ( \3370 , \876 );
or \U$3028 ( \3371 , \3369 , \3370 );
nand \U$3029 ( \3372 , \3364 , \3371 );
not \U$3030 ( \3373 , \3372 );
not \U$3031 ( \3374 , \3287 );
nand \U$3032 ( \3375 , \3374 , \1136 );
and \U$3033 ( \3376 , \1275 , RI98718c0_129);
not \U$3034 ( \3377 , \1275 );
and \U$3035 ( \3378 , \3377 , \1111 );
nor \U$3036 ( \3379 , \3376 , \3378 );
nand \U$3037 ( \3380 , \3379 , \1083 );
and \U$3038 ( \3381 , \3375 , \3380 );
not \U$3039 ( \3382 , \3381 );
or \U$3040 ( \3383 , \3373 , \3382 );
or \U$3041 ( \3384 , \3381 , \3372 );
nand \U$3042 ( \3385 , \3383 , \3384 );
not \U$3043 ( \3386 , \3385 );
or \U$3044 ( \3387 , \3363 , \3386 );
not \U$3045 ( \3388 , \3381 );
nand \U$3046 ( \3389 , \3388 , \3372 );
nand \U$3047 ( \3390 , \3387 , \3389 );
not \U$3048 ( \3391 , \3390 );
or \U$3049 ( \3392 , \3356 , \3391 );
not \U$3050 ( \3393 , \1382 );
not \U$3051 ( \3394 , \1189 );
not \U$3052 ( \3395 , \3394 );
not \U$3053 ( \3396 , \3395 );
xnor \U$3054 ( \3397 , \3396 , RI9871e60_141);
not \U$3055 ( \3398 , \3397 );
or \U$3056 ( \3399 , \3393 , \3398 );
not \U$3057 ( \3400 , \3132 );
nand \U$3058 ( \3401 , \3400 , \1353 );
nand \U$3059 ( \3402 , \3399 , \3401 );
not \U$3060 ( \3403 , \832 );
not \U$3061 ( \3404 , \3116 );
or \U$3062 ( \3405 , \3403 , \3404 );
not \U$3063 ( \3406 , \1047 );
xor \U$3064 ( \3407 , RI9871d70_139, \3406 );
or \U$3065 ( \3408 , \3407 , \860 );
nand \U$3066 ( \3409 , \3405 , \3408 );
and \U$3067 ( \3410 , \3402 , \3409 );
not \U$3068 ( \3411 , \3402 );
not \U$3069 ( \3412 , \3409 );
and \U$3070 ( \3413 , \3411 , \3412 );
nor \U$3071 ( \3414 , \3410 , \3413 );
and \U$3072 ( \3415 , \3303 , \2087 );
xor \U$3073 ( \3416 , \1106 , RI9871aa0_133);
and \U$3074 ( \3417 , \3416 , \2074 );
nor \U$3075 ( \3418 , \3415 , \3417 );
not \U$3076 ( \3419 , \3418 );
and \U$3077 ( \3420 , \3414 , \3419 );
and \U$3078 ( \3421 , \3402 , \3409 );
nor \U$3079 ( \3422 , \3420 , \3421 );
not \U$3080 ( \3423 , \3422 );
not \U$3081 ( \3424 , \3390 );
not \U$3082 ( \3425 , \3172 );
and \U$3083 ( \3426 , \3424 , \3425 );
and \U$3084 ( \3427 , \3390 , \3172 );
nor \U$3085 ( \3428 , \3426 , \3427 );
not \U$3086 ( \3429 , \3428 );
nand \U$3087 ( \3430 , \3423 , \3429 );
nand \U$3088 ( \3431 , \3392 , \3430 );
not \U$3089 ( \3432 , \3431 );
or \U$3090 ( \3433 , \3355 , \3432 );
not \U$3091 ( \3434 , \3348 );
nand \U$3092 ( \3435 , \3434 , \3350 );
nand \U$3093 ( \3436 , \3433 , \3435 );
not \U$3094 ( \3437 , \3436 );
xnor \U$3095 ( \3438 , \3063 , \3018 );
not \U$3096 ( \3439 , \3438 );
xor \U$3097 ( \3440 , \3100 , \3094 );
xor \U$3098 ( \3441 , \3440 , \3182 );
not \U$3099 ( \3442 , \3441 );
or \U$3100 ( \3443 , \3439 , \3442 );
or \U$3101 ( \3444 , \3441 , \3438 );
nand \U$3102 ( \3445 , \3443 , \3444 );
not \U$3103 ( \3446 , \3445 );
or \U$3104 ( \3447 , \3437 , \3446 );
not \U$3105 ( \3448 , \3438 );
nand \U$3106 ( \3449 , \3448 , \3441 );
nand \U$3107 ( \3450 , \3447 , \3449 );
xor \U$3108 ( \3451 , \3450 , \3203 );
xnor \U$3109 ( \3452 , \3451 , \3329 );
not \U$3110 ( \3453 , \3452 );
not \U$3111 ( \3454 , RI98725e0_157);
not \U$3112 ( \3455 , RI9872658_158);
nand \U$3113 ( \3456 , \3454 , \3455 );
nand \U$3114 ( \3457 , RI98725e0_157, RI9872658_158);
and \U$3115 ( \3458 , \3456 , \3457 );
not \U$3116 ( \3459 , \3458 );
and \U$3117 ( \3460 , RI98726d0_159, RI9872658_158);
not \U$3118 ( \3461 , RI98726d0_159);
and \U$3119 ( \3462 , \3461 , \3455 );
nor \U$3120 ( \3463 , \3460 , \3462 );
and \U$3121 ( \3464 , \3459 , \3463 );
buf \U$3122 ( \3465 , \3464 );
buf \U$3123 ( \3466 , \3465 );
buf \U$3124 ( \3467 , \3458 );
or \U$3125 ( \3468 , \3466 , \3467 );
nand \U$3126 ( \3469 , \3468 , RI98726d0_159);
not \U$3127 ( \3470 , \3164 );
xor \U$3128 ( \3471 , RI9872310_151, \1394 );
not \U$3129 ( \3472 , \3471 );
or \U$3130 ( \3473 , \3470 , \3472 );
nand \U$3131 ( \3474 , \3166 , \3170 );
nand \U$3132 ( \3475 , \3473 , \3474 );
xor \U$3133 ( \3476 , \3469 , \3475 );
not \U$3134 ( \3477 , \794 );
xnor \U$3135 ( \3478 , \1799 , RI98719b0_131);
not \U$3136 ( \3479 , \3478 );
or \U$3137 ( \3480 , \3477 , \3479 );
or \U$3138 ( \3481 , \3248 , \3244 );
nand \U$3139 ( \3482 , \3480 , \3481 );
xor \U$3140 ( \3483 , \3476 , \3482 );
not \U$3141 ( \3484 , \1431 );
not \U$3142 ( \3485 , \3107 );
or \U$3143 ( \3486 , \3484 , \3485 );
not \U$3144 ( \3487 , RI9871c08_136);
and \U$3145 ( \3488 , \894 , \3487 );
not \U$3146 ( \3489 , \894 );
and \U$3147 ( \3490 , \3489 , RI9871c08_136);
nor \U$3148 ( \3491 , \3488 , \3490 );
nand \U$3149 ( \3492 , \3491 , \1456 );
nand \U$3150 ( \3493 , \3486 , \3492 );
not \U$3151 ( \3494 , \1162 );
xor \U$3152 ( \3495 , \1200 , \3240 );
not \U$3153 ( \3496 , \3495 );
or \U$3154 ( \3497 , \3494 , \3496 );
nand \U$3155 ( \3498 , \3255 , \1220 );
nand \U$3156 ( \3499 , \3497 , \3498 );
not \U$3157 ( \3500 , \1018 );
and \U$3158 ( \3501 , \3271 , \2962 );
not \U$3159 ( \3502 , \3271 );
and \U$3160 ( \3503 , \3502 , \2111 );
nor \U$3161 ( \3504 , \3501 , \3503 );
not \U$3162 ( \3505 , \3504 );
or \U$3163 ( \3506 , \3500 , \3505 );
or \U$3164 ( \3507 , \3277 , \1068 );
nand \U$3165 ( \3508 , \3506 , \3507 );
xor \U$3166 ( \3509 , \3499 , \3508 );
xor \U$3167 ( \3510 , \3493 , \3509 );
xor \U$3168 ( \3511 , \3483 , \3510 );
and \U$3169 ( \3512 , \3414 , \3419 );
not \U$3170 ( \3513 , \3414 );
and \U$3171 ( \3514 , \3513 , \3418 );
nor \U$3172 ( \3515 , \3512 , \3514 );
and \U$3173 ( \3516 , \3511 , \3515 );
and \U$3174 ( \3517 , \3483 , \3510 );
nor \U$3175 ( \3518 , \3516 , \3517 );
not \U$3176 ( \3519 , \3518 );
not \U$3177 ( \3520 , \3519 );
xnor \U$3178 ( \3521 , \3362 , \3385 );
not \U$3179 ( \3522 , \3521 );
not \U$3180 ( \3523 , \3522 );
not \U$3181 ( \3524 , \1220 );
not \U$3182 ( \3525 , \3495 );
or \U$3183 ( \3526 , \3524 , \3525 );
nand \U$3184 ( \3527 , \3229 , \434 );
not \U$3185 ( \3528 , \3527 );
not \U$3186 ( \3529 , \3528 );
not \U$3187 ( \3530 , \1177 );
not \U$3188 ( \3531 , \3530 );
or \U$3189 ( \3532 , \3529 , \3531 );
not \U$3190 ( \3533 , \3530 );
nand \U$3191 ( \3534 , \3533 , \3527 );
nand \U$3192 ( \3535 , \3532 , \3534 );
buf \U$3193 ( \3536 , \3535 );
buf \U$3194 ( \3537 , \3536 );
not \U$3195 ( \3538 , \3537 );
not \U$3196 ( \3539 , \1716 );
and \U$3197 ( \3540 , \3538 , \3539 );
not \U$3198 ( \3541 , \3536 );
buf \U$3199 ( \3542 , \3541 );
not \U$3200 ( \3543 , \3542 );
and \U$3201 ( \3544 , \3543 , \1716 );
nor \U$3202 ( \3545 , \3540 , \3544 );
not \U$3203 ( \3546 , \3545 );
nand \U$3204 ( \3547 , \3546 , \1162 );
nand \U$3205 ( \3548 , \3526 , \3547 );
buf \U$3206 ( \3549 , \411 );
and \U$3207 ( \3550 , \409 , \3549 , \414 );
not \U$3208 ( \3551 , \3550 );
not \U$3209 ( \3552 , \690 );
not \U$3210 ( \3553 , \687 );
or \U$3211 ( \3554 , \3552 , \3553 );
not \U$3212 ( \3555 , \408 );
nand \U$3213 ( \3556 , \3554 , \3555 );
not \U$3214 ( \3557 , \3556 );
or \U$3215 ( \3558 , \3551 , \3557 );
not \U$3216 ( \3559 , \426 );
nand \U$3217 ( \3560 , \3558 , \3559 );
not \U$3218 ( \3561 , \3560 );
nand \U$3219 ( \3562 , \410 , \428 );
not \U$3220 ( \3563 , \3562 );
and \U$3221 ( \3564 , \3561 , \3563 );
and \U$3222 ( \3565 , \3560 , \3562 );
nor \U$3223 ( \3566 , \3564 , \3565 );
buf \U$3224 ( \3567 , \3566 );
buf \U$3225 ( \3568 , \3567 );
not \U$3226 ( \3569 , \3568 );
nand \U$3227 ( \3570 , \3569 , \1165 );
xnor \U$3228 ( \3571 , \3548 , \3570 );
not \U$3229 ( \3572 , \2087 );
not \U$3230 ( \3573 , \3416 );
or \U$3231 ( \3574 , \3572 , \3573 );
and \U$3232 ( \3575 , RI9871aa0_133, \1417 );
not \U$3233 ( \3576 , RI9871aa0_133);
and \U$3234 ( \3577 , \3576 , \1418 );
nor \U$3235 ( \3578 , \3575 , \3577 );
nand \U$3236 ( \3579 , \3578 , \2074 );
nand \U$3237 ( \3580 , \3574 , \3579 );
and \U$3238 ( \3581 , \3571 , \3580 );
not \U$3239 ( \3582 , \3570 );
and \U$3240 ( \3583 , \3548 , \3582 );
nor \U$3241 ( \3584 , \3581 , \3583 );
not \U$3242 ( \3585 , \3584 );
or \U$3243 ( \3586 , \3264 , \1543 );
xor \U$3244 ( \3587 , RI9871b18_134, \2211 );
or \U$3245 ( \3588 , \3587 , \1293 );
nand \U$3246 ( \3589 , \3586 , \3588 );
nand \U$3247 ( \3590 , \3543 , \1165 );
not \U$3248 ( \3591 , \3467 );
not \U$3249 ( \3592 , \3591 );
not \U$3250 ( \3593 , RI98726d0_159);
not \U$3251 ( \3594 , \3593 );
and \U$3252 ( \3595 , \3592 , \3594 );
and \U$3253 ( \3596 , RI98726d0_159, \1693 );
not \U$3254 ( \3597 , RI98726d0_159);
and \U$3255 ( \3598 , \3597 , \1692 );
or \U$3256 ( \3599 , \3596 , \3598 );
buf \U$3257 ( \3600 , \3465 );
and \U$3258 ( \3601 , \3599 , \3600 );
nor \U$3259 ( \3602 , \3595 , \3601 );
not \U$3260 ( \3603 , \3602 );
and \U$3261 ( \3604 , \3590 , \3603 );
not \U$3262 ( \3605 , \3590 );
and \U$3263 ( \3606 , \3605 , \3602 );
nor \U$3264 ( \3607 , \3604 , \3606 );
and \U$3265 ( \3608 , \3589 , \3607 );
not \U$3266 ( \3609 , \3589 );
not \U$3267 ( \3610 , \3607 );
and \U$3268 ( \3611 , \3609 , \3610 );
or \U$3269 ( \3612 , \3608 , \3611 );
not \U$3270 ( \3613 , \3612 );
or \U$3271 ( \3614 , \3585 , \3613 );
or \U$3272 ( \3615 , \3612 , \3584 );
nand \U$3273 ( \3616 , \3614 , \3615 );
not \U$3274 ( \3617 , \3616 );
or \U$3275 ( \3618 , \3523 , \3617 );
not \U$3276 ( \3619 , \3584 );
nand \U$3277 ( \3620 , \3619 , \3612 );
nand \U$3278 ( \3621 , \3618 , \3620 );
not \U$3279 ( \3622 , \3621 );
xor \U$3280 ( \3623 , \3469 , \3475 );
and \U$3281 ( \3624 , \3623 , \3482 );
and \U$3282 ( \3625 , \3469 , \3475 );
nor \U$3283 ( \3626 , \3624 , \3625 );
not \U$3284 ( \3627 , \3508 );
not \U$3285 ( \3628 , \3499 );
or \U$3286 ( \3629 , \3627 , \3628 );
nand \U$3287 ( \3630 , \3493 , \3509 );
nand \U$3288 ( \3631 , \3629 , \3630 );
and \U$3289 ( \3632 , \3626 , \3631 );
not \U$3290 ( \3633 , \3626 );
not \U$3291 ( \3634 , \3631 );
and \U$3292 ( \3635 , \3633 , \3634 );
or \U$3293 ( \3636 , \3632 , \3635 );
xor \U$3294 ( \3637 , \3226 , \3241 );
xor \U$3295 ( \3638 , \3637 , \3250 );
not \U$3296 ( \3639 , \3638 );
xor \U$3297 ( \3640 , \3636 , \3639 );
not \U$3298 ( \3641 , \3640 );
or \U$3299 ( \3642 , \3622 , \3641 );
or \U$3300 ( \3643 , \3621 , \3640 );
nand \U$3301 ( \3644 , \3642 , \3643 );
not \U$3302 ( \3645 , \3644 );
or \U$3303 ( \3646 , \3520 , \3645 );
not \U$3304 ( \3647 , \3640 );
nand \U$3305 ( \3648 , \3647 , \3621 );
nand \U$3306 ( \3649 , \3646 , \3648 );
not \U$3307 ( \3650 , \3649 );
xor \U$3308 ( \3651 , \3215 , \3205 );
not \U$3309 ( \3652 , \3651 );
not \U$3310 ( \3653 , \3589 );
not \U$3311 ( \3654 , \3610 );
or \U$3312 ( \3655 , \3653 , \3654 );
or \U$3313 ( \3656 , \3602 , \3590 );
nand \U$3314 ( \3657 , \3655 , \3656 );
or \U$3315 ( \3658 , \3360 , \1746 );
and \U$3316 ( \3659 , \1800 , \1949 );
not \U$3317 ( \3660 , \1800 );
and \U$3318 ( \3661 , \3660 , \1344 );
nor \U$3319 ( \3662 , \3659 , \3661 );
or \U$3320 ( \3663 , \3662 , \1591 );
nand \U$3321 ( \3664 , \3658 , \3663 );
not \U$3322 ( \3665 , \797 );
not \U$3323 ( \3666 , \3478 );
or \U$3324 ( \3667 , \3665 , \3666 );
and \U$3325 ( \3668 , RI98719b0_131, \1320 );
not \U$3326 ( \3669 , RI98719b0_131);
and \U$3327 ( \3670 , \3669 , \1309 );
nor \U$3328 ( \3671 , \3668 , \3670 );
not \U$3329 ( \3672 , \3671 );
nand \U$3330 ( \3673 , \3672 , \794 );
nand \U$3331 ( \3674 , \3667 , \3673 );
not \U$3332 ( \3675 , \3164 );
xnor \U$3333 ( \3676 , \2399 , RI9872310_151);
not \U$3334 ( \3677 , \3676 );
or \U$3335 ( \3678 , \3675 , \3677 );
nand \U$3336 ( \3679 , \3471 , \3170 );
nand \U$3337 ( \3680 , \3678 , \3679 );
and \U$3338 ( \3681 , \3674 , \3680 );
not \U$3339 ( \3682 , \3674 );
not \U$3340 ( \3683 , \3680 );
and \U$3341 ( \3684 , \3682 , \3683 );
nor \U$3342 ( \3685 , \3681 , \3684 );
nand \U$3343 ( \3686 , \3664 , \3685 );
nand \U$3344 ( \3687 , \3674 , \3680 );
and \U$3345 ( \3688 , \3686 , \3687 );
not \U$3346 ( \3689 , \3688 );
not \U$3347 ( \3690 , \3689 );
buf \U$3348 ( \3691 , \2947 );
and \U$3349 ( \3692 , \3691 , \1044 );
not \U$3350 ( \3693 , \3691 );
and \U$3351 ( \3694 , \3693 , \1043 );
nor \U$3352 ( \3695 , \3692 , \3694 );
or \U$3353 ( \3696 , \3695 , \1612 );
not \U$3354 ( \3697 , \3504 );
or \U$3355 ( \3698 , \3697 , \1068 );
nand \U$3356 ( \3699 , \3696 , \3698 );
not \U$3357 ( \3700 , \1353 );
not \U$3358 ( \3701 , \3397 );
or \U$3359 ( \3702 , \3700 , \3701 );
and \U$3360 ( \3703 , RI9871e60_141, \1487 );
not \U$3361 ( \3704 , RI9871e60_141);
and \U$3362 ( \3705 , \3704 , \1486 );
nor \U$3363 ( \3706 , \3703 , \3705 );
not \U$3364 ( \3707 , \3706 );
nand \U$3365 ( \3708 , \3707 , \1382 );
nand \U$3366 ( \3709 , \3702 , \3708 );
xor \U$3367 ( \3710 , \3699 , \3709 );
not \U$3368 ( \3711 , \3491 );
or \U$3369 ( \3712 , \3711 , \1432 );
xor \U$3370 ( \3713 , RI9871c08_136, \824 );
or \U$3371 ( \3714 , \3713 , \1457 );
nand \U$3372 ( \3715 , \3712 , \3714 );
and \U$3373 ( \3716 , \3710 , \3715 );
and \U$3374 ( \3717 , \3699 , \3709 );
or \U$3375 ( \3718 , \3716 , \3717 );
not \U$3376 ( \3719 , \3718 );
not \U$3377 ( \3720 , \1083 );
xnor \U$3378 ( \3721 , \916 , RI98718c0_129);
not \U$3379 ( \3722 , \3721 );
or \U$3380 ( \3723 , \3720 , \3722 );
nand \U$3381 ( \3724 , \1136 , \3379 );
nand \U$3382 ( \3725 , \3723 , \3724 );
or \U$3383 ( \3726 , \3407 , \932 );
and \U$3384 ( \3727 , \3130 , RI9871d70_139);
and \U$3385 ( \3728 , \1212 , \1347 );
nor \U$3386 ( \3729 , \3727 , \3728 );
or \U$3387 ( \3730 , \3729 , \860 );
nand \U$3388 ( \3731 , \3726 , \3730 );
xor \U$3389 ( \3732 , \3725 , \3731 );
or \U$3390 ( \3733 , \3369 , \1470 );
and \U$3391 ( \3734 , \1714 , RI9872130_147);
and \U$3392 ( \3735 , \1713 , \919 );
nor \U$3393 ( \3736 , \3734 , \3735 );
or \U$3394 ( \3737 , \1942 , \3736 );
nand \U$3395 ( \3738 , \3733 , \3737 );
and \U$3396 ( \3739 , \3732 , \3738 );
and \U$3397 ( \3740 , \3725 , \3731 );
nor \U$3398 ( \3741 , \3739 , \3740 );
not \U$3399 ( \3742 , \3741 );
or \U$3400 ( \3743 , \3719 , \3742 );
or \U$3401 ( \3744 , \3718 , \3741 );
nand \U$3402 ( \3745 , \3743 , \3744 );
not \U$3403 ( \3746 , \3745 );
or \U$3404 ( \3747 , \3690 , \3746 );
not \U$3405 ( \3748 , \3741 );
nand \U$3406 ( \3749 , \3748 , \3718 );
nand \U$3407 ( \3750 , \3747 , \3749 );
xor \U$3408 ( \3751 , \3657 , \3750 );
and \U$3409 ( \3752 , \3422 , \3429 );
not \U$3410 ( \3753 , \3422 );
and \U$3411 ( \3754 , \3753 , \3428 );
or \U$3412 ( \3755 , \3752 , \3754 );
and \U$3413 ( \3756 , \3751 , \3755 );
and \U$3414 ( \3757 , \3657 , \3750 );
nor \U$3415 ( \3758 , \3756 , \3757 );
not \U$3416 ( \3759 , \3758 );
or \U$3417 ( \3760 , \3652 , \3759 );
or \U$3418 ( \3761 , \3758 , \3651 );
nand \U$3419 ( \3762 , \3760 , \3761 );
not \U$3420 ( \3763 , \3762 );
or \U$3421 ( \3764 , \3650 , \3763 );
not \U$3422 ( \3765 , \3758 );
nand \U$3423 ( \3766 , \3765 , \3651 );
nand \U$3424 ( \3767 , \3764 , \3766 );
not \U$3425 ( \3768 , \3767 );
xor \U$3426 ( \3769 , \3314 , \3253 );
not \U$3427 ( \3770 , \3769 );
not \U$3428 ( \3771 , \3770 );
not \U$3429 ( \3772 , \3639 );
not \U$3430 ( \3773 , \3772 );
not \U$3431 ( \3774 , \3636 );
or \U$3432 ( \3775 , \3773 , \3774 );
or \U$3433 ( \3776 , \3634 , \3626 );
nand \U$3434 ( \3777 , \3775 , \3776 );
not \U$3435 ( \3778 , \3777 );
xor \U$3436 ( \3779 , \3305 , \3297 );
not \U$3437 ( \3780 , \3779 );
and \U$3438 ( \3781 , \3138 , \3109 );
not \U$3439 ( \3782 , \3138 );
and \U$3440 ( \3783 , \3782 , \3110 );
nor \U$3441 ( \3784 , \3781 , \3783 );
not \U$3442 ( \3785 , \3784 );
xnor \U$3443 ( \3786 , \3267 , \3279 );
not \U$3444 ( \3787 , \3786 );
not \U$3445 ( \3788 , \3787 );
or \U$3446 ( \3789 , \3785 , \3788 );
not \U$3447 ( \3790 , \3784 );
nand \U$3448 ( \3791 , \3790 , \3786 );
nand \U$3449 ( \3792 , \3789 , \3791 );
not \U$3450 ( \3793 , \3792 );
or \U$3451 ( \3794 , \3780 , \3793 );
not \U$3452 ( \3795 , \3784 );
nand \U$3453 ( \3796 , \3795 , \3787 );
nand \U$3454 ( \3797 , \3794 , \3796 );
not \U$3455 ( \3798 , \3797 );
not \U$3456 ( \3799 , \3798 );
or \U$3457 ( \3800 , \3778 , \3799 );
not \U$3458 ( \3801 , \3777 );
nand \U$3459 ( \3802 , \3801 , \3797 );
nand \U$3460 ( \3803 , \3800 , \3802 );
not \U$3461 ( \3804 , \3803 );
or \U$3462 ( \3805 , \3771 , \3804 );
nand \U$3463 ( \3806 , \3797 , \3777 );
nand \U$3464 ( \3807 , \3805 , \3806 );
xor \U$3465 ( \3808 , \3220 , \3318 );
xor \U$3466 ( \3809 , \3808 , \3320 );
xor \U$3467 ( \3810 , \3807 , \3809 );
not \U$3468 ( \3811 , \3810 );
or \U$3469 ( \3812 , \3768 , \3811 );
nand \U$3470 ( \3813 , \3807 , \3809 );
nand \U$3471 ( \3814 , \3812 , \3813 );
not \U$3472 ( \3815 , \3814 );
not \U$3473 ( \3816 , \3815 );
and \U$3474 ( \3817 , \3453 , \3816 );
and \U$3475 ( \3818 , \3452 , \3815 );
nor \U$3476 ( \3819 , \3817 , \3818 );
xor \U$3477 ( \3820 , \3445 , \3436 );
xor \U$3478 ( \3821 , \3657 , \3750 );
xor \U$3479 ( \3822 , \3821 , \3755 );
not \U$3480 ( \3823 , \3822 );
and \U$3481 ( \3824 , \3745 , \3689 );
not \U$3482 ( \3825 , \3745 );
and \U$3483 ( \3826 , \3825 , \3688 );
nor \U$3484 ( \3827 , \3824 , \3826 );
not \U$3485 ( \3828 , \3827 );
not \U$3486 ( \3829 , \3587 );
not \U$3487 ( \3830 , \1543 );
and \U$3488 ( \3831 , \3829 , \3830 );
not \U$3489 ( \3832 , \944 );
and \U$3490 ( \3833 , \1283 , \3832 );
not \U$3491 ( \3834 , \1283 );
not \U$3492 ( \3835 , \943 );
not \U$3493 ( \3836 , \3835 );
and \U$3494 ( \3837 , \3834 , \3836 );
nor \U$3495 ( \3838 , \3833 , \3837 );
and \U$3496 ( \3839 , \3838 , \1292 );
nor \U$3497 ( \3840 , \3831 , \3839 );
and \U$3498 ( \3841 , \3840 , \3603 );
not \U$3499 ( \3842 , \3840 );
and \U$3500 ( \3843 , \3842 , \3602 );
nor \U$3501 ( \3844 , \3841 , \3843 );
not \U$3502 ( \3845 , \3844 );
or \U$3503 ( \3846 , \3706 , \1989 );
and \U$3504 ( \3847 , RI9871e60_141, \2962 );
not \U$3505 ( \3848 , RI9871e60_141);
and \U$3506 ( \3849 , \3848 , \2111 );
nor \U$3507 ( \3850 , \3847 , \3849 );
or \U$3508 ( \3851 , \3850 , \1558 );
nand \U$3509 ( \3852 , \3846 , \3851 );
and \U$3510 ( \3853 , \1045 , \3240 );
not \U$3511 ( \3854 , \1045 );
and \U$3512 ( \3855 , \3234 , \3227 );
not \U$3513 ( \3856 , \3234 );
and \U$3514 ( \3857 , \3856 , \3237 );
nor \U$3515 ( \3858 , \3855 , \3857 );
buf \U$3516 ( \3859 , \3858 );
not \U$3517 ( \3860 , \3859 );
not \U$3518 ( \3861 , \3860 );
and \U$3519 ( \3862 , \3854 , \3861 );
nor \U$3520 ( \3863 , \3853 , \3862 );
or \U$3521 ( \3864 , \3863 , \1612 );
or \U$3522 ( \3865 , \3695 , \1068 );
nand \U$3523 ( \3866 , \3864 , \3865 );
xor \U$3524 ( \3867 , \3852 , \3866 );
not \U$3525 ( \3868 , \1136 );
not \U$3526 ( \3869 , \3721 );
or \U$3527 ( \3870 , \3868 , \3869 );
not \U$3528 ( \3871 , \894 );
and \U$3529 ( \3872 , RI98718c0_129, \3871 );
not \U$3530 ( \3873 , RI98718c0_129);
and \U$3531 ( \3874 , \3873 , \894 );
nor \U$3532 ( \3875 , \3872 , \3874 );
nand \U$3533 ( \3876 , \3875 , \1083 );
nand \U$3534 ( \3877 , \3870 , \3876 );
and \U$3535 ( \3878 , \3867 , \3877 );
and \U$3536 ( \3879 , \3852 , \3866 );
or \U$3537 ( \3880 , \3878 , \3879 );
not \U$3538 ( \3881 , \3880 );
or \U$3539 ( \3882 , \3845 , \3881 );
or \U$3540 ( \3883 , \3840 , \3603 );
nand \U$3541 ( \3884 , \3882 , \3883 );
not \U$3542 ( \3885 , \1501 );
not \U$3543 ( \3886 , \1371 );
and \U$3544 ( \3887 , RI9871c80_137, \3886 );
not \U$3545 ( \3888 , RI9871c80_137);
and \U$3546 ( \3889 , \3888 , \1371 );
or \U$3547 ( \3890 , \3887 , \3889 );
not \U$3548 ( \3891 , \3890 );
or \U$3549 ( \3892 , \3885 , \3891 );
or \U$3550 ( \3893 , \3662 , \1746 );
nand \U$3551 ( \3894 , \3892 , \3893 );
not \U$3552 ( \3895 , \1323 );
not \U$3553 ( \3896 , \3838 );
or \U$3554 ( \3897 , \3895 , \3896 );
and \U$3555 ( \3898 , RI9871b18_134, \1257 );
not \U$3556 ( \3899 , RI9871b18_134);
and \U$3557 ( \3900 , \3899 , \1659 );
nor \U$3558 ( \3901 , \3898 , \3900 );
or \U$3559 ( \3902 , \3901 , \1293 );
nand \U$3560 ( \3903 , \3897 , \3902 );
xor \U$3561 ( \3904 , \3894 , \3903 );
or \U$3562 ( \3905 , \3671 , \3244 );
and \U$3563 ( \3906 , \1078 , \1275 );
not \U$3564 ( \3907 , \1078 );
and \U$3565 ( \3908 , \3907 , \1583 );
nor \U$3566 ( \3909 , \3906 , \3908 );
or \U$3567 ( \3910 , \3909 , \792 );
nand \U$3568 ( \3911 , \3905 , \3910 );
and \U$3569 ( \3912 , \3904 , \3911 );
and \U$3570 ( \3913 , \3894 , \3903 );
or \U$3571 ( \3914 , \3912 , \3913 );
not \U$3572 ( \3915 , \2087 );
not \U$3573 ( \3916 , \3578 );
or \U$3574 ( \3917 , \3915 , \3916 );
and \U$3575 ( \3918 , \2076 , \2680 );
not \U$3576 ( \3919 , \2076 );
and \U$3577 ( \3920 , \3919 , \1799 );
nor \U$3578 ( \3921 , \3918 , \3920 );
or \U$3579 ( \3922 , \3921 , \2073 );
nand \U$3580 ( \3923 , \3917 , \3922 );
not \U$3581 ( \3924 , \3923 );
and \U$3582 ( \3925 , RI9872388_152, RI98727c0_161);
nor \U$3583 ( \3926 , \3925 , \3454 );
not \U$3584 ( \3927 , \3926 );
not \U$3585 ( \3928 , \3467 );
not \U$3586 ( \3929 , \3599 );
or \U$3587 ( \3930 , \3928 , \3929 );
not \U$3588 ( \3931 , \1393 );
not \U$3589 ( \3932 , \3593 );
and \U$3590 ( \3933 , \3931 , \3932 );
and \U$3591 ( \3934 , \1394 , \3593 );
nor \U$3592 ( \3935 , \3933 , \3934 );
not \U$3593 ( \3936 , \3935 );
nand \U$3594 ( \3937 , \3936 , \3600 );
nand \U$3595 ( \3938 , \3930 , \3937 );
not \U$3596 ( \3939 , \3938 );
or \U$3597 ( \3940 , \3927 , \3939 );
or \U$3598 ( \3941 , \3938 , \3926 );
nand \U$3599 ( \3942 , \3940 , \3941 );
not \U$3600 ( \3943 , \3942 );
or \U$3601 ( \3944 , \3924 , \3943 );
not \U$3602 ( \3945 , \3926 );
nand \U$3603 ( \3946 , \3945 , \3938 );
nand \U$3604 ( \3947 , \3944 , \3946 );
xor \U$3605 ( \3948 , \3914 , \3947 );
or \U$3606 ( \3949 , \3736 , \1470 );
and \U$3607 ( \3950 , RI9872130_147, \1041 );
not \U$3608 ( \3951 , RI9872130_147);
and \U$3609 ( \3952 , \3951 , \1595 );
nor \U$3610 ( \3953 , \3950 , \3952 );
or \U$3611 ( \3954 , \1942 , \3953 );
nand \U$3612 ( \3955 , \3949 , \3954 );
not \U$3613 ( \3956 , \3170 );
not \U$3614 ( \3957 , \3676 );
or \U$3615 ( \3958 , \3956 , \3957 );
and \U$3616 ( \3959 , \1097 , RI9872310_151);
and \U$3617 ( \3960 , \1106 , \3154 );
nor \U$3618 ( \3961 , \3959 , \3960 );
not \U$3619 ( \3962 , \3163 );
or \U$3620 ( \3963 , \3961 , \3962 );
nand \U$3621 ( \3964 , \3958 , \3963 );
xor \U$3622 ( \3965 , \3955 , \3964 );
or \U$3623 ( \3966 , \3729 , \932 );
and \U$3624 ( \3967 , RI9871d70_139, \1191 );
not \U$3625 ( \3968 , RI9871d70_139);
not \U$3626 ( \3969 , \3396 );
and \U$3627 ( \3970 , \3968 , \3969 );
nor \U$3628 ( \3971 , \3967 , \3970 );
or \U$3629 ( \3972 , \3971 , \860 );
nand \U$3630 ( \3973 , \3966 , \3972 );
and \U$3631 ( \3974 , \3965 , \3973 );
and \U$3632 ( \3975 , \3955 , \3964 );
or \U$3633 ( \3976 , \3974 , \3975 );
and \U$3634 ( \3977 , \3948 , \3976 );
and \U$3635 ( \3978 , \3914 , \3947 );
or \U$3636 ( \3979 , \3977 , \3978 );
xor \U$3637 ( \3980 , \3884 , \3979 );
not \U$3638 ( \3981 , \3980 );
or \U$3639 ( \3982 , \3828 , \3981 );
nand \U$3640 ( \3983 , \3979 , \3884 );
nand \U$3641 ( \3984 , \3982 , \3983 );
not \U$3642 ( \3985 , \3984 );
not \U$3643 ( \3986 , \3779 );
and \U$3644 ( \3987 , \3792 , \3986 );
not \U$3645 ( \3988 , \3792 );
and \U$3646 ( \3989 , \3988 , \3779 );
nor \U$3647 ( \3990 , \3987 , \3989 );
not \U$3648 ( \3991 , \3990 );
or \U$3649 ( \3992 , \3985 , \3991 );
or \U$3650 ( \3993 , \3990 , \3984 );
nand \U$3651 ( \3994 , \3992 , \3993 );
not \U$3652 ( \3995 , \3994 );
or \U$3653 ( \3996 , \3823 , \3995 );
not \U$3654 ( \3997 , \3990 );
nand \U$3655 ( \3998 , \3997 , \3984 );
nand \U$3656 ( \3999 , \3996 , \3998 );
not \U$3657 ( \4000 , \3999 );
not \U$3658 ( \4001 , \3354 );
not \U$3659 ( \4002 , \3431 );
not \U$3660 ( \4003 , \4002 );
or \U$3661 ( \4004 , \4001 , \4003 );
not \U$3662 ( \4005 , \3354 );
nand \U$3663 ( \4006 , \4005 , \3431 );
nand \U$3664 ( \4007 , \4004 , \4006 );
xor \U$3665 ( \4008 , \3769 , \4007 );
xnor \U$3666 ( \4009 , \4008 , \3803 );
not \U$3667 ( \4010 , \4009 );
or \U$3668 ( \4011 , \4000 , \4010 );
and \U$3669 ( \4012 , \3803 , \3769 );
not \U$3670 ( \4013 , \3803 );
and \U$3671 ( \4014 , \4013 , \3770 );
or \U$3672 ( \4015 , \4012 , \4014 );
nand \U$3673 ( \4016 , \4015 , \4007 );
nand \U$3674 ( \4017 , \4011 , \4016 );
xor \U$3675 ( \4018 , \3820 , \4017 );
not \U$3676 ( \4019 , \3810 );
not \U$3677 ( \4020 , \3767 );
not \U$3678 ( \4021 , \4020 );
and \U$3679 ( \4022 , \4019 , \4021 );
and \U$3680 ( \4023 , \3810 , \4020 );
nor \U$3681 ( \4024 , \4022 , \4023 );
not \U$3682 ( \4025 , \4024 );
and \U$3683 ( \4026 , \4018 , \4025 );
and \U$3684 ( \4027 , \3820 , \4017 );
nor \U$3685 ( \4028 , \4026 , \4027 );
nand \U$3686 ( \4029 , \3819 , \4028 );
nand \U$3687 ( \4030 , \3452 , \3814 );
not \U$3688 ( \4031 , \3335 );
and \U$3689 ( \4032 , \3201 , \4031 );
not \U$3690 ( \4033 , \3201 );
and \U$3691 ( \4034 , \4033 , \3335 );
nor \U$3692 ( \4035 , \4032 , \4034 );
and \U$3693 ( \4036 , \3203 , \3329 );
not \U$3694 ( \4037 , \3203 );
and \U$3695 ( \4038 , \4037 , \3330 );
or \U$3696 ( \4039 , \4036 , \4038 );
nand \U$3697 ( \4040 , \4039 , \3450 );
nand \U$3698 ( \4041 , \4030 , \4035 , \4040 );
nand \U$3699 ( \4042 , \3345 , \4029 , \4041 );
not \U$3700 ( \4043 , \4042 );
not \U$3701 ( \4044 , RI9871b18_134);
and \U$3702 ( \4045 , \1344 , \4044 );
not \U$3703 ( \4046 , \1344 );
and \U$3704 ( \4047 , \4046 , RI9871b18_134);
nor \U$3705 ( \4048 , \4045 , \4047 );
not \U$3706 ( \4049 , \4048 );
not \U$3707 ( \4050 , \1292 );
or \U$3708 ( \4051 , \4049 , \4050 );
or \U$3709 ( \4052 , \3901 , \1543 );
nand \U$3710 ( \4053 , \4051 , \4052 );
not \U$3711 ( \4054 , \4053 );
not \U$3712 ( \4055 , \2074 );
xor \U$3713 ( \4056 , \1309 , RI9871aa0_133);
not \U$3714 ( \4057 , \4056 );
or \U$3715 ( \4058 , \4055 , \4057 );
not \U$3716 ( \4059 , \3921 );
nand \U$3717 ( \4060 , \4059 , \2087 );
nand \U$3718 ( \4061 , \4058 , \4060 );
not \U$3719 ( \4062 , \3466 );
not \U$3720 ( \4063 , RI98726d0_159);
and \U$3721 ( \4064 , \1725 , \4063 );
not \U$3722 ( \4065 , \1725 );
and \U$3723 ( \4066 , \4065 , RI98726d0_159);
nor \U$3724 ( \4067 , \4064 , \4066 );
not \U$3725 ( \4068 , \4067 );
or \U$3726 ( \4069 , \4062 , \4068 );
or \U$3727 ( \4070 , \3935 , \3591 );
nand \U$3728 ( \4071 , \4069 , \4070 );
xor \U$3729 ( \4072 , \4061 , \4071 );
not \U$3730 ( \4073 , \4072 );
or \U$3731 ( \4074 , \4054 , \4073 );
nand \U$3732 ( \4075 , \4061 , \4071 );
nand \U$3733 ( \4076 , \4074 , \4075 );
not \U$3734 ( \4077 , \4076 );
not \U$3735 ( \4078 , RI98725e0_157);
and \U$3736 ( \4079 , RI9872388_152, RI98727c0_161);
not \U$3737 ( \4080 , RI9872388_152);
not \U$3738 ( \4081 , RI98727c0_161);
and \U$3739 ( \4082 , \4080 , \4081 );
nor \U$3740 ( \4083 , \4079 , \4082 );
buf \U$3741 ( \4084 , \4083 );
buf \U$3742 ( \4085 , \4084 );
not \U$3743 ( \4086 , \4085 );
or \U$3744 ( \4087 , \4078 , \4086 );
not \U$3745 ( \4088 , RI98725e0_157);
not \U$3746 ( \4089 , \4088 );
not \U$3747 ( \4090 , \1692 );
or \U$3748 ( \4091 , \4089 , \4090 );
not \U$3749 ( \4092 , RI98725e0_157);
or \U$3750 ( \4093 , \780 , \4092 );
nand \U$3751 ( \4094 , \4091 , \4093 );
not \U$3752 ( \4095 , \4083 );
and \U$3753 ( \4096 , RI98725e0_157, RI98727c0_161);
not \U$3754 ( \4097 , RI98725e0_157);
and \U$3755 ( \4098 , \4097 , \4081 );
nor \U$3756 ( \4099 , \4096 , \4098 );
nand \U$3757 ( \4100 , \4095 , \4099 );
not \U$3758 ( \4101 , \4100 );
not \U$3759 ( \4102 , \4101 );
not \U$3760 ( \4103 , \4102 );
nand \U$3761 ( \4104 , \4094 , \4103 );
nand \U$3762 ( \4105 , \4087 , \4104 );
not \U$3763 ( \4106 , \4105 );
not \U$3764 ( \4107 , \4106 );
not \U$3765 ( \4108 , \3890 );
or \U$3766 ( \4109 , \4108 , \1746 );
and \U$3767 ( \4110 , \2842 , RI9871c80_137);
and \U$3768 ( \4111 , \1062 , \1584 );
nor \U$3769 ( \4112 , \4110 , \4111 );
or \U$3770 ( \4113 , \4112 , \1591 );
nand \U$3771 ( \4114 , \4109 , \4113 );
or \U$3772 ( \4115 , \1470 , \3953 );
not \U$3773 ( \4116 , RI9872130_147);
and \U$3774 ( \4117 , \4116 , \1212 );
not \U$3775 ( \4118 , \4116 );
and \U$3776 ( \4119 , \4118 , \3130 );
nor \U$3777 ( \4120 , \4117 , \4119 );
or \U$3778 ( \4121 , \3370 , \4120 );
nand \U$3779 ( \4122 , \4115 , \4121 );
xor \U$3780 ( \4123 , \4114 , \4122 );
or \U$3781 ( \4124 , \3909 , \3244 );
xor \U$3782 ( \4125 , \918 , RI98719b0_131);
or \U$3783 ( \4126 , \4125 , \792 );
nand \U$3784 ( \4127 , \4124 , \4126 );
and \U$3785 ( \4128 , \4123 , \4127 );
and \U$3786 ( \4129 , \4114 , \4122 );
or \U$3787 ( \4130 , \4128 , \4129 );
not \U$3788 ( \4131 , \4130 );
or \U$3789 ( \4132 , \4107 , \4131 );
or \U$3790 ( \4133 , \4130 , \4106 );
nand \U$3791 ( \4134 , \4132 , \4133 );
not \U$3792 ( \4135 , \4134 );
or \U$3793 ( \4136 , \4077 , \4135 );
nand \U$3794 ( \4137 , \4130 , \4105 );
nand \U$3795 ( \4138 , \4136 , \4137 );
xnor \U$3796 ( \4139 , \3732 , \3738 );
not \U$3797 ( \4140 , \4139 );
xor \U$3798 ( \4141 , \3699 , \3709 );
xor \U$3799 ( \4142 , \4141 , \3715 );
not \U$3800 ( \4143 , \4142 );
or \U$3801 ( \4144 , \4140 , \4143 );
or \U$3802 ( \4145 , \4142 , \4139 );
nand \U$3803 ( \4146 , \4144 , \4145 );
nand \U$3804 ( \4147 , \4138 , \4146 );
not \U$3805 ( \4148 , \4139 );
nand \U$3806 ( \4149 , \4148 , \4142 );
and \U$3807 ( \4150 , \4147 , \4149 );
xor \U$3808 ( \4151 , \3980 , \3827 );
xor \U$3809 ( \4152 , \4150 , \4151 );
not \U$3810 ( \4153 , \3567 );
not \U$3811 ( \4154 , \4153 );
not \U$3812 ( \4155 , \4154 );
and \U$3813 ( \4156 , \1716 , \4155 );
not \U$3814 ( \4157 , \1716 );
and \U$3815 ( \4158 , \4157 , \3568 );
nor \U$3816 ( \4159 , \4156 , \4158 );
or \U$3817 ( \4160 , \4159 , \1809 );
or \U$3818 ( \4161 , \3545 , \1719 );
nand \U$3819 ( \4162 , \4160 , \4161 );
not \U$3820 ( \4163 , \3549 );
and \U$3821 ( \4164 , \3556 , \414 );
not \U$3822 ( \4165 , \4164 );
or \U$3823 ( \4166 , \4163 , \4165 );
not \U$3824 ( \4167 , \422 );
nand \U$3825 ( \4168 , \4166 , \4167 );
nand \U$3826 ( \4169 , \409 , \425 );
not \U$3827 ( \4170 , \4169 );
and \U$3828 ( \4171 , \4168 , \4170 );
not \U$3829 ( \4172 , \4168 );
and \U$3830 ( \4173 , \4172 , \4169 );
nor \U$3831 ( \4174 , \4171 , \4173 );
not \U$3832 ( \4175 , \4174 );
buf \U$3833 ( \4176 , \4175 );
not \U$3834 ( \4177 , \4176 );
and \U$3835 ( \4178 , \4177 , \1165 );
xor \U$3836 ( \4179 , \4162 , \4178 );
not \U$3837 ( \4180 , \1431 );
not \U$3838 ( \4181 , \3713 );
not \U$3839 ( \4182 , \4181 );
or \U$3840 ( \4183 , \4180 , \4182 );
and \U$3841 ( \4184 , RI9871c08_136, \848 );
not \U$3842 ( \4185 , RI9871c08_136);
and \U$3843 ( \4186 , \4185 , \847 );
nor \U$3844 ( \4187 , \4184 , \4186 );
or \U$3845 ( \4188 , \4187 , \1457 );
nand \U$3846 ( \4189 , \4183 , \4188 );
xor \U$3847 ( \4190 , \4179 , \4189 );
not \U$3848 ( \4191 , \4190 );
xor \U$3849 ( \4192 , \3852 , \3866 );
xor \U$3850 ( \4193 , \4192 , \3877 );
xor \U$3851 ( \4194 , \3923 , \3942 );
or \U$3852 ( \4195 , \4193 , \4194 );
not \U$3853 ( \4196 , \4195 );
or \U$3854 ( \4197 , \4191 , \4196 );
nand \U$3855 ( \4198 , \4193 , \4194 );
nand \U$3856 ( \4199 , \4197 , \4198 );
not \U$3857 ( \4200 , \4199 );
not \U$3858 ( \4201 , \3880 );
xor \U$3859 ( \4202 , \3844 , \4201 );
not \U$3860 ( \4203 , \4202 );
xor \U$3861 ( \4204 , \3914 , \3947 );
xor \U$3862 ( \4205 , \4204 , \3976 );
not \U$3863 ( \4206 , \4205 );
or \U$3864 ( \4207 , \4203 , \4206 );
or \U$3865 ( \4208 , \4202 , \4205 );
nand \U$3866 ( \4209 , \4207 , \4208 );
not \U$3867 ( \4210 , \4209 );
or \U$3868 ( \4211 , \4200 , \4210 );
not \U$3869 ( \4212 , \4202 );
nand \U$3870 ( \4213 , \4212 , \4205 );
nand \U$3871 ( \4214 , \4211 , \4213 );
xnor \U$3872 ( \4215 , \4152 , \4214 );
xnor \U$3873 ( \4216 , \3521 , \3616 );
not \U$3874 ( \4217 , \4216 );
xor \U$3875 ( \4218 , \3685 , \3664 );
not \U$3876 ( \4219 , \4218 );
not \U$3877 ( \4220 , \4178 );
not \U$3878 ( \4221 , \4162 );
or \U$3879 ( \4222 , \4220 , \4221 );
nand \U$3880 ( \4223 , \4189 , \4179 );
nand \U$3881 ( \4224 , \4222 , \4223 );
xnor \U$3882 ( \4225 , \3571 , \3580 );
and \U$3883 ( \4226 , \4224 , \4225 );
not \U$3884 ( \4227 , \4224 );
not \U$3885 ( \4228 , \4225 );
and \U$3886 ( \4229 , \4227 , \4228 );
or \U$3887 ( \4230 , \4226 , \4229 );
not \U$3888 ( \4231 , \4230 );
or \U$3889 ( \4232 , \4219 , \4231 );
nand \U$3890 ( \4233 , \4228 , \4224 );
nand \U$3891 ( \4234 , \4232 , \4233 );
not \U$3892 ( \4235 , \4234 );
not \U$3893 ( \4236 , \4235 );
and \U$3894 ( \4237 , \4217 , \4236 );
and \U$3895 ( \4238 , \4216 , \4235 );
nor \U$3896 ( \4239 , \4237 , \4238 );
not \U$3897 ( \4240 , \4239 );
xor \U$3898 ( \4241 , \3483 , \3510 );
xor \U$3899 ( \4242 , \4241 , \3515 );
not \U$3900 ( \4243 , \4242 );
and \U$3901 ( \4244 , \4240 , \4243 );
and \U$3902 ( \4245 , \4239 , \4242 );
nor \U$3903 ( \4246 , \4244 , \4245 );
not \U$3904 ( \4247 , \4246 );
xnor \U$3905 ( \4248 , \4230 , \4218 );
not \U$3906 ( \4249 , \4248 );
not \U$3907 ( \4250 , \4249 );
xor \U$3908 ( \4251 , \3894 , \3903 );
xor \U$3909 ( \4252 , \4251 , \3911 );
not \U$3910 ( \4253 , \4252 );
not \U$3911 ( \4254 , \3164 );
and \U$3912 ( \4255 , \1418 , \3154 );
not \U$3913 ( \4256 , \1418 );
and \U$3914 ( \4257 , \4256 , RI9872310_151);
nor \U$3915 ( \4258 , \4255 , \4257 );
not \U$3916 ( \4259 , \4258 );
or \U$3917 ( \4260 , \4254 , \4259 );
not \U$3918 ( \4261 , \3170 );
or \U$3919 ( \4262 , \3961 , \4261 );
nand \U$3920 ( \4263 , \4260 , \4262 );
or \U$3921 ( \4264 , \3971 , \932 );
and \U$3922 ( \4265 , RI9871d70_139, \2116 );
not \U$3923 ( \4266 , RI9871d70_139);
and \U$3924 ( \4267 , \4266 , \1486 );
nor \U$3925 ( \4268 , \4265 , \4267 );
or \U$3926 ( \4269 , \4268 , \860 );
nand \U$3927 ( \4270 , \4264 , \4269 );
xor \U$3928 ( \4271 , \4263 , \4270 );
not \U$3929 ( \4272 , \3875 );
or \U$3930 ( \4273 , \4272 , \1137 );
xor \U$3931 ( \4274 , RI98718c0_129, \824 );
or \U$3932 ( \4275 , \4274 , \1676 );
nand \U$3933 ( \4276 , \4273 , \4275 );
and \U$3934 ( \4277 , \4271 , \4276 );
and \U$3935 ( \4278 , \4263 , \4270 );
or \U$3936 ( \4279 , \4277 , \4278 );
and \U$3937 ( \4280 , \3542 , \1044 );
and \U$3938 ( \4281 , \3543 , \3271 );
nor \U$3939 ( \4282 , \4280 , \4281 );
or \U$3940 ( \4283 , \4282 , \1612 );
or \U$3941 ( \4284 , \3863 , \1068 );
nand \U$3942 ( \4285 , \4283 , \4284 );
not \U$3943 ( \4286 , \1381 );
not \U$3944 ( \4287 , \2948 );
and \U$3945 ( \4288 , RI9871e60_141, \4287 );
not \U$3946 ( \4289 , RI9871e60_141);
and \U$3947 ( \4290 , \4289 , \2948 );
or \U$3948 ( \4291 , \4288 , \4290 );
not \U$3949 ( \4292 , \4291 );
or \U$3950 ( \4293 , \4286 , \4292 );
or \U$3951 ( \4294 , \3850 , \2595 );
nand \U$3952 ( \4295 , \4293 , \4294 );
xor \U$3953 ( \4296 , \4285 , \4295 );
not \U$3954 ( \4297 , \1456 );
xor \U$3955 ( \4298 , \944 , RI9871c08_136);
not \U$3956 ( \4299 , \4298 );
or \U$3957 ( \4300 , \4297 , \4299 );
or \U$3958 ( \4301 , \4187 , \1432 );
nand \U$3959 ( \4302 , \4300 , \4301 );
and \U$3960 ( \4303 , \4296 , \4302 );
and \U$3961 ( \4304 , \4295 , \4285 );
nor \U$3962 ( \4305 , \4303 , \4304 );
not \U$3963 ( \4306 , \4305 );
and \U$3964 ( \4307 , \4279 , \4306 );
not \U$3965 ( \4308 , \4279 );
and \U$3966 ( \4309 , \4308 , \4305 );
nor \U$3967 ( \4310 , \4307 , \4309 );
not \U$3968 ( \4311 , \4310 );
or \U$3969 ( \4312 , \4253 , \4311 );
nand \U$3970 ( \4313 , \4306 , \4279 );
nand \U$3971 ( \4314 , \4312 , \4313 );
not \U$3972 ( \4315 , \4314 );
not \U$3973 ( \4316 , \4315 );
or \U$3974 ( \4317 , \4250 , \4316 );
nand \U$3975 ( \4318 , \4314 , \4248 );
nand \U$3976 ( \4319 , \4317 , \4318 );
not \U$3977 ( \4320 , \4319 );
xor \U$3978 ( \4321 , \4146 , \4138 );
not \U$3979 ( \4322 , \4321 );
or \U$3980 ( \4323 , \4320 , \4322 );
nand \U$3981 ( \4324 , \4314 , \4249 );
nand \U$3982 ( \4325 , \4323 , \4324 );
not \U$3983 ( \4326 , \4325 );
or \U$3984 ( \4327 , \4247 , \4326 );
or \U$3985 ( \4328 , \4325 , \4246 );
nand \U$3986 ( \4329 , \4327 , \4328 );
and \U$3987 ( \4330 , \4215 , \4329 );
not \U$3988 ( \4331 , \4215 );
not \U$3989 ( \4332 , \4329 );
and \U$3990 ( \4333 , \4331 , \4332 );
nor \U$3991 ( \4334 , \4330 , \4333 );
not \U$3992 ( \4335 , \4334 );
xor \U$3993 ( \4336 , \4310 , \4252 );
not \U$3994 ( \4337 , \4336 );
or \U$3995 ( \4338 , \4268 , \932 );
and \U$3996 ( \4339 , RI9871d70_139, \2962 );
not \U$3997 ( \4340 , RI9871d70_139);
and \U$3998 ( \4341 , \4340 , \2111 );
nor \U$3999 ( \4342 , \4339 , \4341 );
or \U$4000 ( \4343 , \4342 , \860 );
nand \U$4001 ( \4344 , \4338 , \4343 );
not \U$4002 ( \4345 , \3467 );
not \U$4003 ( \4346 , \4067 );
or \U$4004 ( \4347 , \4345 , \4346 );
and \U$4005 ( \4348 , \1106 , RI98726d0_159);
not \U$4006 ( \4349 , \1106 );
and \U$4007 ( \4350 , \4349 , \3593 );
nor \U$4008 ( \4351 , \4348 , \4350 );
nand \U$4009 ( \4352 , \4351 , \3466 );
nand \U$4010 ( \4353 , \4347 , \4352 );
xor \U$4011 ( \4354 , \4344 , \4353 );
not \U$4012 ( \4355 , \793 );
and \U$4013 ( \4356 , RI98719b0_131, \895 );
not \U$4014 ( \4357 , RI98719b0_131);
and \U$4015 ( \4358 , \4357 , \1506 );
nor \U$4016 ( \4359 , \4356 , \4358 );
not \U$4017 ( \4360 , \4359 );
or \U$4018 ( \4361 , \4355 , \4360 );
not \U$4019 ( \4362 , \4125 );
nand \U$4020 ( \4363 , \4362 , \797 );
nand \U$4021 ( \4364 , \4361 , \4363 );
and \U$4022 ( \4365 , \4354 , \4364 );
and \U$4023 ( \4366 , \4344 , \4353 );
or \U$4024 ( \4367 , \4365 , \4366 );
not \U$4025 ( \4368 , \1382 );
not \U$4026 ( \4369 , \3859 );
not \U$4027 ( \4370 , \4369 );
xnor \U$4028 ( \4371 , \4370 , RI9871e60_141);
not \U$4029 ( \4372 , \4371 );
or \U$4030 ( \4373 , \4368 , \4372 );
nand \U$4031 ( \4374 , \4291 , \1353 );
nand \U$4032 ( \4375 , \4373 , \4374 );
and \U$4033 ( \4376 , \1044 , \4154 );
not \U$4034 ( \4377 , \1044 );
and \U$4035 ( \4378 , \4377 , \3569 );
nor \U$4036 ( \4379 , \4376 , \4378 );
or \U$4037 ( \4380 , \4379 , \1612 );
or \U$4038 ( \4381 , \4282 , \1068 );
nand \U$4039 ( \4382 , \4380 , \4381 );
xor \U$4040 ( \4383 , \4375 , \4382 );
not \U$4041 ( \4384 , \4383 );
not \U$4042 ( \4385 , \1083 );
xnor \U$4043 ( \4386 , \2211 , RI98718c0_129);
not \U$4044 ( \4387 , \4386 );
or \U$4045 ( \4388 , \4385 , \4387 );
not \U$4046 ( \4389 , \4274 );
nand \U$4047 ( \4390 , \4389 , \1136 );
nand \U$4048 ( \4391 , \4388 , \4390 );
not \U$4049 ( \4392 , \4391 );
or \U$4050 ( \4393 , \4384 , \4392 );
nand \U$4051 ( \4394 , \4375 , \4382 );
nand \U$4052 ( \4395 , \4393 , \4394 );
xor \U$4053 ( \4396 , \4367 , \4395 );
not \U$4054 ( \4397 , \414 );
not \U$4055 ( \4398 , \3556 );
or \U$4056 ( \4399 , \4397 , \4398 );
nand \U$4057 ( \4400 , \4399 , \419 );
not \U$4058 ( \4401 , \4400 );
nand \U$4059 ( \4402 , \3549 , \421 );
not \U$4060 ( \4403 , \4402 );
and \U$4061 ( \4404 , \4401 , \4403 );
and \U$4062 ( \4405 , \4400 , \4402 );
nor \U$4063 ( \4406 , \4404 , \4405 );
not \U$4064 ( \4407 , \4406 );
not \U$4065 ( \4408 , \4407 );
not \U$4066 ( \4409 , \4408 );
not \U$4067 ( \4410 , \4409 );
nor \U$4068 ( \4411 , \4410 , \1716 );
not \U$4069 ( \4412 , \4411 );
not \U$4070 ( \4413 , \4105 );
or \U$4071 ( \4414 , \4412 , \4413 );
or \U$4072 ( \4415 , \4105 , \4411 );
nand \U$4073 ( \4416 , \4414 , \4415 );
and \U$4074 ( \4417 , \4177 , \1716 );
not \U$4075 ( \4418 , \4177 );
and \U$4076 ( \4419 , \4418 , \1165 );
nor \U$4077 ( \4420 , \4417 , \4419 );
or \U$4078 ( \4421 , \4420 , \1809 );
or \U$4079 ( \4422 , \1719 , \4159 );
nand \U$4080 ( \4423 , \4421 , \4422 );
xor \U$4081 ( \4424 , \4416 , \4423 );
and \U$4082 ( \4425 , \4396 , \4424 );
and \U$4083 ( \4426 , \4367 , \4395 );
nor \U$4084 ( \4427 , \4425 , \4426 );
not \U$4085 ( \4428 , \4427 );
xor \U$4086 ( \4429 , \4134 , \4076 );
not \U$4087 ( \4430 , \4429 );
or \U$4088 ( \4431 , \4428 , \4430 );
or \U$4089 ( \4432 , \4427 , \4429 );
nand \U$4090 ( \4433 , \4431 , \4432 );
not \U$4091 ( \4434 , \4433 );
or \U$4092 ( \4435 , \4337 , \4434 );
not \U$4093 ( \4436 , \4427 );
nand \U$4094 ( \4437 , \4436 , \4429 );
nand \U$4095 ( \4438 , \4435 , \4437 );
buf \U$4096 ( \4439 , \4438 );
xor \U$4097 ( \4440 , \3955 , \3964 );
xor \U$4098 ( \4441 , \4440 , \3973 );
and \U$4099 ( \4442 , \4416 , \4423 );
and \U$4100 ( \4443 , \4106 , \4411 );
nor \U$4101 ( \4444 , \4442 , \4443 );
not \U$4102 ( \4445 , \4444 );
and \U$4103 ( \4446 , \4441 , \4445 );
not \U$4104 ( \4447 , \4441 );
and \U$4105 ( \4448 , \4447 , \4444 );
nor \U$4106 ( \4449 , \4446 , \4448 );
not \U$4107 ( \4450 , \4449 );
not \U$4108 ( \4451 , \1323 );
not \U$4109 ( \4452 , \4048 );
or \U$4110 ( \4453 , \4451 , \4452 );
not \U$4111 ( \4454 , \1369 );
not \U$4112 ( \4455 , \4454 );
and \U$4113 ( \4456 , RI9871b18_134, \4455 );
not \U$4114 ( \4457 , RI9871b18_134);
and \U$4115 ( \4458 , \4457 , \3365 );
nor \U$4116 ( \4459 , \4456 , \4458 );
not \U$4117 ( \4460 , \4459 );
nand \U$4118 ( \4461 , \4460 , \1292 );
nand \U$4119 ( \4462 , \4453 , \4461 );
buf \U$4120 ( \4463 , \3556 );
not \U$4121 ( \4464 , \4463 );
nand \U$4122 ( \4465 , \414 , \419 );
not \U$4123 ( \4466 , \4465 );
and \U$4124 ( \4467 , \4464 , \4466 );
and \U$4125 ( \4468 , \4463 , \4465 );
nor \U$4126 ( \4469 , \4467 , \4468 );
buf \U$4127 ( \4470 , \4469 );
buf \U$4128 ( \4471 , \4470 );
not \U$4129 ( \4472 , \4471 );
and \U$4130 ( \4473 , \4472 , \1165 );
xnor \U$4131 ( \4474 , \4462 , \4473 );
not \U$4132 ( \4475 , \4474 );
and \U$4133 ( \4476 , \4298 , \1431 );
and \U$4134 ( \4477 , \1257 , \1619 );
and \U$4135 ( \4478 , \1659 , RI9871c08_136);
nor \U$4136 ( \4479 , \4477 , \4478 );
and \U$4137 ( \4480 , \4479 , \1456 );
nor \U$4138 ( \4481 , \4476 , \4480 );
not \U$4139 ( \4482 , \4481 );
and \U$4140 ( \4483 , \4475 , \4482 );
and \U$4141 ( \4484 , \4462 , \4473 );
nor \U$4142 ( \4485 , \4483 , \4484 );
not \U$4143 ( \4486 , \4485 );
not \U$4144 ( \4487 , \1518 );
not \U$4145 ( \4488 , \4112 );
not \U$4146 ( \4489 , \4488 );
or \U$4147 ( \4490 , \4487 , \4489 );
and \U$4148 ( \4491 , RI9871c80_137, \1595 );
not \U$4149 ( \4492 , RI9871c80_137);
and \U$4150 ( \4493 , \4492 , \1041 );
nor \U$4151 ( \4494 , \4491 , \4493 );
nand \U$4152 ( \4495 , \4494 , \1501 );
nand \U$4153 ( \4496 , \4490 , \4495 );
not \U$4154 ( \4497 , \2087 );
not \U$4155 ( \4498 , \4056 );
or \U$4156 ( \4499 , \4497 , \4498 );
and \U$4157 ( \4500 , RI9871aa0_133, \1838 );
not \U$4158 ( \4501 , RI9871aa0_133);
and \U$4159 ( \4502 , \4501 , \1275 );
nor \U$4160 ( \4503 , \4500 , \4502 );
or \U$4161 ( \4504 , \4503 , \2073 );
nand \U$4162 ( \4505 , \4499 , \4504 );
xor \U$4163 ( \4506 , \4496 , \4505 );
or \U$4164 ( \4507 , \4120 , \1470 );
and \U$4165 ( \4508 , \919 , \3969 );
not \U$4166 ( \4509 , \919 );
and \U$4167 ( \4510 , \4509 , \1191 );
nor \U$4168 ( \4511 , \4508 , \4510 );
or \U$4169 ( \4512 , \4511 , \1942 );
nand \U$4170 ( \4513 , \4507 , \4512 );
and \U$4171 ( \4514 , \4506 , \4513 );
and \U$4172 ( \4515 , \4496 , \4505 );
or \U$4173 ( \4516 , \4514 , \4515 );
not \U$4174 ( \4517 , \4516 );
not \U$4175 ( \4518 , \4103 );
not \U$4176 ( \4519 , \4088 );
not \U$4177 ( \4520 , \2982 );
or \U$4178 ( \4521 , \4519 , \4520 );
or \U$4179 ( \4522 , \1394 , \4088 );
nand \U$4180 ( \4523 , \4521 , \4522 );
not \U$4181 ( \4524 , \4523 );
or \U$4182 ( \4525 , \4518 , \4524 );
nand \U$4183 ( \4526 , \4094 , \4085 );
nand \U$4184 ( \4527 , \4525 , \4526 );
not \U$4185 ( \4528 , \4527 );
not \U$4186 ( \4529 , \4528 );
nand \U$4187 ( \4530 , RI9872400_153, RI9872478_154);
and \U$4188 ( \4531 , \4530 , RI9872388_152);
not \U$4189 ( \4532 , \4531 );
and \U$4190 ( \4533 , \4529 , \4532 );
not \U$4191 ( \4534 , \4527 );
not \U$4192 ( \4535 , \4531 );
and \U$4193 ( \4536 , \4534 , \4535 );
and \U$4194 ( \4537 , \4527 , \4531 );
nor \U$4195 ( \4538 , \4536 , \4537 );
not \U$4196 ( \4539 , \4538 );
not \U$4197 ( \4540 , \3164 );
and \U$4198 ( \4541 , \1799 , \3154 );
not \U$4199 ( \4542 , \1799 );
and \U$4200 ( \4543 , \4542 , RI9872310_151);
nor \U$4201 ( \4544 , \4541 , \4543 );
not \U$4202 ( \4545 , \4544 );
or \U$4203 ( \4546 , \4540 , \4545 );
nand \U$4204 ( \4547 , \4258 , \3170 );
nand \U$4205 ( \4548 , \4546 , \4547 );
and \U$4206 ( \4549 , \4539 , \4548 );
nor \U$4207 ( \4550 , \4533 , \4549 );
nand \U$4208 ( \4551 , \4517 , \4550 );
nand \U$4209 ( \4552 , \4486 , \4551 );
not \U$4210 ( \4553 , \4550 );
nand \U$4211 ( \4554 , \4553 , \4516 );
and \U$4212 ( \4555 , \4552 , \4554 );
not \U$4213 ( \4556 , \4555 );
not \U$4214 ( \4557 , \4556 );
or \U$4215 ( \4558 , \4450 , \4557 );
nand \U$4216 ( \4559 , \4441 , \4445 );
nand \U$4217 ( \4560 , \4558 , \4559 );
and \U$4218 ( \4561 , \4209 , \4199 );
not \U$4219 ( \4562 , \4209 );
not \U$4220 ( \4563 , \4199 );
and \U$4221 ( \4564 , \4562 , \4563 );
nor \U$4222 ( \4565 , \4561 , \4564 );
xor \U$4223 ( \4566 , \4560 , \4565 );
and \U$4224 ( \4567 , \4439 , \4566 );
and \U$4225 ( \4568 , \4560 , \4565 );
nor \U$4226 ( \4569 , \4567 , \4568 );
not \U$4227 ( \4570 , \4321 );
not \U$4228 ( \4571 , \4570 );
not \U$4229 ( \4572 , \4319 );
or \U$4230 ( \4573 , \4571 , \4572 );
or \U$4231 ( \4574 , \4570 , \4319 );
nand \U$4232 ( \4575 , \4573 , \4574 );
not \U$4233 ( \4576 , \4575 );
and \U$4234 ( \4577 , \4449 , \4556 );
not \U$4235 ( \4578 , \4449 );
and \U$4236 ( \4579 , \4578 , \4555 );
nor \U$4237 ( \4580 , \4577 , \4579 );
not \U$4238 ( \4581 , \4580 );
xor \U$4239 ( \4582 , \4053 , \4071 );
xor \U$4240 ( \4583 , \4582 , \4061 );
xor \U$4241 ( \4584 , \4114 , \4122 );
xor \U$4242 ( \4585 , \4584 , \4127 );
or \U$4243 ( \4586 , \4583 , \4585 );
not \U$4244 ( \4587 , \4586 );
xnor \U$4245 ( \4588 , \4296 , \4302 );
or \U$4246 ( \4589 , \4587 , \4588 );
nand \U$4247 ( \4590 , \4583 , \4585 );
nand \U$4248 ( \4591 , \4589 , \4590 );
xor \U$4249 ( \4592 , \4194 , \4190 );
xor \U$4250 ( \4593 , \4592 , \4193 );
xor \U$4251 ( \4594 , \4591 , \4593 );
not \U$4252 ( \4595 , \4594 );
or \U$4253 ( \4596 , \4581 , \4595 );
nand \U$4254 ( \4597 , \4593 , \4591 );
nand \U$4255 ( \4598 , \4596 , \4597 );
not \U$4256 ( \4599 , \4598 );
not \U$4257 ( \4600 , \4599 );
or \U$4258 ( \4601 , \4576 , \4600 );
or \U$4259 ( \4602 , \4599 , \4575 );
nand \U$4260 ( \4603 , \4601 , \4602 );
not \U$4261 ( \4604 , \4603 );
not \U$4262 ( \4605 , \4438 );
not \U$4263 ( \4606 , \4566 );
not \U$4264 ( \4607 , \4606 );
or \U$4265 ( \4608 , \4605 , \4607 );
not \U$4266 ( \4609 , \4438 );
nand \U$4267 ( \4610 , \4609 , \4566 );
nand \U$4268 ( \4611 , \4608 , \4610 );
not \U$4269 ( \4612 , \4611 );
or \U$4270 ( \4613 , \4604 , \4612 );
nand \U$4271 ( \4614 , \4575 , \4598 );
nand \U$4272 ( \4615 , \4613 , \4614 );
xnor \U$4273 ( \4616 , \4569 , \4615 );
not \U$4274 ( \4617 , \4616 );
or \U$4275 ( \4618 , \4335 , \4617 );
not \U$4276 ( \4619 , \4569 );
buf \U$4277 ( \4620 , \4615 );
nand \U$4278 ( \4621 , \4619 , \4620 );
nand \U$4279 ( \4622 , \4618 , \4621 );
not \U$4280 ( \4623 , \4622 );
xor \U$4281 ( \4624 , \3994 , \3822 );
not \U$4282 ( \4625 , \4624 );
not \U$4283 ( \4626 , \4329 );
not \U$4284 ( \4627 , \4215 );
or \U$4285 ( \4628 , \4626 , \4627 );
not \U$4286 ( \4629 , \4246 );
nand \U$4287 ( \4630 , \4629 , \4325 );
nand \U$4288 ( \4631 , \4628 , \4630 );
not \U$4289 ( \4632 , \4631 );
not \U$4290 ( \4633 , \4632 );
or \U$4291 ( \4634 , \4625 , \4633 );
not \U$4292 ( \4635 , \4624 );
nand \U$4293 ( \4636 , \4635 , \4631 );
nand \U$4294 ( \4637 , \4634 , \4636 );
not \U$4295 ( \4638 , \4637 );
not \U$4296 ( \4639 , \4214 );
nand \U$4297 ( \4640 , \4639 , \4150 );
not \U$4298 ( \4641 , \4640 );
not \U$4299 ( \4642 , \4151 );
or \U$4300 ( \4643 , \4641 , \4642 );
not \U$4301 ( \4644 , \4150 );
nand \U$4302 ( \4645 , \4644 , \4214 );
nand \U$4303 ( \4646 , \4643 , \4645 );
not \U$4304 ( \4647 , \3644 );
not \U$4305 ( \4648 , \4647 );
not \U$4306 ( \4649 , \3519 );
or \U$4307 ( \4650 , \4648 , \4649 );
nand \U$4308 ( \4651 , \3644 , \3518 );
nand \U$4309 ( \4652 , \4650 , \4651 );
not \U$4310 ( \4653 , \4242 );
not \U$4311 ( \4654 , \4239 );
not \U$4312 ( \4655 , \4654 );
or \U$4313 ( \4656 , \4653 , \4655 );
not \U$4314 ( \4657 , \4235 );
nand \U$4315 ( \4658 , \4657 , \4216 );
nand \U$4316 ( \4659 , \4656 , \4658 );
xor \U$4317 ( \4660 , \4652 , \4659 );
buf \U$4318 ( \4661 , \4660 );
xor \U$4319 ( \4662 , \4646 , \4661 );
not \U$4320 ( \4663 , \4662 );
not \U$4321 ( \4664 , \4663 );
and \U$4322 ( \4665 , \4638 , \4664 );
and \U$4323 ( \4666 , \4637 , \4663 );
nor \U$4324 ( \4667 , \4665 , \4666 );
and \U$4325 ( \4668 , \4623 , \4667 );
not \U$4326 ( \4669 , \4637 );
not \U$4327 ( \4670 , \4662 );
or \U$4328 ( \4671 , \4669 , \4670 );
nand \U$4329 ( \4672 , \4631 , \4624 );
nand \U$4330 ( \4673 , \4671 , \4672 );
not \U$4331 ( \4674 , \3762 );
not \U$4332 ( \4675 , \3649 );
not \U$4333 ( \4676 , \4675 );
and \U$4334 ( \4677 , \4674 , \4676 );
and \U$4335 ( \4678 , \3762 , \4675 );
nor \U$4336 ( \4679 , \4677 , \4678 );
not \U$4337 ( \4680 , \4646 );
not \U$4338 ( \4681 , \4660 );
or \U$4339 ( \4682 , \4680 , \4681 );
nand \U$4340 ( \4683 , \4652 , \4659 );
nand \U$4341 ( \4684 , \4682 , \4683 );
xor \U$4342 ( \4685 , \4679 , \4684 );
xor \U$4343 ( \4686 , \4007 , \3999 );
xnor \U$4344 ( \4687 , \4686 , \4015 );
xor \U$4345 ( \4688 , \4685 , \4687 );
nor \U$4346 ( \4689 , \4673 , \4688 );
nor \U$4347 ( \4690 , \4668 , \4689 );
not \U$4348 ( \4691 , \4018 );
not \U$4349 ( \4692 , \4024 );
and \U$4350 ( \4693 , \4691 , \4692 );
and \U$4351 ( \4694 , \4018 , \4024 );
nor \U$4352 ( \4695 , \4693 , \4694 );
nand \U$4353 ( \4696 , \4687 , \4679 );
and \U$4354 ( \4697 , \4696 , \4684 );
nor \U$4355 ( \4698 , \4687 , \4679 );
nor \U$4356 ( \4699 , \4697 , \4698 );
nand \U$4357 ( \4700 , \4695 , \4699 );
xor \U$4358 ( \4701 , \4594 , \4580 );
xnor \U$4359 ( \4702 , \4474 , \4481 );
not \U$4360 ( \4703 , \4702 );
not \U$4361 ( \4704 , \4703 );
xor \U$4362 ( \4705 , \4538 , \4548 );
not \U$4363 ( \4706 , \4705 );
not \U$4364 ( \4707 , \1162 );
not \U$4365 ( \4708 , \1716 );
and \U$4366 ( \4709 , \4471 , \4708 );
not \U$4367 ( \4710 , \4469 );
not \U$4368 ( \4711 , \4710 );
not \U$4369 ( \4712 , \4711 );
and \U$4370 ( \4713 , \4712 , \1199 );
nor \U$4371 ( \4714 , \4709 , \4713 );
not \U$4372 ( \4715 , \4714 );
not \U$4373 ( \4716 , \4715 );
or \U$4374 ( \4717 , \4707 , \4716 );
and \U$4375 ( \4718 , \4410 , \1165 );
and \U$4376 ( \4719 , \4409 , \1199 );
nor \U$4377 ( \4720 , \4718 , \4719 );
or \U$4378 ( \4721 , \1719 , \4720 );
nand \U$4379 ( \4722 , \4717 , \4721 );
not \U$4380 ( \4723 , \4722 );
not \U$4381 ( \4724 , \1018 );
not \U$4382 ( \4725 , \1045 );
not \U$4383 ( \4726 , \4177 );
or \U$4384 ( \4727 , \4725 , \4726 );
or \U$4385 ( \4728 , \4177 , \1045 );
nand \U$4386 ( \4729 , \4727 , \4728 );
not \U$4387 ( \4730 , \4729 );
or \U$4388 ( \4731 , \4724 , \4730 );
or \U$4389 ( \4732 , \4379 , \1068 );
nand \U$4390 ( \4733 , \4731 , \4732 );
not \U$4391 ( \4734 , \4733 );
not \U$4392 ( \4735 , \1136 );
not \U$4393 ( \4736 , \4386 );
or \U$4394 ( \4737 , \4735 , \4736 );
not \U$4395 ( \4738 , \1550 );
not \U$4396 ( \4739 , \1111 );
and \U$4397 ( \4740 , \4738 , \4739 );
and \U$4398 ( \4741 , \3836 , \1111 );
nor \U$4399 ( \4742 , \4740 , \4741 );
not \U$4400 ( \4743 , \4742 );
nand \U$4401 ( \4744 , \4743 , \1083 );
nand \U$4402 ( \4745 , \4737 , \4744 );
not \U$4403 ( \4746 , \4745 );
not \U$4404 ( \4747 , \4746 );
or \U$4405 ( \4748 , \4734 , \4747 );
or \U$4406 ( \4749 , \4746 , \4733 );
nand \U$4407 ( \4750 , \4748 , \4749 );
not \U$4408 ( \4751 , \4750 );
or \U$4409 ( \4752 , \4723 , \4751 );
nand \U$4410 ( \4753 , \4745 , \4733 );
nand \U$4411 ( \4754 , \4752 , \4753 );
not \U$4412 ( \4755 , \4754 );
or \U$4413 ( \4756 , \4706 , \4755 );
or \U$4414 ( \4757 , \4754 , \4705 );
nand \U$4415 ( \4758 , \4756 , \4757 );
not \U$4416 ( \4759 , \4758 );
or \U$4417 ( \4760 , \4704 , \4759 );
not \U$4418 ( \4761 , \4705 );
nand \U$4419 ( \4762 , \4761 , \4754 );
nand \U$4420 ( \4763 , \4760 , \4762 );
not \U$4421 ( \4764 , \4763 );
not \U$4422 ( \4765 , \4588 );
nand \U$4423 ( \4766 , \4586 , \4590 );
not \U$4424 ( \4767 , \4766 );
or \U$4425 ( \4768 , \4765 , \4767 );
or \U$4426 ( \4769 , \4766 , \4588 );
nand \U$4427 ( \4770 , \4768 , \4769 );
not \U$4428 ( \4771 , \4770 );
not \U$4429 ( \4772 , \4771 );
or \U$4430 ( \4773 , \4764 , \4772 );
not \U$4431 ( \4774 , \4085 );
and \U$4432 ( \4775 , RI98725e0_157, \2605 );
not \U$4433 ( \4776 , RI98725e0_157);
and \U$4434 ( \4777 , \4776 , \1725 );
nor \U$4435 ( \4778 , \4775 , \4777 );
not \U$4436 ( \4779 , \4778 );
or \U$4437 ( \4780 , \4774 , \4779 );
and \U$4438 ( \4781 , \1098 , \4088 );
not \U$4439 ( \4782 , \1098 );
and \U$4440 ( \4783 , \4782 , RI98725e0_157);
nor \U$4441 ( \4784 , \4781 , \4783 );
nand \U$4442 ( \4785 , \4784 , \4103 );
nand \U$4443 ( \4786 , \4780 , \4785 );
not \U$4444 ( \4787 , \2074 );
and \U$4445 ( \4788 , RI9871aa0_133, \895 );
not \U$4446 ( \4789 , RI9871aa0_133);
and \U$4447 ( \4790 , \4789 , \1506 );
nor \U$4448 ( \4791 , \4788 , \4790 );
not \U$4449 ( \4792 , \4791 );
or \U$4450 ( \4793 , \4787 , \4792 );
and \U$4451 ( \4794 , RI9871aa0_133, \918 );
not \U$4452 ( \4795 , RI9871aa0_133);
and \U$4453 ( \4796 , \4795 , \1513 );
nor \U$4454 ( \4797 , \4794 , \4796 );
not \U$4455 ( \4798 , \4797 );
nand \U$4456 ( \4799 , \4798 , \2087 );
nand \U$4457 ( \4800 , \4793 , \4799 );
xor \U$4458 ( \4801 , \4786 , \4800 );
not \U$4459 ( \4802 , \1501 );
and \U$4460 ( \4803 , \1584 , \1191 );
not \U$4461 ( \4804 , \1584 );
and \U$4462 ( \4805 , \4804 , \3969 );
nor \U$4463 ( \4806 , \4803 , \4805 );
not \U$4464 ( \4807 , \4806 );
or \U$4465 ( \4808 , \4802 , \4807 );
xor \U$4466 ( \4809 , \1212 , RI9871c80_137);
nand \U$4467 ( \4810 , \4809 , \1518 );
nand \U$4468 ( \4811 , \4808 , \4810 );
and \U$4469 ( \4812 , \4801 , \4811 );
and \U$4470 ( \4813 , \4786 , \4800 );
nor \U$4471 ( \4814 , \4812 , \4813 );
not \U$4472 ( \4815 , \4814 );
not \U$4473 ( \4816 , \4815 );
and \U$4474 ( \4817 , RI9871d70_139, \3691 );
not \U$4475 ( \4818 , RI9871d70_139);
and \U$4476 ( \4819 , \4818 , \3693 );
nor \U$4477 ( \4820 , \4817 , \4819 );
or \U$4478 ( \4821 , \4820 , \932 );
and \U$4479 ( \4822 , RI9871d70_139, \3861 );
not \U$4480 ( \4823 , RI9871d70_139);
and \U$4481 ( \4824 , \4823 , \3240 );
nor \U$4482 ( \4825 , \4822 , \4824 );
or \U$4483 ( \4826 , \4825 , \860 );
nand \U$4484 ( \4827 , \4821 , \4826 );
xnor \U$4485 ( \4828 , \3275 , RI9872130_147);
or \U$4486 ( \4829 , \4828 , \1470 );
and \U$4487 ( \4830 , \2111 , \919 );
not \U$4488 ( \4831 , \2111 );
and \U$4489 ( \4832 , \4831 , RI9872130_147);
nor \U$4490 ( \4833 , \4830 , \4832 );
or \U$4491 ( \4834 , \4833 , \1942 );
nand \U$4492 ( \4835 , \4829 , \4834 );
xor \U$4493 ( \4836 , \4827 , \4835 );
not \U$4494 ( \4837 , \794 );
and \U$4495 ( \4838 , RI98719b0_131, \847 );
not \U$4496 ( \4839 , RI98719b0_131);
and \U$4497 ( \4840 , \4839 , \2216 );
nor \U$4498 ( \4841 , \4838 , \4840 );
not \U$4499 ( \4842 , \4841 );
or \U$4500 ( \4843 , \4837 , \4842 );
and \U$4501 ( \4844 , RI98719b0_131, \824 );
not \U$4502 ( \4845 , RI98719b0_131);
and \U$4503 ( \4846 , \4845 , \821 );
nor \U$4504 ( \4847 , \4844 , \4846 );
or \U$4505 ( \4848 , \4847 , \3244 );
nand \U$4506 ( \4849 , \4843 , \4848 );
and \U$4507 ( \4850 , \4836 , \4849 );
and \U$4508 ( \4851 , \4827 , \4835 );
or \U$4509 ( \4852 , \4850 , \4851 );
not \U$4510 ( \4853 , \4852 );
not \U$4511 ( \4854 , \1455 );
xor \U$4512 ( \4855 , \1371 , RI9871c08_136);
not \U$4513 ( \4856 , \4855 );
or \U$4514 ( \4857 , \4854 , \4856 );
and \U$4515 ( \4858 , \1949 , RI9871c08_136);
not \U$4516 ( \4859 , \1949 );
and \U$4517 ( \4860 , \4859 , \1850 );
nor \U$4518 ( \4861 , \4858 , \4860 );
nand \U$4519 ( \4862 , \4861 , \1431 );
nand \U$4520 ( \4863 , \4857 , \4862 );
not \U$4521 ( \4864 , \3164 );
and \U$4522 ( \4865 , RI9872310_151, \1838 );
not \U$4523 ( \4866 , RI9872310_151);
and \U$4524 ( \4867 , \4866 , \1275 );
or \U$4525 ( \4868 , \4865 , \4867 );
not \U$4526 ( \4869 , \4868 );
or \U$4527 ( \4870 , \4864 , \4869 );
and \U$4528 ( \4871 , \2038 , \3154 );
not \U$4529 ( \4872 , \2038 );
and \U$4530 ( \4873 , \4872 , RI9872310_151);
nor \U$4531 ( \4874 , \4871 , \4873 );
nand \U$4532 ( \4875 , \4874 , \3170 );
nand \U$4533 ( \4876 , \4870 , \4875 );
xor \U$4534 ( \4877 , \4863 , \4876 );
and \U$4535 ( \4878 , \2842 , RI9871b18_134);
and \U$4536 ( \4879 , \1062 , \2479 );
nor \U$4537 ( \4880 , \4878 , \4879 );
or \U$4538 ( \4881 , \4880 , \1543 );
not \U$4539 ( \4882 , \1041 );
not \U$4540 ( \4883 , RI9871b18_134);
and \U$4541 ( \4884 , \4882 , \4883 );
and \U$4542 ( \4885 , \1041 , RI9871b18_134);
nor \U$4543 ( \4886 , \4884 , \4885 );
or \U$4544 ( \4887 , \4886 , \1293 );
nand \U$4545 ( \4888 , \4881 , \4887 );
and \U$4546 ( \4889 , \4877 , \4888 );
and \U$4547 ( \4890 , \4863 , \4876 );
nor \U$4548 ( \4891 , \4889 , \4890 );
not \U$4549 ( \4892 , \4891 );
or \U$4550 ( \4893 , \4853 , \4892 );
or \U$4551 ( \4894 , \4852 , \4891 );
nand \U$4552 ( \4895 , \4893 , \4894 );
not \U$4553 ( \4896 , \4895 );
or \U$4554 ( \4897 , \4816 , \4896 );
not \U$4555 ( \4898 , \4891 );
nand \U$4556 ( \4899 , \4898 , \4852 );
nand \U$4557 ( \4900 , \4897 , \4899 );
not \U$4558 ( \4901 , \4900 );
not \U$4559 ( \4902 , RI9872388_152);
not \U$4560 ( \4903 , \4902 );
not \U$4561 ( \4904 , \780 );
or \U$4562 ( \4905 , \4903 , \4904 );
or \U$4563 ( \4906 , \780 , \4902 );
nand \U$4564 ( \4907 , \4905 , \4906 );
not \U$4565 ( \4908 , RI9872400_153);
and \U$4566 ( \4909 , \4902 , \4908 );
and \U$4567 ( \4910 , RI9872388_152, RI9872400_153);
and \U$4568 ( \4911 , RI9872478_154, \4908 );
not \U$4569 ( \4912 , RI9872478_154);
and \U$4570 ( \4913 , \4912 , RI9872400_153);
or \U$4571 ( \4914 , \4911 , \4913 );
nor \U$4572 ( \4915 , \4909 , \4910 , \4914 );
buf \U$4573 ( \4916 , \4915 );
not \U$4574 ( \4917 , \4916 );
not \U$4575 ( \4918 , \4917 );
buf \U$4576 ( \4919 , \4918 );
buf \U$4577 ( \4920 , \4919 );
and \U$4578 ( \4921 , \4907 , \4920 );
buf \U$4579 ( \4922 , \4914 );
buf \U$4580 ( \4923 , \4922 );
not \U$4581 ( \4924 , \4923 );
not \U$4582 ( \4925 , \4924 );
and \U$4583 ( \4926 , \4925 , RI9872388_152);
nor \U$4584 ( \4927 , \4921 , \4926 );
not \U$4585 ( \4928 , \4927 );
or \U$4586 ( \4929 , \4720 , \1809 );
or \U$4587 ( \4930 , \4420 , \1719 );
nand \U$4588 ( \4931 , \4929 , \4930 );
not \U$4589 ( \4932 , \4931 );
or \U$4590 ( \4933 , \4928 , \4932 );
or \U$4591 ( \4934 , \4927 , \4931 );
nand \U$4592 ( \4935 , \4933 , \4934 );
not \U$4593 ( \4936 , \4874 );
not \U$4594 ( \4937 , \4936 );
not \U$4595 ( \4938 , \3962 );
and \U$4596 ( \4939 , \4937 , \4938 );
and \U$4597 ( \4940 , \4544 , \3170 );
nor \U$4598 ( \4941 , \4939 , \4940 );
not \U$4599 ( \4942 , \4941 );
not \U$4600 ( \4943 , \4942 );
not \U$4601 ( \4944 , \405 );
not \U$4602 ( \4945 , \4944 );
not \U$4603 ( \4946 , \689 );
not \U$4604 ( \4947 , \687 );
or \U$4605 ( \4948 , \4946 , \4947 );
not \U$4606 ( \4949 , \398 );
nand \U$4607 ( \4950 , \4948 , \4949 );
not \U$4608 ( \4951 , \4950 );
or \U$4609 ( \4952 , \4945 , \4951 );
nand \U$4610 ( \4953 , \4952 , \399 );
xor \U$4611 ( \4954 , RI986e878_26, RI986e800_25);
and \U$4612 ( \4955 , \4953 , \4954 );
not \U$4613 ( \4956 , \4953 );
not \U$4614 ( \4957 , \4954 );
and \U$4615 ( \4958 , \4956 , \4957 );
nor \U$4616 ( \4959 , \4955 , \4958 );
buf \U$4617 ( \4960 , \4959 );
nand \U$4618 ( \4961 , \4960 , \1165 );
not \U$4619 ( \4962 , \4961 );
not \U$4620 ( \4963 , \4103 );
not \U$4621 ( \4964 , \4778 );
or \U$4622 ( \4965 , \4963 , \4964 );
nand \U$4623 ( \4966 , \4523 , \4085 );
nand \U$4624 ( \4967 , \4965 , \4966 );
not \U$4625 ( \4968 , \4967 );
or \U$4626 ( \4969 , \4962 , \4968 );
or \U$4627 ( \4970 , \4967 , \4961 );
nand \U$4628 ( \4971 , \4969 , \4970 );
not \U$4629 ( \4972 , \4971 );
or \U$4630 ( \4973 , \4943 , \4972 );
not \U$4631 ( \4974 , \4961 );
nand \U$4632 ( \4975 , \4974 , \4967 );
nand \U$4633 ( \4976 , \4973 , \4975 );
xor \U$4634 ( \4977 , \4935 , \4976 );
buf \U$4635 ( \4978 , \4950 );
not \U$4636 ( \4979 , \4978 );
or \U$4637 ( \4980 , \400 , \405 );
not \U$4638 ( \4981 , \4980 );
and \U$4639 ( \4982 , \4979 , \4981 );
and \U$4640 ( \4983 , \4978 , \4980 );
nor \U$4641 ( \4984 , \4982 , \4983 );
buf \U$4642 ( \4985 , \4984 );
buf \U$4643 ( \4986 , \4985 );
nor \U$4644 ( \4987 , \4986 , \1716 );
not \U$4645 ( \4988 , \4959 );
not \U$4646 ( \4989 , \4988 );
not \U$4647 ( \4990 , \4989 );
and \U$4648 ( \4991 , \1165 , \4990 );
not \U$4649 ( \4992 , \1165 );
and \U$4650 ( \4993 , \4992 , \4960 );
nor \U$4651 ( \4994 , \4991 , \4993 );
or \U$4652 ( \4995 , \4994 , \1809 );
or \U$4653 ( \4996 , \4714 , \1719 );
nand \U$4654 ( \4997 , \4995 , \4996 );
xor \U$4655 ( \4998 , \4987 , \4997 );
or \U$4656 ( \4999 , \4742 , \1137 );
and \U$4657 ( \5000 , \1257 , RI98718c0_129);
and \U$4658 ( \5001 , \1254 , \1111 );
nor \U$4659 ( \5002 , \5000 , \5001 );
or \U$4660 ( \5003 , \5002 , \1676 );
nand \U$4661 ( \5004 , \4999 , \5003 );
and \U$4662 ( \5005 , \4998 , \5004 );
and \U$4663 ( \5006 , \4987 , \4997 );
nor \U$4664 ( \5007 , \5005 , \5006 );
not \U$4665 ( \5008 , \5007 );
not \U$4666 ( \5009 , \5008 );
not \U$4667 ( \5010 , \3466 );
and \U$4668 ( \5011 , \4063 , \2492 );
not \U$4669 ( \5012 , \4063 );
not \U$4670 ( \5013 , \1799 );
and \U$4671 ( \5014 , \5012 , \5013 );
nor \U$4672 ( \5015 , \5011 , \5014 );
not \U$4673 ( \5016 , \5015 );
or \U$4674 ( \5017 , \5010 , \5016 );
and \U$4675 ( \5018 , \1417 , \4063 );
not \U$4676 ( \5019 , \1417 );
and \U$4677 ( \5020 , \5019 , RI98726d0_159);
nor \U$4678 ( \5021 , \5018 , \5020 );
or \U$4679 ( \5022 , \5021 , \3591 );
nand \U$4680 ( \5023 , \5017 , \5022 );
not \U$4681 ( \5024 , \5023 );
not \U$4682 ( \5025 , RI9872478_154);
not \U$4683 ( \5026 , RI98724f0_155);
and \U$4684 ( \5027 , \5025 , \5026 );
and \U$4685 ( \5028 , RI9872478_154, RI98724f0_155);
and \U$4686 ( \5029 , RI9872568_156, \5026 );
not \U$4687 ( \5030 , RI9872568_156);
and \U$4688 ( \5031 , \5030 , RI98724f0_155);
or \U$4689 ( \5032 , \5029 , \5031 );
nor \U$4690 ( \5033 , \5027 , \5028 , \5032 );
buf \U$4691 ( \5034 , \5033 );
buf \U$4692 ( \5035 , \5032 );
buf \U$4693 ( \5036 , \5035 );
or \U$4694 ( \5037 , \5034 , \5036 );
nand \U$4695 ( \5038 , \5037 , RI9872478_154);
not \U$4696 ( \5039 , \4920 );
not \U$4697 ( \5040 , \4902 );
not \U$4698 ( \5041 , \1393 );
or \U$4699 ( \5042 , \5040 , \5041 );
or \U$4700 ( \5043 , \1394 , \4902 );
nand \U$4701 ( \5044 , \5042 , \5043 );
not \U$4702 ( \5045 , \5044 );
or \U$4703 ( \5046 , \5039 , \5045 );
buf \U$4704 ( \5047 , \4923 );
buf \U$4705 ( \5048 , \5047 );
nand \U$4706 ( \5049 , \4907 , \5048 );
nand \U$4707 ( \5050 , \5046 , \5049 );
xor \U$4708 ( \5051 , \5038 , \5050 );
not \U$4709 ( \5052 , \5051 );
or \U$4710 ( \5053 , \5024 , \5052 );
nand \U$4711 ( \5054 , \5050 , \5038 );
nand \U$4712 ( \5055 , \5053 , \5054 );
or \U$4713 ( \5056 , \4927 , \5055 );
not \U$4714 ( \5057 , \5056 );
or \U$4715 ( \5058 , \5009 , \5057 );
nand \U$4716 ( \5059 , \5055 , \4927 );
nand \U$4717 ( \5060 , \5058 , \5059 );
xor \U$4718 ( \5061 , \4977 , \5060 );
not \U$4719 ( \5062 , \5061 );
or \U$4720 ( \5063 , \4901 , \5062 );
nand \U$4721 ( \5064 , \5060 , \4977 );
nand \U$4722 ( \5065 , \5063 , \5064 );
not \U$4723 ( \5066 , \4763 );
nand \U$4724 ( \5067 , \5066 , \4770 );
nand \U$4725 ( \5068 , \5065 , \5067 );
nand \U$4726 ( \5069 , \4773 , \5068 );
xor \U$4727 ( \5070 , \4701 , \5069 );
not \U$4728 ( \5071 , \1353 );
not \U$4729 ( \5072 , \4371 );
or \U$4730 ( \5073 , \5071 , \5072 );
and \U$4731 ( \5074 , \1367 , \3537 );
not \U$4732 ( \5075 , \1367 );
and \U$4733 ( \5076 , \5075 , \3542 );
nor \U$4734 ( \5077 , \5074 , \5076 );
not \U$4735 ( \5078 , \1381 );
or \U$4736 ( \5079 , \5077 , \5078 );
nand \U$4737 ( \5080 , \5073 , \5079 );
not \U$4738 ( \5081 , \5080 );
or \U$4739 ( \5082 , \4342 , \932 );
or \U$4740 ( \5083 , \4820 , \860 );
nand \U$4741 ( \5084 , \5082 , \5083 );
not \U$4742 ( \5085 , \5084 );
not \U$4743 ( \5086 , \5085 );
not \U$4744 ( \5087 , \797 );
not \U$4745 ( \5088 , \4359 );
or \U$4746 ( \5089 , \5087 , \5088 );
not \U$4747 ( \5090 , \4847 );
nand \U$4748 ( \5091 , \5090 , \793 );
nand \U$4749 ( \5092 , \5089 , \5091 );
not \U$4750 ( \5093 , \5092 );
or \U$4751 ( \5094 , \5086 , \5093 );
or \U$4752 ( \5095 , \5092 , \5085 );
nand \U$4753 ( \5096 , \5094 , \5095 );
not \U$4754 ( \5097 , \5096 );
or \U$4755 ( \5098 , \5081 , \5097 );
nand \U$4756 ( \5099 , \5092 , \5084 );
nand \U$4757 ( \5100 , \5098 , \5099 );
not \U$4758 ( \5101 , \5100 );
not \U$4759 ( \5102 , \1518 );
not \U$4760 ( \5103 , \4494 );
or \U$4761 ( \5104 , \5102 , \5103 );
nand \U$4762 ( \5105 , \4809 , \1501 );
nand \U$4763 ( \5106 , \5104 , \5105 );
not \U$4764 ( \5107 , \5106 );
not \U$4765 ( \5108 , \5021 );
nand \U$4766 ( \5109 , \5108 , \3466 );
nand \U$4767 ( \5110 , \4351 , \3467 );
and \U$4768 ( \5111 , \5109 , \5110 );
not \U$4769 ( \5112 , \5111 );
or \U$4770 ( \5113 , \5107 , \5112 );
or \U$4771 ( \5114 , \5111 , \5106 );
nand \U$4772 ( \5115 , \5113 , \5114 );
or \U$4773 ( \5116 , \4511 , \1470 );
or \U$4774 ( \5117 , \4828 , \1942 );
nand \U$4775 ( \5118 , \5116 , \5117 );
nand \U$4776 ( \5119 , \5115 , \5118 );
not \U$4777 ( \5120 , \5111 );
nand \U$4778 ( \5121 , \5120 , \5106 );
and \U$4779 ( \5122 , \5119 , \5121 );
or \U$4780 ( \5123 , \4459 , \1543 );
or \U$4781 ( \5124 , \4880 , \1293 );
nand \U$4782 ( \5125 , \5123 , \5124 );
or \U$4783 ( \5126 , \4503 , \2086 );
or \U$4784 ( \5127 , \4797 , \2073 );
nand \U$4785 ( \5128 , \5126 , \5127 );
xor \U$4786 ( \5129 , \5125 , \5128 );
and \U$4787 ( \5130 , \4479 , \1431 );
and \U$4788 ( \5131 , \4861 , \1456 );
nor \U$4789 ( \5132 , \5130 , \5131 );
not \U$4790 ( \5133 , \5132 );
and \U$4791 ( \5134 , \5129 , \5133 );
and \U$4792 ( \5135 , \5125 , \5128 );
nor \U$4793 ( \5136 , \5134 , \5135 );
and \U$4794 ( \5137 , \5122 , \5136 );
not \U$4795 ( \5138 , \5122 );
not \U$4796 ( \5139 , \5136 );
and \U$4797 ( \5140 , \5138 , \5139 );
nor \U$4798 ( \5141 , \5137 , \5140 );
not \U$4799 ( \5142 , \5141 );
or \U$4800 ( \5143 , \5101 , \5142 );
not \U$4801 ( \5144 , \5122 );
nand \U$4802 ( \5145 , \5144 , \5139 );
nand \U$4803 ( \5146 , \5143 , \5145 );
not \U$4804 ( \5147 , \5146 );
not \U$4805 ( \5148 , \4935 );
not \U$4806 ( \5149 , \4976 );
or \U$4807 ( \5150 , \5148 , \5149 );
not \U$4808 ( \5151 , \4927 );
nand \U$4809 ( \5152 , \5151 , \4931 );
nand \U$4810 ( \5153 , \5150 , \5152 );
xor \U$4811 ( \5154 , \4263 , \4270 );
xor \U$4812 ( \5155 , \5154 , \4276 );
xnor \U$4813 ( \5156 , \5153 , \5155 );
not \U$4814 ( \5157 , \5156 );
or \U$4815 ( \5158 , \5147 , \5157 );
or \U$4816 ( \5159 , \5156 , \5146 );
nand \U$4817 ( \5160 , \5158 , \5159 );
xor \U$4818 ( \5161 , \4383 , \4391 );
xor \U$4819 ( \5162 , \4344 , \4353 );
xor \U$4820 ( \5163 , \5162 , \4364 );
xor \U$4821 ( \5164 , \5161 , \5163 );
xor \U$4822 ( \5165 , \4496 , \4505 );
xor \U$4823 ( \5166 , \5165 , \4513 );
and \U$4824 ( \5167 , \5164 , \5166 );
and \U$4825 ( \5168 , \5161 , \5163 );
or \U$4826 ( \5169 , \5167 , \5168 );
xor \U$4827 ( \5170 , \4485 , \4516 );
xor \U$4828 ( \5171 , \5170 , \4550 );
xor \U$4829 ( \5172 , \5169 , \5171 );
xor \U$4830 ( \5173 , \4367 , \4395 );
xor \U$4831 ( \5174 , \5173 , \4424 );
xor \U$4832 ( \5175 , \5172 , \5174 );
xor \U$4833 ( \5176 , \5160 , \5175 );
xor \U$4834 ( \5177 , \5118 , \5115 );
not \U$4835 ( \5178 , \5177 );
not \U$4836 ( \5179 , \1353 );
not \U$4837 ( \5180 , \5077 );
not \U$4838 ( \5181 , \5180 );
or \U$4839 ( \5182 , \5179 , \5181 );
and \U$4840 ( \5183 , RI9871e60_141, \4154 );
not \U$4841 ( \5184 , RI9871e60_141);
and \U$4842 ( \5185 , \5184 , \4155 );
nor \U$4843 ( \5186 , \5183 , \5185 );
or \U$4844 ( \5187 , \5186 , \5078 );
nand \U$4845 ( \5188 , \5182 , \5187 );
not \U$4846 ( \5189 , \5188 );
not \U$4847 ( \5190 , \5034 );
not \U$4848 ( \5191 , \5025 );
not \U$4849 ( \5192 , \2361 );
or \U$4850 ( \5193 , \5191 , \5192 );
or \U$4851 ( \5194 , \780 , \5025 );
nand \U$4852 ( \5195 , \5193 , \5194 );
not \U$4853 ( \5196 , \5195 );
or \U$4854 ( \5197 , \5190 , \5196 );
nand \U$4855 ( \5198 , \5036 , RI9872478_154);
nand \U$4856 ( \5199 , \5197 , \5198 );
not \U$4857 ( \5200 , \5199 );
not \U$4858 ( \5201 , \5200 );
or \U$4859 ( \5202 , \5189 , \5201 );
or \U$4860 ( \5203 , \5200 , \5188 );
nand \U$4861 ( \5204 , \5202 , \5203 );
buf \U$4862 ( \5205 , \4406 );
buf \U$4863 ( \5206 , \5205 );
and \U$4864 ( \5207 , \5206 , \1044 );
not \U$4865 ( \5208 , \5205 );
and \U$4866 ( \5209 , \5208 , \1045 );
nor \U$4867 ( \5210 , \5207 , \5209 );
not \U$4868 ( \5211 , \5210 );
not \U$4869 ( \5212 , \1612 );
and \U$4870 ( \5213 , \5211 , \5212 );
and \U$4871 ( \5214 , \4729 , \1067 );
nor \U$4872 ( \5215 , \5213 , \5214 );
not \U$4873 ( \5216 , \5215 );
and \U$4874 ( \5217 , \5204 , \5216 );
and \U$4875 ( \5218 , \5199 , \5188 );
nor \U$4876 ( \5219 , \5217 , \5218 );
not \U$4877 ( \5220 , \5219 );
xor \U$4878 ( \5221 , \5080 , \5085 );
xnor \U$4879 ( \5222 , \5221 , \5092 );
not \U$4880 ( \5223 , \5222 );
or \U$4881 ( \5224 , \5220 , \5223 );
or \U$4882 ( \5225 , \5222 , \5219 );
nand \U$4883 ( \5226 , \5224 , \5225 );
not \U$4884 ( \5227 , \5226 );
or \U$4885 ( \5228 , \5178 , \5227 );
not \U$4886 ( \5229 , \5219 );
nand \U$4887 ( \5230 , \5229 , \5222 );
nand \U$4888 ( \5231 , \5228 , \5230 );
not \U$4889 ( \5232 , \5141 );
not \U$4890 ( \5233 , \5100 );
not \U$4891 ( \5234 , \5233 );
and \U$4892 ( \5235 , \5232 , \5234 );
and \U$4893 ( \5236 , \5141 , \5233 );
nor \U$4894 ( \5237 , \5235 , \5236 );
xor \U$4895 ( \5238 , \5231 , \5237 );
and \U$4896 ( \5239 , \5129 , \5133 );
not \U$4897 ( \5240 , \5129 );
and \U$4898 ( \5241 , \5240 , \5132 );
nor \U$4899 ( \5242 , \5239 , \5241 );
not \U$4900 ( \5243 , \5242 );
not \U$4901 ( \5244 , \4722 );
not \U$4902 ( \5245 , \5244 );
not \U$4903 ( \5246 , \4750 );
or \U$4904 ( \5247 , \5245 , \5246 );
or \U$4905 ( \5248 , \5244 , \4750 );
nand \U$4906 ( \5249 , \5247 , \5248 );
not \U$4907 ( \5250 , \4971 );
not \U$4908 ( \5251 , \4941 );
and \U$4909 ( \5252 , \5250 , \5251 );
and \U$4910 ( \5253 , \4971 , \4941 );
nor \U$4911 ( \5254 , \5252 , \5253 );
xnor \U$4912 ( \5255 , \5249 , \5254 );
not \U$4913 ( \5256 , \5255 );
or \U$4914 ( \5257 , \5243 , \5256 );
not \U$4915 ( \5258 , \5254 );
nand \U$4916 ( \5259 , \5258 , \5249 );
nand \U$4917 ( \5260 , \5257 , \5259 );
not \U$4918 ( \5261 , \5260 );
or \U$4919 ( \5262 , \5238 , \5261 );
not \U$4920 ( \5263 , \5237 );
nand \U$4921 ( \5264 , \5231 , \5263 );
nand \U$4922 ( \5265 , \5262 , \5264 );
and \U$4923 ( \5266 , \5176 , \5265 );
and \U$4924 ( \5267 , \5160 , \5175 );
or \U$4925 ( \5268 , \5266 , \5267 );
and \U$4926 ( \5269 , \5070 , \5268 );
and \U$4927 ( \5270 , \4701 , \5069 );
or \U$4928 ( \5271 , \5269 , \5270 );
not \U$4929 ( \5272 , \5271 );
not \U$4930 ( \5273 , \5156 );
nand \U$4931 ( \5274 , \5273 , \5146 );
nand \U$4932 ( \5275 , \5153 , \5155 );
and \U$4933 ( \5276 , \5274 , \5275 );
not \U$4934 ( \5277 , \5276 );
xor \U$4935 ( \5278 , \4336 , \4433 );
xor \U$4936 ( \5279 , \5277 , \5278 );
xor \U$4937 ( \5280 , \5169 , \5171 );
and \U$4938 ( \5281 , \5280 , \5174 );
and \U$4939 ( \5282 , \5169 , \5171 );
or \U$4940 ( \5283 , \5281 , \5282 );
and \U$4941 ( \5284 , \5279 , \5283 );
and \U$4942 ( \5285 , \5277 , \5278 );
nor \U$4943 ( \5286 , \5284 , \5285 );
not \U$4944 ( \5287 , \5286 );
xor \U$4945 ( \5288 , \4611 , \4603 );
not \U$4946 ( \5289 , \5288 );
or \U$4947 ( \5290 , \5287 , \5289 );
or \U$4948 ( \5291 , \5288 , \5286 );
nand \U$4949 ( \5292 , \5290 , \5291 );
not \U$4950 ( \5293 , \5292 );
or \U$4951 ( \5294 , \5272 , \5293 );
not \U$4952 ( \5295 , \5286 );
nand \U$4953 ( \5296 , \5295 , \5288 );
nand \U$4954 ( \5297 , \5294 , \5296 );
not \U$4955 ( \5298 , \5297 );
xor \U$4956 ( \5299 , \4569 , \4334 );
xnor \U$4957 ( \5300 , \5299 , \4620 );
not \U$4958 ( \5301 , \5300 );
nand \U$4959 ( \5302 , \5298 , \5301 );
nand \U$4960 ( \5303 , \4690 , \4700 , \5302 );
not \U$4961 ( \5304 , \5303 );
xor \U$4962 ( \5305 , \4927 , \5007 );
xnor \U$4963 ( \5306 , \5305 , \5055 );
not \U$4964 ( \5307 , \4814 );
not \U$4965 ( \5308 , \4895 );
or \U$4966 ( \5309 , \5307 , \5308 );
or \U$4967 ( \5310 , \4814 , \4895 );
nand \U$4968 ( \5311 , \5309 , \5310 );
xor \U$4969 ( \5312 , \5306 , \5311 );
not \U$4970 ( \5313 , \4920 );
not \U$4971 ( \5314 , RI9872388_152);
not \U$4972 ( \5315 , \2399 );
or \U$4973 ( \5316 , \5314 , \5315 );
or \U$4974 ( \5317 , \1128 , RI9872388_152);
nand \U$4975 ( \5318 , \5316 , \5317 );
not \U$4976 ( \5319 , \5318 );
or \U$4977 ( \5320 , \5313 , \5319 );
not \U$4978 ( \5321 , \5044 );
or \U$4979 ( \5322 , \5321 , \4924 );
nand \U$4980 ( \5323 , \5320 , \5322 );
and \U$4981 ( \5324 , \4986 , \1165 );
not \U$4982 ( \5325 , \4986 );
and \U$4983 ( \5326 , \5325 , \1199 );
nor \U$4984 ( \5327 , \5324 , \5326 );
or \U$4985 ( \5328 , \5327 , \1809 );
or \U$4986 ( \5329 , \4994 , \1719 );
nand \U$4987 ( \5330 , \5328 , \5329 );
and \U$4988 ( \5331 , \5323 , \5330 );
not \U$4989 ( \5332 , \5323 );
not \U$4990 ( \5333 , \5330 );
and \U$4991 ( \5334 , \5332 , \5333 );
nor \U$4992 ( \5335 , \5331 , \5334 );
or \U$4993 ( \5336 , \5002 , \1137 );
xor \U$4994 ( \5337 , \1344 , RI98718c0_129);
or \U$4995 ( \5338 , \5337 , \1688 );
nand \U$4996 ( \5339 , \5336 , \5338 );
nand \U$4997 ( \5340 , \5335 , \5339 );
nand \U$4998 ( \5341 , \5323 , \5330 );
and \U$4999 ( \5342 , \5340 , \5341 );
not \U$5000 ( \5343 , \5342 );
not \U$5001 ( \5344 , \5343 );
or \U$5002 ( \5345 , \4825 , \932 );
and \U$5003 ( \5346 , RI9871d70_139, \3542 );
not \U$5004 ( \5347 , RI9871d70_139);
and \U$5005 ( \5348 , \5347 , \3537 );
nor \U$5006 ( \5349 , \5346 , \5348 );
buf \U$5007 ( \5350 , \859 );
not \U$5008 ( \5351 , \5350 );
or \U$5009 ( \5352 , \5349 , \5351 );
nand \U$5010 ( \5353 , \5345 , \5352 );
not \U$5011 ( \5354 , \1382 );
not \U$5012 ( \5355 , \1367 );
not \U$5013 ( \5356 , \4177 );
or \U$5014 ( \5357 , \5355 , \5356 );
nand \U$5015 ( \5358 , \4176 , RI9871e60_141);
nand \U$5016 ( \5359 , \5357 , \5358 );
not \U$5017 ( \5360 , \5359 );
or \U$5018 ( \5361 , \5354 , \5360 );
or \U$5019 ( \5362 , \5186 , \2595 );
nand \U$5020 ( \5363 , \5361 , \5362 );
xor \U$5021 ( \5364 , \5353 , \5363 );
not \U$5022 ( \5365 , \4841 );
or \U$5023 ( \5366 , \5365 , \3244 );
not \U$5024 ( \5367 , RI98719b0_131);
not \U$5025 ( \5368 , \5367 );
not \U$5026 ( \5369 , \943 );
or \U$5027 ( \5370 , \5368 , \5369 );
not \U$5028 ( \5371 , \3835 );
or \U$5029 ( \5372 , \5371 , \5367 );
nand \U$5030 ( \5373 , \5370 , \5372 );
not \U$5031 ( \5374 , \5373 );
or \U$5032 ( \5375 , \5374 , \1398 );
nand \U$5033 ( \5376 , \5366 , \5375 );
and \U$5034 ( \5377 , \5364 , \5376 );
and \U$5035 ( \5378 , \5353 , \5363 );
or \U$5036 ( \5379 , \5377 , \5378 );
not \U$5037 ( \5380 , \5379 );
not \U$5038 ( \5381 , \688 );
not \U$5039 ( \5382 , \5381 );
not \U$5040 ( \5383 , \1020 );
or \U$5041 ( \5384 , \5382 , \5383 );
nand \U$5042 ( \5385 , \5384 , \395 );
not \U$5043 ( \5386 , \394 );
nand \U$5044 ( \5387 , \5386 , \397 );
not \U$5045 ( \5388 , \5387 );
and \U$5046 ( \5389 , \5385 , \5388 );
not \U$5047 ( \5390 , \5385 );
and \U$5048 ( \5391 , \5390 , \5387 );
nor \U$5049 ( \5392 , \5389 , \5391 );
buf \U$5050 ( \5393 , \5392 );
and \U$5051 ( \5394 , \5393 , \1200 );
not \U$5052 ( \5395 , \3467 );
not \U$5053 ( \5396 , \5015 );
or \U$5054 ( \5397 , \5395 , \5396 );
and \U$5055 ( \5398 , RI98726d0_159, \1320 );
not \U$5056 ( \5399 , RI98726d0_159);
and \U$5057 ( \5400 , \5399 , \1740 );
or \U$5058 ( \5401 , \5398 , \5400 );
nand \U$5059 ( \5402 , \5401 , \3466 );
nand \U$5060 ( \5403 , \5397 , \5402 );
xor \U$5061 ( \5404 , \5394 , \5403 );
not \U$5062 ( \5405 , \1431 );
not \U$5063 ( \5406 , \4855 );
or \U$5064 ( \5407 , \5405 , \5406 );
and \U$5065 ( \5408 , \2842 , RI9871c08_136);
and \U$5066 ( \5409 , \1062 , \1619 );
nor \U$5067 ( \5410 , \5408 , \5409 );
not \U$5068 ( \5411 , \1455 );
or \U$5069 ( \5412 , \5410 , \5411 );
nand \U$5070 ( \5413 , \5407 , \5412 );
and \U$5071 ( \5414 , \5404 , \5413 );
and \U$5072 ( \5415 , \5394 , \5403 );
nor \U$5073 ( \5416 , \5414 , \5415 );
not \U$5074 ( \5417 , \5416 );
or \U$5075 ( \5418 , \5380 , \5417 );
or \U$5076 ( \5419 , \5416 , \5379 );
nand \U$5077 ( \5420 , \5418 , \5419 );
not \U$5078 ( \5421 , \5420 );
or \U$5079 ( \5422 , \5344 , \5421 );
not \U$5080 ( \5423 , \5416 );
nand \U$5081 ( \5424 , \5423 , \5379 );
nand \U$5082 ( \5425 , \5422 , \5424 );
and \U$5083 ( \5426 , \5312 , \5425 );
and \U$5084 ( \5427 , \5306 , \5311 );
or \U$5085 ( \5428 , \5426 , \5427 );
not \U$5086 ( \5429 , \5428 );
xor \U$5087 ( \5430 , \5161 , \5163 );
xor \U$5088 ( \5431 , \5430 , \5166 );
not \U$5089 ( \5432 , \5431 );
not \U$5090 ( \5433 , \4758 );
not \U$5091 ( \5434 , \4702 );
and \U$5092 ( \5435 , \5433 , \5434 );
and \U$5093 ( \5436 , \4758 , \4702 );
nor \U$5094 ( \5437 , \5435 , \5436 );
not \U$5095 ( \5438 , \5437 );
or \U$5096 ( \5439 , \5432 , \5438 );
or \U$5097 ( \5440 , \5437 , \5431 );
nand \U$5098 ( \5441 , \5439 , \5440 );
not \U$5099 ( \5442 , \5441 );
or \U$5100 ( \5443 , \5429 , \5442 );
not \U$5101 ( \5444 , \5437 );
nand \U$5102 ( \5445 , \5444 , \5431 );
nand \U$5103 ( \5446 , \5443 , \5445 );
not \U$5104 ( \5447 , \5446 );
not \U$5105 ( \5448 , \4763 );
not \U$5106 ( \5449 , \4770 );
or \U$5107 ( \5450 , \5448 , \5449 );
or \U$5108 ( \5451 , \4763 , \4770 );
nand \U$5109 ( \5452 , \5450 , \5451 );
not \U$5110 ( \5453 , \5452 );
not \U$5111 ( \5454 , \5065 );
or \U$5112 ( \5455 , \5453 , \5454 );
or \U$5113 ( \5456 , \5065 , \5452 );
nand \U$5114 ( \5457 , \5455 , \5456 );
nand \U$5115 ( \5458 , \5447 , \5457 );
not \U$5116 ( \5459 , \5458 );
xor \U$5117 ( \5460 , \5260 , \5263 );
xnor \U$5118 ( \5461 , \5460 , \5231 );
not \U$5119 ( \5462 , \5461 );
not \U$5120 ( \5463 , \5462 );
and \U$5121 ( \5464 , \5204 , \5215 );
not \U$5122 ( \5465 , \5204 );
and \U$5123 ( \5466 , \5465 , \5216 );
or \U$5124 ( \5467 , \5464 , \5466 );
xor \U$5125 ( \5468 , \5023 , \5051 );
xor \U$5126 ( \5469 , \5467 , \5468 );
xor \U$5127 ( \5470 , \4863 , \4876 );
xor \U$5128 ( \5471 , \5470 , \4888 );
and \U$5129 ( \5472 , \5469 , \5471 );
and \U$5130 ( \5473 , \5467 , \5468 );
nor \U$5131 ( \5474 , \5472 , \5473 );
not \U$5132 ( \5475 , \5474 );
xor \U$5133 ( \5476 , \4987 , \4997 );
xor \U$5134 ( \5477 , \5476 , \5004 );
not \U$5135 ( \5478 , \5477 );
not \U$5136 ( \5479 , \915 );
not \U$5137 ( \5480 , \5479 );
xor \U$5138 ( \5481 , RI9872310_151, \5480 );
not \U$5139 ( \5482 , \5481 );
not \U$5140 ( \5483 , \3962 );
and \U$5141 ( \5484 , \5482 , \5483 );
and \U$5142 ( \5485 , \4868 , \3170 );
nor \U$5143 ( \5486 , \5484 , \5485 );
not \U$5144 ( \5487 , \5486 );
not \U$5145 ( \5488 , \5487 );
or \U$5146 ( \5489 , \4886 , \1543 );
and \U$5147 ( \5490 , RI9871b18_134, \1212 );
not \U$5148 ( \5491 , RI9871b18_134);
and \U$5149 ( \5492 , \5491 , \3129 );
nor \U$5150 ( \5493 , \5490 , \5492 );
not \U$5151 ( \5494 , \5493 );
or \U$5152 ( \5495 , \5494 , \1293 );
nand \U$5153 ( \5496 , \5489 , \5495 );
not \U$5154 ( \5497 , \5496 );
not \U$5155 ( \5498 , \1518 );
not \U$5156 ( \5499 , \4806 );
or \U$5157 ( \5500 , \5498 , \5499 );
xor \U$5158 ( \5501 , \3275 , RI9871c80_137);
nand \U$5159 ( \5502 , \5501 , \1501 );
nand \U$5160 ( \5503 , \5500 , \5502 );
not \U$5161 ( \5504 , \5503 );
not \U$5162 ( \5505 , \5504 );
or \U$5163 ( \5506 , \5497 , \5505 );
not \U$5164 ( \5507 , \5496 );
nand \U$5165 ( \5508 , \5507 , \5503 );
nand \U$5166 ( \5509 , \5506 , \5508 );
not \U$5167 ( \5510 , \5509 );
or \U$5168 ( \5511 , \5488 , \5510 );
nand \U$5169 ( \5512 , \5503 , \5496 );
nand \U$5170 ( \5513 , \5511 , \5512 );
not \U$5171 ( \5514 , \876 );
and \U$5172 ( \5515 , RI9872130_147, \2948 );
not \U$5173 ( \5516 , RI9872130_147);
and \U$5174 ( \5517 , \5516 , \3691 );
nor \U$5175 ( \5518 , \5515 , \5517 );
not \U$5176 ( \5519 , \5518 );
or \U$5177 ( \5520 , \5514 , \5519 );
or \U$5178 ( \5521 , \4833 , \1470 );
nand \U$5179 ( \5522 , \5520 , \5521 );
not \U$5180 ( \5523 , \4085 );
not \U$5181 ( \5524 , \4784 );
or \U$5182 ( \5525 , \5523 , \5524 );
and \U$5183 ( \5526 , RI98725e0_157, \1417 );
not \U$5184 ( \5527 , RI98725e0_157);
and \U$5185 ( \5528 , \5527 , \1416 );
nor \U$5186 ( \5529 , \5526 , \5528 );
not \U$5187 ( \5530 , \4102 );
nand \U$5188 ( \5531 , \5529 , \5530 );
nand \U$5189 ( \5532 , \5525 , \5531 );
xor \U$5190 ( \5533 , \5522 , \5532 );
not \U$5191 ( \5534 , \2087 );
not \U$5192 ( \5535 , \4791 );
or \U$5193 ( \5536 , \5534 , \5535 );
xor \U$5194 ( \5537 , RI9871aa0_133, \821 );
nand \U$5195 ( \5538 , \5537 , \2074 );
nand \U$5196 ( \5539 , \5536 , \5538 );
and \U$5197 ( \5540 , \5533 , \5539 );
and \U$5198 ( \5541 , \5522 , \5532 );
or \U$5199 ( \5542 , \5540 , \5541 );
or \U$5200 ( \5543 , \5513 , \5542 );
not \U$5201 ( \5544 , \5543 );
or \U$5202 ( \5545 , \5478 , \5544 );
nand \U$5203 ( \5546 , \5513 , \5542 );
nand \U$5204 ( \5547 , \5545 , \5546 );
xor \U$5205 ( \5548 , \5475 , \5547 );
not \U$5206 ( \5549 , \5242 );
not \U$5207 ( \5550 , \5255 );
not \U$5208 ( \5551 , \5550 );
or \U$5209 ( \5552 , \5549 , \5551 );
not \U$5210 ( \5553 , \5242 );
nand \U$5211 ( \5554 , \5553 , \5255 );
nand \U$5212 ( \5555 , \5552 , \5554 );
and \U$5213 ( \5556 , \5548 , \5555 );
and \U$5214 ( \5557 , \5475 , \5547 );
nor \U$5215 ( \5558 , \5556 , \5557 );
not \U$5216 ( \5559 , \4900 );
and \U$5217 ( \5560 , \5061 , \5559 );
not \U$5218 ( \5561 , \5061 );
and \U$5219 ( \5562 , \5561 , \4900 );
nor \U$5220 ( \5563 , \5560 , \5562 );
and \U$5221 ( \5564 , \5558 , \5563 );
not \U$5222 ( \5565 , \5558 );
not \U$5223 ( \5566 , \5563 );
and \U$5224 ( \5567 , \5565 , \5566 );
nor \U$5225 ( \5568 , \5564 , \5567 );
not \U$5226 ( \5569 , \5568 );
or \U$5227 ( \5570 , \5463 , \5569 );
not \U$5228 ( \5571 , \5558 );
nand \U$5229 ( \5572 , \5571 , \5566 );
nand \U$5230 ( \5573 , \5570 , \5572 );
not \U$5231 ( \5574 , \5573 );
or \U$5232 ( \5575 , \5459 , \5574 );
not \U$5233 ( \5576 , \5457 );
nand \U$5234 ( \5577 , \5576 , \5446 );
nand \U$5235 ( \5578 , \5575 , \5577 );
not \U$5236 ( \5579 , \5578 );
xor \U$5237 ( \5580 , \4701 , \5069 );
xor \U$5238 ( \5581 , \5580 , \5268 );
xor \U$5239 ( \5582 , \5276 , \5283 );
xnor \U$5240 ( \5583 , \5582 , \5278 );
or \U$5241 ( \5584 , \5581 , \5583 );
not \U$5242 ( \5585 , \5584 );
or \U$5243 ( \5586 , \5579 , \5585 );
nand \U$5244 ( \5587 , \5581 , \5583 );
nand \U$5245 ( \5588 , \5586 , \5587 );
not \U$5246 ( \5589 , \5588 );
xnor \U$5247 ( \5590 , \5292 , \5271 );
nand \U$5248 ( \5591 , \5589 , \5590 );
and \U$5249 ( \5592 , \4043 , \5304 , \5591 );
not \U$5250 ( \5593 , \859 );
buf \U$5251 ( \5594 , \4174 );
not \U$5252 ( \5595 , \5594 );
buf \U$5253 ( \5596 , \5595 );
and \U$5254 ( \5597 , RI9871d70_139, \5596 );
not \U$5255 ( \5598 , RI9871d70_139);
not \U$5256 ( \5599 , \4176 );
and \U$5257 ( \5600 , \5598 , \5599 );
or \U$5258 ( \5601 , \5597 , \5600 );
not \U$5259 ( \5602 , \5601 );
or \U$5260 ( \5603 , \5593 , \5602 );
and \U$5261 ( \5604 , \4154 , RI9871d70_139);
and \U$5262 ( \5605 , \3569 , \1347 );
nor \U$5263 ( \5606 , \5604 , \5605 );
or \U$5264 ( \5607 , \5606 , \932 );
nand \U$5265 ( \5608 , \5603 , \5607 );
not \U$5266 ( \5609 , \1353 );
not \U$5267 ( \5610 , \1367 );
not \U$5268 ( \5611 , \5205 );
not \U$5269 ( \5612 , \5611 );
or \U$5270 ( \5613 , \5610 , \5612 );
not \U$5271 ( \5614 , \4407 );
not \U$5272 ( \5615 , \5614 );
not \U$5273 ( \5616 , RI9871e60_141);
or \U$5274 ( \5617 , \5615 , \5616 );
nand \U$5275 ( \5618 , \5613 , \5617 );
not \U$5276 ( \5619 , \5618 );
or \U$5277 ( \5620 , \5609 , \5619 );
not \U$5278 ( \5621 , RI9871e60_141);
not \U$5279 ( \5622 , \5621 );
not \U$5280 ( \5623 , \4470 );
not \U$5281 ( \5624 , \5623 );
or \U$5282 ( \5625 , \5622 , \5624 );
or \U$5283 ( \5626 , \4712 , \5616 );
nand \U$5284 ( \5627 , \5625 , \5626 );
nand \U$5285 ( \5628 , \5627 , \1381 );
nand \U$5286 ( \5629 , \5620 , \5628 );
not \U$5287 ( \5630 , \5629 );
not \U$5288 ( \5631 , RI9872838_162);
not \U$5289 ( \5632 , RI98728b0_163);
nand \U$5290 ( \5633 , \5631 , \5632 );
nand \U$5291 ( \5634 , RI9872838_162, RI98728b0_163);
and \U$5292 ( \5635 , \5633 , \5634 );
not \U$5293 ( \5636 , \5635 );
and \U$5294 ( \5637 , RI9872568_156, RI9872838_162);
not \U$5295 ( \5638 , RI9872568_156);
and \U$5296 ( \5639 , \5638 , \5631 );
nor \U$5297 ( \5640 , \5637 , \5639 );
and \U$5298 ( \5641 , \5636 , \5640 );
buf \U$5299 ( \5642 , \5641 );
not \U$5300 ( \5643 , \5642 );
not \U$5301 ( \5644 , RI9872568_156);
not \U$5302 ( \5645 , \5644 );
not \U$5303 ( \5646 , \2361 );
or \U$5304 ( \5647 , \5645 , \5646 );
not \U$5305 ( \5648 , RI9872568_156);
or \U$5306 ( \5649 , \780 , \5648 );
nand \U$5307 ( \5650 , \5647 , \5649 );
not \U$5308 ( \5651 , \5650 );
or \U$5309 ( \5652 , \5643 , \5651 );
buf \U$5310 ( \5653 , \5635 );
nand \U$5311 ( \5654 , \5653 , RI9872568_156);
nand \U$5312 ( \5655 , \5652 , \5654 );
not \U$5313 ( \5656 , \5655 );
or \U$5314 ( \5657 , \5630 , \5656 );
or \U$5315 ( \5658 , \5655 , \5629 );
nand \U$5316 ( \5659 , \5657 , \5658 );
xor \U$5317 ( \5660 , \5608 , \5659 );
not \U$5318 ( \5661 , \5660 );
not \U$5319 ( \5662 , \5661 );
not \U$5320 ( \5663 , \654 );
not \U$5321 ( \5664 , \564 );
not \U$5322 ( \5665 , \638 );
nor \U$5323 ( \5666 , \5664 , \5665 );
not \U$5324 ( \5667 , \5666 );
not \U$5325 ( \5668 , \548 );
not \U$5326 ( \5669 , \536 );
buf \U$5327 ( \5670 , \614 );
not \U$5328 ( \5671 , \5670 );
nand \U$5329 ( \5672 , \5669 , \5671 );
not \U$5330 ( \5673 , \5672 );
or \U$5331 ( \5674 , \5668 , \5673 );
not \U$5332 ( \5675 , \547 );
not \U$5333 ( \5676 , \649 );
or \U$5334 ( \5677 , \5675 , \5676 );
buf \U$5335 ( \5678 , \651 );
nand \U$5336 ( \5679 , \5677 , \5678 );
not \U$5337 ( \5680 , \5679 );
nand \U$5338 ( \5681 , \5680 , \634 );
not \U$5339 ( \5682 , \5681 );
nand \U$5340 ( \5683 , \5674 , \5682 );
not \U$5341 ( \5684 , \5683 );
or \U$5342 ( \5685 , \5667 , \5684 );
not \U$5343 ( \5686 , \560 );
not \U$5344 ( \5687 , \678 );
or \U$5345 ( \5688 , \5686 , \5687 );
buf \U$5346 ( \5689 , \682 );
nand \U$5347 ( \5690 , \5688 , \5689 );
nand \U$5348 ( \5691 , \5690 , \564 );
nand \U$5349 ( \5692 , \5685 , \5691 );
not \U$5350 ( \5693 , \5692 );
or \U$5351 ( \5694 , \5663 , \5693 );
not \U$5352 ( \5695 , \664 );
nand \U$5353 ( \5696 , \5694 , \5695 );
nand \U$5354 ( \5697 , \665 , \684 );
not \U$5355 ( \5698 , \5697 );
and \U$5356 ( \5699 , \5696 , \5698 );
not \U$5357 ( \5700 , \5696 );
and \U$5358 ( \5701 , \5700 , \5697 );
nor \U$5359 ( \5702 , \5699 , \5701 );
buf \U$5360 ( \5703 , \5702 );
not \U$5361 ( \5704 , \5703 );
buf \U$5362 ( \5705 , \5704 );
not \U$5363 ( \5706 , \5705 );
not \U$5364 ( \5707 , \5706 );
buf \U$5365 ( \5708 , \5707 );
not \U$5366 ( \5709 , \5708 );
nand \U$5367 ( \5710 , \5709 , \1200 );
not \U$5368 ( \5711 , \793 );
not \U$5369 ( \5712 , \1340 );
and \U$5370 ( \5713 , RI98719b0_131, \5712 );
not \U$5371 ( \5714 , RI98719b0_131);
and \U$5372 ( \5715 , \5714 , \1344 );
nor \U$5373 ( \5716 , \5713 , \5715 );
not \U$5374 ( \5717 , \5716 );
or \U$5375 ( \5718 , \5711 , \5717 );
not \U$5376 ( \5719 , \1252 );
not \U$5377 ( \5720 , \5719 );
not \U$5378 ( \5721 , \5720 );
and \U$5379 ( \5722 , RI98719b0_131, \5721 );
not \U$5380 ( \5723 , RI98719b0_131);
and \U$5381 ( \5724 , \5723 , \5720 );
nor \U$5382 ( \5725 , \5722 , \5724 );
nand \U$5383 ( \5726 , \5725 , \796 );
nand \U$5384 ( \5727 , \5718 , \5726 );
xor \U$5385 ( \5728 , \5710 , \5727 );
not \U$5386 ( \5729 , \1067 );
and \U$5387 ( \5730 , \4990 , \1043 );
not \U$5388 ( \5731 , \4990 );
and \U$5389 ( \5732 , \5731 , \1044 );
nor \U$5390 ( \5733 , \5730 , \5732 );
not \U$5391 ( \5734 , \5733 );
or \U$5392 ( \5735 , \5729 , \5734 );
buf \U$5393 ( \5736 , \4984 );
and \U$5394 ( \5737 , \3271 , \5736 );
not \U$5395 ( \5738 , \3271 );
not \U$5396 ( \5739 , \5736 );
and \U$5397 ( \5740 , \5738 , \5739 );
nor \U$5398 ( \5741 , \5737 , \5740 );
not \U$5399 ( \5742 , \5741 );
or \U$5400 ( \5743 , \5742 , \1612 );
nand \U$5401 ( \5744 , \5735 , \5743 );
xor \U$5402 ( \5745 , \5728 , \5744 );
not \U$5403 ( \5746 , \5745 );
and \U$5404 ( \5747 , \5662 , \5746 );
not \U$5405 ( \5748 , \5745 );
not \U$5406 ( \5749 , \5660 );
or \U$5407 ( \5750 , \5748 , \5749 );
or \U$5408 ( \5751 , \5660 , \5745 );
nand \U$5409 ( \5752 , \5750 , \5751 );
not \U$5410 ( \5753 , \1164 );
buf \U$5411 ( \5754 , \1020 );
nand \U$5412 ( \5755 , \5381 , \395 );
and \U$5413 ( \5756 , \5754 , \5755 );
not \U$5414 ( \5757 , \5754 );
not \U$5415 ( \5758 , \5755 );
and \U$5416 ( \5759 , \5757 , \5758 );
nor \U$5417 ( \5760 , \5756 , \5759 );
buf \U$5418 ( \5761 , \5760 );
not \U$5419 ( \5762 , \5761 );
not \U$5420 ( \5763 , \5762 );
and \U$5421 ( \5764 , \5753 , \5763 );
not \U$5422 ( \5765 , \5753 );
not \U$5423 ( \5766 , \5761 );
and \U$5424 ( \5767 , \5765 , \5766 );
nor \U$5425 ( \5768 , \5764 , \5767 );
or \U$5426 ( \5769 , \5768 , \1809 );
not \U$5427 ( \5770 , \5385 );
not \U$5428 ( \5771 , \5387 );
and \U$5429 ( \5772 , \5770 , \5771 );
and \U$5430 ( \5773 , \5385 , \5387 );
nor \U$5431 ( \5774 , \5772 , \5773 );
buf \U$5432 ( \5775 , \5774 );
buf \U$5433 ( \5776 , \5775 );
and \U$5434 ( \5777 , \5776 , \1165 );
and \U$5435 ( \5778 , \5393 , \1199 );
nor \U$5436 ( \5779 , \5777 , \5778 );
or \U$5437 ( \5780 , \5779 , \1719 );
nand \U$5438 ( \5781 , \5769 , \5780 );
not \U$5439 ( \5782 , \5034 );
not \U$5440 ( \5783 , RI9872478_154);
not \U$5441 ( \5784 , \1127 );
or \U$5442 ( \5785 , \5783 , \5784 );
or \U$5443 ( \5786 , \1725 , RI9872478_154);
nand \U$5444 ( \5787 , \5785 , \5786 );
not \U$5445 ( \5788 , \5787 );
or \U$5446 ( \5789 , \5782 , \5788 );
not \U$5447 ( \5790 , \5025 );
not \U$5448 ( \5791 , \1393 );
or \U$5449 ( \5792 , \5790 , \5791 );
or \U$5450 ( \5793 , \2982 , \5025 );
nand \U$5451 ( \5794 , \5792 , \5793 );
not \U$5452 ( \5795 , \5035 );
not \U$5453 ( \5796 , \5795 );
nand \U$5454 ( \5797 , \5794 , \5796 );
nand \U$5455 ( \5798 , \5789 , \5797 );
xor \U$5456 ( \5799 , \5781 , \5798 );
and \U$5457 ( \5800 , \1111 , \1605 );
not \U$5458 ( \5801 , \1111 );
and \U$5459 ( \5802 , \5801 , \1606 );
nor \U$5460 ( \5803 , \5800 , \5802 );
or \U$5461 ( \5804 , \5803 , \1137 );
and \U$5462 ( \5805 , RI98718c0_129, \1062 );
not \U$5463 ( \5806 , RI98718c0_129);
and \U$5464 ( \5807 , \5806 , \2842 );
nor \U$5465 ( \5808 , \5805 , \5807 );
not \U$5466 ( \5809 , \5808 );
or \U$5467 ( \5810 , \5809 , \1676 );
nand \U$5468 ( \5811 , \5804 , \5810 );
not \U$5469 ( \5812 , \5811 );
and \U$5470 ( \5813 , \5799 , \5812 );
not \U$5471 ( \5814 , \5799 );
and \U$5472 ( \5815 , \5814 , \5811 );
nor \U$5473 ( \5816 , \5813 , \5815 );
not \U$5474 ( \5817 , \5816 );
and \U$5475 ( \5818 , \5752 , \5817 );
nor \U$5476 ( \5819 , \5747 , \5818 );
not \U$5477 ( \5820 , \1018 );
not \U$5478 ( \5821 , \5733 );
or \U$5479 ( \5822 , \5820 , \5821 );
and \U$5480 ( \5823 , \4471 , \3272 );
and \U$5481 ( \5824 , \4712 , \1045 );
nor \U$5482 ( \5825 , \5823 , \5824 );
or \U$5483 ( \5826 , \5825 , \1068 );
nand \U$5484 ( \5827 , \5822 , \5826 );
not \U$5485 ( \5828 , \797 );
not \U$5486 ( \5829 , \5373 );
or \U$5487 ( \5830 , \5828 , \5829 );
nand \U$5488 ( \5831 , \793 , \5725 );
nand \U$5489 ( \5832 , \5830 , \5831 );
xor \U$5490 ( \5833 , \5827 , \5832 );
or \U$5491 ( \5834 , \5779 , \1809 );
or \U$5492 ( \5835 , \5327 , \1719 );
nand \U$5493 ( \5836 , \5834 , \5835 );
xor \U$5494 ( \5837 , \5833 , \5836 );
not \U$5495 ( \5838 , \3467 );
not \U$5496 ( \5839 , \5401 );
or \U$5497 ( \5840 , \5838 , \5839 );
and \U$5498 ( \5841 , RI98726d0_159, \1583 );
not \U$5499 ( \5842 , RI98726d0_159);
and \U$5500 ( \5843 , \5842 , \1275 );
or \U$5501 ( \5844 , \5841 , \5843 );
nand \U$5502 ( \5845 , \5844 , \3600 );
nand \U$5503 ( \5846 , \5840 , \5845 );
buf \U$5504 ( \5847 , \4084 );
not \U$5505 ( \5848 , \5847 );
not \U$5506 ( \5849 , \5529 );
or \U$5507 ( \5850 , \5848 , \5849 );
and \U$5508 ( \5851 , RI98725e0_157, \2680 );
not \U$5509 ( \5852 , RI98725e0_157);
and \U$5510 ( \5853 , \5852 , \1447 );
nor \U$5511 ( \5854 , \5851 , \5853 );
nand \U$5512 ( \5855 , \5854 , \5530 );
nand \U$5513 ( \5856 , \5850 , \5855 );
xor \U$5514 ( \5857 , \5846 , \5856 );
not \U$5515 ( \5858 , \5857 );
or \U$5516 ( \5859 , \5337 , \1137 );
or \U$5517 ( \5860 , \5803 , \1676 );
nand \U$5518 ( \5861 , \5859 , \5860 );
not \U$5519 ( \5862 , \5861 );
not \U$5520 ( \5863 , \5862 );
and \U$5521 ( \5864 , \5858 , \5863 );
and \U$5522 ( \5865 , \5857 , \5862 );
nor \U$5523 ( \5866 , \5864 , \5865 );
xor \U$5524 ( \5867 , \5837 , \5866 );
and \U$5525 ( \5868 , \4370 , \919 );
not \U$5526 ( \5869 , \4370 );
and \U$5527 ( \5870 , \5869 , RI9872130_147);
nor \U$5528 ( \5871 , \5868 , \5870 );
not \U$5529 ( \5872 , \5871 );
or \U$5530 ( \5873 , \5872 , \1470 );
not \U$5531 ( \5874 , \919 );
not \U$5532 ( \5875 , \3543 );
or \U$5533 ( \5876 , \5874 , \5875 );
not \U$5534 ( \5877 , RI9872130_147);
or \U$5535 ( \5878 , \3537 , \5877 );
nand \U$5536 ( \5879 , \5876 , \5878 );
not \U$5537 ( \5880 , \5879 );
or \U$5538 ( \5881 , \5880 , \1942 );
nand \U$5539 ( \5882 , \5873 , \5881 );
not \U$5540 ( \5883 , \5882 );
not \U$5541 ( \5884 , \2947 );
not \U$5542 ( \5885 , \5884 );
and \U$5543 ( \5886 , \5885 , \1584 );
not \U$5544 ( \5887 , \5885 );
and \U$5545 ( \5888 , \5887 , RI9871c80_137);
nor \U$5546 ( \5889 , \5886 , \5888 );
not \U$5547 ( \5890 , \5889 );
not \U$5548 ( \5891 , \1501 );
or \U$5549 ( \5892 , \5890 , \5891 );
not \U$5550 ( \5893 , RI9871c80_137);
xor \U$5551 ( \5894 , \2962 , \5893 );
not \U$5552 ( \5895 , \5894 );
or \U$5553 ( \5896 , \5895 , \1746 );
nand \U$5554 ( \5897 , \5892 , \5896 );
not \U$5555 ( \5898 , \2087 );
not \U$5556 ( \5899 , \2076 );
not \U$5557 ( \5900 , \2216 );
not \U$5558 ( \5901 , \5900 );
or \U$5559 ( \5902 , \5899 , \5901 );
nand \U$5560 ( \5903 , \848 , RI9871aa0_133);
nand \U$5561 ( \5904 , \5902 , \5903 );
not \U$5562 ( \5905 , \5904 );
or \U$5563 ( \5906 , \5898 , \5905 );
buf \U$5564 ( \5907 , \941 );
not \U$5565 ( \5908 , \5907 );
not \U$5566 ( \5909 , \5908 );
not \U$5567 ( \5910 , \2076 );
and \U$5568 ( \5911 , \5909 , \5910 );
and \U$5569 ( \5912 , \5371 , \2080 );
nor \U$5570 ( \5913 , \5911 , \5912 );
not \U$5571 ( \5914 , \5913 );
nand \U$5572 ( \5915 , \5914 , \2074 );
nand \U$5573 ( \5916 , \5906 , \5915 );
xor \U$5574 ( \5917 , \5897 , \5916 );
not \U$5575 ( \5918 , \5917 );
or \U$5576 ( \5919 , \5883 , \5918 );
nand \U$5577 ( \5920 , \5916 , \5897 );
nand \U$5578 ( \5921 , \5919 , \5920 );
xor \U$5579 ( \5922 , \5867 , \5921 );
xor \U$5580 ( \5923 , \5819 , \5922 );
and \U$5581 ( \5924 , \5608 , \5659 );
not \U$5582 ( \5925 , \5655 );
and \U$5583 ( \5926 , \5925 , \5629 );
nor \U$5584 ( \5927 , \5924 , \5926 );
not \U$5585 ( \5928 , \1456 );
and \U$5586 ( \5929 , RI9871c08_136, \1047 );
not \U$5587 ( \5930 , RI9871c08_136);
and \U$5588 ( \5931 , \5930 , \1041 );
nor \U$5589 ( \5932 , \5929 , \5931 );
not \U$5590 ( \5933 , \5932 );
or \U$5591 ( \5934 , \5928 , \5933 );
or \U$5592 ( \5935 , \5410 , \1432 );
nand \U$5593 ( \5936 , \5934 , \5935 );
buf \U$5594 ( \5937 , \4925 );
not \U$5595 ( \5938 , \5937 );
not \U$5596 ( \5939 , \5318 );
or \U$5597 ( \5940 , \5938 , \5939 );
xnor \U$5598 ( \5941 , RI9872388_152, \1097 );
buf \U$5599 ( \5942 , \4919 );
nand \U$5600 ( \5943 , \5941 , \5942 );
nand \U$5601 ( \5944 , \5940 , \5943 );
not \U$5602 ( \5945 , \1292 );
buf \U$5603 ( \5946 , \3394 );
not \U$5604 ( \5947 , \5946 );
not \U$5605 ( \5948 , \5947 );
not \U$5606 ( \5949 , \5948 );
xor \U$5607 ( \5950 , RI9871b18_134, \5949 );
not \U$5608 ( \5951 , \5950 );
or \U$5609 ( \5952 , \5945 , \5951 );
nand \U$5610 ( \5953 , \5493 , \1323 );
nand \U$5611 ( \5954 , \5952 , \5953 );
xor \U$5612 ( \5955 , \5944 , \5954 );
xor \U$5613 ( \5956 , \5936 , \5955 );
xnor \U$5614 ( \5957 , \5927 , \5956 );
or \U$5615 ( \5958 , \5349 , \932 );
or \U$5616 ( \5959 , \5606 , \5351 );
nand \U$5617 ( \5960 , \5958 , \5959 );
and \U$5618 ( \5961 , \5359 , \1353 );
and \U$5619 ( \5962 , \5618 , \1381 );
nor \U$5620 ( \5963 , \5961 , \5962 );
not \U$5621 ( \5964 , \5963 );
xor \U$5622 ( \5965 , \5960 , \5964 );
not \U$5623 ( \5966 , \2087 );
not \U$5624 ( \5967 , \5537 );
or \U$5625 ( \5968 , \5966 , \5967 );
nand \U$5626 ( \5969 , \5904 , \2074 );
nand \U$5627 ( \5970 , \5968 , \5969 );
xnor \U$5628 ( \5971 , \5965 , \5970 );
xor \U$5629 ( \5972 , \5957 , \5971 );
and \U$5630 ( \5973 , \5923 , \5972 );
and \U$5631 ( \5974 , \5819 , \5922 );
or \U$5632 ( \5975 , \5973 , \5974 );
not \U$5633 ( \5976 , \5339 );
xor \U$5634 ( \5977 , \5335 , \5976 );
not \U$5635 ( \5978 , \5977 );
not \U$5636 ( \5979 , \5936 );
not \U$5637 ( \5980 , \5955 );
or \U$5638 ( \5981 , \5979 , \5980 );
nand \U$5639 ( \5982 , \5954 , \5944 );
nand \U$5640 ( \5983 , \5981 , \5982 );
not \U$5641 ( \5984 , \5960 );
not \U$5642 ( \5985 , \5963 );
not \U$5643 ( \5986 , \5970 );
or \U$5644 ( \5987 , \5985 , \5986 );
or \U$5645 ( \5988 , \5970 , \5963 );
nand \U$5646 ( \5989 , \5987 , \5988 );
not \U$5647 ( \5990 , \5989 );
or \U$5648 ( \5991 , \5984 , \5990 );
nand \U$5649 ( \5992 , \5970 , \5964 );
nand \U$5650 ( \5993 , \5991 , \5992 );
xor \U$5651 ( \5994 , \5983 , \5993 );
not \U$5652 ( \5995 , \5994 );
or \U$5653 ( \5996 , \5978 , \5995 );
or \U$5654 ( \5997 , \5994 , \5977 );
nand \U$5655 ( \5998 , \5996 , \5997 );
not \U$5656 ( \5999 , \5998 );
not \U$5657 ( \6000 , \5744 );
not \U$5658 ( \6001 , \5728 );
not \U$5659 ( \6002 , \6001 );
or \U$5660 ( \6003 , \6000 , \6002 );
not \U$5661 ( \6004 , \5710 );
nand \U$5662 ( \6005 , \6004 , \5727 );
nand \U$5663 ( \6006 , \6003 , \6005 );
not \U$5664 ( \6007 , \6006 );
not \U$5665 ( \6008 , \6007 );
not \U$5666 ( \6009 , \5811 );
not \U$5667 ( \6010 , \5799 );
or \U$5668 ( \6011 , \6009 , \6010 );
nand \U$5669 ( \6012 , \5798 , \5781 );
nand \U$5670 ( \6013 , \6011 , \6012 );
not \U$5671 ( \6014 , \6013 );
not \U$5672 ( \6015 , \6014 );
or \U$5673 ( \6016 , \6008 , \6015 );
not \U$5674 ( \6017 , \1431 );
not \U$5675 ( \6018 , \5932 );
or \U$5676 ( \6019 , \6017 , \6018 );
not \U$5677 ( \6020 , \1209 );
not \U$5678 ( \6021 , \6020 );
and \U$5679 ( \6022 , RI9871c08_136, \6021 );
not \U$5680 ( \6023 , RI9871c08_136);
and \U$5681 ( \6024 , \6023 , \3128 );
or \U$5682 ( \6025 , \6022 , \6024 );
nand \U$5683 ( \6026 , \6025 , \1456 );
nand \U$5684 ( \6027 , \6019 , \6026 );
not \U$5685 ( \6028 , \3467 );
not \U$5686 ( \6029 , \5844 );
or \U$5687 ( \6030 , \6028 , \6029 );
not \U$5688 ( \6031 , RI98726d0_159);
not \U$5689 ( \6032 , \5480 );
or \U$5690 ( \6033 , \6031 , \6032 );
or \U$5691 ( \6034 , \916 , RI98726d0_159);
nand \U$5692 ( \6035 , \6033 , \6034 );
nand \U$5693 ( \6036 , \6035 , \3600 );
nand \U$5694 ( \6037 , \6030 , \6036 );
xor \U$5695 ( \6038 , \6027 , \6037 );
not \U$5696 ( \6039 , \5530 );
and \U$5697 ( \6040 , \1309 , RI98725e0_157);
not \U$5698 ( \6041 , \1309 );
not \U$5699 ( \6042 , RI98725e0_157);
and \U$5700 ( \6043 , \6041 , \6042 );
nor \U$5701 ( \6044 , \6040 , \6043 );
not \U$5702 ( \6045 , \6044 );
or \U$5703 ( \6046 , \6039 , \6045 );
not \U$5704 ( \6047 , \5854 );
not \U$5705 ( \6048 , \5847 );
or \U$5706 ( \6049 , \6047 , \6048 );
nand \U$5707 ( \6050 , \6046 , \6049 );
and \U$5708 ( \6051 , \6038 , \6050 );
and \U$5709 ( \6052 , \6027 , \6037 );
or \U$5710 ( \6053 , \6051 , \6052 );
nand \U$5711 ( \6054 , \6016 , \6053 );
nand \U$5712 ( \6055 , \6013 , \6006 );
nand \U$5713 ( \6056 , \6054 , \6055 );
not \U$5714 ( \6057 , \6056 );
not \U$5715 ( \6058 , \5760 );
not \U$5716 ( \6059 , \6058 );
not \U$5717 ( \6060 , \6059 );
nand \U$5718 ( \6061 , \6060 , \1165 );
not \U$5719 ( \6062 , \6061 );
buf \U$5720 ( \6063 , \5641 );
or \U$5721 ( \6064 , \6063 , \5653 );
nand \U$5722 ( \6065 , \6064 , RI9872568_156);
not \U$5723 ( \6066 , \6065 );
and \U$5724 ( \6067 , \6062 , \6066 );
and \U$5725 ( \6068 , \6061 , \6065 );
nor \U$5726 ( \6069 , \6067 , \6068 );
not \U$5727 ( \6070 , \6069 );
not \U$5728 ( \6071 , \6070 );
not \U$5729 ( \6072 , \5034 );
not \U$5730 ( \6073 , \5794 );
or \U$5731 ( \6074 , \6072 , \6073 );
nand \U$5732 ( \6075 , \5195 , \5796 );
nand \U$5733 ( \6076 , \6074 , \6075 );
not \U$5734 ( \6077 , \6076 );
or \U$5735 ( \6078 , \6071 , \6077 );
not \U$5736 ( \6079 , \6061 );
nand \U$5737 ( \6080 , \6079 , \6065 );
nand \U$5738 ( \6081 , \6078 , \6080 );
not \U$5739 ( \6082 , \6081 );
xor \U$5740 ( \6083 , \5827 , \5832 );
and \U$5741 ( \6084 , \6083 , \5836 );
and \U$5742 ( \6085 , \5827 , \5832 );
nor \U$5743 ( \6086 , \6084 , \6085 );
xor \U$5744 ( \6087 , \6082 , \6086 );
not \U$5745 ( \6088 , \5861 );
not \U$5746 ( \6089 , \5857 );
or \U$5747 ( \6090 , \6088 , \6089 );
nand \U$5748 ( \6091 , \5856 , \5846 );
nand \U$5749 ( \6092 , \6090 , \6091 );
xnor \U$5750 ( \6093 , \6087 , \6092 );
not \U$5751 ( \6094 , \6093 );
or \U$5752 ( \6095 , \6057 , \6094 );
or \U$5753 ( \6096 , \6093 , \6056 );
nand \U$5754 ( \6097 , \6095 , \6096 );
not \U$5755 ( \6098 , \6097 );
not \U$5756 ( \6099 , \6098 );
or \U$5757 ( \6100 , \5999 , \6099 );
not \U$5758 ( \6101 , \5998 );
nand \U$5759 ( \6102 , \6101 , \6097 );
nand \U$5760 ( \6103 , \6100 , \6102 );
xnor \U$5761 ( \6104 , \5975 , \6103 );
xor \U$5762 ( \6105 , \5394 , \5413 );
xnor \U$5763 ( \6106 , \6105 , \5403 );
not \U$5764 ( \6107 , \6106 );
not \U$5765 ( \6108 , \5486 );
not \U$5766 ( \6109 , \5509 );
or \U$5767 ( \6110 , \6108 , \6109 );
or \U$5768 ( \6111 , \5509 , \5486 );
nand \U$5769 ( \6112 , \6110 , \6111 );
not \U$5770 ( \6113 , \6112 );
or \U$5771 ( \6114 , \6107 , \6113 );
or \U$5772 ( \6115 , \6106 , \6112 );
nand \U$5773 ( \6116 , \6114 , \6115 );
xor \U$5774 ( \6117 , \5353 , \5363 );
xor \U$5775 ( \6118 , \6117 , \5376 );
xnor \U$5776 ( \6119 , \6116 , \6118 );
not \U$5777 ( \6120 , \6119 );
not \U$5778 ( \6121 , \5971 );
not \U$5779 ( \6122 , \6121 );
not \U$5780 ( \6123 , \5957 );
or \U$5781 ( \6124 , \6122 , \6123 );
not \U$5782 ( \6125 , \5927 );
nand \U$5783 ( \6126 , \6125 , \5956 );
nand \U$5784 ( \6127 , \6124 , \6126 );
not \U$5785 ( \6128 , \5921 );
nand \U$5786 ( \6129 , \6128 , \5866 );
not \U$5787 ( \6130 , \6129 );
not \U$5788 ( \6131 , \5837 );
or \U$5789 ( \6132 , \6130 , \6131 );
not \U$5790 ( \6133 , \5866 );
nand \U$5791 ( \6134 , \6133 , \5921 );
nand \U$5792 ( \6135 , \6132 , \6134 );
xor \U$5793 ( \6136 , \6127 , \6135 );
not \U$5794 ( \6137 , \6136 );
or \U$5795 ( \6138 , \6120 , \6137 );
or \U$5796 ( \6139 , \6136 , \6119 );
nand \U$5797 ( \6140 , \6138 , \6139 );
xnor \U$5798 ( \6141 , \6104 , \6140 );
not \U$5799 ( \6142 , \6141 );
not \U$5800 ( \6143 , \6142 );
buf \U$5801 ( \6144 , \796 );
buf \U$5802 ( \6145 , \6144 );
not \U$5803 ( \6146 , \6145 );
not \U$5804 ( \6147 , \5716 );
or \U$5805 ( \6148 , \6146 , \6147 );
xnor \U$5806 ( \6149 , RI98719b0_131, \1366 );
nand \U$5807 ( \6150 , \6149 , \793 );
nand \U$5808 ( \6151 , \6148 , \6150 );
not \U$5809 ( \6152 , \5642 );
not \U$5810 ( \6153 , \5644 );
not \U$5811 ( \6154 , \2982 );
or \U$5812 ( \6155 , \6153 , \6154 );
or \U$5813 ( \6156 , \1394 , \5644 );
nand \U$5814 ( \6157 , \6155 , \6156 );
not \U$5815 ( \6158 , \6157 );
or \U$5816 ( \6159 , \6152 , \6158 );
nand \U$5817 ( \6160 , \5650 , \5653 );
nand \U$5818 ( \6161 , \6159 , \6160 );
xor \U$5819 ( \6162 , \6151 , \6161 );
not \U$5820 ( \6163 , \4902 );
not \U$5821 ( \6164 , \1446 );
buf \U$5822 ( \6165 , \6164 );
not \U$5823 ( \6166 , \6165 );
or \U$5824 ( \6167 , \6163 , \6166 );
nand \U$5825 ( \6168 , \2492 , RI9872388_152);
nand \U$5826 ( \6169 , \6167 , \6168 );
not \U$5827 ( \6170 , \6169 );
not \U$5828 ( \6171 , \5942 );
or \U$5829 ( \6172 , \6170 , \6171 );
not \U$5830 ( \6173 , RI9872388_152);
not \U$5831 ( \6174 , \1415 );
not \U$5832 ( \6175 , \6174 );
or \U$5833 ( \6176 , \6173 , \6175 );
or \U$5834 ( \6177 , \1418 , RI9872388_152);
nand \U$5835 ( \6178 , \6176 , \6177 );
nand \U$5836 ( \6179 , \6178 , \5048 );
nand \U$5837 ( \6180 , \6172 , \6179 );
xor \U$5838 ( \6181 , \6162 , \6180 );
not \U$5839 ( \6182 , \1018 );
not \U$5840 ( \6183 , \3271 );
not \U$5841 ( \6184 , \5392 );
not \U$5842 ( \6185 , \6184 );
not \U$5843 ( \6186 , \6185 );
or \U$5844 ( \6187 , \6183 , \6186 );
or \U$5845 ( \6188 , \6185 , \3271 );
nand \U$5846 ( \6189 , \6187 , \6188 );
not \U$5847 ( \6190 , \6189 );
or \U$5848 ( \6191 , \6182 , \6190 );
nand \U$5849 ( \6192 , \5741 , \1013 );
nand \U$5850 ( \6193 , \6191 , \6192 );
not \U$5851 ( \6194 , \1380 );
not \U$5852 ( \6195 , \6194 );
not \U$5853 ( \6196 , \6195 );
not \U$5854 ( \6197 , RI9871e60_141);
not \U$5855 ( \6198 , \4990 );
or \U$5856 ( \6199 , \6197 , \6198 );
or \U$5857 ( \6200 , \4990 , RI9871e60_141);
nand \U$5858 ( \6201 , \6199 , \6200 );
not \U$5859 ( \6202 , \6201 );
or \U$5860 ( \6203 , \6196 , \6202 );
nand \U$5861 ( \6204 , \5627 , \1353 );
nand \U$5862 ( \6205 , \6203 , \6204 );
xor \U$5863 ( \6206 , \6193 , \6205 );
or \U$5864 ( \6207 , \5913 , \2086 );
and \U$5865 ( \6208 , RI9871aa0_133, \1658 );
not \U$5866 ( \6209 , RI9871aa0_133);
and \U$5867 ( \6210 , \6209 , \5719 );
nor \U$5868 ( \6211 , \6208 , \6210 );
or \U$5869 ( \6212 , \6211 , \2073 );
nand \U$5870 ( \6213 , \6207 , \6212 );
xor \U$5871 ( \6214 , \6206 , \6213 );
xor \U$5872 ( \6215 , \6181 , \6214 );
not \U$5873 ( \6216 , \3170 );
and \U$5874 ( \6217 , RI9872310_151, \820 );
not \U$5875 ( \6218 , RI9872310_151);
not \U$5876 ( \6219 , \820 );
and \U$5877 ( \6220 , \6218 , \6219 );
or \U$5878 ( \6221 , \6217 , \6220 );
not \U$5879 ( \6222 , \6221 );
or \U$5880 ( \6223 , \6216 , \6222 );
not \U$5881 ( \6224 , \846 );
buf \U$5882 ( \6225 , \6224 );
and \U$5883 ( \6226 , RI9872310_151, \6225 );
not \U$5884 ( \6227 , RI9872310_151);
and \U$5885 ( \6228 , \6227 , \847 );
or \U$5886 ( \6229 , \6226 , \6228 );
nand \U$5887 ( \6230 , \6229 , \3164 );
nand \U$5888 ( \6231 , \6223 , \6230 );
not \U$5889 ( \6232 , \1518 );
not \U$5890 ( \6233 , \5889 );
or \U$5891 ( \6234 , \6232 , \6233 );
not \U$5892 ( \6235 , \1800 );
not \U$5893 ( \6236 , \3240 );
or \U$5894 ( \6237 , \6235 , \6236 );
nand \U$5895 ( \6238 , \4370 , RI9871c80_137);
nand \U$5896 ( \6239 , \6237 , \6238 );
nand \U$5897 ( \6240 , \6239 , \1501 );
nand \U$5898 ( \6241 , \6234 , \6240 );
not \U$5899 ( \6242 , \876 );
xor \U$5900 ( \6243 , \4153 , RI9872130_147);
not \U$5901 ( \6244 , \6243 );
or \U$5902 ( \6245 , \6242 , \6244 );
nand \U$5903 ( \6246 , \5879 , \924 );
nand \U$5904 ( \6247 , \6245 , \6246 );
and \U$5905 ( \6248 , \6241 , \6247 );
not \U$5906 ( \6249 , \6241 );
not \U$5907 ( \6250 , \6247 );
and \U$5908 ( \6251 , \6249 , \6250 );
nor \U$5909 ( \6252 , \6248 , \6251 );
xor \U$5910 ( \6253 , \6231 , \6252 );
and \U$5911 ( \6254 , \6215 , \6253 );
and \U$5912 ( \6255 , \6181 , \6214 );
nor \U$5913 ( \6256 , \6254 , \6255 );
not \U$5914 ( \6257 , \6256 );
not \U$5915 ( \6258 , \6257 );
not \U$5916 ( \6259 , \6151 );
not \U$5917 ( \6260 , \6161 );
not \U$5918 ( \6261 , \6260 );
not \U$5919 ( \6262 , \6180 );
or \U$5920 ( \6263 , \6261 , \6262 );
or \U$5921 ( \6264 , \6180 , \6260 );
nand \U$5922 ( \6265 , \6263 , \6264 );
not \U$5923 ( \6266 , \6265 );
or \U$5924 ( \6267 , \6259 , \6266 );
nand \U$5925 ( \6268 , \6180 , \6161 );
nand \U$5926 ( \6269 , \6267 , \6268 );
not \U$5927 ( \6270 , \6269 );
xor \U$5928 ( \6271 , \6193 , \6205 );
and \U$5929 ( \6272 , \6271 , \6213 );
and \U$5930 ( \6273 , \6193 , \6205 );
or \U$5931 ( \6274 , \6272 , \6273 );
xor \U$5932 ( \6275 , RI9872928_164, RI98729a0_165);
not \U$5933 ( \6276 , \6275 );
and \U$5934 ( \6277 , RI98728b0_163, RI9872928_164);
not \U$5935 ( \6278 , RI98728b0_163);
not \U$5936 ( \6279 , RI9872928_164);
and \U$5937 ( \6280 , \6278 , \6279 );
nor \U$5938 ( \6281 , \6277 , \6280 );
and \U$5939 ( \6282 , \6276 , \6281 );
not \U$5940 ( \6283 , \6282 );
not \U$5941 ( \6284 , \6283 );
buf \U$5942 ( \6285 , \6275 );
buf \U$5943 ( \6286 , \6285 );
or \U$5944 ( \6287 , \6284 , \6286 );
nand \U$5945 ( \6288 , \6287 , RI98728b0_163);
buf \U$5946 ( \6289 , \660 );
nor \U$5947 ( \6290 , \5692 , \6289 );
nand \U$5948 ( \6291 , \654 , \663 );
and \U$5949 ( \6292 , \6290 , \6291 );
not \U$5950 ( \6293 , \6290 );
not \U$5951 ( \6294 , \6291 );
and \U$5952 ( \6295 , \6293 , \6294 );
nor \U$5953 ( \6296 , \6292 , \6295 );
not \U$5954 ( \6297 , \6296 );
not \U$5955 ( \6298 , \6297 );
and \U$5956 ( \6299 , \4708 , \6298 );
xor \U$5957 ( \6300 , \6288 , \6299 );
not \U$5958 ( \6301 , \1162 );
not \U$5959 ( \6302 , \4708 );
buf \U$5960 ( \6303 , \5703 );
buf \U$5961 ( \6304 , \6303 );
not \U$5962 ( \6305 , \6304 );
not \U$5963 ( \6306 , \6305 );
or \U$5964 ( \6307 , \6302 , \6306 );
buf \U$5965 ( \6308 , \5704 );
not \U$5966 ( \6309 , \6308 );
nand \U$5967 ( \6310 , \6309 , \1199 );
nand \U$5968 ( \6311 , \6307 , \6310 );
not \U$5969 ( \6312 , \6311 );
or \U$5970 ( \6313 , \6301 , \6312 );
not \U$5971 ( \6314 , \5768 );
not \U$5972 ( \6315 , \1219 );
buf \U$5973 ( \6316 , \6315 );
nand \U$5974 ( \6317 , \6314 , \6316 );
nand \U$5975 ( \6318 , \6313 , \6317 );
and \U$5976 ( \6319 , \6300 , \6318 );
and \U$5977 ( \6320 , \6288 , \6299 );
or \U$5978 ( \6321 , \6319 , \6320 );
not \U$5979 ( \6322 , \6321 );
xor \U$5980 ( \6323 , \6274 , \6322 );
not \U$5981 ( \6324 , \6323 );
and \U$5982 ( \6325 , \6270 , \6324 );
and \U$5983 ( \6326 , \6269 , \6323 );
nor \U$5984 ( \6327 , \6325 , \6326 );
not \U$5985 ( \6328 , \6327 );
not \U$5986 ( \6329 , \1083 );
not \U$5987 ( \6330 , \1038 );
and \U$5988 ( \6331 , RI98718c0_129, \6330 );
not \U$5989 ( \6332 , RI98718c0_129);
not \U$5990 ( \6333 , \1037 );
not \U$5991 ( \6334 , \6333 );
and \U$5992 ( \6335 , \6332 , \6334 );
or \U$5993 ( \6336 , \6331 , \6335 );
not \U$5994 ( \6337 , \6336 );
or \U$5995 ( \6338 , \6329 , \6337 );
nand \U$5996 ( \6339 , \5808 , \1136 );
nand \U$5997 ( \6340 , \6338 , \6339 );
not \U$5998 ( \6341 , \6340 );
not \U$5999 ( \6342 , \1455 );
and \U$6000 ( \6343 , RI9871c08_136, \3396 );
not \U$6001 ( \6344 , RI9871c08_136);
and \U$6002 ( \6345 , \6344 , \5947 );
or \U$6003 ( \6346 , \6343 , \6345 );
not \U$6004 ( \6347 , \6346 );
or \U$6005 ( \6348 , \6342 , \6347 );
nand \U$6006 ( \6349 , \6025 , \1430 );
nand \U$6007 ( \6350 , \6348 , \6349 );
not \U$6008 ( \6351 , \6350 );
or \U$6009 ( \6352 , \6341 , \6351 );
or \U$6010 ( \6353 , \6340 , \6350 );
not \U$6011 ( \6354 , \5847 );
not \U$6012 ( \6355 , \6044 );
or \U$6013 ( \6356 , \6354 , \6355 );
and \U$6014 ( \6357 , RI98725e0_157, \1834 );
not \U$6015 ( \6358 , RI98725e0_157);
and \U$6016 ( \6359 , \6358 , \1275 );
or \U$6017 ( \6360 , \6357 , \6359 );
nand \U$6018 ( \6361 , \6360 , \4103 );
nand \U$6019 ( \6362 , \6356 , \6361 );
nand \U$6020 ( \6363 , \6353 , \6362 );
nand \U$6021 ( \6364 , \6352 , \6363 );
not \U$6022 ( \6365 , \6241 );
nand \U$6023 ( \6366 , \6365 , \6250 );
not \U$6024 ( \6367 , \6366 );
not \U$6025 ( \6368 , \6231 );
or \U$6026 ( \6369 , \6367 , \6368 );
nand \U$6027 ( \6370 , \6241 , \6247 );
nand \U$6028 ( \6371 , \6369 , \6370 );
and \U$6029 ( \6372 , \6364 , \6371 );
not \U$6030 ( \6373 , \6364 );
not \U$6031 ( \6374 , \6371 );
and \U$6032 ( \6375 , \6373 , \6374 );
nor \U$6033 ( \6376 , \6372 , \6375 );
not \U$6034 ( \6377 , \1292 );
not \U$6035 ( \6378 , \2110 );
xnor \U$6036 ( \6379 , \6378 , RI9871b18_134);
not \U$6037 ( \6380 , \6379 );
or \U$6038 ( \6381 , \6377 , \6380 );
not \U$6039 ( \6382 , \1485 );
and \U$6040 ( \6383 , RI9871b18_134, \6382 );
not \U$6041 ( \6384 , RI9871b18_134);
and \U$6042 ( \6385 , \6384 , \1485 );
nor \U$6043 ( \6386 , \6383 , \6385 );
nand \U$6044 ( \6387 , \6386 , \1323 );
nand \U$6045 ( \6388 , \6381 , \6387 );
not \U$6046 ( \6389 , \5796 );
not \U$6047 ( \6390 , \5787 );
or \U$6048 ( \6391 , \6389 , \6390 );
and \U$6049 ( \6392 , RI9872478_154, \1097 );
not \U$6050 ( \6393 , RI9872478_154);
and \U$6051 ( \6394 , \6393 , \1106 );
or \U$6052 ( \6395 , \6392 , \6394 );
nand \U$6053 ( \6396 , \6395 , \5034 );
nand \U$6054 ( \6397 , \6391 , \6396 );
xor \U$6055 ( \6398 , \6388 , \6397 );
not \U$6056 ( \6399 , \3600 );
not \U$6057 ( \6400 , \1505 );
and \U$6058 ( \6401 , \6400 , RI98726d0_159);
not \U$6059 ( \6402 , \6400 );
and \U$6060 ( \6403 , \6402 , \4063 );
nor \U$6061 ( \6404 , \6401 , \6403 );
not \U$6062 ( \6405 , \6404 );
or \U$6063 ( \6406 , \6399 , \6405 );
nand \U$6064 ( \6407 , \6035 , \3467 );
nand \U$6065 ( \6408 , \6406 , \6407 );
and \U$6066 ( \6409 , \6398 , \6408 );
and \U$6067 ( \6410 , \6388 , \6397 );
or \U$6068 ( \6411 , \6409 , \6410 );
buf \U$6069 ( \6412 , \6411 );
and \U$6070 ( \6413 , \6376 , \6412 );
not \U$6071 ( \6414 , \6376 );
not \U$6072 ( \6415 , \6412 );
and \U$6073 ( \6416 , \6414 , \6415 );
nor \U$6074 ( \6417 , \6413 , \6416 );
not \U$6075 ( \6418 , \6417 );
or \U$6076 ( \6419 , \6328 , \6418 );
or \U$6077 ( \6420 , \6417 , \6327 );
nand \U$6078 ( \6421 , \6419 , \6420 );
not \U$6079 ( \6422 , \6421 );
or \U$6080 ( \6423 , \6258 , \6422 );
not \U$6081 ( \6424 , \6327 );
nand \U$6082 ( \6425 , \6424 , \6417 );
nand \U$6083 ( \6426 , \6423 , \6425 );
not \U$6084 ( \6427 , \6426 );
not \U$6085 ( \6428 , \924 );
not \U$6086 ( \6429 , \5518 );
or \U$6087 ( \6430 , \6428 , \6429 );
buf \U$6088 ( \6431 , \875 );
nand \U$6089 ( \6432 , \5871 , \6431 );
nand \U$6090 ( \6433 , \6430 , \6432 );
not \U$6091 ( \6434 , \1518 );
not \U$6092 ( \6435 , \5501 );
or \U$6093 ( \6436 , \6434 , \6435 );
nand \U$6094 ( \6437 , \5894 , \1501 );
nand \U$6095 ( \6438 , \6436 , \6437 );
xor \U$6096 ( \6439 , \6433 , \6438 );
not \U$6097 ( \6440 , \3164 );
not \U$6098 ( \6441 , \3154 );
not \U$6099 ( \6442 , \891 );
buf \U$6100 ( \6443 , \6442 );
not \U$6101 ( \6444 , \6443 );
not \U$6102 ( \6445 , \6444 );
or \U$6103 ( \6446 , \6441 , \6445 );
nand \U$6104 ( \6447 , \893 , RI9872310_151);
nand \U$6105 ( \6448 , \6446 , \6447 );
not \U$6106 ( \6449 , \6448 );
or \U$6107 ( \6450 , \6440 , \6449 );
not \U$6108 ( \6451 , \5481 );
nand \U$6109 ( \6452 , \6451 , \3170 );
nand \U$6110 ( \6453 , \6450 , \6452 );
xor \U$6111 ( \6454 , \6439 , \6453 );
not \U$6112 ( \6455 , \6364 );
not \U$6113 ( \6456 , \6411 );
or \U$6114 ( \6457 , \6455 , \6456 );
or \U$6115 ( \6458 , \6411 , \6364 );
nand \U$6116 ( \6459 , \6458 , \6371 );
nand \U$6117 ( \6460 , \6457 , \6459 );
and \U$6118 ( \6461 , \6454 , \6460 );
not \U$6119 ( \6462 , \6454 );
not \U$6120 ( \6463 , \6460 );
and \U$6121 ( \6464 , \6462 , \6463 );
nor \U$6122 ( \6465 , \6461 , \6464 );
not \U$6123 ( \6466 , \6323 );
not \U$6124 ( \6467 , \6466 );
not \U$6125 ( \6468 , \6269 );
or \U$6126 ( \6469 , \6467 , \6468 );
not \U$6127 ( \6470 , \6322 );
nand \U$6128 ( \6471 , \6470 , \6274 );
nand \U$6129 ( \6472 , \6469 , \6471 );
xnor \U$6130 ( \6473 , \6465 , \6472 );
not \U$6131 ( \6474 , \6473 );
not \U$6132 ( \6475 , \1013 );
not \U$6133 ( \6476 , \6189 );
or \U$6134 ( \6477 , \6475 , \6476 );
and \U$6135 ( \6478 , \1043 , \6060 );
not \U$6136 ( \6479 , \1043 );
not \U$6137 ( \6480 , \5760 );
not \U$6138 ( \6481 , \6480 );
and \U$6139 ( \6482 , \6479 , \6481 );
nor \U$6140 ( \6483 , \6478 , \6482 );
or \U$6141 ( \6484 , \6483 , \1612 );
nand \U$6142 ( \6485 , \6477 , \6484 );
not \U$6143 ( \6486 , \1353 );
not \U$6144 ( \6487 , \6201 );
or \U$6145 ( \6488 , \6486 , \6487 );
and \U$6146 ( \6489 , RI9871e60_141, \5736 );
not \U$6147 ( \6490 , RI9871e60_141);
and \U$6148 ( \6491 , \6490 , \5739 );
or \U$6149 ( \6492 , \6489 , \6491 );
nand \U$6150 ( \6493 , \6492 , \6195 );
nand \U$6151 ( \6494 , \6488 , \6493 );
xor \U$6152 ( \6495 , \6485 , \6494 );
not \U$6153 ( \6496 , \5642 );
not \U$6154 ( \6497 , RI9872568_156);
not \U$6155 ( \6498 , \1127 );
or \U$6156 ( \6499 , \6497 , \6498 );
or \U$6157 ( \6500 , \1725 , RI9872568_156);
nand \U$6158 ( \6501 , \6499 , \6500 );
not \U$6159 ( \6502 , \6501 );
or \U$6160 ( \6503 , \6496 , \6502 );
nand \U$6161 ( \6504 , \6157 , \5653 );
nand \U$6162 ( \6505 , \6503 , \6504 );
and \U$6163 ( \6506 , \6495 , \6505 );
and \U$6164 ( \6507 , \6485 , \6494 );
or \U$6165 ( \6508 , \6506 , \6507 );
not \U$6166 ( \6509 , \6508 );
not \U$6167 ( \6510 , \562 );
not \U$6168 ( \6511 , \6510 );
not \U$6169 ( \6512 , \5665 );
not \U$6170 ( \6513 , \6512 );
not \U$6171 ( \6514 , \5683 );
or \U$6172 ( \6515 , \6513 , \6514 );
not \U$6173 ( \6516 , \5690 );
nand \U$6174 ( \6517 , \6515 , \6516 );
not \U$6175 ( \6518 , \6517 );
or \U$6176 ( \6519 , \6511 , \6518 );
buf \U$6177 ( \6520 , \657 );
nand \U$6178 ( \6521 , \6519 , \6520 );
xor \U$6179 ( \6522 , RI98717d0_127, RI9871848_128);
and \U$6180 ( \6523 , \6521 , \6522 );
not \U$6181 ( \6524 , \6521 );
not \U$6182 ( \6525 , \6522 );
and \U$6183 ( \6526 , \6524 , \6525 );
nor \U$6184 ( \6527 , \6523 , \6526 );
buf \U$6185 ( \6528 , \6527 );
not \U$6186 ( \6529 , \6528 );
not \U$6187 ( \6530 , \6529 );
and \U$6188 ( \6531 , \4708 , \6530 );
not \U$6189 ( \6532 , \1220 );
not \U$6190 ( \6533 , \6311 );
or \U$6191 ( \6534 , \6532 , \6533 );
xor \U$6192 ( \6535 , \4708 , \6298 );
nand \U$6193 ( \6536 , \6535 , \1162 );
nand \U$6194 ( \6537 , \6534 , \6536 );
xor \U$6195 ( \6538 , \6531 , \6537 );
not \U$6196 ( \6539 , \6538 );
not \U$6197 ( \6540 , \2074 );
xnor \U$6198 ( \6541 , RI9871aa0_133, \1344 );
not \U$6199 ( \6542 , \6541 );
or \U$6200 ( \6543 , \6540 , \6542 );
not \U$6201 ( \6544 , \6211 );
nand \U$6202 ( \6545 , \6544 , \2087 );
nand \U$6203 ( \6546 , \6543 , \6545 );
not \U$6204 ( \6547 , \6546 );
or \U$6205 ( \6548 , \6539 , \6547 );
nand \U$6206 ( \6549 , \6537 , \6531 );
nand \U$6207 ( \6550 , \6548 , \6549 );
not \U$6208 ( \6551 , \6550 );
not \U$6209 ( \6552 , \6551 );
buf \U$6210 ( \6553 , \4919 );
not \U$6211 ( \6554 , \6553 );
not \U$6212 ( \6555 , RI9872388_152);
not \U$6213 ( \6556 , \2038 );
or \U$6214 ( \6557 , \6555 , \6556 );
not \U$6215 ( \6558 , RI9872388_152);
nand \U$6216 ( \6559 , \6558 , \1740 );
nand \U$6217 ( \6560 , \6557 , \6559 );
not \U$6218 ( \6561 , \6560 );
or \U$6219 ( \6562 , \6554 , \6561 );
nand \U$6220 ( \6563 , \6169 , \5048 );
nand \U$6221 ( \6564 , \6562 , \6563 );
not \U$6222 ( \6565 , \6145 );
not \U$6223 ( \6566 , \6149 );
or \U$6224 ( \6567 , \6565 , \6566 );
not \U$6225 ( \6568 , RI98719b0_131);
not \U$6226 ( \6569 , \6568 );
not \U$6227 ( \6570 , \1713 );
or \U$6228 ( \6571 , \6569 , \6570 );
not \U$6229 ( \6572 , \1060 );
not \U$6230 ( \6573 , \6572 );
not \U$6231 ( \6574 , RI98719b0_131);
or \U$6232 ( \6575 , \6573 , \6574 );
nand \U$6233 ( \6576 , \6571 , \6575 );
nand \U$6234 ( \6577 , \6576 , \793 );
nand \U$6235 ( \6578 , \6567 , \6577 );
or \U$6236 ( \6579 , \6564 , \6578 );
not \U$6237 ( \6580 , \4085 );
not \U$6238 ( \6581 , \6360 );
or \U$6239 ( \6582 , \6580 , \6581 );
and \U$6240 ( \6583 , RI98725e0_157, \917 );
not \U$6241 ( \6584 , RI98725e0_157);
buf \U$6242 ( \6585 , \914 );
and \U$6243 ( \6586 , \6584 , \6585 );
nor \U$6244 ( \6587 , \6583 , \6586 );
nand \U$6245 ( \6588 , \6587 , \4103 );
nand \U$6246 ( \6589 , \6582 , \6588 );
nand \U$6247 ( \6590 , \6579 , \6589 );
nand \U$6248 ( \6591 , \6564 , \6578 );
nand \U$6249 ( \6592 , \6590 , \6591 );
not \U$6250 ( \6593 , \6592 );
or \U$6251 ( \6594 , \6552 , \6593 );
nand \U$6252 ( \6595 , \6550 , \6590 , \6591 );
nand \U$6253 ( \6596 , \6594 , \6595 );
not \U$6254 ( \6597 , \6596 );
or \U$6255 ( \6598 , \6509 , \6597 );
nand \U$6256 ( \6599 , \6592 , \6550 );
nand \U$6257 ( \6600 , \6598 , \6599 );
not \U$6258 ( \6601 , \6600 );
not \U$6259 ( \6602 , \6284 );
and \U$6260 ( \6603 , RI98728b0_163, \1690 );
not \U$6261 ( \6604 , RI98728b0_163);
and \U$6262 ( \6605 , \6604 , \779 );
nor \U$6263 ( \6606 , \6603 , \6605 );
not \U$6264 ( \6607 , \6606 );
or \U$6265 ( \6608 , \6602 , \6607 );
not \U$6266 ( \6609 , \6285 );
not \U$6267 ( \6610 , \6609 );
buf \U$6268 ( \6611 , \6610 );
nand \U$6269 ( \6612 , \6611 , RI98728b0_163);
nand \U$6270 ( \6613 , \6608 , \6612 );
not \U$6271 ( \6614 , \832 );
not \U$6272 ( \6615 , \5601 );
or \U$6273 ( \6616 , \6614 , \6615 );
not \U$6274 ( \6617 , \5208 );
and \U$6275 ( \6618 , RI9871d70_139, \6617 );
not \U$6276 ( \6619 , RI9871d70_139);
and \U$6277 ( \6620 , \6619 , \4409 );
or \U$6278 ( \6621 , \6618 , \6620 );
nand \U$6279 ( \6622 , \6621 , \859 );
nand \U$6280 ( \6623 , \6616 , \6622 );
xor \U$6281 ( \6624 , \6613 , \6623 );
xor \U$6282 ( \6625 , \6288 , \6299 );
xor \U$6283 ( \6626 , \6625 , \6318 );
and \U$6284 ( \6627 , \6624 , \6626 );
and \U$6285 ( \6628 , \6613 , \6623 );
nor \U$6286 ( \6629 , \6627 , \6628 );
not \U$6287 ( \6630 , \6629 );
not \U$6288 ( \6631 , \832 );
not \U$6289 ( \6632 , \6621 );
or \U$6290 ( \6633 , \6631 , \6632 );
xor \U$6291 ( \6634 , \4472 , RI9871d70_139);
not \U$6292 ( \6635 , \5351 );
nand \U$6293 ( \6636 , \6634 , \6635 );
nand \U$6294 ( \6637 , \6633 , \6636 );
not \U$6295 ( \6638 , \876 );
and \U$6296 ( \6639 , \5596 , \919 );
not \U$6297 ( \6640 , \5596 );
and \U$6298 ( \6641 , \6640 , RI9872130_147);
nor \U$6299 ( \6642 , \6639 , \6641 );
not \U$6300 ( \6643 , \6642 );
or \U$6301 ( \6644 , \6638 , \6643 );
nand \U$6302 ( \6645 , \6243 , \924 );
nand \U$6303 ( \6646 , \6644 , \6645 );
xor \U$6304 ( \6647 , \6637 , \6646 );
not \U$6305 ( \6648 , \3170 );
not \U$6306 ( \6649 , \6229 );
or \U$6307 ( \6650 , \6648 , \6649 );
not \U$6308 ( \6651 , \5907 );
xor \U$6309 ( \6652 , RI9872310_151, \6651 );
buf \U$6310 ( \6653 , \3163 );
nand \U$6311 ( \6654 , \6652 , \6653 );
nand \U$6312 ( \6655 , \6650 , \6654 );
and \U$6313 ( \6656 , \6647 , \6655 );
and \U$6314 ( \6657 , \6637 , \6646 );
or \U$6315 ( \6658 , \6656 , \6657 );
not \U$6316 ( \6659 , \6658 );
not \U$6317 ( \6660 , \1430 );
not \U$6318 ( \6661 , \6346 );
or \U$6319 ( \6662 , \6660 , \6661 );
not \U$6320 ( \6663 , \1850 );
not \U$6321 ( \6664 , \1486 );
or \U$6322 ( \6665 , \6663 , \6664 );
or \U$6323 ( \6666 , \2118 , \1850 );
nand \U$6324 ( \6667 , \6665 , \6666 );
nand \U$6325 ( \6668 , \6667 , \1456 );
nand \U$6326 ( \6669 , \6662 , \6668 );
not \U$6327 ( \6670 , \6669 );
not \U$6328 ( \6671 , \1134 );
not \U$6329 ( \6672 , \6671 );
buf \U$6330 ( \6673 , \6672 );
not \U$6331 ( \6674 , \6673 );
not \U$6332 ( \6675 , \6336 );
or \U$6333 ( \6676 , \6674 , \6675 );
not \U$6334 ( \6677 , RI98718c0_129);
not \U$6335 ( \6678 , \3126 );
not \U$6336 ( \6679 , \6678 );
or \U$6337 ( \6680 , \6677 , \6679 );
nand \U$6338 ( \6681 , \6020 , \1111 );
nand \U$6339 ( \6682 , \6680 , \6681 );
nand \U$6340 ( \6683 , \6682 , \1083 );
nand \U$6341 ( \6684 , \6676 , \6683 );
not \U$6342 ( \6685 , \6684 );
or \U$6343 ( \6686 , \6670 , \6685 );
or \U$6344 ( \6687 , \6669 , \6684 );
not \U$6345 ( \6688 , \5034 );
not \U$6346 ( \6689 , RI9872478_154);
not \U$6347 ( \6690 , \6174 );
or \U$6348 ( \6691 , \6689 , \6690 );
not \U$6349 ( \6692 , \1415 );
not \U$6350 ( \6693 , \6692 );
nand \U$6351 ( \6694 , \6693 , \5025 );
nand \U$6352 ( \6695 , \6691 , \6694 );
not \U$6353 ( \6696 , \6695 );
or \U$6354 ( \6697 , \6688 , \6696 );
buf \U$6355 ( \6698 , \5036 );
nand \U$6356 ( \6699 , \6395 , \6698 );
nand \U$6357 ( \6700 , \6697 , \6699 );
nand \U$6358 ( \6701 , \6687 , \6700 );
nand \U$6359 ( \6702 , \6686 , \6701 );
not \U$6360 ( \6703 , \1323 );
not \U$6361 ( \6704 , \6379 );
or \U$6362 ( \6705 , \6703 , \6704 );
and \U$6363 ( \6706 , RI9871b18_134, \3691 );
not \U$6364 ( \6707 , RI9871b18_134);
and \U$6365 ( \6708 , \6707 , \5884 );
or \U$6366 ( \6709 , \6706 , \6708 );
nand \U$6367 ( \6710 , \6709 , \1292 );
nand \U$6368 ( \6711 , \6705 , \6710 );
not \U$6369 ( \6712 , \1518 );
not \U$6370 ( \6713 , \6239 );
or \U$6371 ( \6714 , \6712 , \6713 );
not \U$6372 ( \6715 , \1584 );
not \U$6373 ( \6716 , \3537 );
or \U$6374 ( \6717 , \6715 , \6716 );
not \U$6375 ( \6718 , \3541 );
or \U$6376 ( \6719 , \6718 , \1584 );
nand \U$6377 ( \6720 , \6717 , \6719 );
nand \U$6378 ( \6721 , \6720 , \1501 );
nand \U$6379 ( \6722 , \6714 , \6721 );
or \U$6380 ( \6723 , \6711 , \6722 );
not \U$6381 ( \6724 , \6723 );
not \U$6382 ( \6725 , \3467 );
not \U$6383 ( \6726 , \6404 );
or \U$6384 ( \6727 , \6725 , \6726 );
xnor \U$6385 ( \6728 , RI98726d0_159, \820 );
nand \U$6386 ( \6729 , \6728 , \3466 );
nand \U$6387 ( \6730 , \6727 , \6729 );
not \U$6388 ( \6731 , \6730 );
or \U$6389 ( \6732 , \6724 , \6731 );
nand \U$6390 ( \6733 , \6711 , \6722 );
nand \U$6391 ( \6734 , \6732 , \6733 );
and \U$6392 ( \6735 , \6702 , \6734 );
not \U$6393 ( \6736 , \6702 );
not \U$6394 ( \6737 , \6734 );
and \U$6395 ( \6738 , \6736 , \6737 );
nor \U$6396 ( \6739 , \6735 , \6738 );
not \U$6397 ( \6740 , \6739 );
or \U$6398 ( \6741 , \6659 , \6740 );
nand \U$6399 ( \6742 , \6734 , \6702 );
nand \U$6400 ( \6743 , \6741 , \6742 );
not \U$6401 ( \6744 , \6743 );
or \U$6402 ( \6745 , \6630 , \6744 );
or \U$6403 ( \6746 , \6743 , \6629 );
nand \U$6404 ( \6747 , \6745 , \6746 );
not \U$6405 ( \6748 , \6747 );
or \U$6406 ( \6749 , \6601 , \6748 );
not \U$6407 ( \6750 , \6629 );
nand \U$6408 ( \6751 , \6750 , \6743 );
nand \U$6409 ( \6752 , \6749 , \6751 );
not \U$6410 ( \6753 , \6752 );
or \U$6411 ( \6754 , \6474 , \6753 );
or \U$6412 ( \6755 , \6752 , \6473 );
nand \U$6413 ( \6756 , \6754 , \6755 );
not \U$6414 ( \6757 , \6756 );
or \U$6415 ( \6758 , \6427 , \6757 );
not \U$6416 ( \6759 , \6473 );
nand \U$6417 ( \6760 , \6759 , \6752 );
nand \U$6418 ( \6761 , \6758 , \6760 );
not \U$6419 ( \6762 , \6761 );
xor \U$6420 ( \6763 , \6027 , \6037 );
xor \U$6421 ( \6764 , \6763 , \6050 );
xor \U$6422 ( \6765 , \5882 , \5917 );
xor \U$6423 ( \6766 , \6764 , \6765 );
not \U$6424 ( \6767 , \4925 );
not \U$6425 ( \6768 , \5941 );
or \U$6426 ( \6769 , \6767 , \6768 );
nand \U$6427 ( \6770 , \4920 , \6178 );
nand \U$6428 ( \6771 , \6769 , \6770 );
not \U$6429 ( \6772 , \6386 );
not \U$6430 ( \6773 , \1292 );
or \U$6431 ( \6774 , \6772 , \6773 );
not \U$6432 ( \6775 , \5950 );
or \U$6433 ( \6776 , \6775 , \1543 );
nand \U$6434 ( \6777 , \6774 , \6776 );
xor \U$6435 ( \6778 , \6771 , \6777 );
not \U$6436 ( \6779 , \3164 );
not \U$6437 ( \6780 , \6221 );
or \U$6438 ( \6781 , \6779 , \6780 );
not \U$6439 ( \6782 , \6448 );
or \U$6440 ( \6783 , \6782 , \4261 );
nand \U$6441 ( \6784 , \6781 , \6783 );
xor \U$6442 ( \6785 , \6778 , \6784 );
and \U$6443 ( \6786 , \6766 , \6785 );
and \U$6444 ( \6787 , \6764 , \6765 );
or \U$6445 ( \6788 , \6786 , \6787 );
not \U$6446 ( \6789 , \6788 );
xor \U$6447 ( \6790 , \6771 , \6777 );
and \U$6448 ( \6791 , \6790 , \6784 );
and \U$6449 ( \6792 , \6771 , \6777 );
or \U$6450 ( \6793 , \6791 , \6792 );
xnor \U$6451 ( \6794 , \6076 , \6069 );
xnor \U$6452 ( \6795 , \5925 , \6794 );
xnor \U$6453 ( \6796 , \6793 , \6795 );
nand \U$6454 ( \6797 , \6789 , \6796 );
not \U$6455 ( \6798 , \6797 );
and \U$6456 ( \6799 , \6053 , \6007 );
not \U$6457 ( \6800 , \6053 );
and \U$6458 ( \6801 , \6800 , \6006 );
or \U$6459 ( \6802 , \6799 , \6801 );
and \U$6460 ( \6803 , \6802 , \6013 );
not \U$6461 ( \6804 , \6802 );
and \U$6462 ( \6805 , \6804 , \6014 );
nor \U$6463 ( \6806 , \6803 , \6805 );
not \U$6464 ( \6807 , \6806 );
or \U$6465 ( \6808 , \6798 , \6807 );
not \U$6466 ( \6809 , \6796 );
nand \U$6467 ( \6810 , \6809 , \6788 );
nand \U$6468 ( \6811 , \6808 , \6810 );
not \U$6469 ( \6812 , \6811 );
not \U$6470 ( \6813 , \6812 );
not \U$6471 ( \6814 , \6472 );
not \U$6472 ( \6815 , \6465 );
or \U$6473 ( \6816 , \6814 , \6815 );
not \U$6474 ( \6817 , \6463 );
nand \U$6475 ( \6818 , \6817 , \6454 );
nand \U$6476 ( \6819 , \6816 , \6818 );
not \U$6477 ( \6820 , \6795 );
not \U$6478 ( \6821 , \6793 );
or \U$6479 ( \6822 , \6820 , \6821 );
nand \U$6480 ( \6823 , \6794 , \5655 );
nand \U$6481 ( \6824 , \6822 , \6823 );
xor \U$6482 ( \6825 , \5522 , \5532 );
xor \U$6483 ( \6826 , \6825 , \5539 );
nor \U$6484 ( \6827 , \6824 , \6826 );
not \U$6485 ( \6828 , \6827 );
nand \U$6486 ( \6829 , \6824 , \6826 );
nand \U$6487 ( \6830 , \6828 , \6829 );
or \U$6488 ( \6831 , \5825 , \1612 );
or \U$6489 ( \6832 , \5210 , \1068 );
nand \U$6490 ( \6833 , \6831 , \6832 );
xor \U$6491 ( \6834 , \6833 , \5200 );
xor \U$6492 ( \6835 , \6433 , \6438 );
and \U$6493 ( \6836 , \6835 , \6453 );
and \U$6494 ( \6837 , \6433 , \6438 );
or \U$6495 ( \6838 , \6836 , \6837 );
xor \U$6496 ( \6839 , \6834 , \6838 );
and \U$6497 ( \6840 , \6830 , \6839 );
not \U$6498 ( \6841 , \6830 );
not \U$6499 ( \6842 , \6839 );
and \U$6500 ( \6843 , \6841 , \6842 );
nor \U$6501 ( \6844 , \6840 , \6843 );
and \U$6502 ( \6845 , \6819 , \6844 );
not \U$6503 ( \6846 , \6819 );
not \U$6504 ( \6847 , \6844 );
and \U$6505 ( \6848 , \6846 , \6847 );
or \U$6506 ( \6849 , \6845 , \6848 );
not \U$6507 ( \6850 , \6849 );
and \U$6508 ( \6851 , \6813 , \6850 );
and \U$6509 ( \6852 , \6849 , \6812 );
nor \U$6510 ( \6853 , \6851 , \6852 );
not \U$6511 ( \6854 , \6853 );
or \U$6512 ( \6855 , \6762 , \6854 );
or \U$6513 ( \6856 , \6761 , \6853 );
nand \U$6514 ( \6857 , \6855 , \6856 );
not \U$6515 ( \6858 , \6857 );
or \U$6516 ( \6859 , \6143 , \6858 );
not \U$6517 ( \6860 , \6853 );
nand \U$6518 ( \6861 , \6860 , \6761 );
nand \U$6519 ( \6862 , \6859 , \6861 );
xor \U$6520 ( \6863 , \5467 , \5468 );
xor \U$6521 ( \6864 , \6863 , \5471 );
not \U$6522 ( \6865 , \6118 );
not \U$6523 ( \6866 , \6116 );
or \U$6524 ( \6867 , \6865 , \6866 );
not \U$6525 ( \6868 , \6106 );
nand \U$6526 ( \6869 , \6868 , \6112 );
nand \U$6527 ( \6870 , \6867 , \6869 );
xor \U$6528 ( \6871 , \6864 , \6870 );
not \U$6529 ( \6872 , \5977 );
not \U$6530 ( \6873 , \6872 );
not \U$6531 ( \6874 , \5994 );
or \U$6532 ( \6875 , \6873 , \6874 );
nand \U$6533 ( \6876 , \5993 , \5983 );
nand \U$6534 ( \6877 , \6875 , \6876 );
not \U$6535 ( \6878 , \6877 );
xnor \U$6536 ( \6879 , \6871 , \6878 );
xor \U$6537 ( \6880 , \6086 , \6082 );
not \U$6538 ( \6881 , \6092 );
and \U$6539 ( \6882 , \6880 , \6881 );
and \U$6540 ( \6883 , \6086 , \6082 );
or \U$6541 ( \6884 , \6882 , \6883 );
not \U$6542 ( \6885 , \6884 );
not \U$6543 ( \6886 , \5342 );
not \U$6544 ( \6887 , \5420 );
or \U$6545 ( \6888 , \6886 , \6887 );
or \U$6546 ( \6889 , \5420 , \5342 );
nand \U$6547 ( \6890 , \6888 , \6889 );
xor \U$6548 ( \6891 , \6885 , \6890 );
xor \U$6549 ( \6892 , \5477 , \5542 );
xor \U$6550 ( \6893 , \6892 , \5513 );
xor \U$6551 ( \6894 , \6891 , \6893 );
xor \U$6552 ( \6895 , \6879 , \6894 );
not \U$6553 ( \6896 , \6119 );
not \U$6554 ( \6897 , \6896 );
not \U$6555 ( \6898 , \6136 );
or \U$6556 ( \6899 , \6897 , \6898 );
nand \U$6557 ( \6900 , \6127 , \6135 );
nand \U$6558 ( \6901 , \6899 , \6900 );
xnor \U$6559 ( \6902 , \6895 , \6901 );
not \U$6560 ( \6903 , \6902 );
or \U$6561 ( \6904 , \6862 , \6903 );
not \U$6562 ( \6905 , \6849 );
not \U$6563 ( \6906 , \6811 );
or \U$6564 ( \6907 , \6905 , \6906 );
nand \U$6565 ( \6908 , \6847 , \6819 );
nand \U$6566 ( \6909 , \6907 , \6908 );
or \U$6567 ( \6910 , \6827 , \6842 );
nand \U$6568 ( \6911 , \6910 , \6829 );
xor \U$6569 ( \6912 , \4827 , \4835 );
xor \U$6570 ( \6913 , \6912 , \4849 );
xor \U$6571 ( \6914 , \6833 , \5200 );
and \U$6572 ( \6915 , \6914 , \6838 );
and \U$6573 ( \6916 , \6833 , \5200 );
or \U$6574 ( \6917 , \6915 , \6916 );
xor \U$6575 ( \6918 , \6913 , \6917 );
xor \U$6576 ( \6919 , \4786 , \4800 );
xor \U$6577 ( \6920 , \6919 , \4811 );
xor \U$6578 ( \6921 , \6918 , \6920 );
xor \U$6579 ( \6922 , \6911 , \6921 );
not \U$6580 ( \6923 , \5998 );
not \U$6581 ( \6924 , \6097 );
or \U$6582 ( \6925 , \6923 , \6924 );
not \U$6583 ( \6926 , \6093 );
nand \U$6584 ( \6927 , \6926 , \6056 );
nand \U$6585 ( \6928 , \6925 , \6927 );
xor \U$6586 ( \6929 , \6922 , \6928 );
xor \U$6587 ( \6930 , \6909 , \6929 );
not \U$6588 ( \6931 , \6140 );
not \U$6589 ( \6932 , \6104 );
or \U$6590 ( \6933 , \6931 , \6932 );
not \U$6591 ( \6934 , \5975 );
nand \U$6592 ( \6935 , \6934 , \6103 );
nand \U$6593 ( \6936 , \6933 , \6935 );
xor \U$6594 ( \6937 , \6930 , \6936 );
nand \U$6595 ( \6938 , \6904 , \6937 );
nand \U$6596 ( \6939 , \6862 , \6903 );
nand \U$6597 ( \6940 , \6938 , \6939 );
not \U$6598 ( \6941 , \6940 );
xor \U$6599 ( \6942 , \5306 , \5311 );
xor \U$6600 ( \6943 , \6942 , \5425 );
not \U$6601 ( \6944 , \6864 );
nand \U$6602 ( \6945 , \6944 , \6878 );
and \U$6603 ( \6946 , \6945 , \6870 );
and \U$6604 ( \6947 , \6877 , \6864 );
nor \U$6605 ( \6948 , \6946 , \6947 );
xor \U$6606 ( \6949 , \6943 , \6948 );
xor \U$6607 ( \6950 , \5474 , \5555 );
xor \U$6608 ( \6951 , \6950 , \5547 );
not \U$6609 ( \6952 , \6951 );
xor \U$6610 ( \6953 , \6949 , \6952 );
not \U$6611 ( \6954 , \6953 );
xor \U$6612 ( \6955 , \6913 , \6917 );
and \U$6613 ( \6956 , \6955 , \6920 );
and \U$6614 ( \6957 , \6913 , \6917 );
or \U$6615 ( \6958 , \6956 , \6957 );
xor \U$6616 ( \6959 , \5219 , \5177 );
xnor \U$6617 ( \6960 , \6959 , \5222 );
xor \U$6618 ( \6961 , \6958 , \6960 );
xor \U$6619 ( \6962 , \6885 , \6890 );
and \U$6620 ( \6963 , \6962 , \6893 );
and \U$6621 ( \6964 , \6885 , \6890 );
or \U$6622 ( \6965 , \6963 , \6964 );
xor \U$6623 ( \6966 , \6961 , \6965 );
xor \U$6624 ( \6967 , \6911 , \6921 );
and \U$6625 ( \6968 , \6967 , \6928 );
and \U$6626 ( \6969 , \6911 , \6921 );
or \U$6627 ( \6970 , \6968 , \6969 );
xor \U$6628 ( \6971 , \6966 , \6970 );
not \U$6629 ( \6972 , \6879 );
not \U$6630 ( \6973 , \6894 );
or \U$6631 ( \6974 , \6972 , \6973 );
or \U$6632 ( \6975 , \6879 , \6894 );
nand \U$6633 ( \6976 , \6975 , \6901 );
nand \U$6634 ( \6977 , \6974 , \6976 );
xor \U$6635 ( \6978 , \6971 , \6977 );
not \U$6636 ( \6979 , \6978 );
or \U$6637 ( \6980 , \6954 , \6979 );
or \U$6638 ( \6981 , \6978 , \6953 );
nand \U$6639 ( \6982 , \6980 , \6981 );
xor \U$6640 ( \6983 , \6909 , \6929 );
and \U$6641 ( \6984 , \6983 , \6936 );
and \U$6642 ( \6985 , \6909 , \6929 );
or \U$6643 ( \6986 , \6984 , \6985 );
xnor \U$6644 ( \6987 , \6982 , \6986 );
nand \U$6645 ( \6988 , \6941 , \6987 );
not \U$6646 ( \6989 , \6142 );
not \U$6647 ( \6990 , \6857 );
not \U$6648 ( \6991 , \6990 );
or \U$6649 ( \6992 , \6989 , \6991 );
nand \U$6650 ( \6993 , \6857 , \6141 );
nand \U$6651 ( \6994 , \6992 , \6993 );
buf \U$6652 ( \6995 , \6517 );
not \U$6653 ( \6996 , \6995 );
nand \U$6654 ( \6997 , \6510 , \657 );
not \U$6655 ( \6998 , \6997 );
and \U$6656 ( \6999 , \6996 , \6998 );
and \U$6657 ( \7000 , \6995 , \6997 );
nor \U$6658 ( \7001 , \6999 , \7000 );
buf \U$6659 ( \7002 , \7001 );
not \U$6660 ( \7003 , \7002 );
buf \U$6661 ( \7004 , \7003 );
and \U$6662 ( \7005 , \5753 , \7004 );
not \U$6663 ( \7006 , \859 );
not \U$6664 ( \7007 , \4960 );
xnor \U$6665 ( \7008 , \7007 , RI9871d70_139);
not \U$6666 ( \7009 , \7008 );
or \U$6667 ( \7010 , \7006 , \7009 );
nand \U$6668 ( \7011 , \6634 , \832 );
nand \U$6669 ( \7012 , \7010 , \7011 );
xor \U$6670 ( \7013 , \7005 , \7012 );
not \U$6671 ( \7014 , \3170 );
not \U$6672 ( \7015 , \6652 );
or \U$6673 ( \7016 , \7014 , \7015 );
and \U$6674 ( \7017 , RI9872310_151, \1659 );
not \U$6675 ( \7018 , RI9872310_151);
not \U$6676 ( \7019 , \5719 );
and \U$6677 ( \7020 , \7018 , \7019 );
nor \U$6678 ( \7021 , \7017 , \7020 );
nand \U$6679 ( \7022 , \7021 , \3163 );
nand \U$6680 ( \7023 , \7016 , \7022 );
and \U$6681 ( \7024 , \7013 , \7023 );
and \U$6682 ( \7025 , \7005 , \7012 );
or \U$6683 ( \7026 , \7024 , \7025 );
not \U$6684 ( \7027 , \6195 );
not \U$6685 ( \7028 , \6184 );
and \U$6686 ( \7029 , RI9871e60_141, \7028 );
not \U$6687 ( \7030 , RI9871e60_141);
and \U$6688 ( \7031 , \7030 , \5776 );
nor \U$6689 ( \7032 , \7029 , \7031 );
not \U$6690 ( \7033 , \7032 );
or \U$6691 ( \7034 , \7027 , \7033 );
nand \U$6692 ( \7035 , \6492 , \1353 );
nand \U$6693 ( \7036 , \7034 , \7035 );
not \U$6694 ( \7037 , \2074 );
not \U$6695 ( \7038 , \2076 );
not \U$6696 ( \7039 , \1371 );
or \U$6697 ( \7040 , \7038 , \7039 );
nand \U$6698 ( \7041 , \4455 , RI9871aa0_133);
nand \U$6699 ( \7042 , \7040 , \7041 );
not \U$6700 ( \7043 , \7042 );
or \U$6701 ( \7044 , \7037 , \7043 );
nand \U$6702 ( \7045 , \6541 , \2087 );
nand \U$6703 ( \7046 , \7044 , \7045 );
xor \U$6704 ( \7047 , \7036 , \7046 );
not \U$6705 ( \7048 , \6284 );
not \U$6706 ( \7049 , RI98728b0_163);
not \U$6707 ( \7050 , \7049 );
not \U$6708 ( \7051 , \2982 );
or \U$6709 ( \7052 , \7050 , \7051 );
or \U$6710 ( \7053 , \1393 , \5632 );
nand \U$6711 ( \7054 , \7052 , \7053 );
not \U$6712 ( \7055 , \7054 );
or \U$6713 ( \7056 , \7048 , \7055 );
nand \U$6714 ( \7057 , \6606 , \6611 );
nand \U$6715 ( \7058 , \7056 , \7057 );
and \U$6716 ( \7059 , \7047 , \7058 );
and \U$6717 ( \7060 , \7036 , \7046 );
or \U$6718 ( \7061 , \7059 , \7060 );
xor \U$6719 ( \7062 , \7026 , \7061 );
not \U$6720 ( \7063 , \4920 );
buf \U$6721 ( \7064 , \1581 );
and \U$6722 ( \7065 , RI9872388_152, \7064 );
not \U$6723 ( \7066 , RI9872388_152);
and \U$6724 ( \7067 , \7066 , \1275 );
or \U$6725 ( \7068 , \7065 , \7067 );
not \U$6726 ( \7069 , \7068 );
or \U$6727 ( \7070 , \7063 , \7069 );
nand \U$6728 ( \7071 , \6560 , \5048 );
nand \U$6729 ( \7072 , \7070 , \7071 );
not \U$6730 ( \7073 , \7072 );
not \U$6731 ( \7074 , \793 );
not \U$6732 ( \7075 , RI98719b0_131);
and \U$6733 ( \7076 , \1040 , \7075 );
not \U$6734 ( \7077 , \1040 );
and \U$6735 ( \7078 , \7077 , RI98719b0_131);
nor \U$6736 ( \7079 , \7076 , \7078 );
not \U$6737 ( \7080 , \7079 );
or \U$6738 ( \7081 , \7074 , \7080 );
nand \U$6739 ( \7082 , \6576 , \6145 );
nand \U$6740 ( \7083 , \7081 , \7082 );
not \U$6741 ( \7084 , \7083 );
or \U$6742 ( \7085 , \7073 , \7084 );
not \U$6743 ( \7086 , \7072 );
not \U$6744 ( \7087 , \7086 );
not \U$6745 ( \7088 , \7083 );
not \U$6746 ( \7089 , \7088 );
or \U$6747 ( \7090 , \7087 , \7089 );
not \U$6748 ( \7091 , \5034 );
not \U$6749 ( \7092 , \6165 );
and \U$6750 ( \7093 , \7092 , \5025 );
not \U$6751 ( \7094 , \7092 );
and \U$6752 ( \7095 , \7094 , RI9872478_154);
nor \U$6753 ( \7096 , \7093 , \7095 );
not \U$6754 ( \7097 , \7096 );
or \U$6755 ( \7098 , \7091 , \7097 );
nand \U$6756 ( \7099 , \6695 , \5796 );
nand \U$6757 ( \7100 , \7098 , \7099 );
nand \U$6758 ( \7101 , \7090 , \7100 );
nand \U$6759 ( \7102 , \7085 , \7101 );
and \U$6760 ( \7103 , \7062 , \7102 );
and \U$6761 ( \7104 , \7026 , \7061 );
or \U$6762 ( \7105 , \7103 , \7104 );
not \U$6763 ( \7106 , \1018 );
not \U$6764 ( \7107 , \3271 );
not \U$6765 ( \7108 , \5705 );
not \U$6766 ( \7109 , \7108 );
or \U$6767 ( \7110 , \7107 , \7109 );
not \U$6768 ( \7111 , \5703 );
not \U$6769 ( \7112 , \7111 );
or \U$6770 ( \7113 , \7112 , \3271 );
nand \U$6771 ( \7114 , \7110 , \7113 );
not \U$6772 ( \7115 , \7114 );
or \U$6773 ( \7116 , \7106 , \7115 );
not \U$6774 ( \7117 , \6483 );
nand \U$6775 ( \7118 , \7117 , \1013 );
nand \U$6776 ( \7119 , \7116 , \7118 );
nand \U$6777 ( \7120 , RI9872a18_166, RI9872a90_167);
and \U$6778 ( \7121 , \7120 , RI98729a0_165);
not \U$6779 ( \7122 , \7121 );
or \U$6780 ( \7123 , \7119 , \7122 );
not \U$6781 ( \7124 , \1162 );
xor \U$6782 ( \7125 , \4708 , \6530 );
not \U$6783 ( \7126 , \7125 );
or \U$6784 ( \7127 , \7124 , \7126 );
nand \U$6785 ( \7128 , \6535 , \1220 );
nand \U$6786 ( \7129 , \7127 , \7128 );
nand \U$6787 ( \7130 , \7123 , \7129 );
nand \U$6788 ( \7131 , \7119 , \7122 );
nand \U$6789 ( \7132 , \7130 , \7131 );
or \U$6790 ( \7133 , \7132 , \6613 );
not \U$6791 ( \7134 , \7131 );
not \U$6792 ( \7135 , \7130 );
or \U$6793 ( \7136 , \7134 , \7135 );
nand \U$6794 ( \7137 , \7136 , \6613 );
nand \U$6795 ( \7138 , \7133 , \7137 );
not \U$6796 ( \7139 , \7138 );
not \U$6797 ( \7140 , \6546 );
and \U$6798 ( \7141 , \6538 , \7140 );
not \U$6799 ( \7142 , \6538 );
and \U$6800 ( \7143 , \7142 , \6546 );
nor \U$6801 ( \7144 , \7141 , \7143 );
not \U$6802 ( \7145 , \7144 );
not \U$6803 ( \7146 , \7145 );
or \U$6804 ( \7147 , \7139 , \7146 );
not \U$6805 ( \7148 , \6613 );
nand \U$6806 ( \7149 , \7148 , \7132 );
nand \U$6807 ( \7150 , \7147 , \7149 );
xor \U$6808 ( \7151 , \7105 , \7150 );
xor \U$6809 ( \7152 , \6637 , \6646 );
xor \U$6810 ( \7153 , \7152 , \6655 );
not \U$6811 ( \7154 , \3467 );
not \U$6812 ( \7155 , \6728 );
or \U$6813 ( \7156 , \7154 , \7155 );
and \U$6814 ( \7157 , RI98726d0_159, \847 );
not \U$6815 ( \7158 , RI98726d0_159);
and \U$6816 ( \7159 , \7158 , \2211 );
nor \U$6817 ( \7160 , \7157 , \7159 );
nand \U$6818 ( \7161 , \7160 , \3600 );
nand \U$6819 ( \7162 , \7156 , \7161 );
not \U$6820 ( \7163 , \1455 );
not \U$6821 ( \7164 , \2111 );
and \U$6822 ( \7165 , \7164 , \1619 );
not \U$6823 ( \7166 , \7164 );
and \U$6824 ( \7167 , \7166 , RI9871c08_136);
nor \U$6825 ( \7168 , \7165 , \7167 );
not \U$6826 ( \7169 , \7168 );
or \U$6827 ( \7170 , \7163 , \7169 );
nand \U$6828 ( \7171 , \6667 , \1430 );
nand \U$6829 ( \7172 , \7170 , \7171 );
or \U$6830 ( \7173 , \7162 , \7172 );
not \U$6831 ( \7174 , \1292 );
not \U$6832 ( \7175 , \3240 );
not \U$6833 ( \7176 , RI9871b18_134);
and \U$6834 ( \7177 , \7175 , \7176 );
and \U$6835 ( \7178 , \3240 , RI9871b18_134);
nor \U$6836 ( \7179 , \7177 , \7178 );
not \U$6837 ( \7180 , \7179 );
or \U$6838 ( \7181 , \7174 , \7180 );
nand \U$6839 ( \7182 , \6709 , \1323 );
nand \U$6840 ( \7183 , \7181 , \7182 );
nand \U$6841 ( \7184 , \7173 , \7183 );
nand \U$6842 ( \7185 , \7162 , \7172 );
nand \U$6843 ( \7186 , \7184 , \7185 );
xor \U$6844 ( \7187 , \7153 , \7186 );
buf \U$6845 ( \7188 , \5653 );
not \U$6846 ( \7189 , \7188 );
not \U$6847 ( \7190 , \6501 );
or \U$6848 ( \7191 , \7189 , \7190 );
not \U$6849 ( \7192 , RI9872568_156);
not \U$6850 ( \7193 , \1097 );
or \U$6851 ( \7194 , \7192 , \7193 );
nand \U$6852 ( \7195 , \1106 , \5648 );
nand \U$6853 ( \7196 , \7194 , \7195 );
nand \U$6854 ( \7197 , \7196 , \5642 );
nand \U$6855 ( \7198 , \7191 , \7197 );
not \U$6856 ( \7199 , \1083 );
and \U$6857 ( \7200 , RI98718c0_129, \3969 );
not \U$6858 ( \7201 , RI98718c0_129);
and \U$6859 ( \7202 , \7201 , \3396 );
nor \U$6860 ( \7203 , \7200 , \7202 );
not \U$6861 ( \7204 , \7203 );
or \U$6862 ( \7205 , \7199 , \7204 );
nand \U$6863 ( \7206 , \6682 , \1136 );
nand \U$6864 ( \7207 , \7205 , \7206 );
xor \U$6865 ( \7208 , \7198 , \7207 );
not \U$6866 ( \7209 , \5530 );
not \U$6867 ( \7210 , RI98725e0_157);
xor \U$6868 ( \7211 , \1506 , \7210 );
not \U$6869 ( \7212 , \7211 );
or \U$6870 ( \7213 , \7209 , \7212 );
nand \U$6871 ( \7214 , \6587 , \4085 );
nand \U$6872 ( \7215 , \7213 , \7214 );
and \U$6873 ( \7216 , \7208 , \7215 );
and \U$6874 ( \7217 , \7198 , \7207 );
or \U$6875 ( \7218 , \7216 , \7217 );
and \U$6876 ( \7219 , \7187 , \7218 );
and \U$6877 ( \7220 , \7153 , \7186 );
or \U$6878 ( \7221 , \7219 , \7220 );
and \U$6879 ( \7222 , \7151 , \7221 );
and \U$6880 ( \7223 , \7105 , \7150 );
or \U$6881 ( \7224 , \7222 , \7223 );
and \U$6882 ( \7225 , \6700 , \6684 );
not \U$6883 ( \7226 , \6700 );
not \U$6884 ( \7227 , \6684 );
and \U$6885 ( \7228 , \7226 , \7227 );
nor \U$6886 ( \7229 , \7225 , \7228 );
and \U$6887 ( \7230 , \7229 , \6669 );
not \U$6888 ( \7231 , \7229 );
not \U$6889 ( \7232 , \6669 );
and \U$6890 ( \7233 , \7231 , \7232 );
nor \U$6891 ( \7234 , \7230 , \7233 );
xor \U$6892 ( \7235 , \6485 , \6494 );
xor \U$6893 ( \7236 , \7235 , \6505 );
xor \U$6894 ( \7237 , \7234 , \7236 );
xor \U$6895 ( \7238 , \6578 , \6589 );
xor \U$6896 ( \7239 , \7238 , \6564 );
and \U$6897 ( \7240 , \7237 , \7239 );
and \U$6898 ( \7241 , \7234 , \7236 );
or \U$6899 ( \7242 , \7240 , \7241 );
not \U$6900 ( \7243 , \6508 );
not \U$6901 ( \7244 , \7243 );
not \U$6902 ( \7245 , \6596 );
or \U$6903 ( \7246 , \7244 , \7245 );
or \U$6904 ( \7247 , \6596 , \7243 );
nand \U$6905 ( \7248 , \7246 , \7247 );
xor \U$6906 ( \7249 , \7242 , \7248 );
not \U$6907 ( \7250 , \6658 );
not \U$6908 ( \7251 , \7250 );
buf \U$6909 ( \7252 , \6739 );
not \U$6910 ( \7253 , \7252 );
or \U$6911 ( \7254 , \7251 , \7253 );
or \U$6912 ( \7255 , \7252 , \7250 );
nand \U$6913 ( \7256 , \7254 , \7255 );
and \U$6914 ( \7257 , \7249 , \7256 );
and \U$6915 ( \7258 , \7242 , \7248 );
or \U$6916 ( \7259 , \7257 , \7258 );
xor \U$6917 ( \7260 , \7224 , \7259 );
and \U$6918 ( \7261 , \6747 , \6600 );
not \U$6919 ( \7262 , \6747 );
not \U$6920 ( \7263 , \6600 );
and \U$6921 ( \7264 , \7262 , \7263 );
nor \U$6922 ( \7265 , \7261 , \7264 );
and \U$6923 ( \7266 , \7260 , \7265 );
and \U$6924 ( \7267 , \7224 , \7259 );
or \U$6925 ( \7268 , \7266 , \7267 );
not \U$6926 ( \7269 , \7268 );
not \U$6927 ( \7270 , \6756 );
not \U$6928 ( \7271 , \6426 );
not \U$6929 ( \7272 , \7271 );
and \U$6930 ( \7273 , \7270 , \7272 );
and \U$6931 ( \7274 , \6756 , \7271 );
nor \U$6932 ( \7275 , \7273 , \7274 );
not \U$6933 ( \7276 , \7275 );
or \U$6934 ( \7277 , \7269 , \7276 );
or \U$6935 ( \7278 , \7268 , \7275 );
nand \U$6936 ( \7279 , \7277 , \7278 );
xor \U$6937 ( \7280 , \6624 , \6626 );
xor \U$6938 ( \7281 , \6388 , \6397 );
xor \U$6939 ( \7282 , \7281 , \6408 );
xor \U$6940 ( \7283 , \7280 , \7282 );
and \U$6941 ( \7284 , \6350 , \6340 );
not \U$6942 ( \7285 , \6350 );
not \U$6943 ( \7286 , \6340 );
and \U$6944 ( \7287 , \7285 , \7286 );
nor \U$6945 ( \7288 , \7284 , \7287 );
xor \U$6946 ( \7289 , \7288 , \6362 );
and \U$6947 ( \7290 , \7283 , \7289 );
and \U$6948 ( \7291 , \7280 , \7282 );
or \U$6949 ( \7292 , \7290 , \7291 );
not \U$6950 ( \7293 , \7292 );
not \U$6951 ( \7294 , \5752 );
not \U$6952 ( \7295 , \5816 );
and \U$6953 ( \7296 , \7294 , \7295 );
and \U$6954 ( \7297 , \5752 , \5816 );
nor \U$6955 ( \7298 , \7296 , \7297 );
not \U$6956 ( \7299 , \7298 );
or \U$6957 ( \7300 , \7293 , \7299 );
or \U$6958 ( \7301 , \7298 , \7292 );
nand \U$6959 ( \7302 , \7300 , \7301 );
xor \U$6960 ( \7303 , \6764 , \6765 );
xor \U$6961 ( \7304 , \7303 , \6785 );
xnor \U$6962 ( \7305 , \7302 , \7304 );
not \U$6963 ( \7306 , \7305 );
not \U$6964 ( \7307 , \7306 );
xor \U$6965 ( \7308 , \6722 , \6711 );
not \U$6966 ( \7309 , \7308 );
not \U$6967 ( \7310 , \6730 );
and \U$6968 ( \7311 , \7309 , \7310 );
and \U$6969 ( \7312 , \6730 , \7308 );
nor \U$6970 ( \7313 , \7311 , \7312 );
and \U$6971 ( \7314 , RI98729a0_165, RI9872a90_167);
not \U$6972 ( \7315 , RI98729a0_165);
not \U$6973 ( \7316 , RI9872a90_167);
and \U$6974 ( \7317 , \7315 , \7316 );
nor \U$6975 ( \7318 , \7314 , \7317 );
not \U$6976 ( \7319 , \7318 );
and \U$6977 ( \7320 , RI9872a18_166, RI9872a90_167);
not \U$6978 ( \7321 , RI9872a18_166);
and \U$6979 ( \7322 , \7321 , \7316 );
nor \U$6980 ( \7323 , \7320 , \7322 );
nor \U$6981 ( \7324 , \7319 , \7323 );
buf \U$6982 ( \7325 , \7324 );
buf \U$6983 ( \7326 , \7325 );
not \U$6984 ( \7327 , \7326 );
not \U$6985 ( \7328 , RI98729a0_165);
not \U$6986 ( \7329 , \7328 );
not \U$6987 ( \7330 , \1691 );
not \U$6988 ( \7331 , \7330 );
or \U$6989 ( \7332 , \7329 , \7331 );
not \U$6990 ( \7333 , RI98729a0_165);
or \U$6991 ( \7334 , \780 , \7333 );
nand \U$6992 ( \7335 , \7332 , \7334 );
not \U$6993 ( \7336 , \7335 );
or \U$6994 ( \7337 , \7327 , \7336 );
buf \U$6995 ( \7338 , \7323 );
nand \U$6996 ( \7339 , \7338 , RI98729a0_165);
nand \U$6997 ( \7340 , \7337 , \7339 );
not \U$6998 ( \7341 , \1501 );
and \U$6999 ( \7342 , RI9871c80_137, \4155 );
not \U$7000 ( \7343 , RI9871c80_137);
and \U$7001 ( \7344 , \7343 , \3568 );
nor \U$7002 ( \7345 , \7342 , \7344 );
not \U$7003 ( \7346 , \7345 );
or \U$7004 ( \7347 , \7341 , \7346 );
nand \U$7005 ( \7348 , \6720 , \1518 );
nand \U$7006 ( \7349 , \7347 , \7348 );
or \U$7007 ( \7350 , \7340 , \7349 );
not \U$7008 ( \7351 , \924 );
not \U$7009 ( \7352 , \6642 );
or \U$7010 ( \7353 , \7351 , \7352 );
not \U$7011 ( \7354 , \919 );
not \U$7012 ( \7355 , \5614 );
not \U$7013 ( \7356 , \7355 );
or \U$7014 ( \7357 , \7354 , \7356 );
nand \U$7015 ( \7358 , \5614 , RI9872130_147);
nand \U$7016 ( \7359 , \7357 , \7358 );
nand \U$7017 ( \7360 , \7359 , \6431 );
nand \U$7018 ( \7361 , \7353 , \7360 );
nand \U$7019 ( \7362 , \7350 , \7361 );
nand \U$7020 ( \7363 , \7340 , \7349 );
nand \U$7021 ( \7364 , \7362 , \7363 );
nor \U$7022 ( \7365 , \7313 , \7364 );
not \U$7023 ( \7366 , \7138 );
not \U$7024 ( \7367 , \7144 );
and \U$7025 ( \7368 , \7366 , \7367 );
and \U$7026 ( \7369 , \7138 , \7144 );
nor \U$7027 ( \7370 , \7368 , \7369 );
or \U$7028 ( \7371 , \7365 , \7370 );
nand \U$7029 ( \7372 , \7313 , \7364 );
nand \U$7030 ( \7373 , \7371 , \7372 );
xor \U$7031 ( \7374 , \7280 , \7282 );
xor \U$7032 ( \7375 , \7374 , \7289 );
xor \U$7033 ( \7376 , \7373 , \7375 );
xor \U$7034 ( \7377 , \6253 , \6214 );
xor \U$7035 ( \7378 , \7377 , \6181 );
and \U$7036 ( \7379 , \7376 , \7378 );
and \U$7037 ( \7380 , \7373 , \7375 );
or \U$7038 ( \7381 , \7379 , \7380 );
not \U$7039 ( \7382 , \7381 );
xor \U$7040 ( \7383 , \6256 , \6421 );
not \U$7041 ( \7384 , \7383 );
or \U$7042 ( \7385 , \7382 , \7384 );
or \U$7043 ( \7386 , \7381 , \7383 );
nand \U$7044 ( \7387 , \7385 , \7386 );
not \U$7045 ( \7388 , \7387 );
or \U$7046 ( \7389 , \7307 , \7388 );
not \U$7047 ( \7390 , \7383 );
nand \U$7048 ( \7391 , \7390 , \7381 );
nand \U$7049 ( \7392 , \7389 , \7391 );
nand \U$7050 ( \7393 , \7279 , \7392 );
not \U$7051 ( \7394 , \7275 );
nand \U$7052 ( \7395 , \7394 , \7268 );
and \U$7053 ( \7396 , \7393 , \7395 );
not \U$7054 ( \7397 , \7304 );
not \U$7055 ( \7398 , \7302 );
or \U$7056 ( \7399 , \7397 , \7398 );
not \U$7057 ( \7400 , \7298 );
nand \U$7058 ( \7401 , \7400 , \7292 );
nand \U$7059 ( \7402 , \7399 , \7401 );
not \U$7060 ( \7403 , \7402 );
xor \U$7061 ( \7404 , \5819 , \5922 );
xor \U$7062 ( \7405 , \7404 , \5972 );
xor \U$7063 ( \7406 , \6796 , \6806 );
xnor \U$7064 ( \7407 , \7406 , \6788 );
xnor \U$7065 ( \7408 , \7405 , \7407 );
not \U$7066 ( \7409 , \7408 );
or \U$7067 ( \7410 , \7403 , \7409 );
not \U$7068 ( \7411 , \7405 );
nand \U$7069 ( \7412 , \7411 , \7407 );
nand \U$7070 ( \7413 , \7410 , \7412 );
not \U$7071 ( \7414 , \7413 );
and \U$7072 ( \7415 , \7396 , \7414 );
not \U$7073 ( \7416 , \7396 );
and \U$7074 ( \7417 , \7416 , \7413 );
nor \U$7075 ( \7418 , \7415 , \7417 );
not \U$7076 ( \7419 , \7418 );
and \U$7077 ( \7420 , \6994 , \7419 );
not \U$7078 ( \7421 , \6994 );
and \U$7079 ( \7422 , \7421 , \7418 );
nor \U$7080 ( \7423 , \7420 , \7422 );
xor \U$7081 ( \7424 , \7279 , \7392 );
not \U$7082 ( \7425 , \7424 );
not \U$7083 ( \7426 , \7408 );
not \U$7084 ( \7427 , \7402 );
not \U$7085 ( \7428 , \7427 );
and \U$7086 ( \7429 , \7426 , \7428 );
and \U$7087 ( \7430 , \7408 , \7427 );
nor \U$7088 ( \7431 , \7429 , \7430 );
not \U$7089 ( \7432 , \7431 );
xor \U$7090 ( \7433 , \7224 , \7259 );
xor \U$7091 ( \7434 , \7433 , \7265 );
and \U$7092 ( \7435 , \6298 , \3272 );
not \U$7093 ( \7436 , \6298 );
and \U$7094 ( \7437 , \7436 , \1043 );
nor \U$7095 ( \7438 , \7435 , \7437 );
not \U$7096 ( \7439 , \7438 );
not \U$7097 ( \7440 , \7439 );
not \U$7098 ( \7441 , \1612 );
and \U$7099 ( \7442 , \7440 , \7441 );
buf \U$7100 ( \7443 , \7114 );
and \U$7101 ( \7444 , \7443 , \1067 );
nor \U$7102 ( \7445 , \7442 , \7444 );
not \U$7103 ( \7446 , \7445 );
not \U$7104 ( \7447 , \7446 );
buf \U$7105 ( \7448 , \554 );
and \U$7106 ( \7449 , \7448 , \557 , \551 );
not \U$7107 ( \7450 , \7449 );
not \U$7108 ( \7451 , \548 );
not \U$7109 ( \7452 , \5672 );
or \U$7110 ( \7453 , \7451 , \7452 );
nand \U$7111 ( \7454 , \7453 , \5682 );
not \U$7112 ( \7455 , \7454 );
or \U$7113 ( \7456 , \7450 , \7455 );
not \U$7114 ( \7457 , \678 );
nand \U$7115 ( \7458 , \7456 , \7457 );
not \U$7116 ( \7459 , \7458 );
nand \U$7117 ( \7460 , \560 , \5689 );
not \U$7118 ( \7461 , \7460 );
and \U$7119 ( \7462 , \7459 , \7461 );
and \U$7120 ( \7463 , \7458 , \7460 );
nor \U$7121 ( \7464 , \7462 , \7463 );
buf \U$7122 ( \7465 , \7464 );
buf \U$7123 ( \7466 , \7465 );
not \U$7124 ( \7467 , \7466 );
and \U$7125 ( \7468 , \4708 , \7467 );
not \U$7126 ( \7469 , \1220 );
not \U$7127 ( \7470 , \7125 );
or \U$7128 ( \7471 , \7469 , \7470 );
xor \U$7129 ( \7472 , \5753 , \7004 );
nand \U$7130 ( \7473 , \7472 , \1162 );
nand \U$7131 ( \7474 , \7471 , \7473 );
xor \U$7132 ( \7475 , \7468 , \7474 );
not \U$7133 ( \7476 , \7475 );
or \U$7134 ( \7477 , \7447 , \7476 );
nand \U$7135 ( \7478 , \7474 , \7468 );
nand \U$7136 ( \7479 , \7477 , \7478 );
buf \U$7137 ( \7480 , \7119 );
xor \U$7138 ( \7481 , \7121 , \7480 );
xnor \U$7139 ( \7482 , \7481 , \7129 );
or \U$7140 ( \7483 , \7479 , \7482 );
not \U$7141 ( \7484 , \1501 );
and \U$7142 ( \7485 , \1584 , \4176 );
not \U$7143 ( \7486 , \1584 );
and \U$7144 ( \7487 , \7486 , \4177 );
nor \U$7145 ( \7488 , \7485 , \7487 );
not \U$7146 ( \7489 , \7488 );
or \U$7147 ( \7490 , \7484 , \7489 );
nand \U$7148 ( \7491 , \7345 , \1518 );
nand \U$7149 ( \7492 , \7490 , \7491 );
not \U$7150 ( \7493 , \7492 );
and \U$7151 ( \7494 , \1283 , \3537 );
not \U$7152 ( \7495 , \1283 );
and \U$7153 ( \7496 , \7495 , \3542 );
nor \U$7154 ( \7497 , \7494 , \7496 );
not \U$7155 ( \7498 , \7497 );
not \U$7156 ( \7499 , \1293 );
and \U$7157 ( \7500 , \7498 , \7499 );
and \U$7158 ( \7501 , \7179 , \1323 );
nor \U$7159 ( \7502 , \7500 , \7501 );
nand \U$7160 ( \7503 , \7493 , \7502 );
not \U$7161 ( \7504 , \7503 );
not \U$7162 ( \7505 , \3467 );
not \U$7163 ( \7506 , \7160 );
or \U$7164 ( \7507 , \7505 , \7506 );
not \U$7165 ( \7508 , \3593 );
not \U$7166 ( \7509 , \944 );
or \U$7167 ( \7510 , \7508 , \7509 );
or \U$7168 ( \7511 , \944 , \4063 );
nand \U$7169 ( \7512 , \7510 , \7511 );
nand \U$7170 ( \7513 , \7512 , \3466 );
nand \U$7171 ( \7514 , \7507 , \7513 );
not \U$7172 ( \7515 , \7514 );
or \U$7173 ( \7516 , \7504 , \7515 );
not \U$7174 ( \7517 , \7502 );
nand \U$7175 ( \7518 , \7517 , \7492 );
nand \U$7176 ( \7519 , \7516 , \7518 );
and \U$7177 ( \7520 , \7483 , \7519 );
and \U$7178 ( \7521 , \7482 , \7479 );
nor \U$7179 ( \7522 , \7520 , \7521 );
not \U$7180 ( \7523 , \7522 );
not \U$7181 ( \7524 , \7523 );
not \U$7182 ( \7525 , \832 );
not \U$7183 ( \7526 , \7008 );
or \U$7184 ( \7527 , \7525 , \7526 );
and \U$7185 ( \7528 , \2312 , \5325 );
not \U$7186 ( \7529 , \2312 );
and \U$7187 ( \7530 , \7529 , \4986 );
nor \U$7188 ( \7531 , \7528 , \7530 );
not \U$7189 ( \7532 , \7531 );
nand \U$7190 ( \7533 , \7532 , \6635 );
nand \U$7191 ( \7534 , \7527 , \7533 );
not \U$7192 ( \7535 , \7534 );
not \U$7193 ( \7536 , \1353 );
not \U$7194 ( \7537 , \7032 );
or \U$7195 ( \7538 , \7536 , \7537 );
and \U$7196 ( \7539 , RI9871e60_141, \5761 );
not \U$7197 ( \7540 , RI9871e60_141);
buf \U$7198 ( \7541 , \6480 );
and \U$7199 ( \7542 , \7540 , \7541 );
nor \U$7200 ( \7543 , \7539 , \7542 );
or \U$7201 ( \7544 , \7543 , \6194 );
nand \U$7202 ( \7545 , \7538 , \7544 );
not \U$7203 ( \7546 , \7545 );
and \U$7204 ( \7547 , \7535 , \7546 );
not \U$7205 ( \7548 , \3164 );
and \U$7206 ( \7549 , RI9872310_151, \1341 );
not \U$7207 ( \7550 , RI9872310_151);
and \U$7208 ( \7551 , \7550 , \1344 );
nor \U$7209 ( \7552 , \7549 , \7551 );
not \U$7210 ( \7553 , \7552 );
or \U$7211 ( \7554 , \7548 , \7553 );
nand \U$7212 ( \7555 , \7021 , \3170 );
nand \U$7213 ( \7556 , \7554 , \7555 );
not \U$7214 ( \7557 , \7556 );
nand \U$7215 ( \7558 , \7534 , \7545 );
and \U$7216 ( \7559 , \7557 , \7558 );
nor \U$7217 ( \7560 , \7547 , \7559 );
not \U$7218 ( \7561 , \2072 );
not \U$7219 ( \7562 , \2076 );
not \U$7220 ( \7563 , \6573 );
or \U$7221 ( \7564 , \7562 , \7563 );
or \U$7222 ( \7565 , \1713 , \2080 );
nand \U$7223 ( \7566 , \7564 , \7565 );
not \U$7224 ( \7567 , \7566 );
or \U$7225 ( \7568 , \7561 , \7567 );
not \U$7226 ( \7569 , \7042 );
or \U$7227 ( \7570 , \7569 , \2086 );
nand \U$7228 ( \7571 , \7568 , \7570 );
not \U$7229 ( \7572 , \6611 );
not \U$7230 ( \7573 , \7054 );
or \U$7231 ( \7574 , \7572 , \7573 );
not \U$7232 ( \7575 , \1725 );
not \U$7233 ( \7576 , RI98728b0_163);
and \U$7234 ( \7577 , \7575 , \7576 );
and \U$7235 ( \7578 , \2399 , RI98728b0_163);
nor \U$7236 ( \7579 , \7577 , \7578 );
or \U$7237 ( \7580 , \7579 , \6283 );
nand \U$7238 ( \7581 , \7574 , \7580 );
xor \U$7239 ( \7582 , \7571 , \7581 );
not \U$7240 ( \7583 , \7096 );
not \U$7241 ( \7584 , \5796 );
or \U$7242 ( \7585 , \7583 , \7584 );
and \U$7243 ( \7586 , RI9872478_154, \1740 );
not \U$7244 ( \7587 , RI9872478_154);
and \U$7245 ( \7588 , \7587 , \1320 );
nor \U$7246 ( \7589 , \7586 , \7588 );
not \U$7247 ( \7590 , \7589 );
not \U$7248 ( \7591 , \5034 );
or \U$7249 ( \7592 , \7590 , \7591 );
nand \U$7250 ( \7593 , \7585 , \7592 );
and \U$7251 ( \7594 , \7582 , \7593 );
and \U$7252 ( \7595 , \7571 , \7581 );
or \U$7253 ( \7596 , \7594 , \7595 );
xor \U$7254 ( \7597 , \7560 , \7596 );
not \U$7255 ( \7598 , \797 );
not \U$7256 ( \7599 , \7079 );
or \U$7257 ( \7600 , \7598 , \7599 );
not \U$7258 ( \7601 , \6568 );
not \U$7259 ( \7602 , \1212 );
or \U$7260 ( \7603 , \7601 , \7602 );
not \U$7261 ( \7604 , \6020 );
not \U$7262 ( \7605 , \7604 );
or \U$7263 ( \7606 , \7605 , \6574 );
nand \U$7264 ( \7607 , \7603 , \7606 );
nand \U$7265 ( \7608 , \7607 , \793 );
nand \U$7266 ( \7609 , \7600 , \7608 );
not \U$7267 ( \7610 , \5048 );
not \U$7268 ( \7611 , \7068 );
or \U$7269 ( \7612 , \7610 , \7611 );
not \U$7270 ( \7613 , RI9872388_152);
not \U$7271 ( \7614 , \5480 );
or \U$7272 ( \7615 , \7613 , \7614 );
or \U$7273 ( \7616 , \916 , RI9872388_152);
nand \U$7274 ( \7617 , \7615 , \7616 );
nand \U$7275 ( \7618 , \7617 , \5942 );
nand \U$7276 ( \7619 , \7612 , \7618 );
xor \U$7277 ( \7620 , \7609 , \7619 );
not \U$7278 ( \7621 , \1136 );
not \U$7279 ( \7622 , \7203 );
or \U$7280 ( \7623 , \7621 , \7622 );
xnor \U$7281 ( \7624 , \2116 , RI98718c0_129);
nand \U$7282 ( \7625 , \7624 , \1083 );
nand \U$7283 ( \7626 , \7623 , \7625 );
and \U$7284 ( \7627 , \7620 , \7626 );
and \U$7285 ( \7628 , \7609 , \7619 );
or \U$7286 ( \7629 , \7627 , \7628 );
and \U$7287 ( \7630 , \7597 , \7629 );
and \U$7288 ( \7631 , \7560 , \7596 );
or \U$7289 ( \7632 , \7630 , \7631 );
not \U$7290 ( \7633 , \7632 );
or \U$7291 ( \7634 , \7524 , \7633 );
not \U$7292 ( \7635 , \7632 );
not \U$7293 ( \7636 , \7522 );
and \U$7294 ( \7637 , \7635 , \7636 );
and \U$7295 ( \7638 , \7632 , \7522 );
nor \U$7296 ( \7639 , \7637 , \7638 );
xor \U$7297 ( \7640 , \7153 , \7186 );
xor \U$7298 ( \7641 , \7640 , \7218 );
not \U$7299 ( \7642 , \7641 );
or \U$7300 ( \7643 , \7639 , \7642 );
nand \U$7301 ( \7644 , \7634 , \7643 );
xor \U$7302 ( \7645 , \7105 , \7150 );
xor \U$7303 ( \7646 , \7645 , \7221 );
xor \U$7304 ( \7647 , \7644 , \7646 );
xor \U$7305 ( \7648 , \7026 , \7061 );
xor \U$7306 ( \7649 , \7648 , \7102 );
xor \U$7307 ( \7650 , \7198 , \7207 );
xor \U$7308 ( \7651 , \7650 , \7215 );
not \U$7309 ( \7652 , \7651 );
xor \U$7310 ( \7653 , \7005 , \7012 );
xor \U$7311 ( \7654 , \7653 , \7023 );
not \U$7312 ( \7655 , \7654 );
xor \U$7313 ( \7656 , \7349 , \7361 );
xnor \U$7314 ( \7657 , \7656 , \7340 );
nand \U$7315 ( \7658 , \7655 , \7657 );
not \U$7316 ( \7659 , \7658 );
or \U$7317 ( \7660 , \7652 , \7659 );
not \U$7318 ( \7661 , \7657 );
nand \U$7319 ( \7662 , \7661 , \7654 );
nand \U$7320 ( \7663 , \7660 , \7662 );
xor \U$7321 ( \7664 , \7649 , \7663 );
xor \U$7322 ( \7665 , \7036 , \7046 );
xor \U$7323 ( \7666 , \7665 , \7058 );
not \U$7324 ( \7667 , \7666 );
not \U$7325 ( \7668 , \1431 );
not \U$7326 ( \7669 , \7168 );
or \U$7327 ( \7670 , \7668 , \7669 );
xnor \U$7328 ( \7671 , \3691 , RI9871c08_136);
nand \U$7329 ( \7672 , \7671 , \1455 );
nand \U$7330 ( \7673 , \7670 , \7672 );
not \U$7331 ( \7674 , \7673 );
not \U$7332 ( \7675 , \7196 );
not \U$7333 ( \7676 , \7675 );
not \U$7334 ( \7677 , \7188 );
not \U$7335 ( \7678 , \7677 );
and \U$7336 ( \7679 , \7676 , \7678 );
not \U$7337 ( \7680 , \1416 );
not \U$7338 ( \7681 , RI9872568_156);
and \U$7339 ( \7682 , \7680 , \7681 );
and \U$7340 ( \7683 , \1416 , RI9872568_156);
nor \U$7341 ( \7684 , \7682 , \7683 );
not \U$7342 ( \7685 , \7684 );
and \U$7343 ( \7686 , \7685 , \5642 );
nor \U$7344 ( \7687 , \7679 , \7686 );
not \U$7345 ( \7688 , \4085 );
not \U$7346 ( \7689 , \7211 );
or \U$7347 ( \7690 , \7688 , \7689 );
not \U$7348 ( \7691 , \820 );
xor \U$7349 ( \7692 , \7691 , RI98725e0_157);
nand \U$7350 ( \7693 , \7692 , \4103 );
nand \U$7351 ( \7694 , \7690 , \7693 );
xnor \U$7352 ( \7695 , \7687 , \7694 );
not \U$7353 ( \7696 , \7695 );
or \U$7354 ( \7697 , \7674 , \7696 );
not \U$7355 ( \7698 , \7687 );
nand \U$7356 ( \7699 , \7694 , \7698 );
nand \U$7357 ( \7700 , \7697 , \7699 );
not \U$7358 ( \7701 , \7700 );
and \U$7359 ( \7702 , \7100 , \7083 );
not \U$7360 ( \7703 , \7100 );
and \U$7361 ( \7704 , \7703 , \7088 );
nor \U$7362 ( \7705 , \7702 , \7704 );
not \U$7363 ( \7706 , \7705 );
not \U$7364 ( \7707 , \7086 );
and \U$7365 ( \7708 , \7706 , \7707 );
and \U$7366 ( \7709 , \7705 , \7086 );
nor \U$7367 ( \7710 , \7708 , \7709 );
nand \U$7368 ( \7711 , \7701 , \7710 );
not \U$7369 ( \7712 , \7711 );
or \U$7370 ( \7713 , \7667 , \7712 );
not \U$7371 ( \7714 , \7710 );
nand \U$7372 ( \7715 , \7714 , \7700 );
nand \U$7373 ( \7716 , \7713 , \7715 );
and \U$7374 ( \7717 , \7664 , \7716 );
and \U$7375 ( \7718 , \7649 , \7663 );
or \U$7376 ( \7719 , \7717 , \7718 );
and \U$7377 ( \7720 , \7647 , \7719 );
and \U$7378 ( \7721 , \7644 , \7646 );
or \U$7379 ( \7722 , \7720 , \7721 );
xor \U$7380 ( \7723 , \7434 , \7722 );
not \U$7381 ( \7724 , \7305 );
not \U$7382 ( \7725 , \7387 );
or \U$7383 ( \7726 , \7724 , \7725 );
or \U$7384 ( \7727 , \7387 , \7305 );
nand \U$7385 ( \7728 , \7726 , \7727 );
and \U$7386 ( \7729 , \7723 , \7728 );
and \U$7387 ( \7730 , \7434 , \7722 );
or \U$7388 ( \7731 , \7729 , \7730 );
not \U$7389 ( \7732 , \7731 );
and \U$7390 ( \7733 , \7432 , \7732 );
and \U$7391 ( \7734 , \7431 , \7731 );
nor \U$7392 ( \7735 , \7733 , \7734 );
not \U$7393 ( \7736 , \7735 );
not \U$7394 ( \7737 , \7736 );
or \U$7395 ( \7738 , \7425 , \7737 );
not \U$7396 ( \7739 , \7431 );
nand \U$7397 ( \7740 , \7739 , \7731 );
nand \U$7398 ( \7741 , \7738 , \7740 );
not \U$7399 ( \7742 , \7741 );
nand \U$7400 ( \7743 , \7423 , \7742 );
buf \U$7401 ( \7744 , \7743 );
not \U$7402 ( \7745 , \6862 );
not \U$7403 ( \7746 , \6902 );
not \U$7404 ( \7747 , \6937 );
or \U$7405 ( \7748 , \7746 , \7747 );
or \U$7406 ( \7749 , \6937 , \6902 );
nand \U$7407 ( \7750 , \7748 , \7749 );
not \U$7408 ( \7751 , \7750 );
or \U$7409 ( \7752 , \7745 , \7751 );
or \U$7410 ( \7753 , \7750 , \6862 );
nand \U$7411 ( \7754 , \7752 , \7753 );
nand \U$7412 ( \7755 , \7418 , \6994 );
not \U$7413 ( \7756 , \7395 );
not \U$7414 ( \7757 , \7393 );
or \U$7415 ( \7758 , \7756 , \7757 );
nand \U$7416 ( \7759 , \7758 , \7413 );
nand \U$7417 ( \7760 , \7754 , \7755 , \7759 );
not \U$7418 ( \7761 , \7424 );
not \U$7419 ( \7762 , \7735 );
or \U$7420 ( \7763 , \7761 , \7762 );
or \U$7421 ( \7764 , \7424 , \7735 );
nand \U$7422 ( \7765 , \7763 , \7764 );
not \U$7423 ( \7766 , \7765 );
xor \U$7424 ( \7767 , \7434 , \7722 );
xor \U$7425 ( \7768 , \7767 , \7728 );
not \U$7426 ( \7769 , \7768 );
xor \U$7427 ( \7770 , \7234 , \7236 );
xor \U$7428 ( \7771 , \7770 , \7239 );
not \U$7429 ( \7772 , \7771 );
not \U$7430 ( \7773 , \7364 );
and \U$7431 ( \7774 , \7313 , \7773 );
not \U$7432 ( \7775 , \7313 );
and \U$7433 ( \7776 , \7775 , \7364 );
nor \U$7434 ( \7777 , \7774 , \7776 );
xnor \U$7435 ( \7778 , \7370 , \7777 );
not \U$7436 ( \7779 , \7778 );
or \U$7437 ( \7780 , \7772 , \7779 );
or \U$7438 ( \7781 , \7771 , \7778 );
nand \U$7439 ( \7782 , \7780 , \7781 );
or \U$7440 ( \7783 , \7531 , \932 );
and \U$7441 ( \7784 , \5776 , RI9871d70_139);
and \U$7442 ( \7785 , \6185 , \1347 );
nor \U$7443 ( \7786 , \7784 , \7785 );
or \U$7444 ( \7787 , \7786 , \860 );
nand \U$7445 ( \7788 , \7783 , \7787 );
not \U$7446 ( \7789 , \876 );
not \U$7447 ( \7790 , RI9872130_147);
buf \U$7448 ( \7791 , \4988 );
not \U$7449 ( \7792 , \7791 );
or \U$7450 ( \7793 , \7790 , \7792 );
or \U$7451 ( \7794 , \7007 , RI9872130_147);
nand \U$7452 ( \7795 , \7793 , \7794 );
not \U$7453 ( \7796 , \7795 );
or \U$7454 ( \7797 , \7789 , \7796 );
and \U$7455 ( \7798 , RI9872130_147, \4471 );
not \U$7456 ( \7799 , RI9872130_147);
and \U$7457 ( \7800 , \7799 , \5623 );
nor \U$7458 ( \7801 , \7798 , \7800 );
or \U$7459 ( \7802 , \7801 , \1470 );
nand \U$7460 ( \7803 , \7797 , \7802 );
xor \U$7461 ( \7804 , \7788 , \7803 );
not \U$7462 ( \7805 , \7326 );
not \U$7463 ( \7806 , \7328 );
not \U$7464 ( \7807 , \1393 );
or \U$7465 ( \7808 , \7806 , \7807 );
or \U$7466 ( \7809 , \2982 , \7333 );
nand \U$7467 ( \7810 , \7808 , \7809 );
not \U$7468 ( \7811 , \7810 );
or \U$7469 ( \7812 , \7805 , \7811 );
nand \U$7470 ( \7813 , \7335 , \7338 );
nand \U$7471 ( \7814 , \7812 , \7813 );
and \U$7472 ( \7815 , \7804 , \7814 );
and \U$7473 ( \7816 , \7788 , \7803 );
or \U$7474 ( \7817 , \7815 , \7816 );
not \U$7475 ( \7818 , \3164 );
not \U$7476 ( \7819 , RI9872310_151);
not \U$7477 ( \7820 , \3886 );
or \U$7478 ( \7821 , \7819 , \7820 );
or \U$7479 ( \7822 , \1366 , RI9872310_151);
nand \U$7480 ( \7823 , \7821 , \7822 );
not \U$7481 ( \7824 , \7823 );
or \U$7482 ( \7825 , \7818 , \7824 );
nand \U$7483 ( \7826 , \7552 , \3170 );
nand \U$7484 ( \7827 , \7825 , \7826 );
not \U$7485 ( \7828 , \2074 );
and \U$7486 ( \7829 , RI9871aa0_133, \1047 );
not \U$7487 ( \7830 , RI9871aa0_133);
and \U$7488 ( \7831 , \7830 , \1041 );
nor \U$7489 ( \7832 , \7829 , \7831 );
not \U$7490 ( \7833 , \7832 );
or \U$7491 ( \7834 , \7828 , \7833 );
nand \U$7492 ( \7835 , \7566 , \2087 );
nand \U$7493 ( \7836 , \7834 , \7835 );
xor \U$7494 ( \7837 , \7827 , \7836 );
or \U$7495 ( \7838 , \7684 , \7677 );
not \U$7496 ( \7839 , \5648 );
not \U$7497 ( \7840 , \2680 );
or \U$7498 ( \7841 , \7839 , \7840 );
nand \U$7499 ( \7842 , \2492 , RI9872568_156);
nand \U$7500 ( \7843 , \7841 , \7842 );
not \U$7501 ( \7844 , \7843 );
not \U$7502 ( \7845 , \5642 );
or \U$7503 ( \7846 , \7844 , \7845 );
nand \U$7504 ( \7847 , \7838 , \7846 );
and \U$7505 ( \7848 , \7837 , \7847 );
and \U$7506 ( \7849 , \7827 , \7836 );
or \U$7507 ( \7850 , \7848 , \7849 );
xor \U$7508 ( \7851 , \7817 , \7850 );
not \U$7509 ( \7852 , \5796 );
not \U$7510 ( \7853 , \7589 );
or \U$7511 ( \7854 , \7852 , \7853 );
not \U$7512 ( \7855 , \5025 );
not \U$7513 ( \7856 , \1275 );
or \U$7514 ( \7857 , \7855 , \7856 );
nand \U$7515 ( \7858 , \7064 , RI9872478_154);
nand \U$7516 ( \7859 , \7857 , \7858 );
nand \U$7517 ( \7860 , \7859 , \5034 );
nand \U$7518 ( \7861 , \7854 , \7860 );
not \U$7519 ( \7862 , \6284 );
not \U$7520 ( \7863 , RI98728b0_163);
not \U$7521 ( \7864 , \1097 );
or \U$7522 ( \7865 , \7863 , \7864 );
or \U$7523 ( \7866 , \1098 , RI98728b0_163);
nand \U$7524 ( \7867 , \7865 , \7866 );
not \U$7525 ( \7868 , \7867 );
or \U$7526 ( \7869 , \7862 , \7868 );
not \U$7527 ( \7870 , \7579 );
nand \U$7528 ( \7871 , \7870 , \6611 );
nand \U$7529 ( \7872 , \7869 , \7871 );
xor \U$7530 ( \7873 , \7861 , \7872 );
not \U$7531 ( \7874 , \794 );
and \U$7532 ( \7875 , RI98719b0_131, \3969 );
not \U$7533 ( \7876 , RI98719b0_131);
and \U$7534 ( \7877 , \7876 , \1191 );
nor \U$7535 ( \7878 , \7875 , \7877 );
not \U$7536 ( \7879 , \7878 );
or \U$7537 ( \7880 , \7874 , \7879 );
nand \U$7538 ( \7881 , \7607 , \797 );
nand \U$7539 ( \7882 , \7880 , \7881 );
and \U$7540 ( \7883 , \7873 , \7882 );
and \U$7541 ( \7884 , \7861 , \7872 );
or \U$7542 ( \7885 , \7883 , \7884 );
and \U$7543 ( \7886 , \7851 , \7885 );
and \U$7544 ( \7887 , \7817 , \7850 );
or \U$7545 ( \7888 , \7886 , \7887 );
not \U$7546 ( \7889 , \7888 );
not \U$7547 ( \7890 , \1381 );
and \U$7548 ( \7891 , \5708 , RI9871e60_141);
not \U$7549 ( \7892 , \5708 );
and \U$7550 ( \7893 , \7892 , \1367 );
or \U$7551 ( \7894 , \7891 , \7893 );
not \U$7552 ( \7895 , \7894 );
or \U$7553 ( \7896 , \7890 , \7895 );
or \U$7554 ( \7897 , \7543 , \2595 );
nand \U$7555 ( \7898 , \7896 , \7897 );
not \U$7556 ( \7899 , \7898 );
and \U$7557 ( \7900 , RI9872b08_168, RI9872b80_169);
not \U$7558 ( \7901 , RI9872a18_166);
nor \U$7559 ( \7902 , \7900 , \7901 );
not \U$7560 ( \7903 , \7902 );
not \U$7561 ( \7904 , \1018 );
buf \U$7562 ( \7905 , \6528 );
and \U$7563 ( \7906 , \7905 , \1044 );
not \U$7564 ( \7907 , \7905 );
and \U$7565 ( \7908 , \7907 , \3271 );
nor \U$7566 ( \7909 , \7906 , \7908 );
not \U$7567 ( \7910 , \7909 );
or \U$7568 ( \7911 , \7904 , \7910 );
nand \U$7569 ( \7912 , \7438 , \1013 );
nand \U$7570 ( \7913 , \7911 , \7912 );
not \U$7571 ( \7914 , \7913 );
or \U$7572 ( \7915 , \7903 , \7914 );
or \U$7573 ( \7916 , \7913 , \7902 );
nand \U$7574 ( \7917 , \7915 , \7916 );
not \U$7575 ( \7918 , \7917 );
or \U$7576 ( \7919 , \7899 , \7918 );
not \U$7577 ( \7920 , \7902 );
nand \U$7578 ( \7921 , \7920 , \7913 );
nand \U$7579 ( \7922 , \7919 , \7921 );
not \U$7580 ( \7923 , \7922 );
not \U$7581 ( \7924 , \924 );
not \U$7582 ( \7925 , \7359 );
or \U$7583 ( \7926 , \7924 , \7925 );
not \U$7584 ( \7927 , \876 );
or \U$7585 ( \7928 , \7801 , \7927 );
nand \U$7586 ( \7929 , \7926 , \7928 );
not \U$7587 ( \7930 , \7929 );
not \U$7588 ( \7931 , \7340 );
or \U$7589 ( \7932 , \7930 , \7931 );
or \U$7590 ( \7933 , \7340 , \7929 );
nand \U$7591 ( \7934 , \7932 , \7933 );
not \U$7592 ( \7935 , \7934 );
or \U$7593 ( \7936 , \7923 , \7935 );
not \U$7594 ( \7937 , \7340 );
nand \U$7595 ( \7938 , \7937 , \7929 );
nand \U$7596 ( \7939 , \7936 , \7938 );
xor \U$7597 ( \7940 , \7183 , \7172 );
xnor \U$7598 ( \7941 , \7940 , \7162 );
xnor \U$7599 ( \7942 , \7939 , \7941 );
not \U$7600 ( \7943 , \7942 );
or \U$7601 ( \7944 , \7889 , \7943 );
not \U$7602 ( \7945 , \7941 );
nand \U$7603 ( \7946 , \7945 , \7939 );
nand \U$7604 ( \7947 , \7944 , \7946 );
xor \U$7605 ( \7948 , \7782 , \7947 );
xor \U$7606 ( \7949 , \7649 , \7663 );
xor \U$7607 ( \7950 , \7949 , \7716 );
xor \U$7608 ( \7951 , \7948 , \7950 );
nand \U$7609 ( \7952 , \7658 , \7662 );
not \U$7610 ( \7953 , \7952 );
not \U$7611 ( \7954 , \7651 );
and \U$7612 ( \7955 , \7953 , \7954 );
and \U$7613 ( \7956 , \7952 , \7651 );
nor \U$7614 ( \7957 , \7955 , \7956 );
not \U$7615 ( \7958 , \7957 );
not \U$7616 ( \7959 , \7958 );
not \U$7617 ( \7960 , \7888 );
xor \U$7618 ( \7961 , \7939 , \7941 );
not \U$7619 ( \7962 , \7961 );
and \U$7620 ( \7963 , \7960 , \7962 );
and \U$7621 ( \7964 , \7961 , \7888 );
nor \U$7622 ( \7965 , \7963 , \7964 );
not \U$7623 ( \7966 , \7965 );
not \U$7624 ( \7967 , \7966 );
or \U$7625 ( \7968 , \7959 , \7967 );
not \U$7626 ( \7969 , \7957 );
not \U$7627 ( \7970 , \7965 );
or \U$7628 ( \7971 , \7969 , \7970 );
not \U$7629 ( \7972 , \6611 );
not \U$7630 ( \7973 , \7867 );
or \U$7631 ( \7974 , \7972 , \7973 );
not \U$7632 ( \7975 , \5632 );
not \U$7633 ( \7976 , \1417 );
or \U$7634 ( \7977 , \7975 , \7976 );
nand \U$7635 ( \7978 , \6174 , RI98728b0_163);
nand \U$7636 ( \7979 , \7977 , \7978 );
nand \U$7637 ( \7980 , \7979 , \6284 );
nand \U$7638 ( \7981 , \7974 , \7980 );
not \U$7639 ( \7982 , \797 );
not \U$7640 ( \7983 , \7878 );
or \U$7641 ( \7984 , \7982 , \7983 );
and \U$7642 ( \7985 , RI98719b0_131, \2116 );
not \U$7643 ( \7986 , RI98719b0_131);
and \U$7644 ( \7987 , \7986 , \1486 );
nor \U$7645 ( \7988 , \7985 , \7987 );
not \U$7646 ( \7989 , \7988 );
nand \U$7647 ( \7990 , \7989 , \793 );
nand \U$7648 ( \7991 , \7984 , \7990 );
xor \U$7649 ( \7992 , \7981 , \7991 );
not \U$7650 ( \7993 , RI9872388_152);
not \U$7651 ( \7994 , \7993 );
not \U$7652 ( \7995 , \2955 );
or \U$7653 ( \7996 , \7994 , \7995 );
nand \U$7654 ( \7997 , \6443 , RI9872388_152);
nand \U$7655 ( \7998 , \7996 , \7997 );
not \U$7656 ( \7999 , \7998 );
or \U$7657 ( \8000 , \7999 , \4924 );
not \U$7658 ( \8001 , RI9872388_152);
not \U$7659 ( \8002 , \820 );
or \U$7660 ( \8003 , \8001 , \8002 );
not \U$7661 ( \8004 , \819 );
buf \U$7662 ( \8005 , \8004 );
not \U$7663 ( \8006 , \8005 );
or \U$7664 ( \8007 , \8006 , RI9872388_152);
nand \U$7665 ( \8008 , \8003 , \8007 );
not \U$7666 ( \8009 , \8008 );
not \U$7667 ( \8010 , \4920 );
or \U$7668 ( \8011 , \8009 , \8010 );
nand \U$7669 ( \8012 , \8000 , \8011 );
and \U$7670 ( \8013 , \7992 , \8012 );
and \U$7671 ( \8014 , \7981 , \7991 );
or \U$7672 ( \8015 , \8013 , \8014 );
not \U$7673 ( \8016 , \8015 );
not \U$7674 ( \8017 , RI9872b08_168);
and \U$7675 ( \8018 , RI9872b80_169, \8017 );
not \U$7676 ( \8019 , RI9872b80_169);
and \U$7677 ( \8020 , \8019 , RI9872b08_168);
nor \U$7678 ( \8021 , \8018 , \8020 );
and \U$7679 ( \8022 , RI9872a18_166, RI9872b08_168);
not \U$7680 ( \8023 , RI9872a18_166);
and \U$7681 ( \8024 , \8023 , \8017 );
nor \U$7682 ( \8025 , \8022 , \8024 );
and \U$7683 ( \8026 , \8021 , \8025 );
buf \U$7684 ( \8027 , \8026 );
buf \U$7685 ( \8028 , \8027 );
buf \U$7686 ( \8029 , \8028 );
not \U$7687 ( \8030 , \8029 );
not \U$7688 ( \8031 , RI9872a18_166);
not \U$7689 ( \8032 , \8031 );
not \U$7690 ( \8033 , \1692 );
or \U$7691 ( \8034 , \8032 , \8033 );
or \U$7692 ( \8035 , \2361 , \8031 );
nand \U$7693 ( \8036 , \8034 , \8035 );
not \U$7694 ( \8037 , \8036 );
or \U$7695 ( \8038 , \8030 , \8037 );
not \U$7696 ( \8039 , \8021 );
not \U$7697 ( \8040 , \8039 );
not \U$7698 ( \8041 , \8040 );
nand \U$7699 ( \8042 , \8041 , RI9872a18_166);
nand \U$7700 ( \8043 , \8038 , \8042 );
not \U$7701 ( \8044 , \8043 );
not \U$7702 ( \8045 , \8044 );
not \U$7703 ( \8046 , \1353 );
not \U$7704 ( \8047 , \7894 );
or \U$7705 ( \8048 , \8046 , \8047 );
and \U$7706 ( \8049 , \6290 , \6294 );
not \U$7707 ( \8050 , \6290 );
and \U$7708 ( \8051 , \8050 , \6291 );
nor \U$7709 ( \8052 , \8049 , \8051 );
buf \U$7710 ( \8053 , \8052 );
buf \U$7711 ( \8054 , \8053 );
and \U$7712 ( \8055 , RI9871e60_141, \8054 );
not \U$7713 ( \8056 , RI9871e60_141);
and \U$7714 ( \8057 , \8056 , \6298 );
or \U$7715 ( \8058 , \8055 , \8057 );
nand \U$7716 ( \8059 , \8058 , \1381 );
nand \U$7717 ( \8060 , \8048 , \8059 );
not \U$7718 ( \8061 , \8060 );
not \U$7719 ( \8062 , \7448 );
not \U$7720 ( \8063 , \5683 );
or \U$7721 ( \8064 , \8062 , \8063 );
buf \U$7722 ( \8065 , \671 );
nand \U$7723 ( \8066 , \8064 , \8065 );
nand \U$7724 ( \8067 , \557 , \673 );
not \U$7725 ( \8068 , \8067 );
and \U$7726 ( \8069 , \8066 , \8068 );
not \U$7727 ( \8070 , \8066 );
and \U$7728 ( \8071 , \8070 , \8067 );
nor \U$7729 ( \8072 , \8069 , \8071 );
not \U$7730 ( \8073 , \8072 );
buf \U$7731 ( \8074 , \8073 );
not \U$7732 ( \8075 , \8074 );
nand \U$7733 ( \8076 , \8075 , \1165 );
not \U$7734 ( \8077 , \8076 );
not \U$7735 ( \8078 , \1067 );
not \U$7736 ( \8079 , \7909 );
or \U$7737 ( \8080 , \8078 , \8079 );
buf \U$7738 ( \8081 , \7002 );
not \U$7739 ( \8082 , \8081 );
and \U$7740 ( \8083 , \8082 , \1044 );
not \U$7741 ( \8084 , \8082 );
not \U$7742 ( \8085 , \1043 );
not \U$7743 ( \8086 , \8085 );
and \U$7744 ( \8087 , \8084 , \8086 );
nor \U$7745 ( \8088 , \8083 , \8087 );
nand \U$7746 ( \8089 , \8088 , \1018 );
nand \U$7747 ( \8090 , \8080 , \8089 );
not \U$7748 ( \8091 , \8090 );
or \U$7749 ( \8092 , \8077 , \8091 );
or \U$7750 ( \8093 , \8090 , \8076 );
nand \U$7751 ( \8094 , \8092 , \8093 );
not \U$7752 ( \8095 , \8094 );
or \U$7753 ( \8096 , \8061 , \8095 );
not \U$7754 ( \8097 , \8076 );
nand \U$7755 ( \8098 , \8097 , \8090 );
nand \U$7756 ( \8099 , \8096 , \8098 );
not \U$7757 ( \8100 , \8099 );
or \U$7758 ( \8101 , \8045 , \8100 );
or \U$7759 ( \8102 , \8044 , \8099 );
nand \U$7760 ( \8103 , \8101 , \8102 );
not \U$7761 ( \8104 , \8103 );
or \U$7762 ( \8105 , \8016 , \8104 );
nand \U$7763 ( \8106 , \8099 , \8043 );
nand \U$7764 ( \8107 , \8105 , \8106 );
xnor \U$7765 ( \8108 , \7922 , \7934 );
xor \U$7766 ( \8109 , \8107 , \8108 );
not \U$7767 ( \8110 , \8109 );
not \U$7768 ( \8111 , \8110 );
or \U$7769 ( \8112 , \7786 , \932 );
and \U$7770 ( \8113 , RI9871d70_139, \5761 );
not \U$7771 ( \8114 , RI9871d70_139);
and \U$7772 ( \8115 , \8114 , \5762 );
nor \U$7773 ( \8116 , \8113 , \8115 );
or \U$7774 ( \8117 , \8116 , \5351 );
nand \U$7775 ( \8118 , \8112 , \8117 );
not \U$7776 ( \8119 , \3170 );
not \U$7777 ( \8120 , \7823 );
or \U$7778 ( \8121 , \8119 , \8120 );
xor \U$7779 ( \8122 , \1062 , RI9872310_151);
nand \U$7780 ( \8123 , \8122 , \3163 );
nand \U$7781 ( \8124 , \8121 , \8123 );
xor \U$7782 ( \8125 , \8118 , \8124 );
not \U$7783 ( \8126 , \7326 );
not \U$7784 ( \8127 , RI98729a0_165);
not \U$7785 ( \8128 , \1725 );
or \U$7786 ( \8129 , \8127 , \8128 );
or \U$7787 ( \8130 , \1725 , RI98729a0_165);
nand \U$7788 ( \8131 , \8129 , \8130 );
not \U$7789 ( \8132 , \8131 );
or \U$7790 ( \8133 , \8126 , \8132 );
nand \U$7791 ( \8134 , \7810 , \7338 );
nand \U$7792 ( \8135 , \8133 , \8134 );
and \U$7793 ( \8136 , \8125 , \8135 );
and \U$7794 ( \8137 , \8118 , \8124 );
or \U$7795 ( \8138 , \8136 , \8137 );
not \U$7796 ( \8139 , \8138 );
not \U$7797 ( \8140 , \1430 );
and \U$7798 ( \8141 , RI9871c08_136, \3861 );
not \U$7799 ( \8142 , RI9871c08_136);
and \U$7800 ( \8143 , \8142 , \3240 );
or \U$7801 ( \8144 , \8141 , \8143 );
not \U$7802 ( \8145 , \8144 );
or \U$7803 ( \8146 , \8140 , \8145 );
xor \U$7804 ( \8147 , RI9871c08_136, \3537 );
nand \U$7805 ( \8148 , \8147 , \1456 );
nand \U$7806 ( \8149 , \8146 , \8148 );
not \U$7807 ( \8150 , \8149 );
not \U$7808 ( \8151 , \6673 );
xnor \U$7809 ( \8152 , \2962 , RI98718c0_129);
not \U$7810 ( \8153 , \8152 );
or \U$7811 ( \8154 , \8151 , \8153 );
and \U$7812 ( \8155 , RI98718c0_129, \4287 );
not \U$7813 ( \8156 , RI98718c0_129);
and \U$7814 ( \8157 , \8156 , \2948 );
or \U$7815 ( \8158 , \8155 , \8157 );
nand \U$7816 ( \8159 , \8158 , \1083 );
nand \U$7817 ( \8160 , \8154 , \8159 );
not \U$7818 ( \8161 , \5847 );
xnor \U$7819 ( \8162 , \6225 , RI98725e0_157);
not \U$7820 ( \8163 , \8162 );
or \U$7821 ( \8164 , \8161 , \8163 );
buf \U$7822 ( \8165 , \5908 );
not \U$7823 ( \8166 , \8165 );
not \U$7824 ( \8167 , \3454 );
and \U$7825 ( \8168 , \8166 , \8167 );
not \U$7826 ( \8169 , \3832 );
and \U$7827 ( \8170 , \8169 , \4088 );
nor \U$7828 ( \8171 , \8168 , \8170 );
not \U$7829 ( \8172 , \8171 );
nand \U$7830 ( \8173 , \8172 , \4101 );
nand \U$7831 ( \8174 , \8164 , \8173 );
xor \U$7832 ( \8175 , \8160 , \8174 );
not \U$7833 ( \8176 , \8175 );
or \U$7834 ( \8177 , \8150 , \8176 );
nand \U$7835 ( \8178 , \8174 , \8160 );
nand \U$7836 ( \8179 , \8177 , \8178 );
not \U$7837 ( \8180 , \8179 );
not \U$7838 ( \8181 , \2087 );
not \U$7839 ( \8182 , \7832 );
or \U$7840 ( \8183 , \8181 , \8182 );
and \U$7841 ( \8184 , RI9871aa0_133, \3129 );
not \U$7842 ( \8185 , RI9871aa0_133);
and \U$7843 ( \8186 , \8185 , \7605 );
or \U$7844 ( \8187 , \8184 , \8186 );
not \U$7845 ( \8188 , \8187 );
or \U$7846 ( \8189 , \8188 , \2073 );
nand \U$7847 ( \8190 , \8183 , \8189 );
not \U$7848 ( \8191 , \8190 );
not \U$7849 ( \8192 , \5796 );
not \U$7850 ( \8193 , \7859 );
or \U$7851 ( \8194 , \8192 , \8193 );
not \U$7852 ( \8195 , RI9872478_154);
not \U$7853 ( \8196 , \5480 );
or \U$7854 ( \8197 , \8195 , \8196 );
or \U$7855 ( \8198 , \918 , RI9872478_154);
nand \U$7856 ( \8199 , \8197 , \8198 );
nand \U$7857 ( \8200 , \8199 , \5034 );
nand \U$7858 ( \8201 , \8194 , \8200 );
not \U$7859 ( \8202 , \5642 );
and \U$7860 ( \8203 , \1309 , RI9872568_156);
not \U$7861 ( \8204 , \1309 );
and \U$7862 ( \8205 , \8204 , \5648 );
nor \U$7863 ( \8206 , \8203 , \8205 );
not \U$7864 ( \8207 , \8206 );
or \U$7865 ( \8208 , \8202 , \8207 );
nand \U$7866 ( \8209 , \7843 , \7188 );
nand \U$7867 ( \8210 , \8208 , \8209 );
and \U$7868 ( \8211 , \8201 , \8210 );
not \U$7869 ( \8212 , \8201 );
not \U$7870 ( \8213 , \8210 );
and \U$7871 ( \8214 , \8212 , \8213 );
nor \U$7872 ( \8215 , \8211 , \8214 );
not \U$7873 ( \8216 , \8215 );
or \U$7874 ( \8217 , \8191 , \8216 );
nand \U$7875 ( \8218 , \8210 , \8201 );
nand \U$7876 ( \8219 , \8217 , \8218 );
not \U$7877 ( \8220 , \8219 );
not \U$7878 ( \8221 , \8220 );
or \U$7879 ( \8222 , \8180 , \8221 );
or \U$7880 ( \8223 , \8220 , \8179 );
nand \U$7881 ( \8224 , \8222 , \8223 );
not \U$7882 ( \8225 , \8224 );
or \U$7883 ( \8226 , \8139 , \8225 );
nand \U$7884 ( \8227 , \8179 , \8219 );
nand \U$7885 ( \8228 , \8226 , \8227 );
not \U$7886 ( \8229 , \8228 );
or \U$7887 ( \8230 , \8111 , \8229 );
not \U$7888 ( \8231 , \8108 );
nand \U$7889 ( \8232 , \8231 , \8107 );
nand \U$7890 ( \8233 , \8230 , \8232 );
nand \U$7891 ( \8234 , \7971 , \8233 );
nand \U$7892 ( \8235 , \7968 , \8234 );
and \U$7893 ( \8236 , \7951 , \8235 );
and \U$7894 ( \8237 , \7948 , \7950 );
or \U$7895 ( \8238 , \8236 , \8237 );
xor \U$7896 ( \8239 , \7644 , \7646 );
xor \U$7897 ( \8240 , \8239 , \7719 );
xor \U$7898 ( \8241 , \8238 , \8240 );
xor \U$7899 ( \8242 , \7482 , \7479 );
xor \U$7900 ( \8243 , \8242 , \7519 );
xor \U$7901 ( \8244 , \7560 , \7596 );
xor \U$7902 ( \8245 , \8244 , \7629 );
xor \U$7903 ( \8246 , \8243 , \8245 );
xor \U$7904 ( \8247 , \7666 , \7710 );
xnor \U$7905 ( \8248 , \8247 , \7700 );
and \U$7906 ( \8249 , \8246 , \8248 );
and \U$7907 ( \8250 , \8243 , \8245 );
or \U$7908 ( \8251 , \8249 , \8250 );
not \U$7909 ( \8252 , \8251 );
xnor \U$7910 ( \8253 , \7639 , \7641 );
not \U$7911 ( \8254 , \8253 );
or \U$7912 ( \8255 , \8252 , \8254 );
not \U$7913 ( \8256 , \8253 );
not \U$7914 ( \8257 , \8251 );
not \U$7915 ( \8258 , \8257 );
or \U$7916 ( \8259 , \8256 , \8258 );
not \U$7917 ( \8260 , \8253 );
nand \U$7918 ( \8261 , \8260 , \8251 );
nand \U$7919 ( \8262 , \8259 , \8261 );
not \U$7920 ( \8263 , \8262 );
xnor \U$7921 ( \8264 , \7556 , \7545 );
not \U$7922 ( \8265 , \8264 );
not \U$7923 ( \8266 , \7534 );
and \U$7924 ( \8267 , \8265 , \8266 );
and \U$7925 ( \8268 , \8264 , \7534 );
nor \U$7926 ( \8269 , \8267 , \8268 );
xor \U$7927 ( \8270 , \7492 , \7502 );
xor \U$7928 ( \8271 , \8270 , \7514 );
xor \U$7929 ( \8272 , \8269 , \8271 );
xor \U$7930 ( \8273 , \7673 , \7698 );
xnor \U$7931 ( \8274 , \8273 , \7694 );
and \U$7932 ( \8275 , \8272 , \8274 );
and \U$7933 ( \8276 , \8269 , \8271 );
or \U$7934 ( \8277 , \8275 , \8276 );
not \U$7935 ( \8278 , \8277 );
not \U$7936 ( \8279 , \8278 );
xor \U$7937 ( \8280 , \7571 , \7581 );
xor \U$7938 ( \8281 , \8280 , \7593 );
not \U$7939 ( \8282 , \8281 );
xor \U$7940 ( \8283 , \7609 , \7619 );
xor \U$7941 ( \8284 , \8283 , \7626 );
and \U$7942 ( \8285 , \4154 , \4044 );
not \U$7943 ( \8286 , \4154 );
and \U$7944 ( \8287 , \8286 , RI9871b18_134);
nor \U$7945 ( \8288 , \8285 , \8287 );
not \U$7946 ( \8289 , \8288 );
not \U$7947 ( \8290 , \1292 );
or \U$7948 ( \8291 , \8289 , \8290 );
or \U$7949 ( \8292 , \7497 , \1543 );
nand \U$7950 ( \8293 , \8291 , \8292 );
not \U$7951 ( \8294 , \1518 );
not \U$7952 ( \8295 , \7488 );
or \U$7953 ( \8296 , \8294 , \8295 );
and \U$7954 ( \8297 , RI9871c80_137, \5208 );
not \U$7955 ( \8298 , RI9871c80_137);
and \U$7956 ( \8299 , \8298 , \4410 );
nor \U$7957 ( \8300 , \8297 , \8299 );
nand \U$7958 ( \8301 , \8300 , \1501 );
nand \U$7959 ( \8302 , \8296 , \8301 );
xor \U$7960 ( \8303 , \8293 , \8302 );
not \U$7961 ( \8304 , \4085 );
not \U$7962 ( \8305 , \7692 );
or \U$7963 ( \8306 , \8304 , \8305 );
nand \U$7964 ( \8307 , \8162 , \4103 );
nand \U$7965 ( \8308 , \8306 , \8307 );
and \U$7966 ( \8309 , \8303 , \8308 );
and \U$7967 ( \8310 , \8293 , \8302 );
or \U$7968 ( \8311 , \8309 , \8310 );
xor \U$7969 ( \8312 , \8284 , \8311 );
not \U$7970 ( \8313 , \8312 );
or \U$7971 ( \8314 , \8282 , \8313 );
nand \U$7972 ( \8315 , \8284 , \8311 );
nand \U$7973 ( \8316 , \8314 , \8315 );
not \U$7974 ( \8317 , \8316 );
xnor \U$7975 ( \8318 , \7445 , \7475 );
not \U$7976 ( \8319 , \8318 );
not \U$7977 ( \8320 , \7448 );
nor \U$7978 ( \8321 , \8320 , \670 );
not \U$7979 ( \8322 , \8321 );
not \U$7980 ( \8323 , \7454 );
or \U$7981 ( \8324 , \8322 , \8323 );
not \U$7982 ( \8325 , \674 );
nand \U$7983 ( \8326 , \8324 , \8325 );
not \U$7984 ( \8327 , \8326 );
nand \U$7985 ( \8328 , \551 , \677 );
not \U$7986 ( \8329 , \8328 );
and \U$7987 ( \8330 , \8327 , \8329 );
and \U$7988 ( \8331 , \8326 , \8328 );
nor \U$7989 ( \8332 , \8330 , \8331 );
buf \U$7990 ( \8333 , \8332 );
buf \U$7991 ( \8334 , \8333 );
not \U$7992 ( \8335 , \8334 );
nand \U$7993 ( \8336 , \4708 , \8335 );
not \U$7994 ( \8337 , \8336 );
not \U$7995 ( \8338 , \1162 );
xor \U$7996 ( \8339 , \4708 , \7467 );
not \U$7997 ( \8340 , \8339 );
or \U$7998 ( \8341 , \8338 , \8340 );
nand \U$7999 ( \8342 , \7472 , \1220 );
nand \U$8000 ( \8343 , \8341 , \8342 );
not \U$8001 ( \8344 , \8343 );
or \U$8002 ( \8345 , \8337 , \8344 );
or \U$8003 ( \8346 , \8343 , \8336 );
nand \U$8004 ( \8347 , \8345 , \8346 );
not \U$8005 ( \8348 , \3467 );
not \U$8006 ( \8349 , \7512 );
or \U$8007 ( \8350 , \8348 , \8349 );
xor \U$8008 ( \8351 , \1658 , RI98726d0_159);
not \U$8009 ( \8352 , \8351 );
nand \U$8010 ( \8353 , \8352 , \3600 );
nand \U$8011 ( \8354 , \8350 , \8353 );
and \U$8012 ( \8355 , \8347 , \8354 );
not \U$8013 ( \8356 , \8343 );
nor \U$8014 ( \8357 , \8356 , \8336 );
nor \U$8015 ( \8358 , \8355 , \8357 );
not \U$8016 ( \8359 , \8358 );
and \U$8017 ( \8360 , \8319 , \8359 );
and \U$8018 ( \8361 , \8318 , \8358 );
nor \U$8019 ( \8362 , \8360 , \8361 );
not \U$8020 ( \8363 , \8362 );
not \U$8021 ( \8364 , \8363 );
not \U$8022 ( \8365 , \1083 );
not \U$8023 ( \8366 , \8152 );
or \U$8024 ( \8367 , \8365 , \8366 );
nand \U$8025 ( \8368 , \7624 , \1136 );
nand \U$8026 ( \8369 , \8367 , \8368 );
not \U$8027 ( \8370 , \8369 );
not \U$8028 ( \8371 , \4920 );
not \U$8029 ( \8372 , \7998 );
or \U$8030 ( \8373 , \8371 , \8372 );
nand \U$8031 ( \8374 , \7617 , \4925 );
nand \U$8032 ( \8375 , \8373 , \8374 );
not \U$8033 ( \8376 , \8375 );
and \U$8034 ( \8377 , \8144 , \1456 );
and \U$8035 ( \8378 , \7671 , \1430 );
nor \U$8036 ( \8379 , \8377 , \8378 );
not \U$8037 ( \8380 , \8379 );
or \U$8038 ( \8381 , \8376 , \8380 );
or \U$8039 ( \8382 , \8375 , \8379 );
nand \U$8040 ( \8383 , \8381 , \8382 );
not \U$8041 ( \8384 , \8383 );
or \U$8042 ( \8385 , \8370 , \8384 );
not \U$8043 ( \8386 , \8379 );
nand \U$8044 ( \8387 , \8386 , \8375 );
nand \U$8045 ( \8388 , \8385 , \8387 );
not \U$8046 ( \8389 , \8388 );
or \U$8047 ( \8390 , \8364 , \8389 );
not \U$8048 ( \8391 , \8358 );
nand \U$8049 ( \8392 , \8391 , \8318 );
nand \U$8050 ( \8393 , \8390 , \8392 );
not \U$8051 ( \8394 , \8393 );
not \U$8052 ( \8395 , \8394 );
or \U$8053 ( \8396 , \8317 , \8395 );
or \U$8054 ( \8397 , \8316 , \8394 );
nand \U$8055 ( \8398 , \8396 , \8397 );
not \U$8056 ( \8399 , \8398 );
or \U$8057 ( \8400 , \8279 , \8399 );
nand \U$8058 ( \8401 , \8316 , \8393 );
nand \U$8059 ( \8402 , \8400 , \8401 );
not \U$8060 ( \8403 , \8402 );
or \U$8061 ( \8404 , \8263 , \8403 );
nand \U$8062 ( \8405 , \8255 , \8404 );
and \U$8063 ( \8406 , \8241 , \8405 );
and \U$8064 ( \8407 , \8238 , \8240 );
or \U$8065 ( \8408 , \8406 , \8407 );
not \U$8066 ( \8409 , \8408 );
or \U$8067 ( \8410 , \7769 , \8409 );
or \U$8068 ( \8411 , \8408 , \7768 );
not \U$8069 ( \8412 , \7947 );
not \U$8070 ( \8413 , \7782 );
or \U$8071 ( \8414 , \8412 , \8413 );
not \U$8072 ( \8415 , \7778 );
nand \U$8073 ( \8416 , \8415 , \7771 );
nand \U$8074 ( \8417 , \8414 , \8416 );
not \U$8075 ( \8418 , \8417 );
xor \U$8076 ( \8419 , \7373 , \7375 );
xor \U$8077 ( \8420 , \8419 , \7378 );
xor \U$8078 ( \8421 , \7242 , \7248 );
xor \U$8079 ( \8422 , \8421 , \7256 );
or \U$8080 ( \8423 , \8420 , \8422 );
not \U$8081 ( \8424 , \8423 );
or \U$8082 ( \8425 , \8418 , \8424 );
nand \U$8083 ( \8426 , \8420 , \8422 );
nand \U$8084 ( \8427 , \8425 , \8426 );
nand \U$8085 ( \8428 , \8411 , \8427 );
nand \U$8086 ( \8429 , \8410 , \8428 );
not \U$8087 ( \8430 , \8429 );
nand \U$8088 ( \8431 , \7766 , \8430 );
and \U$8089 ( \8432 , \6988 , \7744 , \7760 , \8431 );
not \U$8090 ( \8433 , \6948 );
not \U$8091 ( \8434 , \6951 );
or \U$8092 ( \8435 , \8433 , \8434 );
nand \U$8093 ( \8436 , \8435 , \6943 );
not \U$8094 ( \8437 , \6948 );
nand \U$8095 ( \8438 , \8437 , \6952 );
nand \U$8096 ( \8439 , \8436 , \8438 );
not \U$8097 ( \8440 , \8439 );
xor \U$8098 ( \8441 , \6958 , \6960 );
and \U$8099 ( \8442 , \8441 , \6965 );
and \U$8100 ( \8443 , \6958 , \6960 );
or \U$8101 ( \8444 , \8442 , \8443 );
not \U$8102 ( \8445 , \8444 );
not \U$8103 ( \8446 , \5428 );
not \U$8104 ( \8447 , \8446 );
not \U$8105 ( \8448 , \5441 );
and \U$8106 ( \8449 , \8447 , \8448 );
and \U$8107 ( \8450 , \5441 , \8446 );
nor \U$8108 ( \8451 , \8449 , \8450 );
not \U$8109 ( \8452 , \8451 );
or \U$8110 ( \8453 , \8445 , \8452 );
or \U$8111 ( \8454 , \8444 , \8451 );
nand \U$8112 ( \8455 , \8453 , \8454 );
not \U$8113 ( \8456 , \8455 );
or \U$8114 ( \8457 , \8440 , \8456 );
not \U$8115 ( \8458 , \8451 );
nand \U$8116 ( \8459 , \8458 , \8444 );
nand \U$8117 ( \8460 , \8457 , \8459 );
not \U$8118 ( \8461 , \8460 );
not \U$8119 ( \8462 , \8461 );
xor \U$8120 ( \8463 , \5160 , \5175 );
xor \U$8121 ( \8464 , \8463 , \5265 );
not \U$8122 ( \8465 , \8464 );
and \U$8123 ( \8466 , \8462 , \8465 );
and \U$8124 ( \8467 , \8461 , \8464 );
nor \U$8125 ( \8468 , \8466 , \8467 );
not \U$8126 ( \8469 , \8468 );
not \U$8127 ( \8470 , \5446 );
not \U$8128 ( \8471 , \5457 );
or \U$8129 ( \8472 , \8470 , \8471 );
or \U$8130 ( \8473 , \5446 , \5457 );
nand \U$8131 ( \8474 , \8472 , \8473 );
not \U$8132 ( \8475 , \8474 );
not \U$8133 ( \8476 , \5573 );
or \U$8134 ( \8477 , \8475 , \8476 );
or \U$8135 ( \8478 , \5573 , \8474 );
nand \U$8136 ( \8479 , \8477 , \8478 );
nand \U$8137 ( \8480 , \8469 , \8479 );
not \U$8138 ( \8481 , \8480 );
not \U$8139 ( \8482 , \8464 );
nand \U$8140 ( \8483 , \8482 , \8461 );
not \U$8141 ( \8484 , \8483 );
or \U$8142 ( \8485 , \8481 , \8484 );
not \U$8143 ( \8486 , \5578 );
not \U$8144 ( \8487 , \8486 );
nand \U$8145 ( \8488 , \5587 , \5584 );
not \U$8146 ( \8489 , \8488 );
or \U$8147 ( \8490 , \8487 , \8489 );
or \U$8148 ( \8491 , \8488 , \8486 );
nand \U$8149 ( \8492 , \8490 , \8491 );
nand \U$8150 ( \8493 , \8485 , \8492 );
xor \U$8151 ( \8494 , \6966 , \6970 );
and \U$8152 ( \8495 , \8494 , \6977 );
and \U$8153 ( \8496 , \6966 , \6970 );
or \U$8154 ( \8497 , \8495 , \8496 );
not \U$8155 ( \8498 , \8497 );
not \U$8156 ( \8499 , \8498 );
xnor \U$8157 ( \8500 , \5568 , \5461 );
not \U$8158 ( \8501 , \8500 );
xor \U$8159 ( \8502 , \8439 , \8455 );
not \U$8160 ( \8503 , \8502 );
not \U$8161 ( \8504 , \8503 );
or \U$8162 ( \8505 , \8501 , \8504 );
not \U$8163 ( \8506 , \8500 );
nand \U$8164 ( \8507 , \8506 , \8502 );
nand \U$8165 ( \8508 , \8505 , \8507 );
not \U$8166 ( \8509 , \8508 );
or \U$8167 ( \8510 , \8499 , \8509 );
or \U$8168 ( \8511 , \8508 , \8498 );
nand \U$8169 ( \8512 , \8510 , \8511 );
not \U$8170 ( \8513 , \6986 );
not \U$8171 ( \8514 , \6982 );
or \U$8172 ( \8515 , \8513 , \8514 );
not \U$8173 ( \8516 , \6953 );
nand \U$8174 ( \8517 , \8516 , \6978 );
nand \U$8175 ( \8518 , \8515 , \8517 );
or \U$8176 ( \8519 , \8512 , \8518 );
not \U$8177 ( \8520 , \8468 );
not \U$8178 ( \8521 , \8479 );
and \U$8179 ( \8522 , \8520 , \8521 );
and \U$8180 ( \8523 , \8468 , \8479 );
nor \U$8181 ( \8524 , \8522 , \8523 );
not \U$8182 ( \8525 , \8497 );
not \U$8183 ( \8526 , \8508 );
or \U$8184 ( \8527 , \8525 , \8526 );
nand \U$8185 ( \8528 , \8502 , \8500 );
nand \U$8186 ( \8529 , \8527 , \8528 );
nor \U$8187 ( \8530 , \8524 , \8529 );
not \U$8188 ( \8531 , \8530 );
and \U$8189 ( \8532 , \8493 , \8519 , \8531 );
nand \U$8190 ( \8533 , \5592 , \8432 , \8532 );
nor \U$8191 ( \8534 , \3089 , \8533 );
not \U$8192 ( \8535 , \8534 );
not \U$8193 ( \8536 , \1018 );
not \U$8194 ( \8537 , \545 );
not \U$8195 ( \8538 , \8537 );
nor \U$8196 ( \8539 , \536 , \5670 );
not \U$8197 ( \8540 , \543 );
or \U$8198 ( \8541 , \8539 , \8540 );
not \U$8199 ( \8542 , \622 );
nand \U$8200 ( \8543 , \8541 , \8542 );
not \U$8201 ( \8544 , \8543 );
or \U$8202 ( \8545 , \8538 , \8544 );
nand \U$8203 ( \8546 , \8545 , \623 );
not \U$8204 ( \8547 , \8546 );
not \U$8205 ( \8548 , \544 );
nand \U$8206 ( \8549 , \8548 , \617 );
not \U$8207 ( \8550 , \8549 );
and \U$8208 ( \8551 , \8547 , \8550 );
and \U$8209 ( \8552 , \8546 , \8549 );
nor \U$8210 ( \8553 , \8551 , \8552 );
buf \U$8211 ( \8554 , \8553 );
buf \U$8212 ( \8555 , \8554 );
and \U$8213 ( \8556 , \8555 , \8086 );
not \U$8214 ( \8557 , \8555 );
and \U$8215 ( \8558 , \8557 , \3272 );
nor \U$8216 ( \8559 , \8556 , \8558 );
not \U$8217 ( \8560 , \8559 );
or \U$8218 ( \8561 , \8536 , \8560 );
not \U$8219 ( \8562 , \538 );
nand \U$8220 ( \8563 , \8562 , \642 );
not \U$8221 ( \8564 , \8563 );
nand \U$8222 ( \8565 , \543 , \546 );
or \U$8223 ( \8566 , \8539 , \8565 );
and \U$8224 ( \8567 , \626 , \617 );
nand \U$8225 ( \8568 , \8566 , \8567 );
buf \U$8226 ( \8569 , \8568 );
not \U$8227 ( \8570 , \8569 );
or \U$8228 ( \8571 , \8564 , \8570 );
or \U$8229 ( \8572 , \8569 , \8563 );
nand \U$8230 ( \8573 , \8571 , \8572 );
buf \U$8231 ( \8574 , \8573 );
buf \U$8232 ( \8575 , \8574 );
not \U$8233 ( \8576 , \8575 );
and \U$8234 ( \8577 , \3271 , \8576 );
not \U$8235 ( \8578 , \3271 );
not \U$8236 ( \8579 , \8574 );
not \U$8237 ( \8580 , \8579 );
and \U$8238 ( \8581 , \8578 , \8580 );
nor \U$8239 ( \8582 , \8577 , \8581 );
nand \U$8240 ( \8583 , \8582 , \1013 );
nand \U$8241 ( \8584 , \8561 , \8583 );
not \U$8242 ( \8585 , \859 );
nand \U$8243 ( \8586 , \547 , \5678 );
not \U$8244 ( \8587 , \8586 );
not \U$8245 ( \8588 , \630 );
not \U$8246 ( \8589 , \8568 );
or \U$8247 ( \8590 , \8588 , \8589 );
not \U$8248 ( \8591 , \649 );
nand \U$8249 ( \8592 , \8590 , \8591 );
not \U$8250 ( \8593 , \8592 );
or \U$8251 ( \8594 , \8587 , \8593 );
or \U$8252 ( \8595 , \8592 , \8586 );
nand \U$8253 ( \8596 , \8594 , \8595 );
buf \U$8254 ( \8597 , \8596 );
and \U$8255 ( \8598 , RI9871d70_139, \8597 );
not \U$8256 ( \8599 , RI9871d70_139);
not \U$8257 ( \8600 , \8592 );
not \U$8258 ( \8601 , \8586 );
and \U$8259 ( \8602 , \8600 , \8601 );
and \U$8260 ( \8603 , \8592 , \8586 );
nor \U$8261 ( \8604 , \8602 , \8603 );
not \U$8262 ( \8605 , \8604 );
buf \U$8263 ( \8606 , \8605 );
not \U$8264 ( \8607 , \8606 );
and \U$8265 ( \8608 , \8599 , \8607 );
nor \U$8266 ( \8609 , \8598 , \8608 );
not \U$8267 ( \8610 , \8609 );
or \U$8268 ( \8611 , \8585 , \8610 );
buf \U$8269 ( \8612 , \7454 );
not \U$8270 ( \8613 , \8612 );
nand \U$8271 ( \8614 , \7448 , \8065 );
not \U$8272 ( \8615 , \8614 );
and \U$8273 ( \8616 , \8613 , \8615 );
and \U$8274 ( \8617 , \8612 , \8614 );
nor \U$8275 ( \8618 , \8616 , \8617 );
not \U$8276 ( \8619 , \8618 );
not \U$8277 ( \8620 , \8619 );
not \U$8278 ( \8621 , \8620 );
and \U$8279 ( \8622 , RI9871d70_139, \8621 );
not \U$8280 ( \8623 , RI9871d70_139);
not \U$8281 ( \8624 , \8621 );
and \U$8282 ( \8625 , \8623 , \8624 );
nor \U$8283 ( \8626 , \8622 , \8625 );
nand \U$8284 ( \8627 , \8626 , \832 );
nand \U$8285 ( \8628 , \8611 , \8627 );
xor \U$8286 ( \8629 , \8584 , \8628 );
not \U$8287 ( \8630 , \1381 );
not \U$8288 ( \8631 , \8562 );
not \U$8289 ( \8632 , \8568 );
or \U$8290 ( \8633 , \8631 , \8632 );
nand \U$8291 ( \8634 , \8633 , \642 );
not \U$8292 ( \8635 , \629 );
nand \U$8293 ( \8636 , \8635 , \644 );
nor \U$8294 ( \8637 , \8634 , \8636 );
not \U$8295 ( \8638 , \8637 );
nand \U$8296 ( \8639 , \8634 , \8636 );
nand \U$8297 ( \8640 , \8638 , \8639 );
not \U$8298 ( \8641 , \8640 );
not \U$8299 ( \8642 , \8641 );
and \U$8300 ( \8643 , RI9871e60_141, \8642 );
not \U$8301 ( \8644 , RI9871e60_141);
not \U$8302 ( \8645 , \8634 );
not \U$8303 ( \8646 , \8636 );
and \U$8304 ( \8647 , \8645 , \8646 );
and \U$8305 ( \8648 , \8634 , \8636 );
nor \U$8306 ( \8649 , \8647 , \8648 );
buf \U$8307 ( \8650 , \8649 );
and \U$8308 ( \8651 , \8644 , \8650 );
nor \U$8309 ( \8652 , \8643 , \8651 );
not \U$8310 ( \8653 , \8652 );
or \U$8311 ( \8654 , \8630 , \8653 );
nor \U$8312 ( \8655 , \629 , \538 );
not \U$8313 ( \8656 , \8655 );
not \U$8314 ( \8657 , \8568 );
or \U$8315 ( \8658 , \8656 , \8657 );
not \U$8316 ( \8659 , \645 );
nand \U$8317 ( \8660 , \8658 , \8659 );
not \U$8318 ( \8661 , \8660 );
nand \U$8319 ( \8662 , \640 , \648 );
not \U$8320 ( \8663 , \8662 );
and \U$8321 ( \8664 , \8661 , \8663 );
and \U$8322 ( \8665 , \8660 , \8662 );
nor \U$8323 ( \8666 , \8664 , \8665 );
buf \U$8324 ( \8667 , \8666 );
buf \U$8325 ( \8668 , \8667 );
and \U$8326 ( \8669 , \8668 , \5616 );
not \U$8327 ( \8670 , \8668 );
and \U$8328 ( \8671 , \8670 , RI9871e60_141);
nor \U$8329 ( \8672 , \8669 , \8671 );
nand \U$8330 ( \8673 , \8672 , \1353 );
nand \U$8331 ( \8674 , \8654 , \8673 );
xor \U$8332 ( \8675 , \8629 , \8674 );
not \U$8333 ( \8676 , \1220 );
not \U$8334 ( \8677 , \1153 );
not \U$8335 ( \8678 , \8677 );
buf \U$8336 ( \8679 , \8678 );
not \U$8337 ( \8680 , \541 );
not \U$8338 ( \8681 , \8680 );
buf \U$8339 ( \8682 , \5672 );
not \U$8340 ( \8683 , \8682 );
or \U$8341 ( \8684 , \8681 , \8683 );
buf \U$8342 ( \8685 , \619 );
nand \U$8343 ( \8686 , \8684 , \8685 );
not \U$8344 ( \8687 , \8686 );
not \U$8345 ( \8688 , \542 );
nand \U$8346 ( \8689 , \8688 , \621 );
not \U$8347 ( \8690 , \8689 );
and \U$8348 ( \8691 , \8687 , \8690 );
and \U$8349 ( \8692 , \8686 , \8689 );
nor \U$8350 ( \8693 , \8691 , \8692 );
not \U$8351 ( \8694 , \8693 );
buf \U$8352 ( \8695 , \8694 );
not \U$8353 ( \8696 , \8695 );
not \U$8354 ( \8697 , \8696 );
xor \U$8355 ( \8698 , \8679 , \8697 );
not \U$8356 ( \8699 , \8698 );
or \U$8357 ( \8700 , \8676 , \8699 );
buf \U$8358 ( \8701 , \8539 );
nand \U$8359 ( \8702 , \8680 , \619 );
and \U$8360 ( \8703 , \8701 , \8702 );
not \U$8361 ( \8704 , \8701 );
not \U$8362 ( \8705 , \8702 );
and \U$8363 ( \8706 , \8704 , \8705 );
nor \U$8364 ( \8707 , \8703 , \8706 );
buf \U$8365 ( \8708 , \8707 );
xor \U$8366 ( \8709 , \5753 , \8708 );
nand \U$8367 ( \8710 , \1162 , \8709 );
nand \U$8368 ( \8711 , \8700 , \8710 );
not \U$8369 ( \8712 , \1013 );
not \U$8370 ( \8713 , \8559 );
or \U$8371 ( \8714 , \8712 , \8713 );
nand \U$8372 ( \8715 , \8537 , \623 );
not \U$8373 ( \8716 , \8715 );
buf \U$8374 ( \8717 , \8543 );
not \U$8375 ( \8718 , \8717 );
or \U$8376 ( \8719 , \8716 , \8718 );
or \U$8377 ( \8720 , \8715 , \8717 );
nand \U$8378 ( \8721 , \8719 , \8720 );
buf \U$8379 ( \8722 , \8721 );
not \U$8380 ( \8723 , \8722 );
and \U$8381 ( \8724 , \3271 , \8723 );
not \U$8382 ( \8725 , \3271 );
and \U$8383 ( \8726 , \8725 , \8722 );
nor \U$8384 ( \8727 , \8724 , \8726 );
nand \U$8385 ( \8728 , \8727 , \1018 );
nand \U$8386 ( \8729 , \8714 , \8728 );
xor \U$8387 ( \8730 , \8711 , \8729 );
not \U$8388 ( \8731 , \8730 );
not \U$8389 ( \8732 , RI9872f40_177);
not \U$8390 ( \8733 , RI9872fb8_178);
and \U$8391 ( \8734 , \8732 , \8733 );
and \U$8392 ( \8735 , RI9872f40_177, RI9872fb8_178);
and \U$8393 ( \8736 , RI9873030_179, RI9872fb8_178);
not \U$8394 ( \8737 , RI9873030_179);
and \U$8395 ( \8738 , \8737 , \8733 );
nor \U$8396 ( \8739 , \8736 , \8738 );
nor \U$8397 ( \8740 , \8734 , \8735 , \8739 );
buf \U$8398 ( \8741 , \8740 );
buf \U$8399 ( \8742 , \8741 );
buf \U$8400 ( \8743 , \8742 );
not \U$8401 ( \8744 , \8743 );
and \U$8402 ( \8745 , RI9872f40_177, \2361 );
not \U$8403 ( \8746 , RI9872f40_177);
and \U$8404 ( \8747 , \8746 , \1691 );
nor \U$8405 ( \8748 , \8745 , \8747 );
not \U$8406 ( \8749 , \8748 );
or \U$8407 ( \8750 , \8744 , \8749 );
buf \U$8408 ( \8751 , \8739 );
buf \U$8409 ( \8752 , \8751 );
nand \U$8410 ( \8753 , \8752 , RI9872f40_177);
nand \U$8411 ( \8754 , \8750 , \8753 );
not \U$8412 ( \8755 , \8754 );
or \U$8413 ( \8756 , \8731 , \8755 );
nand \U$8414 ( \8757 , \8729 , \8711 );
nand \U$8415 ( \8758 , \8756 , \8757 );
xor \U$8416 ( \8759 , \8675 , \8758 );
not \U$8417 ( \8760 , \8759 );
not \U$8418 ( \8761 , \4925 );
and \U$8419 ( \8762 , \3396 , \7993 );
not \U$8420 ( \8763 , \3396 );
and \U$8421 ( \8764 , \8763 , RI9872388_152);
nor \U$8422 ( \8765 , \8762 , \8764 );
not \U$8423 ( \8766 , \8765 );
or \U$8424 ( \8767 , \8761 , \8766 );
not \U$8425 ( \8768 , RI9872388_152);
not \U$8426 ( \8769 , \1485 );
or \U$8427 ( \8770 , \8768 , \8769 );
or \U$8428 ( \8771 , \1485 , RI9872388_152);
nand \U$8429 ( \8772 , \8770 , \8771 );
nand \U$8430 ( \8773 , \8772 , \5942 );
nand \U$8431 ( \8774 , \8767 , \8773 );
not \U$8432 ( \8775 , \8774 );
not \U$8433 ( \8776 , \4085 );
not \U$8434 ( \8777 , RI98725e0_157);
not \U$8435 ( \8778 , \6378 );
or \U$8436 ( \8779 , \8777 , \8778 );
nand \U$8437 ( \8780 , \2110 , \4088 );
nand \U$8438 ( \8781 , \8779 , \8780 );
not \U$8439 ( \8782 , \8781 );
or \U$8440 ( \8783 , \8776 , \8782 );
not \U$8441 ( \8784 , \4088 );
not \U$8442 ( \8785 , \2947 );
not \U$8443 ( \8786 , \8785 );
or \U$8444 ( \8787 , \8784 , \8786 );
nand \U$8445 ( \8788 , \2947 , RI98725e0_157);
nand \U$8446 ( \8789 , \8787 , \8788 );
buf \U$8447 ( \8790 , \4101 );
nand \U$8448 ( \8791 , \8789 , \8790 );
nand \U$8449 ( \8792 , \8783 , \8791 );
not \U$8450 ( \8793 , \8792 );
not \U$8451 ( \8794 , \8793 );
and \U$8452 ( \8795 , RI9872e50_175, RI9872dd8_174);
not \U$8453 ( \8796 , RI9872e50_175);
not \U$8454 ( \8797 , RI9872dd8_174);
and \U$8455 ( \8798 , \8796 , \8797 );
nor \U$8456 ( \8799 , \8795 , \8798 );
buf \U$8457 ( \8800 , \8799 );
buf \U$8458 ( \8801 , \8800 );
buf \U$8459 ( \8802 , \8801 );
not \U$8460 ( \8803 , \8802 );
xor \U$8461 ( \8804 , RI9872d60_173, \1105 );
not \U$8462 ( \8805 , \8804 );
or \U$8463 ( \8806 , \8803 , \8805 );
not \U$8464 ( \8807 , RI9872d60_173);
not \U$8465 ( \8808 , \8807 );
not \U$8466 ( \8809 , \1415 );
or \U$8467 ( \8810 , \8808 , \8809 );
not \U$8468 ( \8811 , RI9872d60_173);
or \U$8469 ( \8812 , \1415 , \8811 );
nand \U$8470 ( \8813 , \8810 , \8812 );
and \U$8471 ( \8814 , \8807 , \8797 );
and \U$8472 ( \8815 , RI9872d60_173, RI9872dd8_174);
nor \U$8473 ( \8816 , \8814 , \8815 , \8799 );
buf \U$8474 ( \8817 , \8816 );
buf \U$8475 ( \8818 , \8817 );
buf \U$8476 ( \8819 , \8818 );
nand \U$8477 ( \8820 , \8813 , \8819 );
nand \U$8478 ( \8821 , \8806 , \8820 );
not \U$8479 ( \8822 , \8821 );
or \U$8480 ( \8823 , \8794 , \8822 );
or \U$8481 ( \8824 , \8821 , \8793 );
nand \U$8482 ( \8825 , \8823 , \8824 );
not \U$8483 ( \8826 , \8825 );
or \U$8484 ( \8827 , \8775 , \8826 );
nand \U$8485 ( \8828 , \8821 , \8792 );
nand \U$8486 ( \8829 , \8827 , \8828 );
not \U$8487 ( \8830 , \8829 );
or \U$8488 ( \8831 , \8760 , \8830 );
nand \U$8489 ( \8832 , \8758 , \8675 );
nand \U$8490 ( \8833 , \8831 , \8832 );
not \U$8491 ( \8834 , \8833 );
not \U$8492 ( \8835 , \8834 );
not \U$8493 ( \8836 , \1353 );
not \U$8494 ( \8837 , \8652 );
or \U$8495 ( \8838 , \8836 , \8837 );
buf \U$8496 ( \8839 , \8573 );
not \U$8497 ( \8840 , \8839 );
buf \U$8498 ( \8841 , \8840 );
buf \U$8499 ( \8842 , \8841 );
and \U$8500 ( \8843 , RI9871e60_141, \8842 );
not \U$8501 ( \8844 , RI9871e60_141);
not \U$8502 ( \8845 , \8841 );
and \U$8503 ( \8846 , \8844 , \8845 );
or \U$8504 ( \8847 , \8843 , \8846 );
nand \U$8505 ( \8848 , \8847 , \1381 );
nand \U$8506 ( \8849 , \8838 , \8848 );
not \U$8507 ( \8850 , \8849 );
not \U$8508 ( \8851 , \832 );
not \U$8509 ( \8852 , \8609 );
or \U$8510 ( \8853 , \8851 , \8852 );
not \U$8511 ( \8854 , RI9871d70_139);
not \U$8512 ( \8855 , \8668 );
or \U$8513 ( \8856 , \8854 , \8855 );
buf \U$8514 ( \8857 , \8667 );
not \U$8515 ( \8858 , \8857 );
not \U$8516 ( \8859 , RI9871d70_139);
nand \U$8517 ( \8860 , \8858 , \8859 );
nand \U$8518 ( \8861 , \8856 , \8860 );
nand \U$8519 ( \8862 , \8861 , \5350 );
nand \U$8520 ( \8863 , \8853 , \8862 );
not \U$8521 ( \8864 , \8863 );
not \U$8522 ( \8865 , \924 );
and \U$8523 ( \8866 , \8074 , \919 );
not \U$8524 ( \8867 , \8074 );
and \U$8525 ( \8868 , \8867 , RI9872130_147);
nor \U$8526 ( \8869 , \8866 , \8868 );
not \U$8527 ( \8870 , \8869 );
or \U$8528 ( \8871 , \8865 , \8870 );
not \U$8529 ( \8872 , RI9872130_147);
not \U$8530 ( \8873 , \8618 );
not \U$8531 ( \8874 , \8873 );
not \U$8532 ( \8875 , \8874 );
or \U$8533 ( \8876 , \8872 , \8875 );
buf \U$8534 ( \8877 , \8619 );
not \U$8535 ( \8878 , \8877 );
or \U$8536 ( \8879 , \8878 , RI9872130_147);
nand \U$8537 ( \8880 , \8876 , \8879 );
nand \U$8538 ( \8881 , \8880 , \876 );
nand \U$8539 ( \8882 , \8871 , \8881 );
not \U$8540 ( \8883 , \8882 );
not \U$8541 ( \8884 , \8883 );
or \U$8542 ( \8885 , \8864 , \8884 );
or \U$8543 ( \8886 , \8863 , \8883 );
nand \U$8544 ( \8887 , \8885 , \8886 );
not \U$8545 ( \8888 , \8887 );
or \U$8546 ( \8889 , \8850 , \8888 );
nand \U$8547 ( \8890 , \8882 , \8863 );
nand \U$8548 ( \8891 , \8889 , \8890 );
not \U$8549 ( \8892 , \8891 );
not \U$8550 ( \8893 , \1430 );
not \U$8551 ( \8894 , RI9871c08_136);
not \U$8552 ( \8895 , \6303 );
not \U$8553 ( \8896 , \8895 );
or \U$8554 ( \8897 , \8894 , \8896 );
or \U$8555 ( \8898 , \6308 , RI9871c08_136);
nand \U$8556 ( \8899 , \8897 , \8898 );
not \U$8557 ( \8900 , \8899 );
or \U$8558 ( \8901 , \8893 , \8900 );
not \U$8559 ( \8902 , RI9871c08_136);
buf \U$8560 ( \8903 , \8052 );
buf \U$8561 ( \8904 , \8903 );
not \U$8562 ( \8905 , \8904 );
or \U$8563 ( \8906 , \8902 , \8905 );
or \U$8564 ( \8907 , \8904 , RI9871c08_136);
nand \U$8565 ( \8908 , \8906 , \8907 );
nand \U$8566 ( \8909 , \8908 , \1455 );
nand \U$8567 ( \8910 , \8901 , \8909 );
not \U$8568 ( \8911 , \8910 );
not \U$8569 ( \8912 , \1501 );
and \U$8570 ( \8913 , RI9871c80_137, \8334 );
not \U$8571 ( \8914 , RI9871c80_137);
buf \U$8572 ( \8915 , \8332 );
not \U$8573 ( \8916 , \8915 );
and \U$8574 ( \8917 , \8914 , \8916 );
or \U$8575 ( \8918 , \8913 , \8917 );
not \U$8576 ( \8919 , \8918 );
or \U$8577 ( \8920 , \8912 , \8919 );
and \U$8578 ( \8921 , RI9871c80_137, \7466 );
not \U$8579 ( \8922 , RI9871c80_137);
not \U$8580 ( \8923 , \7465 );
not \U$8581 ( \8924 , \8923 );
not \U$8582 ( \8925 , \8924 );
and \U$8583 ( \8926 , \8922 , \8925 );
or \U$8584 ( \8927 , \8921 , \8926 );
nand \U$8585 ( \8928 , \8927 , \1518 );
nand \U$8586 ( \8929 , \8920 , \8928 );
not \U$8587 ( \8930 , \8929 );
or \U$8588 ( \8931 , \8911 , \8930 );
or \U$8589 ( \8932 , \8910 , \8929 );
not \U$8590 ( \8933 , \1323 );
not \U$8591 ( \8934 , \6529 );
and \U$8592 ( \8935 , \8934 , RI9871b18_134);
not \U$8593 ( \8936 , \8934 );
and \U$8594 ( \8937 , \8936 , \2479 );
nor \U$8595 ( \8938 , \8935 , \8937 );
not \U$8596 ( \8939 , \8938 );
or \U$8597 ( \8940 , \8933 , \8939 );
not \U$8598 ( \8941 , \4044 );
not \U$8599 ( \8942 , \7002 );
not \U$8600 ( \8943 , \8942 );
not \U$8601 ( \8944 , \8943 );
not \U$8602 ( \8945 , \8944 );
or \U$8603 ( \8946 , \8941 , \8945 );
not \U$8604 ( \8947 , \7002 );
not \U$8605 ( \8948 , \8947 );
nand \U$8606 ( \8949 , \8948 , RI9871b18_134);
nand \U$8607 ( \8950 , \8946 , \8949 );
nand \U$8608 ( \8951 , \8950 , \1292 );
nand \U$8609 ( \8952 , \8940 , \8951 );
nand \U$8610 ( \8953 , \8932 , \8952 );
nand \U$8611 ( \8954 , \8931 , \8953 );
and \U$8612 ( \8955 , RI9872fb8_178, RI9873030_179);
nor \U$8613 ( \8956 , \8955 , \8732 );
not \U$8614 ( \8957 , \8956 );
and \U$8615 ( \8958 , \5753 , \8708 );
not \U$8616 ( \8959 , \8958 );
or \U$8617 ( \8960 , \8957 , \8959 );
or \U$8618 ( \8961 , \8958 , \8956 );
nand \U$8619 ( \8962 , \8960 , \8961 );
not \U$8620 ( \8963 , \1455 );
not \U$8621 ( \8964 , \8899 );
or \U$8622 ( \8965 , \8963 , \8964 );
and \U$8623 ( \8966 , \6481 , \1850 );
not \U$8624 ( \8967 , \6481 );
and \U$8625 ( \8968 , \8967 , RI9871c08_136);
nor \U$8626 ( \8969 , \8966 , \8968 );
nand \U$8627 ( \8970 , \8969 , \1430 );
nand \U$8628 ( \8971 , \8965 , \8970 );
xor \U$8629 ( \8972 , \8962 , \8971 );
buf \U$8630 ( \8973 , \8972 );
xor \U$8631 ( \8974 , \8954 , \8973 );
not \U$8632 ( \8975 , \8974 );
or \U$8633 ( \8976 , \8892 , \8975 );
nand \U$8634 ( \8977 , \8954 , \8973 );
nand \U$8635 ( \8978 , \8976 , \8977 );
not \U$8636 ( \8979 , \8978 );
not \U$8637 ( \8980 , \1323 );
and \U$8638 ( \8981 , \5707 , \1283 );
not \U$8639 ( \8982 , \5707 );
and \U$8640 ( \8983 , \8982 , RI9871b18_134);
nor \U$8641 ( \8984 , \8981 , \8983 );
not \U$8642 ( \8985 , \8984 );
or \U$8643 ( \8986 , \8980 , \8985 );
and \U$8644 ( \8987 , RI9871b18_134, \8054 );
not \U$8645 ( \8988 , RI9871b18_134);
and \U$8646 ( \8989 , \8988 , \6298 );
or \U$8647 ( \8990 , \8987 , \8989 );
nand \U$8648 ( \8991 , \8990 , \1292 );
nand \U$8649 ( \8992 , \8986 , \8991 );
not \U$8650 ( \8993 , \8992 );
not \U$8651 ( \8994 , \8962 );
not \U$8652 ( \8995 , \8971 );
or \U$8653 ( \8996 , \8994 , \8995 );
not \U$8654 ( \8997 , \8956 );
nand \U$8655 ( \8998 , \8997 , \8958 );
nand \U$8656 ( \8999 , \8996 , \8998 );
xor \U$8657 ( \9000 , \8993 , \8999 );
not \U$8658 ( \9001 , \1518 );
not \U$8659 ( \9002 , \1584 );
not \U$8660 ( \9003 , \7004 );
or \U$8661 ( \9004 , \9002 , \9003 );
nand \U$8662 ( \9005 , \8081 , RI9871c80_137);
nand \U$8663 ( \9006 , \9004 , \9005 );
not \U$8664 ( \9007 , \9006 );
or \U$8665 ( \9008 , \9001 , \9007 );
nand \U$8666 ( \9009 , \8927 , \1501 );
nand \U$8667 ( \9010 , \9008 , \9009 );
not \U$8668 ( \9011 , \876 );
not \U$8669 ( \9012 , \8869 );
or \U$8670 ( \9013 , \9011 , \9012 );
not \U$8671 ( \9014 , \919 );
not \U$8672 ( \9015 , \8335 );
or \U$8673 ( \9016 , \9014 , \9015 );
nand \U$8674 ( \9017 , \8334 , RI9872130_147);
nand \U$8675 ( \9018 , \9016 , \9017 );
nand \U$8676 ( \9019 , \9018 , \924 );
nand \U$8677 ( \9020 , \9013 , \9019 );
xor \U$8678 ( \9021 , \9010 , \9020 );
not \U$8679 ( \9022 , \1292 );
not \U$8680 ( \9023 , \8938 );
or \U$8681 ( \9024 , \9022 , \9023 );
nand \U$8682 ( \9025 , \8990 , \1323 );
nand \U$8683 ( \9026 , \9024 , \9025 );
and \U$8684 ( \9027 , \9021 , \9026 );
and \U$8685 ( \9028 , \9010 , \9020 );
or \U$8686 ( \9029 , \9027 , \9028 );
not \U$8687 ( \9030 , \9029 );
and \U$8688 ( \9031 , \9000 , \9030 );
not \U$8689 ( \9032 , \9000 );
and \U$8690 ( \9033 , \9032 , \9029 );
nor \U$8691 ( \9034 , \9031 , \9033 );
not \U$8692 ( \9035 , \9034 );
and \U$8693 ( \9036 , \8979 , \9035 );
and \U$8694 ( \9037 , \8978 , \9034 );
nor \U$8695 ( \9038 , \9036 , \9037 );
not \U$8696 ( \9039 , \9038 );
not \U$8697 ( \9040 , \9039 );
or \U$8698 ( \9041 , \8835 , \9040 );
nand \U$8699 ( \9042 , \9038 , \8833 );
nand \U$8700 ( \9043 , \9041 , \9042 );
not \U$8701 ( \9044 , \9043 );
xor \U$8702 ( \9045 , \8730 , \8754 );
not \U$8703 ( \9046 , \9045 );
not \U$8704 ( \9047 , \9046 );
xor \U$8705 ( \9048 , \8929 , \8910 );
xnor \U$8706 ( \9049 , \9048 , \8952 );
not \U$8707 ( \9050 , \9049 );
not \U$8708 ( \9051 , \9050 );
or \U$8709 ( \9052 , \9047 , \9051 );
nand \U$8710 ( \9053 , \9049 , \9045 );
nand \U$8711 ( \9054 , \9052 , \9053 );
not \U$8712 ( \9055 , \9054 );
not \U$8713 ( \9056 , \3467 );
xor \U$8714 ( \9057 , RI98726d0_159, \3543 );
not \U$8715 ( \9058 , \9057 );
or \U$8716 ( \9059 , \9056 , \9058 );
and \U$8717 ( \9060 , \3568 , \4063 );
not \U$8718 ( \9061 , \3568 );
and \U$8719 ( \9062 , \9061 , RI98726d0_159);
nor \U$8720 ( \9063 , \9060 , \9062 );
nand \U$8721 ( \9064 , \9063 , \3466 );
nand \U$8722 ( \9065 , \9059 , \9064 );
not \U$8723 ( \9066 , \9065 );
and \U$8724 ( \9067 , RI9872a18_166, \820 );
not \U$8725 ( \9068 , RI9872a18_166);
and \U$8726 ( \9069 , \9068 , \6219 );
or \U$8727 ( \9070 , \9067 , \9069 );
buf \U$8728 ( \9071 , \8039 );
buf \U$8729 ( \9072 , \9071 );
nand \U$8730 ( \9073 , \9070 , \9072 );
not \U$8731 ( \9074 , RI9872a18_166);
not \U$8732 ( \9075 , \6224 );
or \U$8733 ( \9076 , \9074 , \9075 );
or \U$8734 ( \9077 , \6224 , RI9872a18_166);
nand \U$8735 ( \9078 , \9076 , \9077 );
buf \U$8736 ( \9079 , \8028 );
nand \U$8737 ( \9080 , \9078 , \9079 );
nand \U$8738 ( \9081 , \9073 , \9080 );
buf \U$8739 ( \9082 , \466 );
not \U$8740 ( \9083 , \9082 );
buf \U$8741 ( \9084 , \460 );
not \U$8742 ( \9085 , \9084 );
nor \U$8743 ( \9086 , \9083 , \9085 , \593 );
not \U$8744 ( \9087 , \9086 );
not \U$8745 ( \9088 , \523 );
not \U$8746 ( \9089 , \534 );
not \U$8747 ( \9090 , \515 );
or \U$8748 ( \9091 , \9089 , \9090 );
not \U$8749 ( \9092 , \587 );
nand \U$8750 ( \9093 , \9091 , \9092 );
not \U$8751 ( \9094 , \9093 );
or \U$8752 ( \9095 , \9088 , \9094 );
not \U$8753 ( \9096 , \493 );
nand \U$8754 ( \9097 , \9095 , \9096 );
not \U$8755 ( \9098 , \9097 );
or \U$8756 ( \9099 , \9087 , \9098 );
not \U$8757 ( \9100 , \463 );
buf \U$8758 ( \9101 , \604 );
not \U$8759 ( \9102 , \9101 );
or \U$8760 ( \9103 , \9100 , \9102 );
nand \U$8761 ( \9104 , \9103 , \607 );
not \U$8762 ( \9105 , \9104 );
nand \U$8763 ( \9106 , \9099 , \9105 );
not \U$8764 ( \9107 , \9106 );
nand \U$8765 ( \9108 , \469 , \609 );
not \U$8766 ( \9109 , \9108 );
and \U$8767 ( \9110 , \9107 , \9109 );
and \U$8768 ( \9111 , \9106 , \9108 );
nor \U$8769 ( \9112 , \9110 , \9111 );
buf \U$8770 ( \9113 , \9112 );
buf \U$8771 ( \9114 , \9113 );
not \U$8772 ( \9115 , \9114 );
not \U$8773 ( \9116 , \9115 );
not \U$8774 ( \9117 , \1166 );
and \U$8775 ( \9118 , \9116 , \9117 );
not \U$8776 ( \9119 , \9113 );
not \U$8777 ( \9120 , \8678 );
and \U$8778 ( \9121 , \9119 , \9120 );
nor \U$8779 ( \9122 , \9118 , \9121 );
not \U$8780 ( \9123 , \9122 );
nand \U$8781 ( \9124 , \9123 , \6316 );
nand \U$8782 ( \9125 , \463 , \607 );
not \U$8783 ( \9126 , \9125 );
not \U$8784 ( \9127 , \9082 );
nor \U$8785 ( \9128 , \9127 , \9085 );
not \U$8786 ( \9129 , \9128 );
not \U$8787 ( \9130 , \9097 );
or \U$8788 ( \9131 , \9129 , \9130 );
not \U$8789 ( \9132 , \9101 );
nand \U$8790 ( \9133 , \9131 , \9132 );
not \U$8791 ( \9134 , \9133 );
or \U$8792 ( \9135 , \9126 , \9134 );
or \U$8793 ( \9136 , \9125 , \9133 );
nand \U$8794 ( \9137 , \9135 , \9136 );
buf \U$8795 ( \9138 , \9137 );
buf \U$8796 ( \9139 , \9138 );
xor \U$8797 ( \9140 , \8679 , \9139 );
nand \U$8798 ( \9141 , \9140 , \1162 );
and \U$8799 ( \9142 , \9124 , \9141 );
and \U$8800 ( \9143 , \9081 , \9142 );
not \U$8801 ( \9144 , \9081 );
not \U$8802 ( \9145 , \9142 );
and \U$8803 ( \9146 , \9144 , \9145 );
or \U$8804 ( \9147 , \9143 , \9146 );
not \U$8805 ( \9148 , \9147 );
or \U$8806 ( \9149 , \9066 , \9148 );
not \U$8807 ( \9150 , \9080 );
not \U$8808 ( \9151 , \9073 );
or \U$8809 ( \9152 , \9150 , \9151 );
nand \U$8810 ( \9153 , \9152 , \9145 );
nand \U$8811 ( \9154 , \9149 , \9153 );
not \U$8812 ( \9155 , \9154 );
or \U$8813 ( \9156 , \9055 , \9155 );
nand \U$8814 ( \9157 , \9050 , \9045 );
nand \U$8815 ( \9158 , \9156 , \9157 );
not \U$8816 ( \9159 , \9158 );
not \U$8817 ( \9160 , \4918 );
not \U$8818 ( \9161 , RI9872388_152);
not \U$8819 ( \9162 , \2110 );
not \U$8820 ( \9163 , \9162 );
or \U$8821 ( \9164 , \9161 , \9163 );
or \U$8822 ( \9165 , \6378 , RI9872388_152);
nand \U$8823 ( \9166 , \9164 , \9165 );
not \U$8824 ( \9167 , \9166 );
or \U$8825 ( \9168 , \9160 , \9167 );
nand \U$8826 ( \9169 , \8772 , \5047 );
nand \U$8827 ( \9170 , \9168 , \9169 );
not \U$8828 ( \9171 , \9170 );
not \U$8829 ( \9172 , \4084 );
not \U$8830 ( \9173 , \8789 );
or \U$8831 ( \9174 , \9172 , \9173 );
not \U$8832 ( \9175 , RI98725e0_157);
not \U$8833 ( \9176 , \4370 );
or \U$8834 ( \9177 , \9175 , \9176 );
nand \U$8835 ( \9178 , \3240 , \3454 );
nand \U$8836 ( \9179 , \9177 , \9178 );
nand \U$8837 ( \9180 , \9179 , \4101 );
nand \U$8838 ( \9181 , \9174 , \9180 );
not \U$8839 ( \9182 , \9181 );
nand \U$8840 ( \9183 , \9171 , \9182 );
not \U$8841 ( \9184 , \9183 );
not \U$8842 ( \9185 , RI9872bf8_170);
not \U$8843 ( \9186 , RI9872c70_171);
nand \U$8844 ( \9187 , \9185 , \9186 );
nand \U$8845 ( \9188 , RI9872bf8_170, RI9872c70_171);
and \U$8846 ( \9189 , \9187 , \9188 );
and \U$8847 ( \9190 , RI9872b80_169, \9186 );
not \U$8848 ( \9191 , RI9872b80_169);
and \U$8849 ( \9192 , \9191 , RI9872c70_171);
nor \U$8850 ( \9193 , \9190 , \9192 );
nor \U$8851 ( \9194 , \9189 , \9193 );
buf \U$8852 ( \9195 , \9194 );
buf \U$8853 ( \9196 , \9195 );
not \U$8854 ( \9197 , \9196 );
not \U$8855 ( \9198 , RI9872b80_169);
not \U$8856 ( \9199 , \9198 );
not \U$8857 ( \9200 , \891 );
or \U$8858 ( \9201 , \9199 , \9200 );
not \U$8859 ( \9202 , \879 );
not \U$8860 ( \9203 , \887 );
or \U$8861 ( \9204 , \9202 , \9203 );
nand \U$8862 ( \9205 , \9204 , \890 );
or \U$8863 ( \9206 , \9205 , \9198 );
nand \U$8864 ( \9207 , \9201 , \9206 );
not \U$8865 ( \9208 , \9207 );
or \U$8866 ( \9209 , \9197 , \9208 );
and \U$8867 ( \9210 , \6585 , \9198 );
not \U$8868 ( \9211 , \6585 );
and \U$8869 ( \9212 , \9211 , RI9872b80_169);
nor \U$8870 ( \9213 , \9210 , \9212 );
buf \U$8871 ( \9214 , \9189 );
nand \U$8872 ( \9215 , \9213 , \9214 );
nand \U$8873 ( \9216 , \9209 , \9215 );
not \U$8874 ( \9217 , \9216 );
or \U$8875 ( \9218 , \9184 , \9217 );
nand \U$8876 ( \9219 , \9181 , \9170 );
nand \U$8877 ( \9220 , \9218 , \9219 );
not \U$8878 ( \9221 , \9220 );
and \U$8879 ( \9222 , RI9872ce8_172, RI9872d60_173);
not \U$8880 ( \9223 , RI9872ce8_172);
and \U$8881 ( \9224 , \9223 , \8807 );
nor \U$8882 ( \9225 , \9222 , \9224 );
buf \U$8883 ( \9226 , \9225 );
buf \U$8884 ( \9227 , \9226 );
not \U$8885 ( \9228 , \9227 );
not \U$8886 ( \9229 , RI9872bf8_170);
buf \U$8887 ( \9230 , \1318 );
not \U$8888 ( \9231 , \9230 );
or \U$8889 ( \9232 , \9229 , \9231 );
or \U$8890 ( \9233 , \1320 , RI9872bf8_170);
nand \U$8891 ( \9234 , \9232 , \9233 );
not \U$8892 ( \9235 , \9234 );
or \U$8893 ( \9236 , \9228 , \9235 );
not \U$8894 ( \9237 , RI9872bf8_170);
not \U$8895 ( \9238 , \1581 );
or \U$8896 ( \9239 , \9237 , \9238 );
or \U$8897 ( \9240 , \1581 , RI9872bf8_170);
nand \U$8898 ( \9241 , \9239 , \9240 );
or \U$8899 ( \9242 , RI9872bf8_170, RI9872ce8_172);
not \U$8900 ( \9243 , RI9872ce8_172);
not \U$8901 ( \9244 , RI9872bf8_170);
or \U$8902 ( \9245 , \9243 , \9244 );
not \U$8903 ( \9246 , \9225 );
nand \U$8904 ( \9247 , \9242 , \9245 , \9246 );
not \U$8905 ( \9248 , \9247 );
buf \U$8906 ( \9249 , \9248 );
nand \U$8907 ( \9250 , \9241 , \9249 );
nand \U$8908 ( \9251 , \9236 , \9250 );
not \U$8909 ( \9252 , \5034 );
not \U$8910 ( \9253 , RI9872478_154);
buf \U$8911 ( \9254 , \3394 );
buf \U$8912 ( \9255 , \9254 );
not \U$8913 ( \9256 , \9255 );
or \U$8914 ( \9257 , \9253 , \9256 );
or \U$8915 ( \9258 , \3396 , RI9872478_154);
nand \U$8916 ( \9259 , \9257 , \9258 );
not \U$8917 ( \9260 , \9259 );
or \U$8918 ( \9261 , \9252 , \9260 );
not \U$8919 ( \9262 , \1208 );
not \U$8920 ( \9263 , \9262 );
and \U$8921 ( \9264 , RI9872478_154, \9263 );
not \U$8922 ( \9265 , RI9872478_154);
and \U$8923 ( \9266 , \9265 , \6020 );
or \U$8924 ( \9267 , \9264 , \9266 );
nand \U$8925 ( \9268 , \9267 , \6698 );
nand \U$8926 ( \9269 , \9261 , \9268 );
or \U$8927 ( \9270 , \9251 , \9269 );
xor \U$8928 ( \9271 , RI9872ec8_176, RI9872f40_177);
buf \U$8929 ( \9272 , \9271 );
buf \U$8930 ( \9273 , \9272 );
not \U$8931 ( \9274 , \9273 );
not \U$8932 ( \9275 , RI9872e50_175);
not \U$8933 ( \9276 , \1126 );
not \U$8934 ( \9277 , \9276 );
or \U$8935 ( \9278 , \9275 , \9277 );
or \U$8936 ( \9279 , \9276 , RI9872e50_175);
nand \U$8937 ( \9280 , \9278 , \9279 );
not \U$8938 ( \9281 , \9280 );
or \U$8939 ( \9282 , \9274 , \9281 );
and \U$8940 ( \9283 , RI9872e50_175, \1106 );
not \U$8941 ( \9284 , RI9872e50_175);
and \U$8942 ( \9285 , \9284 , \1097 );
nor \U$8943 ( \9286 , \9283 , \9285 );
not \U$8944 ( \9287 , \9271 );
and \U$8945 ( \9288 , RI9872e50_175, RI9872ec8_176);
not \U$8946 ( \9289 , RI9872e50_175);
not \U$8947 ( \9290 , RI9872ec8_176);
and \U$8948 ( \9291 , \9289 , \9290 );
nor \U$8949 ( \9292 , \9288 , \9291 );
and \U$8950 ( \9293 , \9287 , \9292 );
buf \U$8951 ( \9294 , \9293 );
nand \U$8952 ( \9295 , \9286 , \9294 );
nand \U$8953 ( \9296 , \9282 , \9295 );
nand \U$8954 ( \9297 , \9270 , \9296 );
nand \U$8955 ( \9298 , \9269 , \9251 );
and \U$8956 ( \9299 , \9221 , \9297 , \9298 );
not \U$8957 ( \9300 , \6284 );
xnor \U$8958 ( \9301 , \1603 , RI98728b0_163);
not \U$8959 ( \9302 , \9301 );
or \U$8960 ( \9303 , \9300 , \9302 );
not \U$8961 ( \9304 , RI98728b0_163);
not \U$8962 ( \9305 , \1340 );
or \U$8963 ( \9306 , \9304 , \9305 );
nand \U$8964 ( \9307 , \5712 , \5632 );
nand \U$8965 ( \9308 , \9306 , \9307 );
nand \U$8966 ( \9309 , \9308 , \6286 );
nand \U$8967 ( \9310 , \9303 , \9309 );
not \U$8968 ( \9311 , \9310 );
buf \U$8969 ( \9312 , \8818 );
not \U$8970 ( \9313 , \9312 );
not \U$8971 ( \9314 , \1446 );
xor \U$8972 ( \9315 , RI9872d60_173, \9314 );
not \U$8973 ( \9316 , \9315 );
or \U$8974 ( \9317 , \9313 , \9316 );
nand \U$8975 ( \9318 , \8813 , \8802 );
nand \U$8976 ( \9319 , \9317 , \9318 );
buf \U$8977 ( \9320 , \5641 );
not \U$8978 ( \9321 , \9320 );
not \U$8979 ( \9322 , RI9872568_156);
not \U$8980 ( \9323 , \1038 );
not \U$8981 ( \9324 , \9323 );
or \U$8982 ( \9325 , \9322 , \9324 );
not \U$8983 ( \9326 , \1038 );
or \U$8984 ( \9327 , \9326 , RI9872568_156);
nand \U$8985 ( \9328 , \9325 , \9327 );
not \U$8986 ( \9329 , \9328 );
or \U$8987 ( \9330 , \9321 , \9329 );
xor \U$8988 ( \9331 , RI9872568_156, \1062 );
nand \U$8989 ( \9332 , \9331 , \7188 );
nand \U$8990 ( \9333 , \9330 , \9332 );
or \U$8991 ( \9334 , \9319 , \9333 );
not \U$8992 ( \9335 , \9334 );
or \U$8993 ( \9336 , \9311 , \9335 );
nand \U$8994 ( \9337 , \9319 , \9333 );
nand \U$8995 ( \9338 , \9336 , \9337 );
not \U$8996 ( \9339 , \9338 );
or \U$8997 ( \9340 , \9299 , \9339 );
not \U$8998 ( \9341 , \9297 );
not \U$8999 ( \9342 , \9298 );
or \U$9000 ( \9343 , \9341 , \9342 );
nand \U$9001 ( \9344 , \9343 , \9220 );
nand \U$9002 ( \9345 , \9340 , \9344 );
not \U$9003 ( \9346 , \9345 );
xor \U$9004 ( \9347 , \8972 , \8954 );
xor \U$9005 ( \9348 , \9347 , \8891 );
buf \U$9006 ( \9349 , \9348 );
not \U$9007 ( \9350 , \9349 );
and \U$9008 ( \9351 , \9346 , \9350 );
not \U$9009 ( \9352 , \9346 );
and \U$9010 ( \9353 , \9352 , \9349 );
nor \U$9011 ( \9354 , \9351 , \9353 );
not \U$9012 ( \9355 , \9354 );
or \U$9013 ( \9356 , \9159 , \9355 );
nand \U$9014 ( \9357 , \9345 , \9349 );
nand \U$9015 ( \9358 , \9356 , \9357 );
not \U$9016 ( \9359 , \9358 );
not \U$9017 ( \9360 , \9359 );
or \U$9018 ( \9361 , \9044 , \9360 );
or \U$9019 ( \9362 , \9359 , \9043 );
nand \U$9020 ( \9363 , \9361 , \9362 );
not \U$9021 ( \9364 , \6145 );
and \U$9022 ( \9365 , RI98719b0_131, \7791 );
not \U$9023 ( \9366 , RI98719b0_131);
not \U$9024 ( \9367 , \7791 );
and \U$9025 ( \9368 , \9366 , \9367 );
or \U$9026 ( \9369 , \9365 , \9368 );
not \U$9027 ( \9370 , \9369 );
or \U$9028 ( \9371 , \9364 , \9370 );
and \U$9029 ( \9372 , RI98719b0_131, \4986 );
not \U$9030 ( \9373 , RI98719b0_131);
not \U$9031 ( \9374 , \4985 );
and \U$9032 ( \9375 , \9373 , \9374 );
nor \U$9033 ( \9376 , \9372 , \9375 );
not \U$9034 ( \9377 , \9376 );
nand \U$9035 ( \9378 , \9377 , \793 );
nand \U$9036 ( \9379 , \9371 , \9378 );
not \U$9037 ( \9380 , \9379 );
not \U$9038 ( \9381 , \6673 );
and \U$9039 ( \9382 , \5776 , \1111 );
not \U$9040 ( \9383 , \5776 );
and \U$9041 ( \9384 , \9383 , RI98718c0_129);
nor \U$9042 ( \9385 , \9382 , \9384 );
not \U$9043 ( \9386 , \9385 );
or \U$9044 ( \9387 , \9381 , \9386 );
xor \U$9045 ( \9388 , \5766 , RI98718c0_129);
nand \U$9046 ( \9389 , \9388 , \1083 );
nand \U$9047 ( \9390 , \9387 , \9389 );
not \U$9048 ( \9391 , \6284 );
not \U$9049 ( \9392 , \9308 );
or \U$9050 ( \9393 , \9391 , \9392 );
and \U$9051 ( \9394 , RI98728b0_163, \5720 );
not \U$9052 ( \9395 , RI98728b0_163);
and \U$9053 ( \9396 , \9395 , \1254 );
or \U$9054 ( \9397 , \9394 , \9396 );
nand \U$9055 ( \9398 , \9397 , \6611 );
nand \U$9056 ( \9399 , \9393 , \9398 );
xor \U$9057 ( \9400 , \9390 , \9399 );
not \U$9058 ( \9401 , \9400 );
or \U$9059 ( \9402 , \9380 , \9401 );
nand \U$9060 ( \9403 , \9399 , \9390 );
nand \U$9061 ( \9404 , \9402 , \9403 );
not \U$9062 ( \9405 , \9404 );
not \U$9063 ( \9406 , \6653 );
not \U$9064 ( \9407 , RI9872310_151);
not \U$9065 ( \9408 , \4176 );
or \U$9066 ( \9409 , \9407 , \9408 );
or \U$9067 ( \9410 , \5596 , RI9872310_151);
nand \U$9068 ( \9411 , \9409 , \9410 );
not \U$9069 ( \9412 , \9411 );
or \U$9070 ( \9413 , \9406 , \9412 );
and \U$9071 ( \9414 , RI9872310_151, \3568 );
not \U$9072 ( \9415 , RI9872310_151);
and \U$9073 ( \9416 , \9415 , \3569 );
or \U$9074 ( \9417 , \9414 , \9416 );
nand \U$9075 ( \9418 , \9417 , \3170 );
nand \U$9076 ( \9419 , \9413 , \9418 );
not \U$9077 ( \9420 , \9419 );
and \U$9078 ( \9421 , RI98730a8_180, RI9873120_181);
not \U$9079 ( \9422 , \9421 );
nand \U$9080 ( \9423 , \9422 , RI9873030_179);
and \U$9081 ( \9424 , \8679 , \9139 );
xor \U$9082 ( \9425 , \9423 , \9424 );
not \U$9083 ( \9426 , \8709 );
not \U$9084 ( \9427 , \6316 );
or \U$9085 ( \9428 , \9426 , \9427 );
buf \U$9086 ( \9429 , \1161 );
not \U$9087 ( \9430 , \9429 );
or \U$9088 ( \9431 , \9122 , \9430 );
nand \U$9089 ( \9432 , \9428 , \9431 );
and \U$9090 ( \9433 , \9425 , \9432 );
and \U$9091 ( \9434 , \9423 , \9424 );
nor \U$9092 ( \9435 , \9433 , \9434 );
buf \U$9093 ( \9436 , \9435 );
not \U$9094 ( \9437 , \2087 );
not \U$9095 ( \9438 , \2076 );
not \U$9096 ( \9439 , \4409 );
or \U$9097 ( \9440 , \9438 , \9439 );
nand \U$9098 ( \9441 , \5205 , RI9871aa0_133);
nand \U$9099 ( \9442 , \9440 , \9441 );
not \U$9100 ( \9443 , \9442 );
or \U$9101 ( \9444 , \9437 , \9443 );
not \U$9102 ( \9445 , \2080 );
not \U$9103 ( \9446 , \4472 );
or \U$9104 ( \9447 , \9445 , \9446 );
nand \U$9105 ( \9448 , \4470 , RI9871aa0_133);
nand \U$9106 ( \9449 , \9447 , \9448 );
nand \U$9107 ( \9450 , \9449 , \2071 );
nand \U$9108 ( \9451 , \9444 , \9450 );
xnor \U$9109 ( \9452 , \9436 , \9451 );
not \U$9110 ( \9453 , \9452 );
or \U$9111 ( \9454 , \9420 , \9453 );
not \U$9112 ( \9455 , \9436 );
nand \U$9113 ( \9456 , \9455 , \9451 );
nand \U$9114 ( \9457 , \9454 , \9456 );
not \U$9115 ( \9458 , \9457 );
xor \U$9116 ( \9459 , \9405 , \9458 );
not \U$9117 ( \9460 , \3467 );
not \U$9118 ( \9461 , \4369 );
and \U$9119 ( \9462 , \9461 , \4063 );
not \U$9120 ( \9463 , \9461 );
and \U$9121 ( \9464 , \9463 , RI98726d0_159);
nor \U$9122 ( \9465 , \9462 , \9464 );
not \U$9123 ( \9466 , \9465 );
or \U$9124 ( \9467 , \9460 , \9466 );
nand \U$9125 ( \9468 , \9057 , \3466 );
nand \U$9126 ( \9469 , \9467 , \9468 );
not \U$9127 ( \9470 , \9469 );
not \U$9128 ( \9471 , \7338 );
not \U$9129 ( \9472 , RI98729a0_165);
not \U$9130 ( \9473 , \6225 );
or \U$9131 ( \9474 , \9472 , \9473 );
or \U$9132 ( \9475 , \2216 , RI98729a0_165);
nand \U$9133 ( \9476 , \9474 , \9475 );
not \U$9134 ( \9477 , \9476 );
or \U$9135 ( \9478 , \9471 , \9477 );
not \U$9136 ( \9479 , \7328 );
not \U$9137 ( \9480 , \1550 );
or \U$9138 ( \9481 , \9479 , \9480 );
or \U$9139 ( \9482 , \7328 , \944 );
nand \U$9140 ( \9483 , \9481 , \9482 );
nand \U$9141 ( \9484 , \9483 , \7325 );
nand \U$9142 ( \9485 , \9478 , \9484 );
not \U$9143 ( \9486 , \9485 );
not \U$9144 ( \9487 , \9486 );
not \U$9145 ( \9488 , \9072 );
and \U$9146 ( \9489 , \893 , \8031 );
not \U$9147 ( \9490 , \893 );
and \U$9148 ( \9491 , \9490 , RI9872a18_166);
nor \U$9149 ( \9492 , \9489 , \9491 );
not \U$9150 ( \9493 , \9492 );
or \U$9151 ( \9494 , \9488 , \9493 );
nand \U$9152 ( \9495 , \9070 , \9079 );
nand \U$9153 ( \9496 , \9494 , \9495 );
not \U$9154 ( \9497 , \9496 );
or \U$9155 ( \9498 , \9487 , \9497 );
or \U$9156 ( \9499 , \9496 , \9486 );
nand \U$9157 ( \9500 , \9498 , \9499 );
not \U$9158 ( \9501 , \9500 );
or \U$9159 ( \9502 , \9470 , \9501 );
nand \U$9160 ( \9503 , \9496 , \9485 );
nand \U$9161 ( \9504 , \9502 , \9503 );
xnor \U$9162 ( \9505 , \9459 , \9504 );
not \U$9163 ( \9506 , \9505 );
not \U$9164 ( \9507 , \9506 );
not \U$9165 ( \9508 , \8829 );
not \U$9166 ( \9509 , \9508 );
not \U$9167 ( \9510 , \8759 );
and \U$9168 ( \9511 , \9509 , \9510 );
and \U$9169 ( \9512 , \9508 , \8759 );
nor \U$9170 ( \9513 , \9511 , \9512 );
not \U$9171 ( \9514 , \9376 );
not \U$9172 ( \9515 , \786 );
and \U$9173 ( \9516 , \9514 , \9515 );
not \U$9174 ( \9517 , RI98719b0_131);
not \U$9175 ( \9518 , \5775 );
or \U$9176 ( \9519 , \9517 , \9518 );
or \U$9177 ( \9520 , \5776 , RI98719b0_131);
nand \U$9178 ( \9521 , \9519 , \9520 );
and \U$9179 ( \9522 , \9521 , \793 );
nor \U$9180 ( \9523 , \9516 , \9522 );
not \U$9181 ( \9524 , \9523 );
buf \U$9182 ( \9525 , \8741 );
buf \U$9183 ( \9526 , \9525 );
buf \U$9184 ( \9527 , \9526 );
not \U$9185 ( \9528 , \9527 );
not \U$9186 ( \9529 , RI9872f40_177);
not \U$9187 ( \9530 , \9529 );
not \U$9188 ( \9531 , \1393 );
or \U$9189 ( \9532 , \9530 , \9531 );
or \U$9190 ( \9533 , \2982 , \8732 );
nand \U$9191 ( \9534 , \9532 , \9533 );
not \U$9192 ( \9535 , \9534 );
or \U$9193 ( \9536 , \9528 , \9535 );
nand \U$9194 ( \9537 , \8748 , \8752 );
nand \U$9195 ( \9538 , \9536 , \9537 );
xor \U$9196 ( \9539 , \9524 , \9538 );
not \U$9197 ( \9540 , \2071 );
and \U$9198 ( \9541 , \9367 , RI9871aa0_133);
not \U$9199 ( \9542 , \9367 );
and \U$9200 ( \9543 , \9542 , \2080 );
nor \U$9201 ( \9544 , \9541 , \9543 );
not \U$9202 ( \9545 , \9544 );
or \U$9203 ( \9546 , \9540 , \9545 );
nand \U$9204 ( \9547 , \9449 , \2085 );
nand \U$9205 ( \9548 , \9546 , \9547 );
and \U$9206 ( \9549 , \9539 , \9548 );
and \U$9207 ( \9550 , \9524 , \9538 );
nor \U$9208 ( \9551 , \9549 , \9550 );
not \U$9209 ( \9552 , \9551 );
not \U$9210 ( \9553 , \9552 );
not \U$9211 ( \9554 , \1083 );
not \U$9212 ( \9555 , RI98718c0_129);
not \U$9213 ( \9556 , \6303 );
not \U$9214 ( \9557 , \9556 );
or \U$9215 ( \9558 , \9555 , \9557 );
or \U$9216 ( \9559 , \8895 , RI98718c0_129);
nand \U$9217 ( \9560 , \9558 , \9559 );
not \U$9218 ( \9561 , \9560 );
or \U$9219 ( \9562 , \9554 , \9561 );
nand \U$9220 ( \9563 , \9388 , \6673 );
nand \U$9221 ( \9564 , \9562 , \9563 );
not \U$9222 ( \9565 , \9564 );
not \U$9223 ( \9566 , \1292 );
and \U$9224 ( \9567 , RI9871b18_134, \7466 );
not \U$9225 ( \9568 , RI9871b18_134);
not \U$9226 ( \9569 , \7465 );
buf \U$9227 ( \9570 , \9569 );
and \U$9228 ( \9571 , \9568 , \9570 );
or \U$9229 ( \9572 , \9567 , \9571 );
not \U$9230 ( \9573 , \9572 );
or \U$9231 ( \9574 , \9566 , \9573 );
nand \U$9232 ( \9575 , \8950 , \1323 );
nand \U$9233 ( \9576 , \9574 , \9575 );
not \U$9234 ( \9577 , \9576 );
not \U$9235 ( \9578 , \9577 );
not \U$9236 ( \9579 , \1455 );
not \U$9237 ( \9580 , \1850 );
not \U$9238 ( \9581 , \7905 );
or \U$9239 ( \9582 , \9580 , \9581 );
or \U$9240 ( \9583 , \8934 , \1850 );
nand \U$9241 ( \9584 , \9582 , \9583 );
not \U$9242 ( \9585 , \9584 );
or \U$9243 ( \9586 , \9579 , \9585 );
nand \U$9244 ( \9587 , \8908 , \1430 );
nand \U$9245 ( \9588 , \9586 , \9587 );
not \U$9246 ( \9589 , \9588 );
or \U$9247 ( \9590 , \9578 , \9589 );
or \U$9248 ( \9591 , \9588 , \9577 );
nand \U$9249 ( \9592 , \9590 , \9591 );
not \U$9250 ( \9593 , \9592 );
or \U$9251 ( \9594 , \9565 , \9593 );
nand \U$9252 ( \9595 , \9588 , \9576 );
nand \U$9253 ( \9596 , \9594 , \9595 );
not \U$9254 ( \9597 , \1501 );
buf \U$9255 ( \9598 , \8072 );
not \U$9256 ( \9599 , \9598 );
xnor \U$9257 ( \9600 , RI9871c80_137, \9599 );
not \U$9258 ( \9601 , \9600 );
or \U$9259 ( \9602 , \9597 , \9601 );
nand \U$9260 ( \9603 , \8918 , \1518 );
nand \U$9261 ( \9604 , \9602 , \9603 );
not \U$9262 ( \9605 , \9604 );
not \U$9263 ( \9606 , \832 );
not \U$9264 ( \9607 , \8861 );
or \U$9265 ( \9608 , \9606 , \9607 );
not \U$9266 ( \9609 , RI9871d70_139);
not \U$9267 ( \9610 , \8650 );
or \U$9268 ( \9611 , \9609 , \9610 );
or \U$9269 ( \9612 , \8650 , RI9871d70_139);
nand \U$9270 ( \9613 , \9611 , \9612 );
nand \U$9271 ( \9614 , \9613 , \859 );
nand \U$9272 ( \9615 , \9608 , \9614 );
not \U$9273 ( \9616 , \9615 );
not \U$9274 ( \9617 , \876 );
not \U$9275 ( \9618 , \919 );
not \U$9276 ( \9619 , \8597 );
or \U$9277 ( \9620 , \9618 , \9619 );
nand \U$9278 ( \9621 , \8607 , RI9872130_147);
nand \U$9279 ( \9622 , \9620 , \9621 );
not \U$9280 ( \9623 , \9622 );
or \U$9281 ( \9624 , \9617 , \9623 );
nand \U$9282 ( \9625 , \8880 , \924 );
nand \U$9283 ( \9626 , \9624 , \9625 );
not \U$9284 ( \9627 , \9626 );
not \U$9285 ( \9628 , \9627 );
or \U$9286 ( \9629 , \9616 , \9628 );
or \U$9287 ( \9630 , \9615 , \9627 );
nand \U$9288 ( \9631 , \9629 , \9630 );
not \U$9289 ( \9632 , \9631 );
or \U$9290 ( \9633 , \9605 , \9632 );
nand \U$9291 ( \9634 , \9626 , \9615 );
nand \U$9292 ( \9635 , \9633 , \9634 );
and \U$9293 ( \9636 , \9596 , \9635 );
not \U$9294 ( \9637 , \9596 );
not \U$9295 ( \9638 , \9635 );
and \U$9296 ( \9639 , \9637 , \9638 );
nor \U$9297 ( \9640 , \9636 , \9639 );
not \U$9298 ( \9641 , \9640 );
or \U$9299 ( \9642 , \9553 , \9641 );
nand \U$9300 ( \9643 , \9596 , \9635 );
nand \U$9301 ( \9644 , \9642 , \9643 );
xnor \U$9302 ( \9645 , \9513 , \9644 );
not \U$9303 ( \9646 , \9645 );
or \U$9304 ( \9647 , \9507 , \9646 );
not \U$9305 ( \9648 , \9513 );
nand \U$9306 ( \9649 , \9648 , \9644 );
nand \U$9307 ( \9650 , \9647 , \9649 );
not \U$9308 ( \9651 , \9650 );
and \U$9309 ( \9652 , \9363 , \9651 );
not \U$9310 ( \9653 , \9363 );
and \U$9311 ( \9654 , \9653 , \9650 );
nor \U$9312 ( \9655 , \9652 , \9654 );
not \U$9313 ( \9656 , \9655 );
not \U$9314 ( \9657 , \9505 );
not \U$9315 ( \9658 , \9645 );
and \U$9316 ( \9659 , \9657 , \9658 );
and \U$9317 ( \9660 , \9505 , \9645 );
nor \U$9318 ( \9661 , \9659 , \9660 );
not \U$9319 ( \9662 , \9661 );
not \U$9320 ( \9663 , \9662 );
and \U$9321 ( \9664 , RI9872bf8_170, \1447 );
not \U$9322 ( \9665 , RI9872bf8_170);
and \U$9323 ( \9666 , \9665 , \6165 );
or \U$9324 ( \9667 , \9664 , \9666 );
buf \U$9325 ( \9668 , \9226 );
and \U$9326 ( \9669 , \9667 , \9668 );
buf \U$9327 ( \9670 , \9249 );
and \U$9328 ( \9671 , \9234 , \9670 );
nor \U$9329 ( \9672 , \9669 , \9671 );
not \U$9330 ( \9673 , \9672 );
not \U$9331 ( \9674 , \9673 );
not \U$9332 ( \9675 , \5653 );
and \U$9333 ( \9676 , \4454 , RI9872568_156);
not \U$9334 ( \9677 , \4454 );
and \U$9335 ( \9678 , \9677 , \5648 );
nor \U$9336 ( \9679 , \9676 , \9678 );
not \U$9337 ( \9680 , \9679 );
or \U$9338 ( \9681 , \9675 , \9680 );
nand \U$9339 ( \9682 , \9331 , \5642 );
nand \U$9340 ( \9683 , \9681 , \9682 );
not \U$9341 ( \9684 , \9683 );
not \U$9342 ( \9685 , \9684 );
buf \U$9343 ( \9686 , \9293 );
not \U$9344 ( \9687 , \9686 );
not \U$9345 ( \9688 , \9280 );
or \U$9346 ( \9689 , \9687 , \9688 );
not \U$9347 ( \9690 , RI9872e50_175);
not \U$9348 ( \9691 , \9690 );
not \U$9349 ( \9692 , \2982 );
or \U$9350 ( \9693 , \9691 , \9692 );
not \U$9351 ( \9694 , RI9872e50_175);
or \U$9352 ( \9695 , \1394 , \9694 );
nand \U$9353 ( \9696 , \9693 , \9695 );
nand \U$9354 ( \9697 , \9696 , \9273 );
nand \U$9355 ( \9698 , \9689 , \9697 );
not \U$9356 ( \9699 , \9698 );
or \U$9357 ( \9700 , \9685 , \9699 );
or \U$9358 ( \9701 , \9698 , \9684 );
nand \U$9359 ( \9702 , \9700 , \9701 );
not \U$9360 ( \9703 , \9702 );
or \U$9361 ( \9704 , \9674 , \9703 );
not \U$9362 ( \9705 , \9684 );
nand \U$9363 ( \9706 , \9705 , \9698 );
nand \U$9364 ( \9707 , \9704 , \9706 );
xor \U$9365 ( \9708 , \9010 , \9020 );
xor \U$9366 ( \9709 , \9708 , \9026 );
not \U$9367 ( \9710 , \5036 );
not \U$9368 ( \9711 , \5025 );
not \U$9369 ( \9712 , \9323 );
not \U$9370 ( \9713 , \9712 );
or \U$9371 ( \9714 , \9711 , \9713 );
nand \U$9372 ( \9715 , \9323 , RI9872478_154);
nand \U$9373 ( \9716 , \9714 , \9715 );
not \U$9374 ( \9717 , \9716 );
or \U$9375 ( \9718 , \9710 , \9717 );
nand \U$9376 ( \9719 , \9267 , \5034 );
nand \U$9377 ( \9720 , \9718 , \9719 );
not \U$9378 ( \9721 , \9720 );
not \U$9379 ( \9722 , \9119 );
not \U$9380 ( \9723 , \8679 );
or \U$9381 ( \9724 , \9722 , \9723 );
not \U$9382 ( \9725 , \9214 );
not \U$9383 ( \9726 , RI9872b80_169);
not \U$9384 ( \9727 , \1581 );
or \U$9385 ( \9728 , \9726 , \9727 );
or \U$9386 ( \9729 , \1581 , RI9872b80_169);
nand \U$9387 ( \9730 , \9728 , \9729 );
not \U$9388 ( \9731 , \9730 );
or \U$9389 ( \9732 , \9725 , \9731 );
nand \U$9390 ( \9733 , \9213 , \9196 );
nand \U$9391 ( \9734 , \9732 , \9733 );
and \U$9392 ( \9735 , \9724 , \9734 );
not \U$9393 ( \9736 , \9724 );
not \U$9394 ( \9737 , \9734 );
and \U$9395 ( \9738 , \9736 , \9737 );
nor \U$9396 ( \9739 , \9735 , \9738 );
not \U$9397 ( \9740 , \9739 );
or \U$9398 ( \9741 , \9721 , \9740 );
nand \U$9399 ( \9742 , \9734 , \9724 );
nand \U$9400 ( \9743 , \9741 , \9742 );
xor \U$9401 ( \9744 , \9709 , \9743 );
xor \U$9402 ( \9745 , \9707 , \9744 );
xor \U$9403 ( \9746 , \9469 , \9486 );
xnor \U$9404 ( \9747 , \9746 , \9496 );
not \U$9405 ( \9748 , \1018 );
not \U$9406 ( \9749 , \8086 );
buf \U$9407 ( \9750 , \8694 );
not \U$9408 ( \9751 , \9750 );
or \U$9409 ( \9752 , \9749 , \9751 );
or \U$9410 ( \9753 , \9750 , \8086 );
nand \U$9411 ( \9754 , \9752 , \9753 );
not \U$9412 ( \9755 , \9754 );
or \U$9413 ( \9756 , \9748 , \9755 );
nand \U$9414 ( \9757 , \8727 , \1013 );
nand \U$9415 ( \9758 , \9756 , \9757 );
not \U$9416 ( \9759 , \1381 );
not \U$9417 ( \9760 , \8554 );
not \U$9418 ( \9761 , \9760 );
and \U$9419 ( \9762 , RI9871e60_141, \9761 );
not \U$9420 ( \9763 , RI9871e60_141);
not \U$9421 ( \9764 , \8555 );
and \U$9422 ( \9765 , \9763 , \9764 );
or \U$9423 ( \9766 , \9762 , \9765 );
not \U$9424 ( \9767 , \9766 );
or \U$9425 ( \9768 , \9759 , \9767 );
nand \U$9426 ( \9769 , \8847 , \1352 );
nand \U$9427 ( \9770 , \9768 , \9769 );
nor \U$9428 ( \9771 , \9758 , \9770 );
not \U$9429 ( \9772 , \9771 );
not \U$9430 ( \9773 , \9772 );
not \U$9431 ( \9774 , \7338 );
not \U$9432 ( \9775 , \9483 );
or \U$9433 ( \9776 , \9774 , \9775 );
xnor \U$9434 ( \9777 , \1253 , RI98729a0_165);
nand \U$9435 ( \9778 , \9777 , \7325 );
nand \U$9436 ( \9779 , \9776 , \9778 );
not \U$9437 ( \9780 , \9779 );
or \U$9438 ( \9781 , \9773 , \9780 );
nand \U$9439 ( \9782 , \9770 , \9758 );
nand \U$9440 ( \9783 , \9781 , \9782 );
not \U$9441 ( \9784 , \8887 );
not \U$9442 ( \9785 , \8849 );
not \U$9443 ( \9786 , \9785 );
and \U$9444 ( \9787 , \9784 , \9786 );
and \U$9445 ( \9788 , \8887 , \9785 );
nor \U$9446 ( \9789 , \9787 , \9788 );
xnor \U$9447 ( \9790 , \9783 , \9789 );
and \U$9448 ( \9791 , \9747 , \9790 );
not \U$9449 ( \9792 , \9747 );
not \U$9450 ( \9793 , \9790 );
and \U$9451 ( \9794 , \9792 , \9793 );
nor \U$9452 ( \9795 , \9791 , \9794 );
and \U$9453 ( \9796 , \9631 , \9604 );
not \U$9454 ( \9797 , \9631 );
not \U$9455 ( \9798 , \9604 );
and \U$9456 ( \9799 , \9797 , \9798 );
nor \U$9457 ( \9800 , \9796 , \9799 );
not \U$9458 ( \9801 , \9782 );
nor \U$9459 ( \9802 , \9801 , \9771 );
not \U$9460 ( \9803 , \9802 );
not \U$9461 ( \9804 , \9779 );
and \U$9462 ( \9805 , \9803 , \9804 );
and \U$9463 ( \9806 , \9779 , \9802 );
nor \U$9464 ( \9807 , \9805 , \9806 );
xor \U$9465 ( \9808 , \9800 , \9807 );
not \U$9466 ( \9809 , \9216 );
not \U$9467 ( \9810 , \9182 );
not \U$9468 ( \9811 , \9170 );
and \U$9469 ( \9812 , \9810 , \9811 );
and \U$9470 ( \9813 , \9182 , \9170 );
nor \U$9471 ( \9814 , \9812 , \9813 );
not \U$9472 ( \9815 , \9814 );
or \U$9473 ( \9816 , \9809 , \9815 );
or \U$9474 ( \9817 , \9814 , \9216 );
nand \U$9475 ( \9818 , \9816 , \9817 );
and \U$9476 ( \9819 , \9808 , \9818 );
and \U$9477 ( \9820 , \9800 , \9807 );
or \U$9478 ( \9821 , \9819 , \9820 );
not \U$9479 ( \9822 , \9821 );
not \U$9480 ( \9823 , \9822 );
not \U$9481 ( \9824 , \2087 );
not \U$9482 ( \9825 , \9544 );
or \U$9483 ( \9826 , \9824 , \9825 );
xnor \U$9484 ( \9827 , \4985 , RI9871aa0_133);
nand \U$9485 ( \9828 , \9827 , \2072 );
nand \U$9486 ( \9829 , \9826 , \9828 );
not \U$9487 ( \9830 , \9829 );
not \U$9488 ( \9831 , \7325 );
and \U$9489 ( \9832 , RI98729a0_165, \1340 );
not \U$9490 ( \9833 , RI98729a0_165);
not \U$9491 ( \9834 , \1340 );
and \U$9492 ( \9835 , \9833 , \9834 );
or \U$9493 ( \9836 , \9832 , \9835 );
not \U$9494 ( \9837 , \9836 );
or \U$9495 ( \9838 , \9831 , \9837 );
nand \U$9496 ( \9839 , \9777 , \7338 );
nand \U$9497 ( \9840 , \9838 , \9839 );
not \U$9498 ( \9841 , \1013 );
not \U$9499 ( \9842 , \9754 );
or \U$9500 ( \9843 , \9841 , \9842 );
and \U$9501 ( \9844 , \8682 , \8702 );
not \U$9502 ( \9845 , \8682 );
and \U$9503 ( \9846 , \9845 , \8705 );
nor \U$9504 ( \9847 , \9844 , \9846 );
not \U$9505 ( \9848 , \9847 );
not \U$9506 ( \9849 , \9848 );
buf \U$9507 ( \9850 , \9849 );
and \U$9508 ( \9851 , \1043 , \9850 );
not \U$9509 ( \9852 , \1043 );
and \U$9510 ( \9853 , \9852 , \8708 );
nor \U$9511 ( \9854 , \9851 , \9853 );
nand \U$9512 ( \9855 , \9854 , \1018 );
nand \U$9513 ( \9856 , \9843 , \9855 );
or \U$9514 ( \9857 , \9840 , \9856 );
not \U$9515 ( \9858 , \9857 );
or \U$9516 ( \9859 , \9830 , \9858 );
nand \U$9517 ( \9860 , \9840 , \9856 );
nand \U$9518 ( \9861 , \9859 , \9860 );
not \U$9519 ( \9862 , \9861 );
not \U$9520 ( \9863 , \1518 );
not \U$9521 ( \9864 , \9600 );
or \U$9522 ( \9865 , \9863 , \9864 );
not \U$9523 ( \9866 , RI9871c80_137);
not \U$9524 ( \9867 , \8874 );
or \U$9525 ( \9868 , \9866 , \9867 );
not \U$9526 ( \9869 , \8620 );
nand \U$9527 ( \9870 , \9869 , \1800 );
nand \U$9528 ( \9871 , \9868 , \9870 );
nand \U$9529 ( \9872 , \9871 , \1501 );
nand \U$9530 ( \9873 , \9865 , \9872 );
not \U$9531 ( \9874 , \9873 );
not \U$9532 ( \9875 , \9874 );
buf \U$9533 ( \9876 , \924 );
not \U$9534 ( \9877 , \9876 );
not \U$9535 ( \9878 , \9622 );
or \U$9536 ( \9879 , \9877 , \9878 );
buf \U$9537 ( \9880 , \8666 );
not \U$9538 ( \9881 , \9880 );
not \U$9539 ( \9882 , \9881 );
and \U$9540 ( \9883 , RI9872130_147, \9882 );
not \U$9541 ( \9884 , RI9872130_147);
not \U$9542 ( \9885 , \8857 );
and \U$9543 ( \9886 , \9884 , \9885 );
or \U$9544 ( \9887 , \9883 , \9886 );
nand \U$9545 ( \9888 , \9887 , \6431 );
nand \U$9546 ( \9889 , \9879 , \9888 );
not \U$9547 ( \9890 , \9889 );
not \U$9548 ( \9891 , \9890 );
or \U$9549 ( \9892 , \9875 , \9891 );
not \U$9550 ( \9893 , \1292 );
not \U$9551 ( \9894 , RI9871b18_134);
buf \U$9552 ( \9895 , \8915 );
not \U$9553 ( \9896 , \9895 );
or \U$9554 ( \9897 , \9894 , \9896 );
not \U$9555 ( \9898 , \8333 );
nand \U$9556 ( \9899 , \9898 , \1283 );
nand \U$9557 ( \9900 , \9897 , \9899 );
not \U$9558 ( \9901 , \9900 );
or \U$9559 ( \9902 , \9893 , \9901 );
nand \U$9560 ( \9903 , \9572 , \1323 );
nand \U$9561 ( \9904 , \9902 , \9903 );
nand \U$9562 ( \9905 , \9892 , \9904 );
nand \U$9563 ( \9906 , \9889 , \9873 );
nand \U$9564 ( \9907 , \9905 , \9906 );
not \U$9565 ( \9908 , \832 );
not \U$9566 ( \9909 , \9613 );
or \U$9567 ( \9910 , \9908 , \9909 );
not \U$9568 ( \9911 , \8574 );
and \U$9569 ( \9912 , RI9871d70_139, \9911 );
not \U$9570 ( \9913 , RI9871d70_139);
and \U$9571 ( \9914 , \9913 , \8575 );
or \U$9572 ( \9915 , \9912 , \9914 );
nand \U$9573 ( \9916 , \9915 , \859 );
nand \U$9574 ( \9917 , \9910 , \9916 );
not \U$9575 ( \9918 , \9917 );
not \U$9576 ( \9919 , \1352 );
not \U$9577 ( \9920 , \9766 );
or \U$9578 ( \9921 , \9919 , \9920 );
not \U$9579 ( \9922 , \1379 );
not \U$9580 ( \9923 , \9922 );
not \U$9581 ( \9924 , \8722 );
and \U$9582 ( \9925 , RI9871e60_141, \9924 );
not \U$9583 ( \9926 , RI9871e60_141);
and \U$9584 ( \9927 , \9926 , \8722 );
or \U$9585 ( \9928 , \9925 , \9927 );
nand \U$9586 ( \9929 , \9923 , \9928 );
nand \U$9587 ( \9930 , \9921 , \9929 );
not \U$9588 ( \9931 , \9930 );
nand \U$9589 ( \9932 , \9918 , \9931 );
not \U$9590 ( \9933 , \9932 );
not \U$9591 ( \9934 , RI9873030_179);
nor \U$9592 ( \9935 , RI98730a8_180, RI9873120_181);
nor \U$9593 ( \9936 , \9421 , \9935 );
buf \U$9594 ( \9937 , \9936 );
not \U$9595 ( \9938 , \9937 );
or \U$9596 ( \9939 , \9934 , \9938 );
not \U$9597 ( \9940 , \779 );
not \U$9598 ( \9941 , RI9873030_179);
and \U$9599 ( \9942 , \9940 , \9941 );
and \U$9600 ( \9943 , \2360 , RI9873030_179);
nor \U$9601 ( \9944 , \9942 , \9943 );
not \U$9602 ( \9945 , \9944 );
not \U$9603 ( \9946 , RI9873030_179);
not \U$9604 ( \9947 , RI9873120_181);
and \U$9605 ( \9948 , \9946 , \9947 );
and \U$9606 ( \9949 , RI9873030_179, RI9873120_181);
nor \U$9607 ( \9950 , \9948 , \9949 , \9936 );
buf \U$9608 ( \9951 , \9950 );
buf \U$9609 ( \9952 , \9951 );
nand \U$9610 ( \9953 , \9945 , \9952 );
nand \U$9611 ( \9954 , \9939 , \9953 );
not \U$9612 ( \9955 , \9954 );
or \U$9613 ( \9956 , \9933 , \9955 );
nand \U$9614 ( \9957 , \9917 , \9930 );
nand \U$9615 ( \9958 , \9956 , \9957 );
xor \U$9616 ( \9959 , \9907 , \9958 );
not \U$9617 ( \9960 , \9959 );
or \U$9618 ( \9961 , \9862 , \9960 );
nand \U$9619 ( \9962 , \9958 , \9907 );
nand \U$9620 ( \9963 , \9961 , \9962 );
not \U$9621 ( \9964 , \9963 );
and \U$9622 ( \9965 , \9823 , \9964 );
and \U$9623 ( \9966 , \9963 , \9822 );
nor \U$9624 ( \9967 , \9965 , \9966 );
not \U$9625 ( \9968 , \9967 );
and \U$9626 ( \9969 , \9795 , \9968 );
not \U$9627 ( \9970 , \9963 );
nor \U$9628 ( \9971 , \9970 , \9822 );
nor \U$9629 ( \9972 , \9969 , \9971 );
not \U$9630 ( \9973 , \9972 );
xor \U$9631 ( \9974 , \9745 , \9973 );
xnor \U$9632 ( \9975 , \9672 , \9702 );
not \U$9633 ( \9976 , \9975 );
and \U$9634 ( \9977 , \8825 , \8774 );
not \U$9635 ( \9978 , \8825 );
not \U$9636 ( \9979 , \8774 );
and \U$9637 ( \9980 , \9978 , \9979 );
nor \U$9638 ( \9981 , \9977 , \9980 );
not \U$9639 ( \9982 , \9981 );
not \U$9640 ( \9983 , \9739 );
not \U$9641 ( \9984 , \9720 );
not \U$9642 ( \9985 , \9984 );
and \U$9643 ( \9986 , \9983 , \9985 );
and \U$9644 ( \9987 , \9739 , \9984 );
nor \U$9645 ( \9988 , \9986 , \9987 );
not \U$9646 ( \9989 , \9988 );
or \U$9647 ( \9990 , \9982 , \9989 );
or \U$9648 ( \9991 , \9988 , \9981 );
nand \U$9649 ( \9992 , \9990 , \9991 );
not \U$9650 ( \9993 , \9992 );
or \U$9651 ( \9994 , \9976 , \9993 );
not \U$9652 ( \9995 , \9988 );
nand \U$9653 ( \9996 , \9995 , \9981 );
nand \U$9654 ( \9997 , \9994 , \9996 );
not \U$9655 ( \9998 , \9747 );
not \U$9656 ( \9999 , \9790 );
or \U$9657 ( \10000 , \9998 , \9999 );
not \U$9658 ( \10001 , \9789 );
nand \U$9659 ( \10002 , \10001 , \9783 );
nand \U$9660 ( \10003 , \10000 , \10002 );
xor \U$9661 ( \10004 , \9997 , \10003 );
not \U$9662 ( \10005 , \10004 );
xnor \U$9663 ( \10006 , \9974 , \10005 );
not \U$9664 ( \10007 , \10006 );
or \U$9665 ( \10008 , \9663 , \10007 );
and \U$9666 ( \10009 , \9745 , \10005 );
not \U$9667 ( \10010 , \9745 );
and \U$9668 ( \10011 , \10010 , \10004 );
or \U$9669 ( \10012 , \10009 , \10011 );
nand \U$9670 ( \10013 , \10012 , \9973 );
nand \U$9671 ( \10014 , \10008 , \10013 );
xor \U$9672 ( \10015 , \9656 , \10014 );
not \U$9673 ( \10016 , \9745 );
not \U$9674 ( \10017 , \10004 );
or \U$9675 ( \10018 , \10016 , \10017 );
nand \U$9676 ( \10019 , \9997 , \10003 );
nand \U$9677 ( \10020 , \10018 , \10019 );
xor \U$9678 ( \10021 , \9390 , \9379 );
xor \U$9679 ( \10022 , \10021 , \9399 );
not \U$9680 ( \10023 , \10022 );
not \U$9681 ( \10024 , \9425 );
and \U$9682 ( \10025 , \9432 , \10024 );
not \U$9683 ( \10026 , \9432 );
and \U$9684 ( \10027 , \10026 , \9425 );
nor \U$9685 ( \10028 , \10025 , \10027 );
not \U$9686 ( \10029 , \3170 );
not \U$9687 ( \10030 , \9411 );
or \U$9688 ( \10031 , \10029 , \10030 );
and \U$9689 ( \10032 , \5614 , \3154 );
not \U$9690 ( \10033 , \5614 );
and \U$9691 ( \10034 , \10033 , RI9872310_151);
nor \U$9692 ( \10035 , \10032 , \10034 );
nand \U$9693 ( \10036 , \10035 , \6653 );
nand \U$9694 ( \10037 , \10031 , \10036 );
not \U$9695 ( \10038 , \10037 );
xor \U$9696 ( \10039 , \10028 , \10038 );
not \U$9697 ( \10040 , \10039 );
not \U$9698 ( \10041 , \1430 );
not \U$9699 ( \10042 , \9584 );
or \U$9700 ( \10043 , \10041 , \10042 );
and \U$9701 ( \10044 , RI9871c08_136, \8081 );
not \U$9702 ( \10045 , RI9871c08_136);
and \U$9703 ( \10046 , \10045 , \7004 );
or \U$9704 ( \10047 , \10044 , \10046 );
nand \U$9705 ( \10048 , \10047 , \1455 );
nand \U$9706 ( \10049 , \10043 , \10048 );
not \U$9707 ( \10050 , \10049 );
not \U$9708 ( \10051 , \9084 );
not \U$9709 ( \10052 , \9097 );
or \U$9710 ( \10053 , \10051 , \10052 );
nand \U$9711 ( \10054 , RI986ff70_75, RI986ffe8_76);
buf \U$9712 ( \10055 , \10054 );
nand \U$9713 ( \10056 , \10053 , \10055 );
not \U$9714 ( \10057 , \10056 );
nand \U$9715 ( \10058 , \9082 , \603 );
not \U$9716 ( \10059 , \10058 );
and \U$9717 ( \10060 , \10057 , \10059 );
and \U$9718 ( \10061 , \10056 , \10058 );
nor \U$9719 ( \10062 , \10060 , \10061 );
buf \U$9720 ( \10063 , \10062 );
buf \U$9721 ( \10064 , \10063 );
or \U$9722 ( \10065 , \10064 , \9723 );
not \U$9723 ( \10066 , \10065 );
not \U$9724 ( \10067 , \6672 );
not \U$9725 ( \10068 , \9560 );
or \U$9726 ( \10069 , \10067 , \10068 );
not \U$9727 ( \10070 , RI98718c0_129);
not \U$9728 ( \10071 , \8053 );
or \U$9729 ( \10072 , \10070 , \10071 );
or \U$9730 ( \10073 , \8904 , RI98718c0_129);
nand \U$9731 ( \10074 , \10072 , \10073 );
nand \U$9732 ( \10075 , \10074 , \1083 );
nand \U$9733 ( \10076 , \10069 , \10075 );
not \U$9734 ( \10077 , \10076 );
or \U$9735 ( \10078 , \10066 , \10077 );
or \U$9736 ( \10079 , \10076 , \10065 );
nand \U$9737 ( \10080 , \10078 , \10079 );
not \U$9738 ( \10081 , \10080 );
or \U$9739 ( \10082 , \10050 , \10081 );
not \U$9740 ( \10083 , \10065 );
nand \U$9741 ( \10084 , \10083 , \10076 );
nand \U$9742 ( \10085 , \10082 , \10084 );
not \U$9743 ( \10086 , \10085 );
or \U$9744 ( \10087 , \10040 , \10086 );
not \U$9745 ( \10088 , \10028 );
nand \U$9746 ( \10089 , \10088 , \10037 );
nand \U$9747 ( \10090 , \10087 , \10089 );
xor \U$9748 ( \10091 , \9435 , \9451 );
xnor \U$9749 ( \10092 , \10091 , \9419 );
xor \U$9750 ( \10093 , \10090 , \10092 );
not \U$9751 ( \10094 , \10093 );
or \U$9752 ( \10095 , \10023 , \10094 );
nand \U$9753 ( \10096 , \10090 , \10092 );
nand \U$9754 ( \10097 , \10095 , \10096 );
not \U$9755 ( \10098 , \6316 );
not \U$9756 ( \10099 , \8723 );
xor \U$9757 ( \10100 , \8679 , \10099 );
not \U$9758 ( \10101 , \10100 );
or \U$9759 ( \10102 , \10098 , \10101 );
nand \U$9760 ( \10103 , \8698 , \1162 );
nand \U$9761 ( \10104 , \10102 , \10103 );
not \U$9762 ( \10105 , \793 );
not \U$9763 ( \10106 , \9369 );
or \U$9764 ( \10107 , \10105 , \10106 );
and \U$9765 ( \10108 , \4471 , \7075 );
not \U$9766 ( \10109 , \4471 );
and \U$9767 ( \10110 , \10109 , RI98719b0_131);
nor \U$9768 ( \10111 , \10108 , \10110 );
nand \U$9769 ( \10112 , \10111 , \796 );
nand \U$9770 ( \10113 , \10107 , \10112 );
xor \U$9771 ( \10114 , \10104 , \10113 );
not \U$9772 ( \10115 , \6286 );
not \U$9773 ( \10116 , \5632 );
not \U$9774 ( \10117 , \943 );
or \U$9775 ( \10118 , \10116 , \10117 );
or \U$9776 ( \10119 , \8165 , \7049 );
nand \U$9777 ( \10120 , \10118 , \10119 );
not \U$9778 ( \10121 , \10120 );
or \U$9779 ( \10122 , \10115 , \10121 );
nand \U$9780 ( \10123 , \9397 , \6284 );
nand \U$9781 ( \10124 , \10122 , \10123 );
xnor \U$9782 ( \10125 , \10114 , \10124 );
not \U$9783 ( \10126 , \5034 );
not \U$9784 ( \10127 , \9716 );
or \U$9785 ( \10128 , \10126 , \10127 );
not \U$9786 ( \10129 , \5025 );
not \U$9787 ( \10130 , \6573 );
or \U$9788 ( \10131 , \10129 , \10130 );
not \U$9789 ( \10132 , \6573 );
not \U$9790 ( \10133 , \10132 );
or \U$9791 ( \10134 , \10133 , \5025 );
nand \U$9792 ( \10135 , \10131 , \10134 );
nand \U$9793 ( \10136 , \10135 , \5036 );
nand \U$9794 ( \10137 , \10128 , \10136 );
not \U$9795 ( \10138 , \9670 );
not \U$9796 ( \10139 , \9667 );
or \U$9797 ( \10140 , \10138 , \10139 );
not \U$9798 ( \10141 , RI9872bf8_170);
not \U$9799 ( \10142 , \1416 );
or \U$9800 ( \10143 , \10141 , \10142 );
buf \U$9801 ( \10144 , \1415 );
not \U$9802 ( \10145 , \10144 );
or \U$9803 ( \10146 , \10145 , RI9872bf8_170);
nand \U$9804 ( \10147 , \10143 , \10146 );
nand \U$9805 ( \10148 , \10147 , \9668 );
nand \U$9806 ( \10149 , \10140 , \10148 );
not \U$9807 ( \10150 , \10149 );
not \U$9808 ( \10151 , \9214 );
not \U$9809 ( \10152 , RI9872b80_169);
not \U$9810 ( \10153 , \9230 );
or \U$9811 ( \10154 , \10152 , \10153 );
or \U$9812 ( \10155 , \1320 , RI9872b80_169);
nand \U$9813 ( \10156 , \10154 , \10155 );
not \U$9814 ( \10157 , \10156 );
or \U$9815 ( \10158 , \10151 , \10157 );
nand \U$9816 ( \10159 , \9730 , \9196 );
nand \U$9817 ( \10160 , \10158 , \10159 );
not \U$9818 ( \10161 , \10160 );
not \U$9819 ( \10162 , \10161 );
or \U$9820 ( \10163 , \10150 , \10162 );
or \U$9821 ( \10164 , \10161 , \10149 );
nand \U$9822 ( \10165 , \10163 , \10164 );
xor \U$9823 ( \10166 , \10137 , \10165 );
xor \U$9824 ( \10167 , \10125 , \10166 );
not \U$9825 ( \10168 , \3164 );
not \U$9826 ( \10169 , \9417 );
or \U$9827 ( \10170 , \10168 , \10169 );
not \U$9828 ( \10171 , \3154 );
not \U$9829 ( \10172 , \3543 );
or \U$9830 ( \10173 , \10171 , \10172 );
or \U$9831 ( \10174 , \3537 , \3154 );
nand \U$9832 ( \10175 , \10173 , \10174 );
nand \U$9833 ( \10176 , \10175 , \3170 );
nand \U$9834 ( \10177 , \10170 , \10176 );
not \U$9835 ( \10178 , \10177 );
not \U$9836 ( \10179 , \2087 );
and \U$9837 ( \10180 , \4176 , \2080 );
not \U$9838 ( \10181 , \4176 );
and \U$9839 ( \10182 , \10181 , RI9871aa0_133);
nor \U$9840 ( \10183 , \10180 , \10182 );
not \U$9841 ( \10184 , \10183 );
or \U$9842 ( \10185 , \10179 , \10184 );
nand \U$9843 ( \10186 , \9442 , \2074 );
nand \U$9844 ( \10187 , \10185 , \10186 );
xor \U$9845 ( \10188 , \10178 , \10187 );
not \U$9846 ( \10189 , \7338 );
and \U$9847 ( \10190 , RI98729a0_165, \8006 );
not \U$9848 ( \10191 , RI98729a0_165);
and \U$9849 ( \10192 , \10191 , \6219 );
or \U$9850 ( \10193 , \10190 , \10192 );
not \U$9851 ( \10194 , \10193 );
or \U$9852 ( \10195 , \10189 , \10194 );
nand \U$9853 ( \10196 , \9476 , \7325 );
nand \U$9854 ( \10197 , \10195 , \10196 );
xnor \U$9855 ( \10198 , \10188 , \10197 );
xnor \U$9856 ( \10199 , \10167 , \10198 );
xor \U$9857 ( \10200 , \10097 , \10199 );
not \U$9858 ( \10201 , \6673 );
and \U$9859 ( \10202 , RI98718c0_129, \4986 );
not \U$9860 ( \10203 , RI98718c0_129);
and \U$9861 ( \10204 , \10203 , \5739 );
or \U$9862 ( \10205 , \10202 , \10204 );
not \U$9863 ( \10206 , \10205 );
or \U$9864 ( \10207 , \10201 , \10206 );
nand \U$9865 ( \10208 , \9385 , \1083 );
nand \U$9866 ( \10209 , \10207 , \10208 );
not \U$9867 ( \10210 , \5642 );
not \U$9868 ( \10211 , \9679 );
or \U$9869 ( \10212 , \10210 , \10211 );
not \U$9870 ( \10213 , RI9872568_156);
not \U$9871 ( \10214 , \1344 );
or \U$9872 ( \10215 , \10213 , \10214 );
nand \U$9873 ( \10216 , \5712 , \5644 );
nand \U$9874 ( \10217 , \10215 , \10216 );
nand \U$9875 ( \10218 , \10217 , \5653 );
nand \U$9876 ( \10219 , \10212 , \10218 );
xor \U$9877 ( \10220 , \10209 , \10219 );
not \U$9878 ( \10221 , \9686 );
not \U$9879 ( \10222 , \9696 );
or \U$9880 ( \10223 , \10221 , \10222 );
not \U$9881 ( \10224 , \9690 );
not \U$9882 ( \10225 , \1692 );
or \U$9883 ( \10226 , \10224 , \10225 );
or \U$9884 ( \10227 , \7330 , \9694 );
nand \U$9885 ( \10228 , \10226 , \10227 );
nand \U$9886 ( \10229 , \10228 , \9273 );
nand \U$9887 ( \10230 , \10223 , \10229 );
xor \U$9888 ( \10231 , \10220 , \10230 );
not \U$9889 ( \10232 , \4085 );
and \U$9890 ( \10233 , RI98725e0_157, \1486 );
not \U$9891 ( \10234 , RI98725e0_157);
not \U$9892 ( \10235 , \3275 );
and \U$9893 ( \10236 , \10234 , \10235 );
nor \U$9894 ( \10237 , \10233 , \10236 );
not \U$9895 ( \10238 , \10237 );
or \U$9896 ( \10239 , \10232 , \10238 );
nand \U$9897 ( \10240 , \8781 , \5530 );
nand \U$9898 ( \10241 , \10239 , \10240 );
buf \U$9899 ( \10242 , \8802 );
not \U$9900 ( \10243 , \10242 );
not \U$9901 ( \10244 , RI9872d60_173);
not \U$9902 ( \10245 , \1127 );
or \U$9903 ( \10246 , \10244 , \10245 );
or \U$9904 ( \10247 , \2399 , RI9872d60_173);
nand \U$9905 ( \10248 , \10246 , \10247 );
not \U$9906 ( \10249 , \10248 );
or \U$9907 ( \10250 , \10243 , \10249 );
buf \U$9908 ( \10251 , \8818 );
nand \U$9909 ( \10252 , \8804 , \10251 );
nand \U$9910 ( \10253 , \10250 , \10252 );
xor \U$9911 ( \10254 , \10241 , \10253 );
not \U$9912 ( \10255 , \5942 );
not \U$9913 ( \10256 , \8765 );
or \U$9914 ( \10257 , \10255 , \10256 );
xnor \U$9915 ( \10258 , \6021 , RI9872388_152);
nand \U$9916 ( \10259 , \10258 , \5937 );
nand \U$9917 ( \10260 , \10257 , \10259 );
xor \U$9918 ( \10261 , \10254 , \10260 );
xor \U$9919 ( \10262 , \10231 , \10261 );
not \U$9920 ( \10263 , \3466 );
not \U$9921 ( \10264 , \9465 );
or \U$9922 ( \10265 , \10263 , \10264 );
xnor \U$9923 ( \10266 , \4287 , RI98726d0_159);
nand \U$9924 ( \10267 , \10266 , \3467 );
nand \U$9925 ( \10268 , \10265 , \10267 );
xor \U$9926 ( \10269 , \9724 , \10268 );
not \U$9927 ( \10270 , \8029 );
not \U$9928 ( \10271 , \9492 );
or \U$9929 ( \10272 , \10270 , \10271 );
not \U$9930 ( \10273 , RI9872a18_166);
not \U$9931 ( \10274 , \916 );
or \U$9932 ( \10275 , \10273 , \10274 );
or \U$9933 ( \10276 , \6585 , RI9872a18_166);
nand \U$9934 ( \10277 , \10275 , \10276 );
nand \U$9935 ( \10278 , \10277 , \8041 );
nand \U$9936 ( \10279 , \10272 , \10278 );
xnor \U$9937 ( \10280 , \10269 , \10279 );
xor \U$9938 ( \10281 , \10262 , \10280 );
and \U$9939 ( \10282 , \10200 , \10281 );
and \U$9940 ( \10283 , \10097 , \10199 );
or \U$9941 ( \10284 , \10282 , \10283 );
xor \U$9942 ( \10285 , \10020 , \10284 );
not \U$9943 ( \10286 , \10187 );
and \U$9944 ( \10287 , \10197 , \10177 );
not \U$9945 ( \10288 , \10197 );
and \U$9946 ( \10289 , \10288 , \10178 );
nor \U$9947 ( \10290 , \10287 , \10289 );
not \U$9948 ( \10291 , \10290 );
or \U$9949 ( \10292 , \10286 , \10291 );
nand \U$9950 ( \10293 , \10197 , \10177 );
nand \U$9951 ( \10294 , \10292 , \10293 );
not \U$9952 ( \10295 , \10113 );
not \U$9953 ( \10296 , \10104 );
not \U$9954 ( \10297 , \10296 );
not \U$9955 ( \10298 , \10124 );
or \U$9956 ( \10299 , \10297 , \10298 );
or \U$9957 ( \10300 , \10296 , \10124 );
nand \U$9958 ( \10301 , \10299 , \10300 );
not \U$9959 ( \10302 , \10301 );
or \U$9960 ( \10303 , \10295 , \10302 );
nand \U$9961 ( \10304 , \10124 , \10104 );
nand \U$9962 ( \10305 , \10303 , \10304 );
not \U$9963 ( \10306 , \10305 );
not \U$9964 ( \10307 , \1353 );
not \U$9965 ( \10308 , \8606 );
buf \U$9966 ( \10309 , \10308 );
and \U$9967 ( \10310 , RI9871e60_141, \10309 );
not \U$9968 ( \10311 , RI9871e60_141);
and \U$9969 ( \10312 , \10311 , \8597 );
or \U$9970 ( \10313 , \10310 , \10312 );
not \U$9971 ( \10314 , \10313 );
or \U$9972 ( \10315 , \10307 , \10314 );
nand \U$9973 ( \10316 , \8672 , \1381 );
nand \U$9974 ( \10317 , \10315 , \10316 );
not \U$9975 ( \10318 , \1067 );
and \U$9976 ( \10319 , \8642 , \3272 );
not \U$9977 ( \10320 , \8642 );
and \U$9978 ( \10321 , \10320 , \8086 );
nor \U$9979 ( \10322 , \10319 , \10321 );
not \U$9980 ( \10323 , \10322 );
or \U$9981 ( \10324 , \10318 , \10323 );
nand \U$9982 ( \10325 , \8582 , \1018 );
nand \U$9983 ( \10326 , \10324 , \10325 );
xor \U$9984 ( \10327 , \10317 , \10326 );
not \U$9985 ( \10328 , \9294 );
not \U$9986 ( \10329 , \10228 );
or \U$9987 ( \10330 , \10328 , \10329 );
buf \U$9988 ( \10331 , \9272 );
buf \U$9989 ( \10332 , \10331 );
buf \U$9990 ( \10333 , \10332 );
nand \U$9991 ( \10334 , \10333 , RI9872e50_175);
nand \U$9992 ( \10335 , \10330 , \10334 );
xnor \U$9993 ( \10336 , \10327 , \10335 );
not \U$9994 ( \10337 , \10336 );
and \U$9995 ( \10338 , \10306 , \10337 );
and \U$9996 ( \10339 , \10305 , \10336 );
nor \U$9997 ( \10340 , \10338 , \10339 );
xnor \U$9998 ( \10341 , \10294 , \10340 );
not \U$9999 ( \10342 , \9458 );
not \U$10000 ( \10343 , \9405 );
or \U$10001 ( \10344 , \10342 , \10343 );
nand \U$10002 ( \10345 , \10344 , \9504 );
nand \U$10003 ( \10346 , \9404 , \9457 );
and \U$10004 ( \10347 , \10345 , \10346 );
xor \U$10005 ( \10348 , \10341 , \10347 );
not \U$10006 ( \10349 , \10198 );
not \U$10007 ( \10350 , \10125 );
and \U$10008 ( \10351 , \10166 , \10350 );
not \U$10009 ( \10352 , \10166 );
and \U$10010 ( \10353 , \10352 , \10125 );
nor \U$10011 ( \10354 , \10351 , \10353 );
not \U$10012 ( \10355 , \10354 );
or \U$10013 ( \10356 , \10349 , \10355 );
nand \U$10014 ( \10357 , \10166 , \10350 );
nand \U$10015 ( \10358 , \10356 , \10357 );
xnor \U$10016 ( \10359 , \10348 , \10358 );
xor \U$10017 ( \10360 , \10285 , \10359 );
buf \U$10018 ( \10361 , \10360 );
and \U$10019 ( \10362 , \10015 , \10361 );
and \U$10020 ( \10363 , \9656 , \10014 );
nor \U$10021 ( \10364 , \10362 , \10363 );
not \U$10022 ( \10365 , \10364 );
and \U$10023 ( \10366 , \8679 , \8697 );
not \U$10024 ( \10367 , \1220 );
not \U$10025 ( \10368 , \5753 );
buf \U$10026 ( \10369 , \8554 );
and \U$10027 ( \10370 , \10368 , \10369 );
not \U$10028 ( \10371 , \10368 );
not \U$10029 ( \10372 , \10369 );
and \U$10030 ( \10373 , \10371 , \10372 );
nor \U$10031 ( \10374 , \10370 , \10373 );
not \U$10032 ( \10375 , \10374 );
or \U$10033 ( \10376 , \10367 , \10375 );
nand \U$10034 ( \10377 , \10100 , \1162 );
nand \U$10035 ( \10378 , \10376 , \10377 );
xor \U$10036 ( \10379 , \10366 , \10378 );
not \U$10037 ( \10380 , \5642 );
not \U$10038 ( \10381 , \10217 );
or \U$10039 ( \10382 , \10380 , \10381 );
and \U$10040 ( \10383 , \1658 , \5648 );
not \U$10041 ( \10384 , \1658 );
and \U$10042 ( \10385 , \10384 , RI9872568_156);
nor \U$10043 ( \10386 , \10383 , \10385 );
nand \U$10044 ( \10387 , \10386 , \5653 );
nand \U$10045 ( \10388 , \10382 , \10387 );
xor \U$10046 ( \10389 , \10379 , \10388 );
not \U$10047 ( \10390 , \832 );
buf \U$10048 ( \10391 , \9598 );
not \U$10049 ( \10392 , \10391 );
xnor \U$10050 ( \10393 , \10392 , RI9871d70_139);
not \U$10051 ( \10394 , \10393 );
or \U$10052 ( \10395 , \10390 , \10394 );
nand \U$10053 ( \10396 , \8626 , \859 );
nand \U$10054 ( \10397 , \10395 , \10396 );
not \U$10055 ( \10398 , \924 );
and \U$10056 ( \10399 , RI9872130_147, \8925 );
not \U$10057 ( \10400 , RI9872130_147);
not \U$10058 ( \10401 , \9570 );
and \U$10059 ( \10402 , \10400 , \10401 );
nor \U$10060 ( \10403 , \10399 , \10402 );
not \U$10061 ( \10404 , \10403 );
or \U$10062 ( \10405 , \10398 , \10404 );
nand \U$10063 ( \10406 , \9018 , \6431 );
nand \U$10064 ( \10407 , \10405 , \10406 );
xor \U$10065 ( \10408 , \10397 , \10407 );
not \U$10066 ( \10409 , \1518 );
not \U$10067 ( \10410 , \1584 );
buf \U$10068 ( \10411 , \6527 );
buf \U$10069 ( \10412 , \10411 );
not \U$10070 ( \10413 , \10412 );
or \U$10071 ( \10414 , \10410 , \10413 );
or \U$10072 ( \10415 , \6530 , \1800 );
nand \U$10073 ( \10416 , \10414 , \10415 );
not \U$10074 ( \10417 , \10416 );
or \U$10075 ( \10418 , \10409 , \10417 );
nand \U$10076 ( \10419 , \9006 , \1501 );
nand \U$10077 ( \10420 , \10418 , \10419 );
xor \U$10078 ( \10421 , \10408 , \10420 );
xor \U$10079 ( \10422 , \10389 , \10421 );
xor \U$10080 ( \10423 , \10241 , \10253 );
and \U$10081 ( \10424 , \10423 , \10260 );
and \U$10082 ( \10425 , \10241 , \10253 );
or \U$10083 ( \10426 , \10424 , \10425 );
and \U$10084 ( \10427 , \10422 , \10426 );
and \U$10085 ( \10428 , \10389 , \10421 );
or \U$10086 ( \10429 , \10427 , \10428 );
not \U$10087 ( \10430 , \10429 );
not \U$10088 ( \10431 , \10305 );
nand \U$10089 ( \10432 , \10431 , \10336 );
not \U$10090 ( \10433 , \10432 );
not \U$10091 ( \10434 , \10294 );
or \U$10092 ( \10435 , \10433 , \10434 );
not \U$10093 ( \10436 , \10336 );
nand \U$10094 ( \10437 , \10436 , \10305 );
nand \U$10095 ( \10438 , \10435 , \10437 );
not \U$10096 ( \10439 , \10438 );
not \U$10097 ( \10440 , \10439 );
or \U$10098 ( \10441 , \10430 , \10440 );
or \U$10099 ( \10442 , \10439 , \10429 );
nand \U$10100 ( \10443 , \10441 , \10442 );
not \U$10101 ( \10444 , \3170 );
and \U$10102 ( \10445 , \9461 , \3154 );
not \U$10103 ( \10446 , \9461 );
and \U$10104 ( \10447 , \10446 , RI9872310_151);
nor \U$10105 ( \10448 , \10445 , \10447 );
not \U$10106 ( \10449 , \10448 );
or \U$10107 ( \10450 , \10444 , \10449 );
nand \U$10108 ( \10451 , \10175 , \3163 );
nand \U$10109 ( \10452 , \10450 , \10451 );
not \U$10110 ( \10453 , \10452 );
not \U$10111 ( \10454 , \3467 );
and \U$10112 ( \10455 , \2111 , RI98726d0_159);
not \U$10113 ( \10456 , \2111 );
and \U$10114 ( \10457 , \10456 , \3593 );
nor \U$10115 ( \10458 , \10455 , \10457 );
not \U$10116 ( \10459 , \10458 );
or \U$10117 ( \10460 , \10454 , \10459 );
nand \U$10118 ( \10461 , \10266 , \3600 );
nand \U$10119 ( \10462 , \10460 , \10461 );
not \U$10120 ( \10463 , \7338 );
xnor \U$10121 ( \10464 , \893 , RI98729a0_165);
not \U$10122 ( \10465 , \10464 );
or \U$10123 ( \10466 , \10463 , \10465 );
nand \U$10124 ( \10467 , \10193 , \7326 );
nand \U$10125 ( \10468 , \10466 , \10467 );
xor \U$10126 ( \10469 , \10462 , \10468 );
not \U$10127 ( \10470 , \10469 );
or \U$10128 ( \10471 , \10453 , \10470 );
nand \U$10129 ( \10472 , \10468 , \10462 );
nand \U$10130 ( \10473 , \10471 , \10472 );
not \U$10131 ( \10474 , \10473 );
not \U$10132 ( \10475 , \4085 );
not \U$10133 ( \10476 , \4088 );
not \U$10134 ( \10477 , \1194 );
or \U$10135 ( \10478 , \10476 , \10477 );
or \U$10136 ( \10479 , \3969 , \4088 );
nand \U$10137 ( \10480 , \10478 , \10479 );
not \U$10138 ( \10481 , \10480 );
or \U$10139 ( \10482 , \10475 , \10481 );
nand \U$10140 ( \10483 , \10237 , \4103 );
nand \U$10141 ( \10484 , \10482 , \10483 );
not \U$10142 ( \10485 , \10484 );
not \U$10143 ( \10486 , \9668 );
not \U$10144 ( \10487 , \10486 );
not \U$10145 ( \10488 , \10487 );
not \U$10146 ( \10489 , RI9872bf8_170);
not \U$10147 ( \10490 , \1097 );
or \U$10148 ( \10491 , \10489 , \10490 );
or \U$10149 ( \10492 , \1097 , RI9872bf8_170);
nand \U$10150 ( \10493 , \10491 , \10492 );
not \U$10151 ( \10494 , \10493 );
or \U$10152 ( \10495 , \10488 , \10494 );
nand \U$10153 ( \10496 , \10147 , \9670 );
nand \U$10154 ( \10497 , \10495 , \10496 );
not \U$10155 ( \10498 , \9072 );
not \U$10156 ( \10499 , RI9872a18_166);
not \U$10157 ( \10500 , \7064 );
or \U$10158 ( \10501 , \10499 , \10500 );
or \U$10159 ( \10502 , \1834 , RI9872a18_166);
nand \U$10160 ( \10503 , \10501 , \10502 );
not \U$10161 ( \10504 , \10503 );
or \U$10162 ( \10505 , \10498 , \10504 );
nand \U$10163 ( \10506 , \10277 , \9079 );
nand \U$10164 ( \10507 , \10505 , \10506 );
xor \U$10165 ( \10508 , \10497 , \10507 );
not \U$10166 ( \10509 , \10508 );
or \U$10167 ( \10510 , \10485 , \10509 );
nand \U$10168 ( \10511 , \10507 , \10497 );
nand \U$10169 ( \10512 , \10510 , \10511 );
not \U$10170 ( \10513 , \10512 );
xor \U$10171 ( \10514 , \10317 , \10335 );
and \U$10172 ( \10515 , \10514 , \10326 );
and \U$10173 ( \10516 , \10317 , \10335 );
nor \U$10174 ( \10517 , \10515 , \10516 );
not \U$10175 ( \10518 , \10517 );
and \U$10176 ( \10519 , \10513 , \10518 );
and \U$10177 ( \10520 , \10512 , \10517 );
nor \U$10178 ( \10521 , \10519 , \10520 );
not \U$10179 ( \10522 , \10521 );
or \U$10180 ( \10523 , \10474 , \10522 );
or \U$10181 ( \10524 , \10521 , \10473 );
nand \U$10182 ( \10525 , \10523 , \10524 );
xnor \U$10183 ( \10526 , \10443 , \10525 );
xor \U$10184 ( \10527 , \8584 , \8628 );
and \U$10185 ( \10528 , \10527 , \8674 );
and \U$10186 ( \10529 , \8584 , \8628 );
or \U$10187 ( \10530 , \10528 , \10529 );
not \U$10188 ( \10531 , \10137 );
not \U$10189 ( \10532 , \10165 );
or \U$10190 ( \10533 , \10531 , \10532 );
nand \U$10191 ( \10534 , \10160 , \10149 );
nand \U$10192 ( \10535 , \10533 , \10534 );
xor \U$10193 ( \10536 , \10530 , \10535 );
not \U$10194 ( \10537 , \10268 );
not \U$10195 ( \10538 , \9724 );
not \U$10196 ( \10539 , \10279 );
or \U$10197 ( \10540 , \10538 , \10539 );
or \U$10198 ( \10541 , \10279 , \9724 );
nand \U$10199 ( \10542 , \10540 , \10541 );
not \U$10200 ( \10543 , \10542 );
or \U$10201 ( \10544 , \10537 , \10543 );
not \U$10202 ( \10545 , \9724 );
nand \U$10203 ( \10546 , \10545 , \10279 );
nand \U$10204 ( \10547 , \10544 , \10546 );
xor \U$10205 ( \10548 , \10536 , \10547 );
xor \U$10206 ( \10549 , \10231 , \10261 );
and \U$10207 ( \10550 , \10549 , \10280 );
and \U$10208 ( \10551 , \10231 , \10261 );
or \U$10209 ( \10552 , \10550 , \10551 );
or \U$10210 ( \10553 , \10548 , \10552 );
not \U$10211 ( \10554 , \10553 );
not \U$10212 ( \10555 , \9707 );
not \U$10213 ( \10556 , \9744 );
or \U$10214 ( \10557 , \10555 , \10556 );
nand \U$10215 ( \10558 , \9743 , \9709 );
nand \U$10216 ( \10559 , \10557 , \10558 );
not \U$10217 ( \10560 , \10559 );
or \U$10218 ( \10561 , \10554 , \10560 );
nand \U$10219 ( \10562 , \10548 , \10552 );
nand \U$10220 ( \10563 , \10561 , \10562 );
xor \U$10221 ( \10564 , \10526 , \10563 );
xor \U$10222 ( \10565 , \10366 , \10378 );
and \U$10223 ( \10566 , \10565 , \10388 );
and \U$10224 ( \10567 , \10366 , \10378 );
or \U$10225 ( \10568 , \10566 , \10567 );
and \U$10226 ( \10569 , \10393 , \6635 );
and \U$10227 ( \10570 , \8335 , RI9871d70_139);
not \U$10228 ( \10571 , \8335 );
and \U$10229 ( \10572 , \10571 , \2243 );
nor \U$10230 ( \10573 , \10570 , \10572 );
and \U$10231 ( \10574 , \10573 , \832 );
nor \U$10232 ( \10575 , \10569 , \10574 );
not \U$10233 ( \10576 , \10575 );
not \U$10234 ( \10577 , \876 );
not \U$10235 ( \10578 , \10403 );
or \U$10236 ( \10579 , \10577 , \10578 );
not \U$10237 ( \10580 , \919 );
not \U$10238 ( \10581 , \7001 );
not \U$10239 ( \10582 , \10581 );
buf \U$10240 ( \10583 , \10582 );
not \U$10241 ( \10584 , \10583 );
not \U$10242 ( \10585 , \10584 );
or \U$10243 ( \10586 , \10580 , \10585 );
not \U$10244 ( \10587 , \7003 );
nand \U$10245 ( \10588 , \10587 , RI9872130_147);
nand \U$10246 ( \10589 , \10586 , \10588 );
nand \U$10247 ( \10590 , \10589 , \9876 );
nand \U$10248 ( \10591 , \10579 , \10590 );
not \U$10249 ( \10592 , \10591 );
not \U$10250 ( \10593 , \1381 );
not \U$10251 ( \10594 , \10313 );
or \U$10252 ( \10595 , \10593 , \10594 );
not \U$10253 ( \10596 , \2595 );
buf \U$10254 ( \10597 , \8877 );
not \U$10255 ( \10598 , \10597 );
and \U$10256 ( \10599 , \3123 , \10598 );
not \U$10257 ( \10600 , \3123 );
not \U$10258 ( \10601 , \8620 );
and \U$10259 ( \10602 , \10600 , \10601 );
nor \U$10260 ( \10603 , \10599 , \10602 );
nand \U$10261 ( \10604 , \10596 , \10603 );
nand \U$10262 ( \10605 , \10595 , \10604 );
not \U$10263 ( \10606 , \10605 );
not \U$10264 ( \10607 , \10606 );
or \U$10265 ( \10608 , \10592 , \10607 );
or \U$10266 ( \10609 , \10591 , \10606 );
nand \U$10267 ( \10610 , \10608 , \10609 );
not \U$10268 ( \10611 , \10610 );
or \U$10269 ( \10612 , \10576 , \10611 );
or \U$10270 ( \10613 , \10610 , \10575 );
nand \U$10271 ( \10614 , \10612 , \10613 );
xor \U$10272 ( \10615 , \10568 , \10614 );
not \U$10273 ( \10616 , \10251 );
not \U$10274 ( \10617 , \10248 );
or \U$10275 ( \10618 , \10616 , \10617 );
not \U$10276 ( \10619 , \8811 );
not \U$10277 ( \10620 , \2982 );
or \U$10278 ( \10621 , \10619 , \10620 );
or \U$10279 ( \10622 , \2982 , \8811 );
nand \U$10280 ( \10623 , \10621 , \10622 );
buf \U$10281 ( \10624 , \8800 );
nand \U$10282 ( \10625 , \10623 , \10624 );
nand \U$10283 ( \10626 , \10618 , \10625 );
not \U$10284 ( \10627 , \1455 );
not \U$10285 ( \10628 , \8969 );
or \U$10286 ( \10629 , \10627 , \10628 );
and \U$10287 ( \10630 , \5776 , \1619 );
not \U$10288 ( \10631 , \5776 );
and \U$10289 ( \10632 , \10631 , RI9871c08_136);
nor \U$10290 ( \10633 , \10630 , \10632 );
nand \U$10291 ( \10634 , \10633 , \1430 );
nand \U$10292 ( \10635 , \10629 , \10634 );
xor \U$10293 ( \10636 , \10626 , \10635 );
and \U$10294 ( \10637 , RI98718c0_129, \7791 );
not \U$10295 ( \10638 , RI98718c0_129);
not \U$10296 ( \10639 , \4990 );
and \U$10297 ( \10640 , \10638 , \10639 );
or \U$10298 ( \10641 , \10637 , \10640 );
and \U$10299 ( \10642 , \10641 , \6673 );
not \U$10300 ( \10643 , \10205 );
nor \U$10301 ( \10644 , \10643 , \1688 );
nor \U$10302 ( \10645 , \10642 , \10644 );
not \U$10303 ( \10646 , \10645 );
and \U$10304 ( \10647 , \10636 , \10646 );
and \U$10305 ( \10648 , \10626 , \10635 );
or \U$10306 ( \10649 , \10647 , \10648 );
xor \U$10307 ( \10650 , \10615 , \10649 );
xor \U$10308 ( \10651 , \10635 , \10645 );
xnor \U$10309 ( \10652 , \10651 , \10626 );
not \U$10310 ( \10653 , \5036 );
xor \U$10311 ( \10654 , \3365 , RI9872478_154);
not \U$10312 ( \10655 , \10654 );
or \U$10313 ( \10656 , \10653 , \10655 );
nand \U$10314 ( \10657 , \10135 , \5034 );
nand \U$10315 ( \10658 , \10656 , \10657 );
not \U$10316 ( \10659 , \5048 );
not \U$10317 ( \10660 , \4902 );
not \U$10318 ( \10661 , \9712 );
or \U$10319 ( \10662 , \10660 , \10661 );
nand \U$10320 ( \10663 , \9323 , RI9872388_152);
nand \U$10321 ( \10664 , \10662 , \10663 );
not \U$10322 ( \10665 , \10664 );
or \U$10323 ( \10666 , \10659 , \10665 );
nand \U$10324 ( \10667 , \10258 , \5942 );
nand \U$10325 ( \10668 , \10666 , \10667 );
xor \U$10326 ( \10669 , \10658 , \10668 );
not \U$10327 ( \10670 , \9214 );
and \U$10328 ( \10671 , RI9872b80_169, \1447 );
not \U$10329 ( \10672 , RI9872b80_169);
not \U$10330 ( \10673 , \1445 );
buf \U$10331 ( \10674 , \10673 );
and \U$10332 ( \10675 , \10672 , \10674 );
or \U$10333 ( \10676 , \10671 , \10675 );
not \U$10334 ( \10677 , \10676 );
or \U$10335 ( \10678 , \10670 , \10677 );
buf \U$10336 ( \10679 , \9196 );
nand \U$10337 ( \10680 , \10156 , \10679 );
nand \U$10338 ( \10681 , \10678 , \10680 );
xor \U$10339 ( \10682 , \10669 , \10681 );
xor \U$10340 ( \10683 , \10652 , \10682 );
not \U$10341 ( \10684 , \6145 );
and \U$10342 ( \10685 , RI98719b0_131, \5206 );
not \U$10343 ( \10686 , RI98719b0_131);
and \U$10344 ( \10687 , \10686 , \5611 );
or \U$10345 ( \10688 , \10685 , \10687 );
not \U$10346 ( \10689 , \10688 );
or \U$10347 ( \10690 , \10684 , \10689 );
nand \U$10348 ( \10691 , \10111 , \793 );
nand \U$10349 ( \10692 , \10690 , \10691 );
not \U$10350 ( \10693 , \2074 );
not \U$10351 ( \10694 , \10183 );
or \U$10352 ( \10695 , \10693 , \10694 );
and \U$10353 ( \10696 , RI9871aa0_133, \3569 );
not \U$10354 ( \10697 , RI9871aa0_133);
not \U$10355 ( \10698 , \3567 );
not \U$10356 ( \10699 , \10698 );
and \U$10357 ( \10700 , \10697 , \10699 );
or \U$10358 ( \10701 , \10696 , \10700 );
not \U$10359 ( \10702 , \10701 );
nand \U$10360 ( \10703 , \10702 , \2087 );
nand \U$10361 ( \10704 , \10695 , \10703 );
xor \U$10362 ( \10705 , \10692 , \10704 );
not \U$10363 ( \10706 , \6611 );
not \U$10364 ( \10707 , RI98728b0_163);
not \U$10365 ( \10708 , \2216 );
or \U$10366 ( \10709 , \10707 , \10708 );
or \U$10367 ( \10710 , \2216 , RI98728b0_163);
nand \U$10368 ( \10711 , \10709 , \10710 );
not \U$10369 ( \10712 , \10711 );
or \U$10370 ( \10713 , \10706 , \10712 );
nand \U$10371 ( \10714 , \10120 , \6284 );
nand \U$10372 ( \10715 , \10713 , \10714 );
xor \U$10373 ( \10716 , \10705 , \10715 );
and \U$10374 ( \10717 , \10683 , \10716 );
and \U$10375 ( \10718 , \10652 , \10682 );
or \U$10376 ( \10719 , \10717 , \10718 );
xor \U$10377 ( \10720 , \10650 , \10719 );
xor \U$10378 ( \10721 , \10209 , \10219 );
and \U$10379 ( \10722 , \10721 , \10230 );
and \U$10380 ( \10723 , \10209 , \10219 );
nor \U$10381 ( \10724 , \10722 , \10723 );
not \U$10382 ( \10725 , \10724 );
xor \U$10383 ( \10726 , \10452 , \10462 );
xnor \U$10384 ( \10727 , \10726 , \10468 );
not \U$10385 ( \10728 , \10727 );
or \U$10386 ( \10729 , \10725 , \10728 );
and \U$10387 ( \10730 , \10508 , \10484 );
not \U$10388 ( \10731 , \10508 );
not \U$10389 ( \10732 , \10484 );
and \U$10390 ( \10733 , \10731 , \10732 );
nor \U$10391 ( \10734 , \10730 , \10733 );
nand \U$10392 ( \10735 , \10729 , \10734 );
not \U$10393 ( \10736 , \10724 );
not \U$10394 ( \10737 , \10727 );
nand \U$10395 ( \10738 , \10736 , \10737 );
and \U$10396 ( \10739 , \10735 , \10738 );
not \U$10397 ( \10740 , \10739 );
xnor \U$10398 ( \10741 , \10720 , \10740 );
not \U$10399 ( \10742 , \10741 );
xnor \U$10400 ( \10743 , \10564 , \10742 );
xor \U$10401 ( \10744 , \10020 , \10284 );
and \U$10402 ( \10745 , \10744 , \10359 );
and \U$10403 ( \10746 , \10020 , \10284 );
or \U$10404 ( \10747 , \10745 , \10746 );
not \U$10405 ( \10748 , \9650 );
not \U$10406 ( \10749 , \9363 );
or \U$10407 ( \10750 , \10748 , \10749 );
not \U$10408 ( \10751 , \9359 );
nand \U$10409 ( \10752 , \10751 , \9043 );
nand \U$10410 ( \10753 , \10750 , \10752 );
and \U$10411 ( \10754 , \10747 , \10753 );
not \U$10412 ( \10755 , \10747 );
not \U$10413 ( \10756 , \10753 );
and \U$10414 ( \10757 , \10755 , \10756 );
nor \U$10415 ( \10758 , \10754 , \10757 );
xor \U$10416 ( \10759 , \10743 , \10758 );
not \U$10417 ( \10760 , \10759 );
xor \U$10418 ( \10761 , \10389 , \10421 );
xor \U$10419 ( \10762 , \10761 , \10426 );
xor \U$10420 ( \10763 , \10652 , \10682 );
xor \U$10421 ( \10764 , \10763 , \10716 );
xor \U$10422 ( \10765 , \10762 , \10764 );
xor \U$10423 ( \10766 , \10734 , \10724 );
xnor \U$10424 ( \10767 , \10766 , \10737 );
and \U$10425 ( \10768 , \10765 , \10767 );
and \U$10426 ( \10769 , \10762 , \10764 );
or \U$10427 ( \10770 , \10768 , \10769 );
not \U$10428 ( \10771 , \10770 );
and \U$10429 ( \10772 , \8679 , \10099 );
not \U$10430 ( \10773 , \1162 );
not \U$10431 ( \10774 , \10374 );
or \U$10432 ( \10775 , \10773 , \10774 );
xor \U$10433 ( \10776 , \1165 , \8575 );
nand \U$10434 ( \10777 , \10776 , \6316 );
nand \U$10435 ( \10778 , \10775 , \10777 );
xor \U$10436 ( \10779 , \10772 , \10778 );
not \U$10437 ( \10780 , \1067 );
and \U$10438 ( \10781 , \8857 , \1043 );
not \U$10439 ( \10782 , \8857 );
and \U$10440 ( \10783 , \10782 , \1044 );
nor \U$10441 ( \10784 , \10781 , \10783 );
not \U$10442 ( \10785 , \10784 );
or \U$10443 ( \10786 , \10780 , \10785 );
nand \U$10444 ( \10787 , \10322 , \1018 );
nand \U$10445 ( \10788 , \10786 , \10787 );
xor \U$10446 ( \10789 , \10779 , \10788 );
not \U$10447 ( \10790 , \10789 );
not \U$10448 ( \10791 , \10790 );
not \U$10449 ( \10792 , \1292 );
not \U$10450 ( \10793 , \8984 );
or \U$10451 ( \10794 , \10792 , \10793 );
not \U$10452 ( \10795 , \7541 );
and \U$10453 ( \10796 , \10795 , RI9871b18_134);
and \U$10454 ( \10797 , \5762 , \4044 );
nor \U$10455 ( \10798 , \10796 , \10797 );
or \U$10456 ( \10799 , \10798 , \1543 );
nand \U$10457 ( \10800 , \10794 , \10799 );
not \U$10458 ( \10801 , \1501 );
not \U$10459 ( \10802 , \10416 );
or \U$10460 ( \10803 , \10801 , \10802 );
not \U$10461 ( \10804 , \1746 );
not \U$10462 ( \10805 , RI9871c80_137);
not \U$10463 ( \10806 , \8054 );
or \U$10464 ( \10807 , \10805 , \10806 );
or \U$10465 ( \10808 , \8054 , RI9871c80_137);
nand \U$10466 ( \10809 , \10807 , \10808 );
nand \U$10467 ( \10810 , \10804 , \10809 );
nand \U$10468 ( \10811 , \10803 , \10810 );
not \U$10469 ( \10812 , \10811 );
nand \U$10470 ( \10813 , RI9872ec8_176, RI9872f40_177);
and \U$10471 ( \10814 , \10813 , RI9872e50_175);
not \U$10472 ( \10815 , \10814 );
and \U$10473 ( \10816 , \10812 , \10815 );
and \U$10474 ( \10817 , \10811 , \10814 );
nor \U$10475 ( \10818 , \10816 , \10817 );
and \U$10476 ( \10819 , \10800 , \10818 );
not \U$10477 ( \10820 , \10800 );
not \U$10478 ( \10821 , \10818 );
and \U$10479 ( \10822 , \10820 , \10821 );
or \U$10480 ( \10823 , \10819 , \10822 );
not \U$10481 ( \10824 , \10823 );
or \U$10482 ( \10825 , \10791 , \10824 );
or \U$10483 ( \10826 , \10823 , \10790 );
nand \U$10484 ( \10827 , \10825 , \10826 );
buf \U$10485 ( \10828 , \10827 );
xor \U$10486 ( \10829 , \10692 , \10704 );
and \U$10487 ( \10830 , \10829 , \10715 );
and \U$10488 ( \10831 , \10692 , \10704 );
or \U$10489 ( \10832 , \10830 , \10831 );
not \U$10490 ( \10833 , \10832 );
and \U$10491 ( \10834 , \10828 , \10833 );
not \U$10492 ( \10835 , \10828 );
and \U$10493 ( \10836 , \10835 , \10832 );
nor \U$10494 ( \10837 , \10834 , \10836 );
not \U$10495 ( \10838 , \5034 );
not \U$10496 ( \10839 , \10654 );
or \U$10497 ( \10840 , \10838 , \10839 );
not \U$10498 ( \10841 , RI9872478_154);
not \U$10499 ( \10842 , \1344 );
or \U$10500 ( \10843 , \10841 , \10842 );
or \U$10501 ( \10844 , \1340 , RI9872478_154);
nand \U$10502 ( \10845 , \10843 , \10844 );
nand \U$10503 ( \10846 , \5036 , \10845 );
nand \U$10504 ( \10847 , \10840 , \10846 );
not \U$10505 ( \10848 , \10251 );
not \U$10506 ( \10849 , \10623 );
or \U$10507 ( \10850 , \10848 , \10849 );
not \U$10508 ( \10851 , \8807 );
not \U$10509 ( \10852 , \780 );
or \U$10510 ( \10853 , \10851 , \10852 );
or \U$10511 ( \10854 , \1692 , \8811 );
nand \U$10512 ( \10855 , \10853 , \10854 );
nand \U$10513 ( \10856 , \10855 , \10624 );
nand \U$10514 ( \10857 , \10850 , \10856 );
xor \U$10515 ( \10858 , \10847 , \10857 );
not \U$10516 ( \10859 , \9214 );
and \U$10517 ( \10860 , \1416 , \9198 );
not \U$10518 ( \10861 , \1416 );
and \U$10519 ( \10862 , \10861 , RI9872b80_169);
nor \U$10520 ( \10863 , \10860 , \10862 );
not \U$10521 ( \10864 , \10863 );
or \U$10522 ( \10865 , \10859 , \10864 );
nand \U$10523 ( \10866 , \10676 , \10679 );
nand \U$10524 ( \10867 , \10865 , \10866 );
and \U$10525 ( \10868 , \10858 , \10867 );
not \U$10526 ( \10869 , \10858 );
not \U$10527 ( \10870 , \10867 );
and \U$10528 ( \10871 , \10869 , \10870 );
nor \U$10529 ( \10872 , \10868 , \10871 );
not \U$10530 ( \10873 , \9374 );
and \U$10531 ( \10874 , RI9871c08_136, \10873 );
not \U$10532 ( \10875 , RI9871c08_136);
and \U$10533 ( \10876 , \10875 , \5739 );
nor \U$10534 ( \10877 , \10874 , \10876 );
not \U$10535 ( \10878 , \1430 );
or \U$10536 ( \10879 , \10877 , \10878 );
not \U$10537 ( \10880 , \10633 );
or \U$10538 ( \10881 , \10880 , \5411 );
nand \U$10539 ( \10882 , \10879 , \10881 );
not \U$10540 ( \10883 , \1083 );
not \U$10541 ( \10884 , \10641 );
or \U$10542 ( \10885 , \10883 , \10884 );
xor \U$10543 ( \10886 , RI98718c0_129, \4712 );
nand \U$10544 ( \10887 , \10886 , \1136 );
nand \U$10545 ( \10888 , \10885 , \10887 );
xor \U$10546 ( \10889 , \10882 , \10888 );
not \U$10547 ( \10890 , \7188 );
not \U$10548 ( \10891 , \5644 );
not \U$10549 ( \10892 , \1550 );
or \U$10550 ( \10893 , \10891 , \10892 );
or \U$10551 ( \10894 , \3836 , \5648 );
nand \U$10552 ( \10895 , \10893 , \10894 );
not \U$10553 ( \10896 , \10895 );
or \U$10554 ( \10897 , \10890 , \10896 );
nand \U$10555 ( \10898 , \10386 , \5642 );
nand \U$10556 ( \10899 , \10897 , \10898 );
xor \U$10557 ( \10900 , \10889 , \10899 );
xor \U$10558 ( \10901 , \10872 , \10900 );
not \U$10559 ( \10902 , \4920 );
not \U$10560 ( \10903 , \10664 );
or \U$10561 ( \10904 , \10902 , \10903 );
not \U$10562 ( \10905 , \4902 );
not \U$10563 ( \10906 , \1062 );
or \U$10564 ( \10907 , \10905 , \10906 );
or \U$10565 ( \10908 , \10133 , \4902 );
nand \U$10566 ( \10909 , \10907 , \10908 );
nand \U$10567 ( \10910 , \4925 , \10909 );
nand \U$10568 ( \10911 , \10904 , \10910 );
not \U$10569 ( \10912 , \8029 );
not \U$10570 ( \10913 , \10503 );
or \U$10571 ( \10914 , \10912 , \10913 );
not \U$10572 ( \10915 , RI9872a18_166);
not \U$10573 ( \10916 , \9230 );
or \U$10574 ( \10917 , \10915 , \10916 );
or \U$10575 ( \10918 , \1320 , RI9872a18_166);
nand \U$10576 ( \10919 , \10917 , \10918 );
nand \U$10577 ( \10920 , \8041 , \10919 );
nand \U$10578 ( \10921 , \10914 , \10920 );
xor \U$10579 ( \10922 , \10911 , \10921 );
not \U$10580 ( \10923 , \4103 );
not \U$10581 ( \10924 , \10480 );
or \U$10582 ( \10925 , \10923 , \10924 );
xor \U$10583 ( \10926 , RI98725e0_157, \7605 );
nand \U$10584 ( \10927 , \10926 , \5847 );
nand \U$10585 ( \10928 , \10925 , \10927 );
xor \U$10586 ( \10929 , \10922 , \10928 );
xnor \U$10587 ( \10930 , \10901 , \10929 );
xor \U$10588 ( \10931 , \10837 , \10930 );
not \U$10589 ( \10932 , \2087 );
not \U$10590 ( \10933 , \2076 );
not \U$10591 ( \10934 , \3537 );
or \U$10592 ( \10935 , \10933 , \10934 );
or \U$10593 ( \10936 , \3543 , \2080 );
nand \U$10594 ( \10937 , \10935 , \10936 );
not \U$10595 ( \10938 , \10937 );
or \U$10596 ( \10939 , \10932 , \10938 );
or \U$10597 ( \10940 , \10701 , \2073 );
nand \U$10598 ( \10941 , \10939 , \10940 );
not \U$10599 ( \10942 , \2947 );
xor \U$10600 ( \10943 , \10942 , RI9872310_151);
not \U$10601 ( \10944 , \10943 );
or \U$10602 ( \10945 , \10944 , \4261 );
not \U$10603 ( \10946 , \10448 );
not \U$10604 ( \10947 , \6653 );
or \U$10605 ( \10948 , \10946 , \10947 );
nand \U$10606 ( \10949 , \10945 , \10948 );
xor \U$10607 ( \10950 , \10941 , \10949 );
not \U$10608 ( \10951 , \6284 );
not \U$10609 ( \10952 , \10711 );
or \U$10610 ( \10953 , \10951 , \10952 );
not \U$10611 ( \10954 , RI98728b0_163);
not \U$10612 ( \10955 , \8006 );
or \U$10613 ( \10956 , \10954 , \10955 );
or \U$10614 ( \10957 , \8006 , RI98728b0_163);
nand \U$10615 ( \10958 , \10956 , \10957 );
not \U$10616 ( \10959 , \10958 );
not \U$10617 ( \10960 , \6611 );
or \U$10618 ( \10961 , \10959 , \10960 );
nand \U$10619 ( \10962 , \10953 , \10961 );
xor \U$10620 ( \10963 , \10950 , \10962 );
xor \U$10621 ( \10964 , \10658 , \10681 );
and \U$10622 ( \10965 , \10964 , \10668 );
and \U$10623 ( \10966 , \10658 , \10681 );
nor \U$10624 ( \10967 , \10965 , \10966 );
xor \U$10625 ( \10968 , \10963 , \10967 );
not \U$10626 ( \10969 , \3466 );
not \U$10627 ( \10970 , \10458 );
or \U$10628 ( \10971 , \10969 , \10970 );
and \U$10629 ( \10972 , \10235 , \4063 );
not \U$10630 ( \10973 , \10235 );
and \U$10631 ( \10974 , \10973 , RI98726d0_159);
nor \U$10632 ( \10975 , \10972 , \10974 );
nand \U$10633 ( \10976 , \10975 , \3467 );
nand \U$10634 ( \10977 , \10971 , \10976 );
not \U$10635 ( \10978 , \10487 );
not \U$10636 ( \10979 , RI9872bf8_170);
not \U$10637 ( \10980 , \2399 );
or \U$10638 ( \10981 , \10979 , \10980 );
or \U$10639 ( \10982 , \2399 , RI9872bf8_170);
nand \U$10640 ( \10983 , \10981 , \10982 );
not \U$10641 ( \10984 , \10983 );
or \U$10642 ( \10985 , \10978 , \10984 );
nand \U$10643 ( \10986 , \10493 , \9670 );
nand \U$10644 ( \10987 , \10985 , \10986 );
not \U$10645 ( \10988 , \10987 );
xor \U$10646 ( \10989 , \10977 , \10988 );
not \U$10647 ( \10990 , \7326 );
not \U$10648 ( \10991 , \10464 );
or \U$10649 ( \10992 , \10990 , \10991 );
and \U$10650 ( \10993 , \916 , \7333 );
not \U$10651 ( \10994 , \916 );
and \U$10652 ( \10995 , \10994 , RI98729a0_165);
nor \U$10653 ( \10996 , \10993 , \10995 );
nand \U$10654 ( \10997 , \10996 , \7338 );
nand \U$10655 ( \10998 , \10992 , \10997 );
xnor \U$10656 ( \10999 , \10989 , \10998 );
xor \U$10657 ( \11000 , \10968 , \10999 );
xor \U$10658 ( \11001 , \10931 , \11000 );
not \U$10659 ( \11002 , \11001 );
or \U$10660 ( \11003 , \10771 , \11002 );
or \U$10661 ( \11004 , \11001 , \10770 );
nand \U$10662 ( \11005 , \11003 , \11004 );
not \U$10663 ( \11006 , \11005 );
not \U$10664 ( \11007 , \10341 );
not \U$10665 ( \11008 , \10347 );
not \U$10666 ( \11009 , \10358 );
or \U$10667 ( \11010 , \11008 , \11009 );
or \U$10668 ( \11011 , \10358 , \10347 );
nand \U$10669 ( \11012 , \11010 , \11011 );
not \U$10670 ( \11013 , \11012 );
or \U$10671 ( \11014 , \11007 , \11013 );
not \U$10672 ( \11015 , \10347 );
nand \U$10673 ( \11016 , \11015 , \10358 );
nand \U$10674 ( \11017 , \11014 , \11016 );
not \U$10675 ( \11018 , \11017 );
xor \U$10676 ( \11019 , \10530 , \10535 );
and \U$10677 ( \11020 , \11019 , \10547 );
and \U$10678 ( \11021 , \10530 , \10535 );
or \U$10679 ( \11022 , \11020 , \11021 );
xor \U$10680 ( \11023 , \10397 , \10407 );
and \U$10681 ( \11024 , \11023 , \10420 );
and \U$10682 ( \11025 , \10397 , \10407 );
or \U$10683 ( \11026 , \11024 , \11025 );
not \U$10684 ( \11027 , \797 );
not \U$10685 ( \11028 , \5594 );
not \U$10686 ( \11029 , \11028 );
xor \U$10687 ( \11030 , \11029 , RI98719b0_131);
not \U$10688 ( \11031 , \11030 );
or \U$10689 ( \11032 , \11027 , \11031 );
nand \U$10690 ( \11033 , \10688 , \793 );
nand \U$10691 ( \11034 , \11032 , \11033 );
xor \U$10692 ( \11035 , \8992 , \11034 );
xor \U$10693 ( \11036 , \11026 , \11035 );
not \U$10694 ( \11037 , \11036 );
and \U$10695 ( \11038 , \9000 , \9029 );
and \U$10696 ( \11039 , \8993 , \8999 );
nor \U$10697 ( \11040 , \11038 , \11039 );
not \U$10698 ( \11041 , \11040 );
or \U$10699 ( \11042 , \11037 , \11041 );
or \U$10700 ( \11043 , \11040 , \11036 );
nand \U$10701 ( \11044 , \11042 , \11043 );
xor \U$10702 ( \11045 , \11022 , \11044 );
not \U$10703 ( \11046 , \11045 );
not \U$10704 ( \11047 , \9038 );
and \U$10705 ( \11048 , \11047 , \8833 );
not \U$10706 ( \11049 , \8978 );
nor \U$10707 ( \11050 , \11049 , \9034 );
nor \U$10708 ( \11051 , \11048 , \11050 );
not \U$10709 ( \11052 , \11051 );
or \U$10710 ( \11053 , \11046 , \11052 );
or \U$10711 ( \11054 , \11051 , \11045 );
nand \U$10712 ( \11055 , \11053 , \11054 );
not \U$10713 ( \11056 , \11055 );
not \U$10714 ( \11057 , \11056 );
and \U$10715 ( \11058 , \11018 , \11057 );
and \U$10716 ( \11059 , \11017 , \11056 );
nor \U$10717 ( \11060 , \11058 , \11059 );
not \U$10718 ( \11061 , \11060 );
and \U$10719 ( \11062 , \11006 , \11061 );
and \U$10720 ( \11063 , \11005 , \11060 );
nor \U$10721 ( \11064 , \11062 , \11063 );
xor \U$10722 ( \11065 , \10762 , \10764 );
xor \U$10723 ( \11066 , \11065 , \10767 );
not \U$10724 ( \11067 , \11066 );
nand \U$10725 ( \11068 , \10553 , \10562 );
xor \U$10726 ( \11069 , \11068 , \10559 );
not \U$10727 ( \11070 , \11069 );
or \U$10728 ( \11071 , \11067 , \11070 );
or \U$10729 ( \11072 , \11066 , \11069 );
nand \U$10730 ( \11073 , \11071 , \11072 );
not \U$10731 ( \11074 , \11073 );
xor \U$10732 ( \11075 , \9154 , \9054 );
not \U$10733 ( \11076 , \11075 );
not \U$10734 ( \11077 , \9299 );
nand \U$10735 ( \11078 , \11077 , \9344 );
and \U$10736 ( \11079 , \11078 , \9338 );
not \U$10737 ( \11080 , \11078 );
and \U$10738 ( \11081 , \11080 , \9339 );
nor \U$10739 ( \11082 , \11079 , \11081 );
not \U$10740 ( \11083 , \11082 );
xor \U$10741 ( \11084 , \9296 , \9251 );
not \U$10742 ( \11085 , \9269 );
xor \U$10743 ( \11086 , \11084 , \11085 );
not \U$10744 ( \11087 , \11086 );
not \U$10745 ( \11088 , \11087 );
xor \U$10746 ( \11089 , \9319 , \9333 );
xor \U$10747 ( \11090 , \11089 , \9310 );
xor \U$10748 ( \11091 , \9523 , \9548 );
xnor \U$10749 ( \11092 , \11091 , \9538 );
xor \U$10750 ( \11093 , \11090 , \11092 );
not \U$10751 ( \11094 , \11093 );
or \U$10752 ( \11095 , \11088 , \11094 );
nand \U$10753 ( \11096 , \11090 , \11092 );
nand \U$10754 ( \11097 , \11095 , \11096 );
not \U$10755 ( \11098 , \11097 );
or \U$10756 ( \11099 , \11083 , \11098 );
or \U$10757 ( \11100 , \11097 , \11082 );
nand \U$10758 ( \11101 , \11099 , \11100 );
not \U$10759 ( \11102 , \11101 );
or \U$10760 ( \11103 , \11076 , \11102 );
not \U$10761 ( \11104 , \11082 );
nand \U$10762 ( \11105 , \11104 , \11097 );
nand \U$10763 ( \11106 , \11103 , \11105 );
not \U$10764 ( \11107 , \11106 );
not \U$10765 ( \11108 , \7188 );
not \U$10766 ( \11109 , \9328 );
or \U$10767 ( \11110 , \11108 , \11109 );
and \U$10768 ( \11111 , RI9872568_156, \3127 );
not \U$10769 ( \11112 , RI9872568_156);
not \U$10770 ( \11113 , \1208 );
buf \U$10771 ( \11114 , \11113 );
and \U$10772 ( \11115 , \11112 , \11114 );
or \U$10773 ( \11116 , \11111 , \11115 );
nand \U$10774 ( \11117 , \11116 , \5642 );
nand \U$10775 ( \11118 , \11110 , \11117 );
not \U$10776 ( \11119 , \11118 );
not \U$10777 ( \11120 , \9668 );
not \U$10778 ( \11121 , \9241 );
or \U$10779 ( \11122 , \11120 , \11121 );
not \U$10780 ( \11123 , RI9872bf8_170);
not \U$10781 ( \11124 , \6585 );
or \U$10782 ( \11125 , \11123 , \11124 );
or \U$10783 ( \11126 , \915 , RI9872bf8_170);
nand \U$10784 ( \11127 , \11125 , \11126 );
nand \U$10785 ( \11128 , \11127 , \9670 );
nand \U$10786 ( \11129 , \11122 , \11128 );
not \U$10787 ( \11130 , \8801 );
not \U$10788 ( \11131 , \9315 );
or \U$10789 ( \11132 , \11130 , \11131 );
not \U$10790 ( \11133 , RI9872d60_173);
not \U$10791 ( \11134 , \1318 );
or \U$10792 ( \11135 , \11133 , \11134 );
or \U$10793 ( \11136 , \1319 , RI9872d60_173);
nand \U$10794 ( \11137 , \11135 , \11136 );
nand \U$10795 ( \11138 , \11137 , \9312 );
nand \U$10796 ( \11139 , \11132 , \11138 );
xor \U$10797 ( \11140 , \11129 , \11139 );
not \U$10798 ( \11141 , \11140 );
or \U$10799 ( \11142 , \11119 , \11141 );
nand \U$10800 ( \11143 , \11139 , \11129 );
nand \U$10801 ( \11144 , \11142 , \11143 );
not \U$10802 ( \11145 , \11144 );
not \U$10803 ( \11146 , \4925 );
not \U$10804 ( \11147 , \9166 );
or \U$10805 ( \11148 , \11146 , \11147 );
and \U$10806 ( \11149 , RI9872388_152, \3691 );
not \U$10807 ( \11150 , RI9872388_152);
and \U$10808 ( \11151 , \11150 , \10942 );
or \U$10809 ( \11152 , \11149 , \11151 );
nand \U$10810 ( \11153 , \11152 , \6553 );
nand \U$10811 ( \11154 , \11148 , \11153 );
not \U$10812 ( \11155 , \11154 );
not \U$10813 ( \11156 , \5796 );
not \U$10814 ( \11157 , \9259 );
or \U$10815 ( \11158 , \11156 , \11157 );
and \U$10816 ( \11159 , \1485 , \5025 );
not \U$10817 ( \11160 , \1485 );
and \U$10818 ( \11161 , \11160 , RI9872478_154);
nor \U$10819 ( \11162 , \11159 , \11161 );
nand \U$10820 ( \11163 , \11162 , \5034 );
nand \U$10821 ( \11164 , \11158 , \11163 );
not \U$10822 ( \11165 , \9273 );
not \U$10823 ( \11166 , \9286 );
or \U$10824 ( \11167 , \11165 , \11166 );
xor \U$10825 ( \11168 , RI9872e50_175, \1415 );
nand \U$10826 ( \11169 , \11168 , \9686 );
nand \U$10827 ( \11170 , \11167 , \11169 );
and \U$10828 ( \11171 , \11164 , \11170 );
not \U$10829 ( \11172 , \11164 );
not \U$10830 ( \11173 , \11170 );
and \U$10831 ( \11174 , \11172 , \11173 );
nor \U$10832 ( \11175 , \11171 , \11174 );
not \U$10833 ( \11176 , \11175 );
or \U$10834 ( \11177 , \11155 , \11176 );
nand \U$10835 ( \11178 , \11164 , \11170 );
nand \U$10836 ( \11179 , \11177 , \11178 );
not \U$10837 ( \11180 , \6611 );
not \U$10838 ( \11181 , \9301 );
or \U$10839 ( \11182 , \11180 , \11181 );
not \U$10840 ( \11183 , \7049 );
not \U$10841 ( \11184 , \10133 );
or \U$10842 ( \11185 , \11183 , \11184 );
or \U$10843 ( \11186 , \1062 , \7049 );
nand \U$10844 ( \11187 , \11185 , \11186 );
nand \U$10845 ( \11188 , \11187 , \6284 );
nand \U$10846 ( \11189 , \11182 , \11188 );
not \U$10847 ( \11190 , \11189 );
not \U$10848 ( \11191 , \8743 );
nor \U$10849 ( \11192 , \1120 , \1112 );
not \U$10850 ( \11193 , \11192 );
nand \U$10851 ( \11194 , \11193 , \1124 );
xor \U$10852 ( \11195 , RI9872f40_177, \11194 );
not \U$10853 ( \11196 , \11195 );
or \U$10854 ( \11197 , \11191 , \11196 );
buf \U$10855 ( \11198 , \8751 );
buf \U$10856 ( \11199 , \11198 );
nand \U$10857 ( \11200 , \9534 , \11199 );
nand \U$10858 ( \11201 , \11197 , \11200 );
not \U$10859 ( \11202 , \6145 );
not \U$10860 ( \11203 , \9521 );
or \U$10861 ( \11204 , \11202 , \11203 );
not \U$10862 ( \11205 , RI98719b0_131);
not \U$10863 ( \11206 , \6481 );
or \U$10864 ( \11207 , \11205 , \11206 );
or \U$10865 ( \11208 , \6059 , RI98719b0_131);
nand \U$10866 ( \11209 , \11207 , \11208 );
nand \U$10867 ( \11210 , \11209 , \793 );
nand \U$10868 ( \11211 , \11204 , \11210 );
xor \U$10869 ( \11212 , \11201 , \11211 );
not \U$10870 ( \11213 , \11212 );
or \U$10871 ( \11214 , \11190 , \11213 );
nand \U$10872 ( \11215 , \11201 , \11211 );
nand \U$10873 ( \11216 , \11214 , \11215 );
and \U$10874 ( \11217 , \11179 , \11216 );
not \U$10875 ( \11218 , \11179 );
not \U$10876 ( \11219 , \11216 );
and \U$10877 ( \11220 , \11218 , \11219 );
nor \U$10878 ( \11221 , \11217 , \11220 );
not \U$10879 ( \11222 , \11221 );
or \U$10880 ( \11223 , \11145 , \11222 );
not \U$10881 ( \11224 , \11219 );
nand \U$10882 ( \11225 , \11224 , \11179 );
nand \U$10883 ( \11226 , \11223 , \11225 );
not \U$10884 ( \11227 , \11226 );
not \U$10885 ( \11228 , \9640 );
not \U$10886 ( \11229 , \9551 );
and \U$10887 ( \11230 , \11228 , \11229 );
and \U$10888 ( \11231 , \9640 , \9551 );
nor \U$10889 ( \11232 , \11230 , \11231 );
not \U$10890 ( \11233 , \11232 );
not \U$10891 ( \11234 , \11233 );
not \U$10892 ( \11235 , \5847 );
not \U$10893 ( \11236 , \9179 );
or \U$10894 ( \11237 , \11235 , \11236 );
and \U$10895 ( \11238 , RI98725e0_157, \3542 );
not \U$10896 ( \11239 , RI98725e0_157);
and \U$10897 ( \11240 , \11239 , \3537 );
or \U$10898 ( \11241 , \11238 , \11240 );
nand \U$10899 ( \11242 , \11241 , \4101 );
nand \U$10900 ( \11243 , \11237 , \11242 );
not \U$10901 ( \11244 , \11243 );
not \U$10902 ( \11245 , \9145 );
not \U$10903 ( \11246 , \9214 );
not \U$10904 ( \11247 , \9207 );
or \U$10905 ( \11248 , \11246 , \11247 );
xor \U$10906 ( \11249 , RI9872b80_169, \8004 );
nand \U$10907 ( \11250 , \11249 , \10679 );
nand \U$10908 ( \11251 , \11248 , \11250 );
not \U$10909 ( \11252 , \11251 );
or \U$10910 ( \11253 , \11245 , \11252 );
or \U$10911 ( \11254 , \11251 , \9145 );
nand \U$10912 ( \11255 , \11253 , \11254 );
not \U$10913 ( \11256 , \11255 );
or \U$10914 ( \11257 , \11244 , \11256 );
nand \U$10915 ( \11258 , \11251 , \9142 );
nand \U$10916 ( \11259 , \11257 , \11258 );
not \U$10917 ( \11260 , \9564 );
and \U$10918 ( \11261 , \9592 , \11260 );
not \U$10919 ( \11262 , \9592 );
and \U$10920 ( \11263 , \11262 , \9564 );
nor \U$10921 ( \11264 , \11261 , \11263 );
not \U$10922 ( \11265 , \11264 );
or \U$10923 ( \11266 , \11259 , \11265 );
not \U$10924 ( \11267 , \3170 );
not \U$10925 ( \11268 , \10035 );
or \U$10926 ( \11269 , \11267 , \11268 );
and \U$10927 ( \11270 , \4471 , \3154 );
not \U$10928 ( \11271 , \4471 );
and \U$10929 ( \11272 , \11271 , RI9872310_151);
nor \U$10930 ( \11273 , \11270 , \11272 );
nand \U$10931 ( \11274 , \11273 , \3164 );
nand \U$10932 ( \11275 , \11269 , \11274 );
not \U$10933 ( \11276 , \11275 );
not \U$10934 ( \11277 , \8041 );
not \U$10935 ( \11278 , \9078 );
or \U$10936 ( \11279 , \11277 , \11278 );
not \U$10937 ( \11280 , \8031 );
not \U$10938 ( \11281 , \943 );
or \U$10939 ( \11282 , \11280 , \11281 );
not \U$10940 ( \11283 , \5907 );
or \U$10941 ( \11284 , \11283 , \8031 );
nand \U$10942 ( \11285 , \11282 , \11284 );
nand \U$10943 ( \11286 , \11285 , \9079 );
nand \U$10944 ( \11287 , \11279 , \11286 );
not \U$10945 ( \11288 , \3465 );
not \U$10946 ( \11289 , RI98726d0_159);
not \U$10947 ( \11290 , \5595 );
or \U$10948 ( \11291 , \11289 , \11290 );
or \U$10949 ( \11292 , \5595 , RI98726d0_159);
nand \U$10950 ( \11293 , \11291 , \11292 );
not \U$10951 ( \11294 , \11293 );
or \U$10952 ( \11295 , \11288 , \11294 );
nand \U$10953 ( \11296 , \9063 , \3467 );
nand \U$10954 ( \11297 , \11295 , \11296 );
xor \U$10955 ( \11298 , \11287 , \11297 );
not \U$10956 ( \11299 , \11298 );
or \U$10957 ( \11300 , \11276 , \11299 );
nand \U$10958 ( \11301 , \11287 , \11297 );
nand \U$10959 ( \11302 , \11300 , \11301 );
nand \U$10960 ( \11303 , \11266 , \11302 );
nand \U$10961 ( \11304 , \11259 , \11265 );
nand \U$10962 ( \11305 , \11303 , \11304 );
not \U$10963 ( \11306 , \11305 );
not \U$10964 ( \11307 , \11306 );
or \U$10965 ( \11308 , \11234 , \11307 );
nand \U$10966 ( \11309 , \11305 , \11232 );
nand \U$10967 ( \11310 , \11308 , \11309 );
not \U$10968 ( \11311 , \11310 );
or \U$10969 ( \11312 , \11227 , \11311 );
nand \U$10970 ( \11313 , \11305 , \11233 );
nand \U$10971 ( \11314 , \11312 , \11313 );
xor \U$10972 ( \11315 , \9348 , \9346 );
xnor \U$10973 ( \11316 , \11315 , \9158 );
xor \U$10974 ( \11317 , \11314 , \11316 );
not \U$10975 ( \11318 , \11317 );
or \U$10976 ( \11319 , \11107 , \11318 );
nand \U$10977 ( \11320 , \11314 , \11316 );
nand \U$10978 ( \11321 , \11319 , \11320 );
not \U$10979 ( \11322 , \11321 );
or \U$10980 ( \11323 , \11074 , \11322 );
not \U$10981 ( \11324 , \11069 );
nand \U$10982 ( \11325 , \11324 , \11066 );
nand \U$10983 ( \11326 , \11323 , \11325 );
xor \U$10984 ( \11327 , \11064 , \11326 );
not \U$10985 ( \11328 , \11327 );
and \U$10986 ( \11329 , \10760 , \11328 );
and \U$10987 ( \11330 , \11327 , \10759 );
nor \U$10988 ( \11331 , \11329 , \11330 );
not \U$10989 ( \11332 , \11331 );
xor \U$10990 ( \11333 , \10365 , \11332 );
xor \U$10991 ( \11334 , \9861 , \9959 );
not \U$10992 ( \11335 , \11334 );
xor \U$10993 ( \11336 , \9065 , \9147 );
and \U$10994 ( \11337 , RI9873210_183, RI9873198_182);
not \U$10995 ( \11338 , RI9873210_183);
not \U$10996 ( \11339 , RI9873198_182);
and \U$10997 ( \11340 , \11338 , \11339 );
nor \U$10998 ( \11341 , \11337 , \11340 );
buf \U$10999 ( \11342 , \11341 );
not \U$11000 ( \11343 , \11342 );
not \U$11001 ( \11344 , \11343 );
not \U$11002 ( \11345 , \11341 );
and \U$11003 ( \11346 , RI98730a8_180, RI9873198_182);
not \U$11004 ( \11347 , RI98730a8_180);
and \U$11005 ( \11348 , \11347 , \11339 );
nor \U$11006 ( \11349 , \11346 , \11348 );
and \U$11007 ( \11350 , \11345 , \11349 );
not \U$11008 ( \11351 , \11350 );
not \U$11009 ( \11352 , \11351 );
or \U$11010 ( \11353 , \11344 , \11352 );
nand \U$11011 ( \11354 , \11353 , RI98730a8_180);
not \U$11012 ( \11355 , \6316 );
not \U$11013 ( \11356 , \9140 );
or \U$11014 ( \11357 , \11355 , \11356 );
not \U$11015 ( \11358 , \10063 );
and \U$11016 ( \11359 , \11358 , \1165 );
not \U$11017 ( \11360 , \11358 );
and \U$11018 ( \11361 , \11360 , \10368 );
nor \U$11019 ( \11362 , \11359 , \11361 );
nand \U$11020 ( \11363 , \11362 , \1162 );
nand \U$11021 ( \11364 , \11357 , \11363 );
xor \U$11022 ( \11365 , \11354 , \11364 );
not \U$11023 ( \11366 , \1018 );
not \U$11024 ( \11367 , \1044 );
not \U$11025 ( \11368 , \9114 );
or \U$11026 ( \11369 , \11367 , \11368 );
not \U$11027 ( \11370 , \9113 );
not \U$11028 ( \11371 , \11370 );
or \U$11029 ( \11372 , \11371 , \8085 );
nand \U$11030 ( \11373 , \11369 , \11372 );
not \U$11031 ( \11374 , \11373 );
or \U$11032 ( \11375 , \11366 , \11374 );
nand \U$11033 ( \11376 , \9854 , \1013 );
nand \U$11034 ( \11377 , \11375 , \11376 );
and \U$11035 ( \11378 , \11365 , \11377 );
and \U$11036 ( \11379 , \11354 , \11364 );
nor \U$11037 ( \11380 , \11378 , \11379 );
buf \U$11038 ( \11381 , \11380 );
not \U$11039 ( \11382 , \11381 );
not \U$11040 ( \11383 , \1380 );
and \U$11041 ( \11384 , RI9871e60_141, \8696 );
not \U$11042 ( \11385 , RI9871e60_141);
and \U$11043 ( \11386 , \11385 , \9750 );
or \U$11044 ( \11387 , \11384 , \11386 );
not \U$11045 ( \11388 , \11387 );
or \U$11046 ( \11389 , \11383 , \11388 );
nand \U$11047 ( \11390 , \9928 , \1352 );
nand \U$11048 ( \11391 , \11389 , \11390 );
not \U$11049 ( \11392 , \5350 );
and \U$11050 ( \11393 , \1347 , \8554 );
not \U$11051 ( \11394 , \1347 );
and \U$11052 ( \11395 , \11394 , \10372 );
nor \U$11053 ( \11396 , \11393 , \11395 );
not \U$11054 ( \11397 , \11396 );
or \U$11055 ( \11398 , \11392 , \11397 );
nand \U$11056 ( \11399 , \9915 , \832 );
nand \U$11057 ( \11400 , \11398 , \11399 );
xor \U$11058 ( \11401 , \11391 , \11400 );
not \U$11059 ( \11402 , \9876 );
not \U$11060 ( \11403 , \9887 );
or \U$11061 ( \11404 , \11402 , \11403 );
not \U$11062 ( \11405 , RI9872130_147);
buf \U$11063 ( \11406 , \8649 );
not \U$11064 ( \11407 , \11406 );
or \U$11065 ( \11408 , \11405 , \11407 );
or \U$11066 ( \11409 , \11406 , RI9872130_147);
nand \U$11067 ( \11410 , \11408 , \11409 );
nand \U$11068 ( \11411 , \11410 , \876 );
nand \U$11069 ( \11412 , \11404 , \11411 );
and \U$11070 ( \11413 , \11401 , \11412 );
and \U$11071 ( \11414 , \11391 , \11400 );
or \U$11072 ( \11415 , \11413 , \11414 );
not \U$11073 ( \11416 , \11415 );
or \U$11074 ( \11417 , \11382 , \11416 );
or \U$11075 ( \11418 , \11381 , \11415 );
nand \U$11076 ( \11419 , \11417 , \11418 );
not \U$11077 ( \11420 , \11419 );
not \U$11078 ( \11421 , \1083 );
not \U$11079 ( \11422 , \1111 );
not \U$11080 ( \11423 , \10412 );
or \U$11081 ( \11424 , \11422 , \11423 );
nand \U$11082 ( \11425 , \6529 , RI98718c0_129);
nand \U$11083 ( \11426 , \11424 , \11425 );
not \U$11084 ( \11427 , \11426 );
or \U$11085 ( \11428 , \11421 , \11427 );
nand \U$11086 ( \11429 , \10074 , \6673 );
nand \U$11087 ( \11430 , \11428 , \11429 );
not \U$11088 ( \11431 , \11430 );
buf \U$11089 ( \11432 , \791 );
buf \U$11090 ( \11433 , \11432 );
not \U$11091 ( \11434 , \11433 );
not \U$11092 ( \11435 , \5703 );
and \U$11093 ( \11436 , RI98719b0_131, \11435 );
not \U$11094 ( \11437 , RI98719b0_131);
not \U$11095 ( \11438 , \7111 );
and \U$11096 ( \11439 , \11437 , \11438 );
or \U$11097 ( \11440 , \11436 , \11439 );
not \U$11098 ( \11441 , \11440 );
or \U$11099 ( \11442 , \11434 , \11441 );
nand \U$11100 ( \11443 , \11209 , \796 );
nand \U$11101 ( \11444 , \11442 , \11443 );
not \U$11102 ( \11445 , \11444 );
buf \U$11103 ( \11446 , \9097 );
not \U$11104 ( \11447 , \11446 );
nand \U$11105 ( \11448 , \9084 , \10054 );
not \U$11106 ( \11449 , \11448 );
and \U$11107 ( \11450 , \11447 , \11449 );
and \U$11108 ( \11451 , \11446 , \11448 );
nor \U$11109 ( \11452 , \11450 , \11451 );
buf \U$11110 ( \11453 , \11452 );
not \U$11111 ( \11454 , \11453 );
not \U$11112 ( \11455 , \11454 );
or \U$11113 ( \11456 , \11455 , \9723 );
and \U$11114 ( \11457 , \11445 , \11456 );
not \U$11115 ( \11458 , \11445 );
not \U$11116 ( \11459 , \11456 );
and \U$11117 ( \11460 , \11458 , \11459 );
nor \U$11118 ( \11461 , \11457 , \11460 );
not \U$11119 ( \11462 , \11461 );
or \U$11120 ( \11463 , \11431 , \11462 );
nand \U$11121 ( \11464 , \11444 , \11459 );
nand \U$11122 ( \11465 , \11463 , \11464 );
not \U$11123 ( \11466 , \11465 );
or \U$11124 ( \11467 , \11420 , \11466 );
not \U$11125 ( \11468 , \11381 );
nand \U$11126 ( \11469 , \11468 , \11415 );
nand \U$11127 ( \11470 , \11467 , \11469 );
xnor \U$11128 ( \11471 , \11336 , \11470 );
not \U$11129 ( \11472 , \11471 );
not \U$11130 ( \11473 , \11472 );
or \U$11131 ( \11474 , \11335 , \11473 );
xor \U$11132 ( \11475 , \9147 , \9065 );
nand \U$11133 ( \11476 , \11475 , \11470 );
nand \U$11134 ( \11477 , \11474 , \11476 );
not \U$11135 ( \11478 , \11477 );
not \U$11136 ( \11479 , \11478 );
xor \U$11137 ( \11480 , \9800 , \9807 );
xor \U$11138 ( \11481 , \11480 , \9818 );
not \U$11139 ( \11482 , \11481 );
xor \U$11140 ( \11483 , \11264 , \11302 );
xor \U$11141 ( \11484 , \11483 , \11259 );
nand \U$11142 ( \11485 , \11482 , \11484 );
not \U$11143 ( \11486 , \11485 );
not \U$11144 ( \11487 , \11144 );
xor \U$11145 ( \11488 , \11216 , \11487 );
xnor \U$11146 ( \11489 , \11488 , \11179 );
not \U$11147 ( \11490 , \11489 );
or \U$11148 ( \11491 , \11486 , \11490 );
not \U$11149 ( \11492 , \11484 );
nand \U$11150 ( \11493 , \11492 , \11481 );
nand \U$11151 ( \11494 , \11491 , \11493 );
not \U$11152 ( \11495 , \11494 );
or \U$11153 ( \11496 , \11479 , \11495 );
or \U$11154 ( \11497 , \11494 , \11478 );
nand \U$11155 ( \11498 , \11496 , \11497 );
not \U$11156 ( \11499 , \11498 );
xor \U$11157 ( \11500 , \9856 , \9829 );
xor \U$11158 ( \11501 , \11500 , \9840 );
not \U$11159 ( \11502 , \11501 );
not \U$11160 ( \11503 , \11189 );
xor \U$11161 ( \11504 , \11211 , \11503 );
xnor \U$11162 ( \11505 , \11504 , \11201 );
not \U$11163 ( \11506 , \11505 );
xor \U$11164 ( \11507 , \11154 , \11170 );
xnor \U$11165 ( \11508 , \11507 , \11164 );
nand \U$11166 ( \11509 , \11506 , \11508 );
not \U$11167 ( \11510 , \11509 );
or \U$11168 ( \11511 , \11502 , \11510 );
not \U$11169 ( \11512 , \11508 );
nand \U$11170 ( \11513 , \11512 , \11505 );
nand \U$11171 ( \11514 , \11511 , \11513 );
not \U$11172 ( \11515 , \11514 );
xor \U$11173 ( \11516 , \11298 , \11275 );
not \U$11174 ( \11517 , \11516 );
and \U$11175 ( \11518 , \11140 , \11118 );
not \U$11176 ( \11519 , \11140 );
not \U$11177 ( \11520 , \11118 );
and \U$11178 ( \11521 , \11519 , \11520 );
nor \U$11179 ( \11522 , \11518 , \11521 );
not \U$11180 ( \11523 , \11522 );
not \U$11181 ( \11524 , \11523 );
xor \U$11182 ( \11525 , \9142 , \11243 );
xnor \U$11183 ( \11526 , \11525 , \11251 );
not \U$11184 ( \11527 , \11526 );
not \U$11185 ( \11528 , \11527 );
or \U$11186 ( \11529 , \11524 , \11528 );
nand \U$11187 ( \11530 , \11526 , \11522 );
nand \U$11188 ( \11531 , \11529 , \11530 );
not \U$11189 ( \11532 , \11531 );
or \U$11190 ( \11533 , \11517 , \11532 );
nand \U$11191 ( \11534 , \11527 , \11522 );
nand \U$11192 ( \11535 , \11533 , \11534 );
not \U$11193 ( \11536 , \2087 );
not \U$11194 ( \11537 , \9827 );
or \U$11195 ( \11538 , \11536 , \11537 );
and \U$11196 ( \11539 , \7028 , RI9871aa0_133);
not \U$11197 ( \11540 , \7028 );
and \U$11198 ( \11541 , \11540 , \2076 );
nor \U$11199 ( \11542 , \11539 , \11541 );
nand \U$11200 ( \11543 , \11542 , \2071 );
nand \U$11201 ( \11544 , \11538 , \11543 );
not \U$11202 ( \11545 , \3170 );
not \U$11203 ( \11546 , \11273 );
or \U$11204 ( \11547 , \11545 , \11546 );
not \U$11205 ( \11548 , \4989 );
and \U$11206 ( \11549 , \3154 , \11548 );
not \U$11207 ( \11550 , \3154 );
and \U$11208 ( \11551 , \11550 , \4960 );
nor \U$11209 ( \11552 , \11549 , \11551 );
nand \U$11210 ( \11553 , \11552 , \6653 );
nand \U$11211 ( \11554 , \11547 , \11553 );
xor \U$11212 ( \11555 , \11544 , \11554 );
not \U$11213 ( \11556 , \8041 );
not \U$11214 ( \11557 , \11285 );
or \U$11215 ( \11558 , \11556 , \11557 );
not \U$11216 ( \11559 , \1252 );
xor \U$11217 ( \11560 , \11559 , RI9872a18_166);
nand \U$11218 ( \11561 , \11560 , \9079 );
nand \U$11219 ( \11562 , \11558 , \11561 );
and \U$11220 ( \11563 , \11555 , \11562 );
and \U$11221 ( \11564 , \11544 , \11554 );
or \U$11222 ( \11565 , \11563 , \11564 );
not \U$11223 ( \11566 , \11565 );
not \U$11224 ( \11567 , \7325 );
and \U$11225 ( \11568 , RI98729a0_165, \1603 );
not \U$11226 ( \11569 , RI98729a0_165);
and \U$11227 ( \11570 , \11569 , \1370 );
or \U$11228 ( \11571 , \11568 , \11570 );
not \U$11229 ( \11572 , \11571 );
or \U$11230 ( \11573 , \11567 , \11572 );
nand \U$11231 ( \11574 , \9836 , \7338 );
nand \U$11232 ( \11575 , \11573 , \11574 );
not \U$11233 ( \11576 , \11575 );
xor \U$11234 ( \11577 , RI9873030_179, \1393 );
not \U$11235 ( \11578 , \11577 );
not \U$11236 ( \11579 , \9952 );
or \U$11237 ( \11580 , \11578 , \11579 );
not \U$11238 ( \11581 , \9937 );
or \U$11239 ( \11582 , \9944 , \11581 );
nand \U$11240 ( \11583 , \11580 , \11582 );
not \U$11241 ( \11584 , \11583 );
not \U$11242 ( \11585 , \9686 );
not \U$11243 ( \11586 , RI9872e50_175);
not \U$11244 ( \11587 , \1446 );
or \U$11245 ( \11588 , \11586 , \11587 );
or \U$11246 ( \11589 , \1446 , RI9872e50_175);
nand \U$11247 ( \11590 , \11588 , \11589 );
not \U$11248 ( \11591 , \11590 );
or \U$11249 ( \11592 , \11585 , \11591 );
nand \U$11250 ( \11593 , \11168 , \10331 );
nand \U$11251 ( \11594 , \11592 , \11593 );
not \U$11252 ( \11595 , \11594 );
not \U$11253 ( \11596 , \11595 );
or \U$11254 ( \11597 , \11584 , \11596 );
not \U$11255 ( \11598 , \11583 );
nand \U$11256 ( \11599 , \11598 , \11594 );
nand \U$11257 ( \11600 , \11597 , \11599 );
not \U$11258 ( \11601 , \11600 );
or \U$11259 ( \11602 , \11576 , \11601 );
nand \U$11260 ( \11603 , \11594 , \11583 );
nand \U$11261 ( \11604 , \11602 , \11603 );
not \U$11262 ( \11605 , \1456 );
and \U$11263 ( \11606 , RI9871c08_136, \9570 );
not \U$11264 ( \11607 , RI9871c08_136);
and \U$11265 ( \11608 , \11607 , \8924 );
nor \U$11266 ( \11609 , \11606 , \11608 );
not \U$11267 ( \11610 , \11609 );
or \U$11268 ( \11611 , \11605 , \11610 );
nand \U$11269 ( \11612 , \10047 , \1429 );
nand \U$11270 ( \11613 , \11611 , \11612 );
not \U$11271 ( \11614 , \11613 );
not \U$11272 ( \11615 , \1501 );
not \U$11273 ( \11616 , RI9871c80_137);
not \U$11274 ( \11617 , \8607 );
or \U$11275 ( \11618 , \11616 , \11617 );
nand \U$11276 ( \11619 , \8597 , \1584 );
nand \U$11277 ( \11620 , \11618 , \11619 );
not \U$11278 ( \11621 , \11620 );
or \U$11279 ( \11622 , \11615 , \11621 );
nand \U$11280 ( \11623 , \9871 , \1518 );
nand \U$11281 ( \11624 , \11622 , \11623 );
not \U$11282 ( \11625 , \1292 );
not \U$11283 ( \11626 , \4044 );
not \U$11284 ( \11627 , \9598 );
buf \U$11285 ( \11628 , \11627 );
not \U$11286 ( \11629 , \11628 );
not \U$11287 ( \11630 , \11629 );
or \U$11288 ( \11631 , \11626 , \11630 );
nand \U$11289 ( \11632 , \10392 , RI9871b18_134);
nand \U$11290 ( \11633 , \11631 , \11632 );
not \U$11291 ( \11634 , \11633 );
or \U$11292 ( \11635 , \11625 , \11634 );
nand \U$11293 ( \11636 , \9900 , \1323 );
nand \U$11294 ( \11637 , \11635 , \11636 );
xor \U$11295 ( \11638 , \11624 , \11637 );
not \U$11296 ( \11639 , \11638 );
or \U$11297 ( \11640 , \11614 , \11639 );
nand \U$11298 ( \11641 , \11637 , \11624 );
nand \U$11299 ( \11642 , \11640 , \11641 );
not \U$11300 ( \11643 , \11642 );
xor \U$11301 ( \11644 , \11604 , \11643 );
not \U$11302 ( \11645 , \11644 );
not \U$11303 ( \11646 , \11645 );
or \U$11304 ( \11647 , \11566 , \11646 );
not \U$11305 ( \11648 , \11643 );
nand \U$11306 ( \11649 , \11648 , \11604 );
nand \U$11307 ( \11650 , \11647 , \11649 );
xor \U$11308 ( \11651 , \11535 , \11650 );
not \U$11309 ( \11652 , \11651 );
or \U$11310 ( \11653 , \11515 , \11652 );
nand \U$11311 ( \11654 , \11535 , \11650 );
nand \U$11312 ( \11655 , \11653 , \11654 );
not \U$11313 ( \11656 , \11655 );
or \U$11314 ( \11657 , \11499 , \11656 );
not \U$11315 ( \11658 , \11478 );
nand \U$11316 ( \11659 , \11658 , \11494 );
nand \U$11317 ( \11660 , \11657 , \11659 );
not \U$11318 ( \11661 , \11660 );
xor \U$11319 ( \11662 , \10097 , \10199 );
xor \U$11320 ( \11663 , \11662 , \10281 );
xor \U$11321 ( \11664 , \9975 , \9992 );
not \U$11322 ( \11665 , \11664 );
xor \U$11323 ( \11666 , \10092 , \10022 );
xor \U$11324 ( \11667 , \11666 , \10090 );
not \U$11325 ( \11668 , \11667 );
nand \U$11326 ( \11669 , \11665 , \11668 );
not \U$11327 ( \11670 , \11669 );
not \U$11328 ( \11671 , \4101 );
not \U$11329 ( \11672 , \4153 );
and \U$11330 ( \11673 , \11672 , \4088 );
not \U$11331 ( \11674 , \11672 );
and \U$11332 ( \11675 , \11674 , RI98725e0_157);
nor \U$11333 ( \11676 , \11673 , \11675 );
not \U$11334 ( \11677 , \11676 );
or \U$11335 ( \11678 , \11671 , \11677 );
nand \U$11336 ( \11679 , \11241 , \4084 );
nand \U$11337 ( \11680 , \11678 , \11679 );
not \U$11338 ( \11681 , \9214 );
not \U$11339 ( \11682 , \11249 );
or \U$11340 ( \11683 , \11681 , \11682 );
not \U$11341 ( \11684 , \9198 );
not \U$11342 ( \11685 , \846 );
or \U$11343 ( \11686 , \11684 , \11685 );
not \U$11344 ( \11687 , \6224 );
not \U$11345 ( \11688 , RI9872b80_169);
or \U$11346 ( \11689 , \11687 , \11688 );
nand \U$11347 ( \11690 , \11686 , \11689 );
not \U$11348 ( \11691 , \9196 );
not \U$11349 ( \11692 , \11691 );
nand \U$11350 ( \11693 , \11690 , \11692 );
nand \U$11351 ( \11694 , \11683 , \11693 );
xor \U$11352 ( \11695 , \11680 , \11694 );
not \U$11353 ( \11696 , \4919 );
xor \U$11354 ( \11697 , \3240 , RI9872388_152);
not \U$11355 ( \11698 , \11697 );
or \U$11356 ( \11699 , \11696 , \11698 );
nand \U$11357 ( \11700 , \11152 , \4925 );
nand \U$11358 ( \11701 , \11699 , \11700 );
and \U$11359 ( \11702 , \11695 , \11701 );
and \U$11360 ( \11703 , \11680 , \11694 );
or \U$11361 ( \11704 , \11702 , \11703 );
not \U$11362 ( \11705 , \11704 );
not \U$11363 ( \11706 , \5034 );
not \U$11364 ( \11707 , \9162 );
xor \U$11365 ( \11708 , RI9872478_154, \11707 );
not \U$11366 ( \11709 , \11708 );
or \U$11367 ( \11710 , \11706 , \11709 );
nand \U$11368 ( \11711 , \11162 , \5036 );
nand \U$11369 ( \11712 , \11710 , \11711 );
not \U$11370 ( \11713 , \11712 );
not \U$11371 ( \11714 , \11198 );
not \U$11372 ( \11715 , \11195 );
or \U$11373 ( \11716 , \11714 , \11715 );
and \U$11374 ( \11717 , RI9872f40_177, \1096 );
not \U$11375 ( \11718 , RI9872f40_177);
and \U$11376 ( \11719 , \11718 , \1105 );
or \U$11377 ( \11720 , \11717 , \11719 );
nand \U$11378 ( \11721 , \11720 , \9526 );
nand \U$11379 ( \11722 , \11716 , \11721 );
not \U$11380 ( \11723 , \11722 );
or \U$11381 ( \11724 , \11713 , \11723 );
not \U$11382 ( \11725 , \11712 );
and \U$11383 ( \11726 , \11722 , \11725 );
not \U$11384 ( \11727 , \11722 );
and \U$11385 ( \11728 , \11727 , \11712 );
nor \U$11386 ( \11729 , \11726 , \11728 );
not \U$11387 ( \11730 , \11729 );
not \U$11388 ( \11731 , \9670 );
not \U$11389 ( \11732 , RI9872bf8_170);
not \U$11390 ( \11733 , \1505 );
or \U$11391 ( \11734 , \11732 , \11733 );
or \U$11392 ( \11735 , \892 , RI9872bf8_170);
nand \U$11393 ( \11736 , \11734 , \11735 );
not \U$11394 ( \11737 , \11736 );
or \U$11395 ( \11738 , \11731 , \11737 );
nand \U$11396 ( \11739 , \11127 , \9227 );
nand \U$11397 ( \11740 , \11738 , \11739 );
nand \U$11398 ( \11741 , \11730 , \11740 );
nand \U$11399 ( \11742 , \11724 , \11741 );
not \U$11400 ( \11743 , \6284 );
not \U$11401 ( \11744 , RI98728b0_163);
not \U$11402 ( \11745 , \6330 );
or \U$11403 ( \11746 , \11744 , \11745 );
or \U$11404 ( \11747 , \9326 , RI98728b0_163);
nand \U$11405 ( \11748 , \11746 , \11747 );
not \U$11406 ( \11749 , \11748 );
or \U$11407 ( \11750 , \11743 , \11749 );
nand \U$11408 ( \11751 , \11187 , \6611 );
nand \U$11409 ( \11752 , \11750 , \11751 );
not \U$11410 ( \11753 , \11752 );
not \U$11411 ( \11754 , \5642 );
not \U$11412 ( \11755 , \1190 );
xor \U$11413 ( \11756 , \11755 , RI9872568_156);
not \U$11414 ( \11757 , \11756 );
or \U$11415 ( \11758 , \11754 , \11757 );
nand \U$11416 ( \11759 , \11116 , \5653 );
nand \U$11417 ( \11760 , \11758 , \11759 );
not \U$11418 ( \11761 , \11760 );
or \U$11419 ( \11762 , \11753 , \11761 );
or \U$11420 ( \11763 , \11760 , \11752 );
not \U$11421 ( \11764 , \9312 );
not \U$11422 ( \11765 , RI9872d60_173);
not \U$11423 ( \11766 , \7064 );
or \U$11424 ( \11767 , \11765 , \11766 );
or \U$11425 ( \11768 , \7064 , RI9872d60_173);
nand \U$11426 ( \11769 , \11767 , \11768 );
not \U$11427 ( \11770 , \11769 );
or \U$11428 ( \11771 , \11764 , \11770 );
nand \U$11429 ( \11772 , \11137 , \10242 );
nand \U$11430 ( \11773 , \11771 , \11772 );
nand \U$11431 ( \11774 , \11763 , \11773 );
nand \U$11432 ( \11775 , \11762 , \11774 );
xor \U$11433 ( \11776 , \11742 , \11775 );
not \U$11434 ( \11777 , \11776 );
or \U$11435 ( \11778 , \11705 , \11777 );
not \U$11436 ( \11779 , \11742 );
not \U$11437 ( \11780 , \11779 );
nand \U$11438 ( \11781 , \11780 , \11775 );
nand \U$11439 ( \11782 , \11778 , \11781 );
not \U$11440 ( \11783 , \11782 );
not \U$11441 ( \11784 , \10039 );
not \U$11442 ( \11785 , \11784 );
not \U$11443 ( \11786 , \10085 );
or \U$11444 ( \11787 , \11785 , \11786 );
or \U$11445 ( \11788 , \10085 , \11784 );
nand \U$11446 ( \11789 , \11787 , \11788 );
xor \U$11447 ( \11790 , \9873 , \9890 );
xnor \U$11448 ( \11791 , \11790 , \9904 );
not \U$11449 ( \11792 , \11791 );
and \U$11450 ( \11793 , \9917 , \9931 );
not \U$11451 ( \11794 , \9917 );
and \U$11452 ( \11795 , \11794 , \9930 );
nor \U$11453 ( \11796 , \11793 , \11795 );
xor \U$11454 ( \11797 , \9954 , \11796 );
not \U$11455 ( \11798 , \11797 );
not \U$11456 ( \11799 , \10076 );
xor \U$11457 ( \11800 , \10065 , \11799 );
xor \U$11458 ( \11801 , \11800 , \10049 );
not \U$11459 ( \11802 , \11801 );
or \U$11460 ( \11803 , \11798 , \11802 );
or \U$11461 ( \11804 , \11801 , \11797 );
nand \U$11462 ( \11805 , \11803 , \11804 );
not \U$11463 ( \11806 , \11805 );
or \U$11464 ( \11807 , \11792 , \11806 );
not \U$11465 ( \11808 , \11801 );
not \U$11466 ( \11809 , \11808 );
not \U$11467 ( \11810 , \11797 );
nand \U$11468 ( \11811 , \11809 , \11810 );
nand \U$11469 ( \11812 , \11807 , \11811 );
xor \U$11470 ( \11813 , \11789 , \11812 );
not \U$11471 ( \11814 , \11813 );
or \U$11472 ( \11815 , \11783 , \11814 );
nand \U$11473 ( \11816 , \11812 , \11789 );
nand \U$11474 ( \11817 , \11815 , \11816 );
not \U$11475 ( \11818 , \11817 );
or \U$11476 ( \11819 , \11670 , \11818 );
nand \U$11477 ( \11820 , \11667 , \11664 );
nand \U$11478 ( \11821 , \11819 , \11820 );
and \U$11479 ( \11822 , \11663 , \11821 );
not \U$11480 ( \11823 , \11663 );
not \U$11481 ( \11824 , \11821 );
and \U$11482 ( \11825 , \11823 , \11824 );
nor \U$11483 ( \11826 , \11822 , \11825 );
not \U$11484 ( \11827 , \11826 );
or \U$11485 ( \11828 , \11661 , \11827 );
nand \U$11486 ( \11829 , \11663 , \11821 );
nand \U$11487 ( \11830 , \11828 , \11829 );
not \U$11488 ( \11831 , \11830 );
not \U$11489 ( \11832 , \11831 );
and \U$11490 ( \11833 , \11073 , \11321 );
not \U$11491 ( \11834 , \11073 );
not \U$11492 ( \11835 , \11321 );
and \U$11493 ( \11836 , \11834 , \11835 );
nor \U$11494 ( \11837 , \11833 , \11836 );
not \U$11495 ( \11838 , \11837 );
or \U$11496 ( \11839 , \11832 , \11838 );
or \U$11497 ( \11840 , \11831 , \11837 );
nand \U$11498 ( \11841 , \11839 , \11840 );
not \U$11499 ( \11842 , \11841 );
xor \U$11500 ( \11843 , \9972 , \9661 );
xnor \U$11501 ( \11844 , \11843 , \10012 );
not \U$11502 ( \11845 , \11844 );
not \U$11503 ( \11846 , \11845 );
not \U$11504 ( \11847 , \9967 );
not \U$11505 ( \11848 , \9795 );
or \U$11506 ( \11849 , \11847 , \11848 );
or \U$11507 ( \11850 , \9967 , \9795 );
nand \U$11508 ( \11851 , \11849 , \11850 );
and \U$11509 ( \11852 , \11310 , \11226 );
not \U$11510 ( \11853 , \11310 );
not \U$11511 ( \11854 , \11226 );
and \U$11512 ( \11855 , \11853 , \11854 );
nor \U$11513 ( \11856 , \11852 , \11855 );
xor \U$11514 ( \11857 , \11851 , \11856 );
xor \U$11515 ( \11858 , \11075 , \11082 );
not \U$11516 ( \11859 , \11097 );
xor \U$11517 ( \11860 , \11858 , \11859 );
and \U$11518 ( \11861 , \11857 , \11860 );
and \U$11519 ( \11862 , \11851 , \11856 );
or \U$11520 ( \11863 , \11861 , \11862 );
not \U$11521 ( \11864 , \11863 );
not \U$11522 ( \11865 , \11864 );
not \U$11523 ( \11866 , \11314 );
xor \U$11524 ( \11867 , \11316 , \11866 );
xnor \U$11525 ( \11868 , \11867 , \11106 );
not \U$11526 ( \11869 , \11868 );
or \U$11527 ( \11870 , \11865 , \11869 );
not \U$11528 ( \11871 , \11863 );
or \U$11529 ( \11872 , \11868 , \11871 );
nand \U$11530 ( \11873 , \11870 , \11872 );
not \U$11531 ( \11874 , \11873 );
or \U$11532 ( \11875 , \11846 , \11874 );
not \U$11533 ( \11876 , \11871 );
nand \U$11534 ( \11877 , \11876 , \11868 );
nand \U$11535 ( \11878 , \11875 , \11877 );
not \U$11536 ( \11879 , \11878 );
or \U$11537 ( \11880 , \11842 , \11879 );
nand \U$11538 ( \11881 , \11830 , \11837 );
nand \U$11539 ( \11882 , \11880 , \11881 );
not \U$11540 ( \11883 , \11882 );
not \U$11541 ( \11884 , \11883 );
and \U$11542 ( \11885 , \11333 , \11884 );
and \U$11543 ( \11886 , \10365 , \11332 );
nor \U$11544 ( \11887 , \11885 , \11886 );
not \U$11545 ( \11888 , \10759 );
not \U$11546 ( \11889 , \11327 );
not \U$11547 ( \11890 , \11889 );
or \U$11548 ( \11891 , \11888 , \11890 );
not \U$11549 ( \11892 , \11064 );
nand \U$11550 ( \11893 , \11892 , \11326 );
nand \U$11551 ( \11894 , \11891 , \11893 );
not \U$11552 ( \11895 , \11894 );
not \U$11553 ( \11896 , \11044 );
not \U$11554 ( \11897 , \11022 );
or \U$11555 ( \11898 , \11896 , \11897 );
not \U$11556 ( \11899 , \11040 );
nand \U$11557 ( \11900 , \11899 , \11036 );
nand \U$11558 ( \11901 , \11898 , \11900 );
and \U$11559 ( \11902 , \11035 , \11026 );
and \U$11560 ( \11903 , \8992 , \11034 );
nor \U$11561 ( \11904 , \11902 , \11903 );
not \U$11562 ( \11905 , \3861 );
not \U$11563 ( \11906 , RI9871aa0_133);
and \U$11564 ( \11907 , \11905 , \11906 );
and \U$11565 ( \11908 , \9461 , RI9871aa0_133);
nor \U$11566 ( \11909 , \11907 , \11908 );
or \U$11567 ( \11910 , \11909 , \2086 );
not \U$11568 ( \11911 , \10937 );
or \U$11569 ( \11912 , \11911 , \2073 );
nand \U$11570 ( \11913 , \11910 , \11912 );
not \U$11571 ( \11914 , \7188 );
not \U$11572 ( \11915 , RI9872568_156);
not \U$11573 ( \11916 , \2216 );
or \U$11574 ( \11917 , \11915 , \11916 );
or \U$11575 ( \11918 , \848 , RI9872568_156);
nand \U$11576 ( \11919 , \11917 , \11918 );
not \U$11577 ( \11920 , \11919 );
or \U$11578 ( \11921 , \11914 , \11920 );
nand \U$11579 ( \11922 , \10895 , \5642 );
nand \U$11580 ( \11923 , \11921 , \11922 );
xor \U$11581 ( \11924 , \11913 , \11923 );
not \U$11582 ( \11925 , \6611 );
not \U$11583 ( \11926 , RI98728b0_163);
not \U$11584 ( \11927 , \893 );
or \U$11585 ( \11928 , \11926 , \11927 );
or \U$11586 ( \11929 , \6443 , RI98728b0_163);
nand \U$11587 ( \11930 , \11928 , \11929 );
not \U$11588 ( \11931 , \11930 );
or \U$11589 ( \11932 , \11925 , \11931 );
nand \U$11590 ( \11933 , \10958 , \6284 );
nand \U$11591 ( \11934 , \11932 , \11933 );
xor \U$11592 ( \11935 , \11924 , \11934 );
xor \U$11593 ( \11936 , \11904 , \11935 );
xor \U$11594 ( \11937 , \10772 , \10778 );
and \U$11595 ( \11938 , \11937 , \10788 );
and \U$11596 ( \11939 , \10772 , \10778 );
nor \U$11597 ( \11940 , \11938 , \11939 );
not \U$11598 ( \11941 , \10575 );
not \U$11599 ( \11942 , \11941 );
not \U$11600 ( \11943 , \10610 );
or \U$11601 ( \11944 , \11942 , \11943 );
nand \U$11602 ( \11945 , \10591 , \10605 );
nand \U$11603 ( \11946 , \11944 , \11945 );
xor \U$11604 ( \11947 , \11940 , \11946 );
not \U$11605 ( \11948 , \10800 );
not \U$11606 ( \11949 , \10821 );
or \U$11607 ( \11950 , \11948 , \11949 );
not \U$11608 ( \11951 , \10814 );
nand \U$11609 ( \11952 , \11951 , \10811 );
nand \U$11610 ( \11953 , \11950 , \11952 );
xnor \U$11611 ( \11954 , \11947 , \11953 );
xnor \U$11612 ( \11955 , \11936 , \11954 );
and \U$11613 ( \11956 , \11901 , \11955 );
not \U$11614 ( \11957 , \11901 );
not \U$11615 ( \11958 , \11955 );
and \U$11616 ( \11959 , \11957 , \11958 );
or \U$11617 ( \11960 , \11956 , \11959 );
not \U$11618 ( \11961 , \10525 );
not \U$11619 ( \11962 , \10443 );
or \U$11620 ( \11963 , \11961 , \11962 );
nand \U$11621 ( \11964 , \10438 , \10429 );
nand \U$11622 ( \11965 , \11963 , \11964 );
not \U$11623 ( \11966 , \11965 );
xor \U$11624 ( \11967 , \11960 , \11966 );
not \U$11625 ( \11968 , \10526 );
not \U$11626 ( \11969 , \10741 );
or \U$11627 ( \11970 , \11968 , \11969 );
nand \U$11628 ( \11971 , \11970 , \10563 );
not \U$11629 ( \11972 , \10526 );
nand \U$11630 ( \11973 , \11972 , \10742 );
nand \U$11631 ( \11974 , \11971 , \11973 );
xor \U$11632 ( \11975 , \11967 , \11974 );
not \U$11633 ( \11976 , \10521 );
not \U$11634 ( \11977 , \11976 );
not \U$11635 ( \11978 , \10473 );
or \U$11636 ( \11979 , \11977 , \11978 );
not \U$11637 ( \11980 , \10517 );
nand \U$11638 ( \11981 , \11980 , \10512 );
nand \U$11639 ( \11982 , \11979 , \11981 );
not \U$11640 ( \11983 , \11982 );
not \U$11641 ( \11984 , \11983 );
not \U$11642 ( \11985 , \10832 );
not \U$11643 ( \11986 , \10827 );
or \U$11644 ( \11987 , \11985 , \11986 );
not \U$11645 ( \11988 , \10790 );
nand \U$11646 ( \11989 , \11988 , \10823 );
nand \U$11647 ( \11990 , \11987 , \11989 );
xor \U$11648 ( \11991 , \10568 , \10614 );
and \U$11649 ( \11992 , \11991 , \10649 );
and \U$11650 ( \11993 , \10568 , \10614 );
or \U$11651 ( \11994 , \11992 , \11993 );
xor \U$11652 ( \11995 , \11990 , \11994 );
not \U$11653 ( \11996 , \11995 );
or \U$11654 ( \11997 , \11984 , \11996 );
or \U$11655 ( \11998 , \11995 , \11983 );
nand \U$11656 ( \11999 , \11997 , \11998 );
not \U$11657 ( \12000 , \10650 );
not \U$11658 ( \12001 , \10740 );
or \U$11659 ( \12002 , \12000 , \12001 );
not \U$11660 ( \12003 , \10650 );
not \U$11661 ( \12004 , \12003 );
not \U$11662 ( \12005 , \10739 );
or \U$11663 ( \12006 , \12004 , \12005 );
nand \U$11664 ( \12007 , \12006 , \10719 );
nand \U$11665 ( \12008 , \12002 , \12007 );
xor \U$11666 ( \12009 , \11999 , \12008 );
not \U$11667 ( \12010 , \10929 );
buf \U$11668 ( \12011 , \10872 );
not \U$11669 ( \12012 , \12011 );
or \U$11670 ( \12013 , \12010 , \12012 );
or \U$11671 ( \12014 , \10929 , \12011 );
nand \U$11672 ( \12015 , \12014 , \10900 );
nand \U$11673 ( \12016 , \12013 , \12015 );
not \U$11674 ( \12017 , \6316 );
xor \U$11675 ( \12018 , \5753 , \8642 );
not \U$11676 ( \12019 , \12018 );
or \U$11677 ( \12020 , \12017 , \12019 );
nand \U$11678 ( \12021 , \10776 , \1162 );
nand \U$11679 ( \12022 , \12020 , \12021 );
not \U$11680 ( \12023 , \1067 );
not \U$11681 ( \12024 , \1044 );
not \U$11682 ( \12025 , \10309 );
or \U$11683 ( \12026 , \12024 , \12025 );
nand \U$11684 ( \12027 , \8597 , \3271 );
nand \U$11685 ( \12028 , \12026 , \12027 );
not \U$11686 ( \12029 , \12028 );
or \U$11687 ( \12030 , \12023 , \12029 );
nand \U$11688 ( \12031 , \10784 , \1018 );
nand \U$11689 ( \12032 , \12030 , \12031 );
xor \U$11690 ( \12033 , \12022 , \12032 );
not \U$11691 ( \12034 , \10251 );
not \U$11692 ( \12035 , \10855 );
or \U$11693 ( \12036 , \12034 , \12035 );
nand \U$11694 ( \12037 , \10242 , RI9872d60_173);
nand \U$11695 ( \12038 , \12036 , \12037 );
xnor \U$11696 ( \12039 , \12033 , \12038 );
not \U$11697 ( \12040 , \12039 );
xor \U$11698 ( \12041 , \10911 , \10921 );
and \U$11699 ( \12042 , \12041 , \10928 );
and \U$11700 ( \12043 , \10911 , \10921 );
or \U$11701 ( \12044 , \12042 , \12043 );
not \U$11702 ( \12045 , \12044 );
or \U$11703 ( \12046 , \12040 , \12045 );
or \U$11704 ( \12047 , \12044 , \12039 );
nand \U$11705 ( \12048 , \12046 , \12047 );
not \U$11706 ( \12049 , \10888 );
not \U$11707 ( \12050 , \10899 );
or \U$11708 ( \12051 , \12049 , \12050 );
xor \U$11709 ( \12052 , \10899 , \10888 );
nand \U$11710 ( \12053 , \12052 , \10882 );
nand \U$11711 ( \12054 , \12051 , \12053 );
not \U$11712 ( \12055 , \12054 );
and \U$11713 ( \12056 , \12048 , \12055 );
not \U$11714 ( \12057 , \12048 );
and \U$11715 ( \12058 , \12057 , \12054 );
nor \U$11716 ( \12059 , \12056 , \12058 );
xor \U$11717 ( \12060 , \12016 , \12059 );
xor \U$11718 ( \12061 , \10999 , \10963 );
not \U$11719 ( \12062 , \10967 );
and \U$11720 ( \12063 , \12061 , \12062 );
and \U$11721 ( \12064 , \10999 , \10963 );
or \U$11722 ( \12065 , \12063 , \12064 );
buf \U$11723 ( \12066 , \12065 );
xnor \U$11724 ( \12067 , \12060 , \12066 );
xor \U$11725 ( \12068 , \12009 , \12067 );
xor \U$11726 ( \12069 , \11975 , \12068 );
not \U$11727 ( \12070 , \12069 );
not \U$11728 ( \12071 , \12070 );
not \U$11729 ( \12072 , \11060 );
not \U$11730 ( \12073 , \12072 );
not \U$11731 ( \12074 , \11005 );
or \U$11732 ( \12075 , \12073 , \12074 );
not \U$11733 ( \12076 , \11001 );
nand \U$11734 ( \12077 , \12076 , \10770 );
nand \U$11735 ( \12078 , \12075 , \12077 );
not \U$11736 ( \12079 , \12078 );
not \U$11737 ( \12080 , \10977 );
not \U$11738 ( \12081 , \10988 );
not \U$11739 ( \12082 , \10998 );
or \U$11740 ( \12083 , \12081 , \12082 );
or \U$11741 ( \12084 , \10998 , \10988 );
nand \U$11742 ( \12085 , \12083 , \12084 );
not \U$11743 ( \12086 , \12085 );
or \U$11744 ( \12087 , \12080 , \12086 );
nand \U$11745 ( \12088 , \10998 , \10987 );
nand \U$11746 ( \12089 , \12087 , \12088 );
not \U$11747 ( \12090 , \12089 );
xor \U$11748 ( \12091 , \10941 , \10949 );
and \U$11749 ( \12092 , \12091 , \10962 );
and \U$11750 ( \12093 , \10941 , \10949 );
or \U$11751 ( \12094 , \12092 , \12093 );
not \U$11752 ( \12095 , \12094 );
not \U$11753 ( \12096 , \9876 );
and \U$11754 ( \12097 , \10412 , RI9872130_147);
not \U$11755 ( \12098 , \10412 );
and \U$11756 ( \12099 , \12098 , \919 );
nor \U$11757 ( \12100 , \12097 , \12099 );
not \U$11758 ( \12101 , \12100 );
or \U$11759 ( \12102 , \12096 , \12101 );
nand \U$11760 ( \12103 , \10589 , \876 );
nand \U$11761 ( \12104 , \12102 , \12103 );
not \U$11762 ( \12105 , \859 );
not \U$11763 ( \12106 , \10573 );
or \U$11764 ( \12107 , \12105 , \12106 );
not \U$11765 ( \12108 , RI9871d70_139);
not \U$11766 ( \12109 , \12108 );
not \U$11767 ( \12110 , \7467 );
or \U$11768 ( \12111 , \12109 , \12110 );
nand \U$11769 ( \12112 , \10401 , RI9871d70_139);
nand \U$11770 ( \12113 , \12111 , \12112 );
nand \U$11771 ( \12114 , \12113 , \832 );
nand \U$11772 ( \12115 , \12107 , \12114 );
and \U$11773 ( \12116 , \12104 , \12115 );
not \U$11774 ( \12117 , \12104 );
not \U$11775 ( \12118 , \12115 );
and \U$11776 ( \12119 , \12117 , \12118 );
nor \U$11777 ( \12120 , \12116 , \12119 );
buf \U$11778 ( \12121 , \12120 );
not \U$11779 ( \12122 , \1353 );
not \U$11780 ( \12123 , \1367 );
not \U$11781 ( \12124 , \9599 );
not \U$11782 ( \12125 , \12124 );
or \U$11783 ( \12126 , \12123 , \12125 );
nand \U$11784 ( \12127 , \8074 , RI9871e60_141);
nand \U$11785 ( \12128 , \12126 , \12127 );
not \U$11786 ( \12129 , \12128 );
or \U$11787 ( \12130 , \12122 , \12129 );
not \U$11788 ( \12131 , \10603 );
or \U$11789 ( \12132 , \12131 , \5078 );
nand \U$11790 ( \12133 , \12130 , \12132 );
xnor \U$11791 ( \12134 , \12121 , \12133 );
not \U$11792 ( \12135 , \12134 );
and \U$11793 ( \12136 , \12095 , \12135 );
and \U$11794 ( \12137 , \12094 , \12134 );
nor \U$11795 ( \12138 , \12136 , \12137 );
not \U$11796 ( \12139 , \12138 );
and \U$11797 ( \12140 , \12090 , \12139 );
and \U$11798 ( \12141 , \12089 , \12138 );
nor \U$11799 ( \12142 , \12140 , \12141 );
not \U$11800 ( \12143 , \12142 );
not \U$11801 ( \12144 , \1136 );
not \U$11802 ( \12145 , \5206 );
xor \U$11803 ( \12146 , RI98718c0_129, \12145 );
not \U$11804 ( \12147 , \12146 );
or \U$11805 ( \12148 , \12144 , \12147 );
nand \U$11806 ( \12149 , \10886 , \1083 );
nand \U$11807 ( \12150 , \12148 , \12149 );
not \U$11808 ( \12151 , \12150 );
not \U$11809 ( \12152 , \12151 );
not \U$11810 ( \12153 , \1518 );
not \U$11811 ( \12154 , \6305 );
not \U$11812 ( \12155 , \12154 );
not \U$11813 ( \12156 , RI9871c80_137);
and \U$11814 ( \12157 , \12155 , \12156 );
not \U$11815 ( \12158 , \5707 );
and \U$11816 ( \12159 , \12158 , RI9871c80_137);
nor \U$11817 ( \12160 , \12157 , \12159 );
not \U$11818 ( \12161 , \12160 );
or \U$11819 ( \12162 , \12153 , \12161 );
nand \U$11820 ( \12163 , \10809 , \1501 );
nand \U$11821 ( \12164 , \12162 , \12163 );
not \U$11822 ( \12165 , \12164 );
not \U$11823 ( \12166 , \12165 );
or \U$11824 ( \12167 , \12152 , \12166 );
nand \U$11825 ( \12168 , \12150 , \12164 );
nand \U$11826 ( \12169 , \12167 , \12168 );
not \U$11827 ( \12170 , \793 );
not \U$11828 ( \12171 , \11030 );
or \U$11829 ( \12172 , \12170 , \12171 );
and \U$11830 ( \12173 , \10699 , \1078 );
not \U$11831 ( \12174 , \10699 );
and \U$11832 ( \12175 , \12174 , RI98719b0_131);
nor \U$11833 ( \12176 , \12173 , \12175 );
nand \U$11834 ( \12177 , \12176 , \6145 );
nand \U$11835 ( \12178 , \12172 , \12177 );
and \U$11836 ( \12179 , \12169 , \12178 );
not \U$11837 ( \12180 , \12169 );
not \U$11838 ( \12181 , \12178 );
and \U$11839 ( \12182 , \12180 , \12181 );
nor \U$11840 ( \12183 , \12179 , \12182 );
not \U$11841 ( \12184 , \10867 );
not \U$11842 ( \12185 , \10858 );
or \U$11843 ( \12186 , \12184 , \12185 );
nand \U$11844 ( \12187 , \10857 , \10847 );
nand \U$11845 ( \12188 , \12186 , \12187 );
not \U$11846 ( \12189 , \12188 );
xor \U$11847 ( \12190 , \12183 , \12189 );
not \U$11848 ( \12191 , \4085 );
and \U$11849 ( \12192 , RI98725e0_157, \1039 );
not \U$11850 ( \12193 , RI98725e0_157);
and \U$11851 ( \12194 , \12193 , \6330 );
nor \U$11852 ( \12195 , \12192 , \12194 );
not \U$11853 ( \12196 , \12195 );
or \U$11854 ( \12197 , \12191 , \12196 );
nand \U$11855 ( \12198 , \4103 , \10926 );
nand \U$11856 ( \12199 , \12197 , \12198 );
not \U$11857 ( \12200 , \9072 );
not \U$11858 ( \12201 , RI9872a18_166);
not \U$11859 ( \12202 , \2492 );
or \U$11860 ( \12203 , \12201 , \12202 );
or \U$11861 ( \12204 , \2492 , RI9872a18_166);
nand \U$11862 ( \12205 , \12203 , \12204 );
not \U$11863 ( \12206 , \12205 );
or \U$11864 ( \12207 , \12200 , \12206 );
nand \U$11865 ( \12208 , \10919 , \9079 );
nand \U$11866 ( \12209 , \12207 , \12208 );
not \U$11867 ( \12210 , \12209 );
not \U$11868 ( \12211 , \7338 );
and \U$11869 ( \12212 , RI98729a0_165, \7064 );
not \U$11870 ( \12213 , RI98729a0_165);
and \U$11871 ( \12214 , \12213 , \1582 );
or \U$11872 ( \12215 , \12212 , \12214 );
not \U$11873 ( \12216 , \12215 );
or \U$11874 ( \12217 , \12211 , \12216 );
nand \U$11875 ( \12218 , \10996 , \7326 );
nand \U$11876 ( \12219 , \12217 , \12218 );
not \U$11877 ( \12220 , \12219 );
not \U$11878 ( \12221 , \12220 );
or \U$11879 ( \12222 , \12210 , \12221 );
or \U$11880 ( \12223 , \12209 , \12220 );
nand \U$11881 ( \12224 , \12222 , \12223 );
xor \U$11882 ( \12225 , \12199 , \12224 );
xnor \U$11883 ( \12226 , \12190 , \12225 );
not \U$11884 ( \12227 , \12226 );
or \U$11885 ( \12228 , \12143 , \12227 );
or \U$11886 ( \12229 , \12226 , \12142 );
nand \U$11887 ( \12230 , \12228 , \12229 );
not \U$11888 ( \12231 , \5034 );
not \U$11889 ( \12232 , \10845 );
or \U$11890 ( \12233 , \12231 , \12232 );
not \U$11891 ( \12234 , RI9872478_154);
not \U$11892 ( \12235 , \7019 );
or \U$11893 ( \12236 , \12234 , \12235 );
or \U$11894 ( \12237 , \7019 , RI9872478_154);
nand \U$11895 ( \12238 , \12236 , \12237 );
nand \U$11896 ( \12239 , \12238 , \5796 );
nand \U$11897 ( \12240 , \12233 , \12239 );
nand \U$11898 ( \12241 , \10372 , \1165 );
xor \U$11899 ( \12242 , \12240 , \12241 );
not \U$11900 ( \12243 , \1430 );
and \U$11901 ( \12244 , RI9871c08_136, \10639 );
not \U$11902 ( \12245 , RI9871c08_136);
and \U$11903 ( \12246 , \12245 , \4990 );
nor \U$11904 ( \12247 , \12244 , \12246 );
not \U$11905 ( \12248 , \12247 );
or \U$11906 ( \12249 , \12243 , \12248 );
or \U$11907 ( \12250 , \10877 , \5411 );
nand \U$11908 ( \12251 , \12249 , \12250 );
xor \U$11909 ( \12252 , \12242 , \12251 );
not \U$11910 ( \12253 , \12252 );
not \U$11911 ( \12254 , \3170 );
and \U$11912 ( \12255 , RI9872310_151, \2111 );
not \U$11913 ( \12256 , RI9872310_151);
and \U$11914 ( \12257 , \12256 , \7164 );
nor \U$11915 ( \12258 , \12255 , \12257 );
not \U$11916 ( \12259 , \12258 );
or \U$11917 ( \12260 , \12254 , \12259 );
nand \U$11918 ( \12261 , \10943 , \3163 );
nand \U$11919 ( \12262 , \12260 , \12261 );
not \U$11920 ( \12263 , \10679 );
not \U$11921 ( \12264 , \10863 );
or \U$11922 ( \12265 , \12263 , \12264 );
and \U$11923 ( \12266 , RI9872b80_169, \1097 );
not \U$11924 ( \12267 , RI9872b80_169);
and \U$11925 ( \12268 , \12267 , \1106 );
or \U$11926 ( \12269 , \12266 , \12268 );
nand \U$11927 ( \12270 , \12269 , \9214 );
nand \U$11928 ( \12271 , \12265 , \12270 );
xor \U$11929 ( \12272 , \12262 , \12271 );
not \U$11930 ( \12273 , \3467 );
and \U$11931 ( \12274 , \1191 , \3593 );
not \U$11932 ( \12275 , \1191 );
and \U$11933 ( \12276 , \12275 , RI98726d0_159);
nor \U$11934 ( \12277 , \12274 , \12276 );
not \U$11935 ( \12278 , \12277 );
or \U$11936 ( \12279 , \12273 , \12278 );
nand \U$11937 ( \12280 , \10975 , \3600 );
nand \U$11938 ( \12281 , \12279 , \12280 );
xor \U$11939 ( \12282 , \12272 , \12281 );
not \U$11940 ( \12283 , \12282 );
or \U$11941 ( \12284 , \12253 , \12283 );
or \U$11942 ( \12285 , \12282 , \12252 );
nand \U$11943 ( \12286 , \12284 , \12285 );
and \U$11944 ( \12287 , RI9871b18_134, \5776 );
not \U$11945 ( \12288 , RI9871b18_134);
and \U$11946 ( \12289 , \12288 , \6185 );
nor \U$11947 ( \12290 , \12287 , \12289 );
or \U$11948 ( \12291 , \12290 , \1543 );
or \U$11949 ( \12292 , \1293 , \10798 );
nand \U$11950 ( \12293 , \12291 , \12292 );
not \U$11951 ( \12294 , \5048 );
not \U$11952 ( \12295 , \1365 );
and \U$11953 ( \12296 , RI9872388_152, \12295 );
not \U$11954 ( \12297 , RI9872388_152);
and \U$11955 ( \12298 , \12297 , \4454 );
or \U$11956 ( \12299 , \12296 , \12298 );
not \U$11957 ( \12300 , \12299 );
or \U$11958 ( \12301 , \12294 , \12300 );
nand \U$11959 ( \12302 , \10909 , \6553 );
nand \U$11960 ( \12303 , \12301 , \12302 );
xor \U$11961 ( \12304 , \12293 , \12303 );
not \U$11962 ( \12305 , \9670 );
not \U$11963 ( \12306 , \10983 );
or \U$11964 ( \12307 , \12305 , \12306 );
not \U$11965 ( \12308 , \9185 );
not \U$11966 ( \12309 , \1393 );
or \U$11967 ( \12310 , \12308 , \12309 );
or \U$11968 ( \12311 , \2982 , \9185 );
nand \U$11969 ( \12312 , \12310 , \12311 );
nand \U$11970 ( \12313 , \12312 , \9668 );
nand \U$11971 ( \12314 , \12307 , \12313 );
xor \U$11972 ( \12315 , \12304 , \12314 );
xor \U$11973 ( \12316 , \12286 , \12315 );
not \U$11974 ( \12317 , \12316 );
and \U$11975 ( \12318 , \12230 , \12317 );
not \U$11976 ( \12319 , \12230 );
and \U$11977 ( \12320 , \12319 , \12316 );
nor \U$11978 ( \12321 , \12318 , \12320 );
not \U$11979 ( \12322 , \12321 );
not \U$11980 ( \12323 , \12322 );
xor \U$11981 ( \12324 , \10837 , \10930 );
and \U$11982 ( \12325 , \12324 , \11000 );
and \U$11983 ( \12326 , \10837 , \10930 );
or \U$11984 ( \12327 , \12325 , \12326 );
not \U$11985 ( \12328 , \12327 );
or \U$11986 ( \12329 , \12323 , \12328 );
not \U$11987 ( \12330 , \12327 );
nand \U$11988 ( \12331 , \12330 , \12321 );
nand \U$11989 ( \12332 , \12329 , \12331 );
not \U$11990 ( \12333 , \11055 );
not \U$11991 ( \12334 , \11017 );
or \U$11992 ( \12335 , \12333 , \12334 );
not \U$11993 ( \12336 , \11051 );
nand \U$11994 ( \12337 , \12336 , \11045 );
nand \U$11995 ( \12338 , \12335 , \12337 );
not \U$11996 ( \12339 , \12338 );
and \U$11997 ( \12340 , \12332 , \12339 );
not \U$11998 ( \12341 , \12332 );
and \U$11999 ( \12342 , \12341 , \12338 );
nor \U$12000 ( \12343 , \12340 , \12342 );
not \U$12001 ( \12344 , \12343 );
and \U$12002 ( \12345 , \12079 , \12344 );
and \U$12003 ( \12346 , \12078 , \12343 );
nor \U$12004 ( \12347 , \12345 , \12346 );
not \U$12005 ( \12348 , \10743 );
not \U$12006 ( \12349 , \10758 );
or \U$12007 ( \12350 , \12348 , \12349 );
nand \U$12008 ( \12351 , \10747 , \10753 );
nand \U$12009 ( \12352 , \12350 , \12351 );
and \U$12010 ( \12353 , \12347 , \12352 );
not \U$12011 ( \12354 , \12347 );
not \U$12012 ( \12355 , \12352 );
and \U$12013 ( \12356 , \12354 , \12355 );
nor \U$12014 ( \12357 , \12353 , \12356 );
not \U$12015 ( \12358 , \12357 );
not \U$12016 ( \12359 , \12358 );
or \U$12017 ( \12360 , \12071 , \12359 );
nand \U$12018 ( \12361 , \12357 , \12069 );
nand \U$12019 ( \12362 , \12360 , \12361 );
not \U$12020 ( \12363 , \12362 );
or \U$12021 ( \12364 , \11895 , \12363 );
or \U$12022 ( \12365 , \12362 , \11894 );
nand \U$12023 ( \12366 , \12364 , \12365 );
nand \U$12024 ( \12367 , \11887 , \12366 );
xor \U$12025 ( \12368 , \9655 , \10360 );
xnor \U$12026 ( \12369 , \12368 , \10014 );
and \U$12027 ( \12370 , \11664 , \11667 );
not \U$12028 ( \12371 , \11664 );
and \U$12029 ( \12372 , \12371 , \11668 );
nor \U$12030 ( \12373 , \12370 , \12372 );
xor \U$12031 ( \12374 , \11817 , \12373 );
xor \U$12032 ( \12375 , \11391 , \11400 );
xor \U$12033 ( \12376 , \12375 , \11412 );
not \U$12034 ( \12377 , \7338 );
not \U$12035 ( \12378 , \11571 );
or \U$12036 ( \12379 , \12377 , \12378 );
not \U$12037 ( \12380 , \7333 );
not \U$12038 ( \12381 , \1062 );
or \U$12039 ( \12382 , \12380 , \12381 );
or \U$12040 ( \12383 , \1061 , \7333 );
nand \U$12041 ( \12384 , \12382 , \12383 );
nand \U$12042 ( \12385 , \7325 , \12384 );
nand \U$12043 ( \12386 , \12379 , \12385 );
not \U$12044 ( \12387 , \6610 );
not \U$12045 ( \12388 , \11748 );
or \U$12046 ( \12389 , \12387 , \12388 );
not \U$12047 ( \12390 , RI98728b0_163);
not \U$12048 ( \12391 , \1210 );
or \U$12049 ( \12392 , \12390 , \12391 );
not \U$12050 ( \12393 , \11114 );
or \U$12051 ( \12394 , \12393 , RI98728b0_163);
nand \U$12052 ( \12395 , \12392 , \12394 );
nand \U$12053 ( \12396 , \12395 , \6284 );
nand \U$12054 ( \12397 , \12389 , \12396 );
xor \U$12055 ( \12398 , \12386 , \12397 );
not \U$12056 ( \12399 , \10333 );
not \U$12057 ( \12400 , \11590 );
or \U$12058 ( \12401 , \12399 , \12400 );
xnor \U$12059 ( \12402 , RI9872e50_175, \1307 );
not \U$12060 ( \12403 , \12402 );
not \U$12061 ( \12404 , \9294 );
or \U$12062 ( \12405 , \12403 , \12404 );
nand \U$12063 ( \12406 , \12401 , \12405 );
and \U$12064 ( \12407 , \12398 , \12406 );
and \U$12065 ( \12408 , \12386 , \12397 );
or \U$12066 ( \12409 , \12407 , \12408 );
xor \U$12067 ( \12410 , \12376 , \12409 );
not \U$12068 ( \12411 , \12410 );
not \U$12069 ( \12412 , \9527 );
and \U$12070 ( \12413 , \6174 , \8732 );
not \U$12071 ( \12414 , \6174 );
and \U$12072 ( \12415 , \12414 , RI9872f40_177);
nor \U$12073 ( \12416 , \12413 , \12415 );
not \U$12074 ( \12417 , \12416 );
or \U$12075 ( \12418 , \12412 , \12417 );
nand \U$12076 ( \12419 , \11720 , \8752 );
nand \U$12077 ( \12420 , \12418 , \12419 );
not \U$12078 ( \12421 , \12420 );
not \U$12079 ( \12422 , \10624 );
not \U$12080 ( \12423 , \11769 );
or \U$12081 ( \12424 , \12422 , \12423 );
not \U$12082 ( \12425 , RI9872d60_173);
not \U$12083 ( \12426 , \915 );
or \U$12084 ( \12427 , \12425 , \12426 );
or \U$12085 ( \12428 , \916 , RI9872d60_173);
nand \U$12086 ( \12429 , \12427 , \12428 );
nand \U$12087 ( \12430 , \12429 , \10251 );
nand \U$12088 ( \12431 , \12424 , \12430 );
not \U$12089 ( \12432 , \12431 );
not \U$12090 ( \12433 , \12432 );
not \U$12091 ( \12434 , \5653 );
not \U$12092 ( \12435 , \11756 );
or \U$12093 ( \12436 , \12434 , \12435 );
not \U$12094 ( \12437 , RI9872568_156);
not \U$12095 ( \12438 , \1485 );
or \U$12096 ( \12439 , \12437 , \12438 );
or \U$12097 ( \12440 , \1485 , RI9872568_156);
nand \U$12098 ( \12441 , \12439 , \12440 );
nand \U$12099 ( \12442 , \5642 , \12441 );
nand \U$12100 ( \12443 , \12436 , \12442 );
not \U$12101 ( \12444 , \12443 );
or \U$12102 ( \12445 , \12433 , \12444 );
or \U$12103 ( \12446 , \12443 , \12432 );
nand \U$12104 ( \12447 , \12445 , \12446 );
not \U$12105 ( \12448 , \12447 );
or \U$12106 ( \12449 , \12421 , \12448 );
nand \U$12107 ( \12450 , \12443 , \12431 );
nand \U$12108 ( \12451 , \12449 , \12450 );
not \U$12109 ( \12452 , \12451 );
or \U$12110 ( \12453 , \12411 , \12452 );
nand \U$12111 ( \12454 , \12409 , \12376 );
nand \U$12112 ( \12455 , \12453 , \12454 );
not \U$12113 ( \12456 , \1352 );
not \U$12114 ( \12457 , \11387 );
or \U$12115 ( \12458 , \12456 , \12457 );
not \U$12116 ( \12459 , RI9871e60_141);
buf \U$12117 ( \12460 , \9847 );
not \U$12118 ( \12461 , \12460 );
or \U$12119 ( \12462 , \12459 , \12461 );
or \U$12120 ( \12463 , \9849 , RI9871e60_141);
nand \U$12121 ( \12464 , \12462 , \12463 );
nand \U$12122 ( \12465 , \12464 , \1380 );
nand \U$12123 ( \12466 , \12458 , \12465 );
not \U$12124 ( \12467 , \832 );
not \U$12125 ( \12468 , \11396 );
or \U$12126 ( \12469 , \12467 , \12468 );
buf \U$12127 ( \12470 , \8722 );
not \U$12128 ( \12471 , \12470 );
and \U$12129 ( \12472 , RI9871d70_139, \12471 );
not \U$12130 ( \12473 , RI9871d70_139);
and \U$12131 ( \12474 , \12473 , \8722 );
or \U$12132 ( \12475 , \12472 , \12474 );
nand \U$12133 ( \12476 , \12475 , \5350 );
nand \U$12134 ( \12477 , \12469 , \12476 );
xor \U$12135 ( \12478 , \12466 , \12477 );
not \U$12136 ( \12479 , \12478 );
not \U$12137 ( \12480 , \9079 );
not \U$12138 ( \12481 , RI9872a18_166);
not \U$12139 ( \12482 , \1340 );
or \U$12140 ( \12483 , \12481 , \12482 );
or \U$12141 ( \12484 , \1340 , RI9872a18_166);
nand \U$12142 ( \12485 , \12483 , \12484 );
not \U$12143 ( \12486 , \12485 );
or \U$12144 ( \12487 , \12480 , \12486 );
nand \U$12145 ( \12488 , \11560 , \8041 );
nand \U$12146 ( \12489 , \12487 , \12488 );
not \U$12147 ( \12490 , \12489 );
or \U$12148 ( \12491 , \12479 , \12490 );
nand \U$12149 ( \12492 , \12477 , \12466 );
nand \U$12150 ( \12493 , \12491 , \12492 );
not \U$12151 ( \12494 , \12493 );
not \U$12152 ( \12495 , \12494 );
not \U$12153 ( \12496 , \2087 );
not \U$12154 ( \12497 , \11542 );
or \U$12155 ( \12498 , \12496 , \12497 );
not \U$12156 ( \12499 , RI9871aa0_133);
not \U$12157 ( \12500 , \5761 );
or \U$12158 ( \12501 , \12499 , \12500 );
or \U$12159 ( \12502 , \6059 , RI9871aa0_133);
nand \U$12160 ( \12503 , \12501 , \12502 );
nand \U$12161 ( \12504 , \12503 , \2071 );
nand \U$12162 ( \12505 , \12498 , \12504 );
not \U$12163 ( \12506 , \12505 );
buf \U$12164 ( \12507 , \9951 );
not \U$12165 ( \12508 , \12507 );
xor \U$12166 ( \12509 , RI9873030_179, \11194 );
not \U$12167 ( \12510 , \12509 );
or \U$12168 ( \12511 , \12508 , \12510 );
nand \U$12169 ( \12512 , \11577 , \9937 );
nand \U$12170 ( \12513 , \12511 , \12512 );
buf \U$12171 ( \12514 , \3169 );
not \U$12172 ( \12515 , \12514 );
not \U$12173 ( \12516 , \11552 );
or \U$12174 ( \12517 , \12515 , \12516 );
and \U$12175 ( \12518 , \3154 , \5736 );
not \U$12176 ( \12519 , \3154 );
and \U$12177 ( \12520 , \12519 , \9374 );
nor \U$12178 ( \12521 , \12518 , \12520 );
nand \U$12179 ( \12522 , \6653 , \12521 );
nand \U$12180 ( \12523 , \12517 , \12522 );
and \U$12181 ( \12524 , \12513 , \12523 );
not \U$12182 ( \12525 , \12513 );
not \U$12183 ( \12526 , \12523 );
and \U$12184 ( \12527 , \12525 , \12526 );
nor \U$12185 ( \12528 , \12524 , \12527 );
not \U$12186 ( \12529 , \12528 );
or \U$12187 ( \12530 , \12506 , \12529 );
nand \U$12188 ( \12531 , \12513 , \12523 );
nand \U$12189 ( \12532 , \12530 , \12531 );
not \U$12190 ( \12533 , \12532 );
or \U$12191 ( \12534 , \12495 , \12533 );
or \U$12192 ( \12535 , \12532 , \12494 );
nand \U$12193 ( \12536 , \12534 , \12535 );
not \U$12194 ( \12537 , \12536 );
not \U$12195 ( \12538 , \5048 );
not \U$12196 ( \12539 , \11697 );
or \U$12197 ( \12540 , \12538 , \12539 );
and \U$12198 ( \12541 , RI9872388_152, \3537 );
not \U$12199 ( \12542 , RI9872388_152);
not \U$12200 ( \12543 , \3536 );
and \U$12201 ( \12544 , \12542 , \12543 );
nor \U$12202 ( \12545 , \12541 , \12544 );
nand \U$12203 ( \12546 , \12545 , \4919 );
nand \U$12204 ( \12547 , \12540 , \12546 );
not \U$12205 ( \12548 , \12547 );
not \U$12206 ( \12549 , RI9872478_154);
not \U$12207 ( \12550 , \2947 );
or \U$12208 ( \12551 , \12549 , \12550 );
or \U$12209 ( \12552 , \2947 , RI9872478_154);
nand \U$12210 ( \12553 , \12551 , \12552 );
not \U$12211 ( \12554 , \12553 );
not \U$12212 ( \12555 , \12554 );
not \U$12213 ( \12556 , \7591 );
and \U$12214 ( \12557 , \12555 , \12556 );
and \U$12215 ( \12558 , \11708 , \6698 );
nor \U$12216 ( \12559 , \12557 , \12558 );
not \U$12217 ( \12560 , \12559 );
not \U$12218 ( \12561 , \9668 );
not \U$12219 ( \12562 , \11736 );
or \U$12220 ( \12563 , \12561 , \12562 );
xnor \U$12221 ( \12564 , \820 , RI9872bf8_170);
nand \U$12222 ( \12565 , \12564 , \9670 );
nand \U$12223 ( \12566 , \12563 , \12565 );
not \U$12224 ( \12567 , \12566 );
or \U$12225 ( \12568 , \12560 , \12567 );
or \U$12226 ( \12569 , \12566 , \12559 );
nand \U$12227 ( \12570 , \12568 , \12569 );
not \U$12228 ( \12571 , \12570 );
or \U$12229 ( \12572 , \12548 , \12571 );
not \U$12230 ( \12573 , \12559 );
nand \U$12231 ( \12574 , \12573 , \12566 );
nand \U$12232 ( \12575 , \12572 , \12574 );
not \U$12233 ( \12576 , \12575 );
or \U$12234 ( \12577 , \12537 , \12576 );
not \U$12235 ( \12578 , \12494 );
nand \U$12236 ( \12579 , \12578 , \12532 );
nand \U$12237 ( \12580 , \12577 , \12579 );
or \U$12238 ( \12581 , \12455 , \12580 );
not \U$12239 ( \12582 , \11613 );
and \U$12240 ( \12583 , \11638 , \12582 );
not \U$12241 ( \12584 , \11638 );
and \U$12242 ( \12585 , \12584 , \11613 );
nor \U$12243 ( \12586 , \12583 , \12585 );
not \U$12244 ( \12587 , \12586 );
not \U$12245 ( \12588 , \12587 );
not \U$12246 ( \12589 , \1013 );
not \U$12247 ( \12590 , \11373 );
or \U$12248 ( \12591 , \12589 , \12590 );
not \U$12249 ( \12592 , \1042 );
not \U$12250 ( \12593 , \12592 );
buf \U$12251 ( \12594 , \9138 );
not \U$12252 ( \12595 , \12594 );
or \U$12253 ( \12596 , \12593 , \12595 );
not \U$12254 ( \12597 , \9138 );
nand \U$12255 ( \12598 , \12597 , \8085 );
nand \U$12256 ( \12599 , \12596 , \12598 );
nand \U$12257 ( \12600 , \12599 , \1018 );
nand \U$12258 ( \12601 , \12591 , \12600 );
not \U$12259 ( \12602 , \12601 );
not \U$12260 ( \12603 , \9214 );
not \U$12261 ( \12604 , \11690 );
or \U$12262 ( \12605 , \12603 , \12604 );
not \U$12263 ( \12606 , \9198 );
not \U$12264 ( \12607 , \943 );
or \U$12265 ( \12608 , \12606 , \12607 );
or \U$12266 ( \12609 , \11283 , \9198 );
nand \U$12267 ( \12610 , \12608 , \12609 );
nand \U$12268 ( \12611 , \12610 , \10679 );
nand \U$12269 ( \12612 , \12605 , \12611 );
xor \U$12270 ( \12613 , \12602 , \12612 );
not \U$12271 ( \12614 , \5530 );
not \U$12272 ( \12615 , RI98725e0_157);
not \U$12273 ( \12616 , \5594 );
not \U$12274 ( \12617 , \12616 );
or \U$12275 ( \12618 , \12615 , \12617 );
or \U$12276 ( \12619 , \11028 , RI98725e0_157);
nand \U$12277 ( \12620 , \12618 , \12619 );
not \U$12278 ( \12621 , \12620 );
or \U$12279 ( \12622 , \12614 , \12621 );
nand \U$12280 ( \12623 , \11676 , \5847 );
nand \U$12281 ( \12624 , \12622 , \12623 );
and \U$12282 ( \12625 , \12613 , \12624 );
and \U$12283 ( \12626 , \12602 , \12612 );
nor \U$12284 ( \12627 , \12625 , \12626 );
xor \U$12285 ( \12628 , \11456 , \11445 );
xor \U$12286 ( \12629 , \12628 , \11430 );
not \U$12287 ( \12630 , \12629 );
and \U$12288 ( \12631 , \12627 , \12630 );
not \U$12289 ( \12632 , \12627 );
and \U$12290 ( \12633 , \12632 , \12629 );
nor \U$12291 ( \12634 , \12631 , \12633 );
not \U$12292 ( \12635 , \12634 );
or \U$12293 ( \12636 , \12588 , \12635 );
not \U$12294 ( \12637 , \12627 );
nand \U$12295 ( \12638 , \12637 , \12629 );
nand \U$12296 ( \12639 , \12636 , \12638 );
nand \U$12297 ( \12640 , \12581 , \12639 );
nand \U$12298 ( \12641 , \12580 , \12455 );
nand \U$12299 ( \12642 , \12640 , \12641 );
not \U$12300 ( \12643 , \12642 );
xor \U$12301 ( \12644 , \11334 , \11471 );
xor \U$12302 ( \12645 , \11092 , \11090 );
xnor \U$12303 ( \12646 , \12645 , \11086 );
xnor \U$12304 ( \12647 , \12644 , \12646 );
not \U$12305 ( \12648 , \12647 );
or \U$12306 ( \12649 , \12643 , \12648 );
xor \U$12307 ( \12650 , \11334 , \11472 );
nand \U$12308 ( \12651 , \12650 , \12646 );
nand \U$12309 ( \12652 , \12649 , \12651 );
xor \U$12310 ( \12653 , \12374 , \12652 );
xor \U$12311 ( \12654 , \11791 , \11810 );
xnor \U$12312 ( \12655 , \12654 , \11808 );
not \U$12313 ( \12656 , \12655 );
not \U$12314 ( \12657 , \12656 );
not \U$12315 ( \12658 , \11565 );
not \U$12316 ( \12659 , \12658 );
not \U$12317 ( \12660 , \11645 );
or \U$12318 ( \12661 , \12659 , \12660 );
nand \U$12319 ( \12662 , \11644 , \11565 );
nand \U$12320 ( \12663 , \12661 , \12662 );
not \U$12321 ( \12664 , \12663 );
or \U$12322 ( \12665 , \12657 , \12664 );
or \U$12323 ( \12666 , \12663 , \12656 );
nand \U$12324 ( \12667 , \12665 , \12666 );
not \U$12325 ( \12668 , \12667 );
and \U$12326 ( \12669 , \11760 , \11752 );
not \U$12327 ( \12670 , \11760 );
not \U$12328 ( \12671 , \11752 );
and \U$12329 ( \12672 , \12670 , \12671 );
nor \U$12330 ( \12673 , \12669 , \12672 );
not \U$12331 ( \12674 , \11773 );
and \U$12332 ( \12675 , \12673 , \12674 );
not \U$12333 ( \12676 , \12673 );
and \U$12334 ( \12677 , \12676 , \11773 );
nor \U$12335 ( \12678 , \12675 , \12677 );
not \U$12336 ( \12679 , \12678 );
xor \U$12337 ( \12680 , \11544 , \11554 );
xnor \U$12338 ( \12681 , \12680 , \11562 );
not \U$12339 ( \12682 , \12681 );
not \U$12340 ( \12683 , \11740 );
not \U$12341 ( \12684 , \11729 );
or \U$12342 ( \12685 , \12683 , \12684 );
or \U$12343 ( \12686 , \11729 , \11740 );
nand \U$12344 ( \12687 , \12685 , \12686 );
not \U$12345 ( \12688 , \12687 );
or \U$12346 ( \12689 , \12682 , \12688 );
or \U$12347 ( \12690 , \12681 , \12687 );
nand \U$12348 ( \12691 , \12689 , \12690 );
nand \U$12349 ( \12692 , \12679 , \12691 );
not \U$12350 ( \12693 , \12681 );
nand \U$12351 ( \12694 , \12693 , \12687 );
nand \U$12352 ( \12695 , \12692 , \12694 );
not \U$12353 ( \12696 , \12695 );
or \U$12354 ( \12697 , \12668 , \12696 );
not \U$12355 ( \12698 , \12656 );
nand \U$12356 ( \12699 , \12698 , \12663 );
nand \U$12357 ( \12700 , \12697 , \12699 );
not \U$12358 ( \12701 , \12700 );
not \U$12359 ( \12702 , \11419 );
not \U$12360 ( \12703 , \12702 );
not \U$12361 ( \12704 , \11465 );
or \U$12362 ( \12705 , \12703 , \12704 );
or \U$12363 ( \12706 , \11465 , \12702 );
nand \U$12364 ( \12707 , \12705 , \12706 );
not \U$12365 ( \12708 , \12707 );
not \U$12366 ( \12709 , \1323 );
not \U$12367 ( \12710 , \11633 );
or \U$12368 ( \12711 , \12709 , \12710 );
not \U$12369 ( \12712 , \8877 );
not \U$12370 ( \12713 , \12712 );
and \U$12371 ( \12714 , RI9871b18_134, \12713 );
not \U$12372 ( \12715 , RI9871b18_134);
not \U$12373 ( \12716 , \8877 );
buf \U$12374 ( \12717 , \12716 );
and \U$12375 ( \12718 , \12715 , \12717 );
nor \U$12376 ( \12719 , \12714 , \12718 );
buf \U$12377 ( \12720 , \1292 );
nand \U$12378 ( \12721 , \12719 , \12720 );
nand \U$12379 ( \12722 , \12711 , \12721 );
not \U$12380 ( \12723 , \1429 );
not \U$12381 ( \12724 , \11609 );
or \U$12382 ( \12725 , \12723 , \12724 );
not \U$12383 ( \12726 , \3487 );
not \U$12384 ( \12727 , \8333 );
not \U$12385 ( \12728 , \12727 );
or \U$12386 ( \12729 , \12726 , \12728 );
nand \U$12387 ( \12730 , \8334 , RI9871c08_136);
nand \U$12388 ( \12731 , \12729 , \12730 );
nand \U$12389 ( \12732 , \12731 , \1455 );
nand \U$12390 ( \12733 , \12725 , \12732 );
xor \U$12391 ( \12734 , \12722 , \12733 );
not \U$12392 ( \12735 , \6673 );
not \U$12393 ( \12736 , \11426 );
or \U$12394 ( \12737 , \12735 , \12736 );
not \U$12395 ( \12738 , \1111 );
not \U$12396 ( \12739 , \8944 );
or \U$12397 ( \12740 , \12738 , \12739 );
nand \U$12398 ( \12741 , \8943 , RI98718c0_129);
nand \U$12399 ( \12742 , \12740 , \12741 );
nand \U$12400 ( \12743 , \12742 , \1083 );
nand \U$12401 ( \12744 , \12737 , \12743 );
and \U$12402 ( \12745 , \12734 , \12744 );
and \U$12403 ( \12746 , \12722 , \12733 );
or \U$12404 ( \12747 , \12745 , \12746 );
not \U$12405 ( \12748 , \12747 );
not \U$12406 ( \12749 , \11377 );
and \U$12407 ( \12750 , \11365 , \12749 );
not \U$12408 ( \12751 , \11365 );
and \U$12409 ( \12752 , \12751 , \11377 );
nor \U$12410 ( \12753 , \12750 , \12752 );
not \U$12411 ( \12754 , \12753 );
not \U$12412 ( \12755 , \478 );
nor \U$12413 ( \12756 , \516 , \518 );
not \U$12414 ( \12757 , \12756 );
not \U$12415 ( \12758 , \9093 );
or \U$12416 ( \12759 , \12757 , \12758 );
not \U$12417 ( \12760 , \485 );
nand \U$12418 ( \12761 , \12759 , \12760 );
not \U$12419 ( \12762 , \12761 );
or \U$12420 ( \12763 , \12755 , \12762 );
nand \U$12421 ( \12764 , \12763 , \488 );
not \U$12422 ( \12765 , \491 );
nand \U$12423 ( \12766 , \12765 , \475 );
and \U$12424 ( \12767 , \12764 , \12766 );
not \U$12425 ( \12768 , \12764 );
not \U$12426 ( \12769 , \12766 );
and \U$12427 ( \12770 , \12768 , \12769 );
nor \U$12428 ( \12771 , \12767 , \12770 );
buf \U$12429 ( \12772 , \12771 );
buf \U$12430 ( \12773 , \12772 );
not \U$12431 ( \12774 , \12773 );
nand \U$12432 ( \12775 , \12774 , \1165 );
not \U$12433 ( \12776 , \12775 );
not \U$12434 ( \12777 , \6316 );
not \U$12435 ( \12778 , \11362 );
or \U$12436 ( \12779 , \12777 , \12778 );
not \U$12437 ( \12780 , \1153 );
not \U$12438 ( \12781 , \12780 );
not \U$12439 ( \12782 , \12781 );
not \U$12440 ( \12783 , \11453 );
not \U$12441 ( \12784 , \12783 );
not \U$12442 ( \12785 , \12784 );
or \U$12443 ( \12786 , \12782 , \12785 );
not \U$12444 ( \12787 , \11453 );
not \U$12445 ( \12788 , \12787 );
or \U$12446 ( \12789 , \12788 , \8679 );
nand \U$12447 ( \12790 , \12786 , \12789 );
nand \U$12448 ( \12791 , \12790 , \9429 );
nand \U$12449 ( \12792 , \12779 , \12791 );
not \U$12450 ( \12793 , \12792 );
or \U$12451 ( \12794 , \12776 , \12793 );
or \U$12452 ( \12795 , \12792 , \12775 );
nand \U$12453 ( \12796 , \12794 , \12795 );
not \U$12454 ( \12797 , \12796 );
not \U$12455 ( \12798 , \796 );
not \U$12456 ( \12799 , \11440 );
or \U$12457 ( \12800 , \12798 , \12799 );
not \U$12458 ( \12801 , \7075 );
not \U$12459 ( \12802 , \6297 );
not \U$12460 ( \12803 , \12802 );
or \U$12461 ( \12804 , \12801 , \12803 );
buf \U$12462 ( \12805 , \8052 );
not \U$12463 ( \12806 , \12805 );
not \U$12464 ( \12807 , \12806 );
nand \U$12465 ( \12808 , \12807 , RI98719b0_131);
nand \U$12466 ( \12809 , \12804 , \12808 );
nand \U$12467 ( \12810 , \12809 , \11433 );
nand \U$12468 ( \12811 , \12800 , \12810 );
not \U$12469 ( \12812 , \12811 );
or \U$12470 ( \12813 , \12797 , \12812 );
not \U$12471 ( \12814 , \12775 );
nand \U$12472 ( \12815 , \12814 , \12792 );
nand \U$12473 ( \12816 , \12813 , \12815 );
not \U$12474 ( \12817 , \12816 );
or \U$12475 ( \12818 , \12754 , \12817 );
or \U$12476 ( \12819 , \12816 , \12753 );
nand \U$12477 ( \12820 , \12818 , \12819 );
not \U$12478 ( \12821 , \12820 );
or \U$12479 ( \12822 , \12748 , \12821 );
not \U$12480 ( \12823 , \12753 );
nand \U$12481 ( \12824 , \12823 , \12816 );
nand \U$12482 ( \12825 , \12822 , \12824 );
not \U$12483 ( \12826 , \3467 );
not \U$12484 ( \12827 , \11293 );
or \U$12485 ( \12828 , \12826 , \12827 );
not \U$12486 ( \12829 , RI98726d0_159);
not \U$12487 ( \12830 , \5205 );
or \U$12488 ( \12831 , \12829 , \12830 );
not \U$12489 ( \12832 , \4407 );
or \U$12490 ( \12833 , \12832 , RI98726d0_159);
nand \U$12491 ( \12834 , \12831 , \12833 );
nand \U$12492 ( \12835 , \12834 , \3465 );
nand \U$12493 ( \12836 , \12828 , \12835 );
not \U$12494 ( \12837 , \12836 );
not \U$12495 ( \12838 , \12602 );
and \U$12496 ( \12839 , \12837 , \12838 );
and \U$12497 ( \12840 , \12836 , \12602 );
nor \U$12498 ( \12841 , \12839 , \12840 );
not \U$12499 ( \12842 , \12841 );
not \U$12500 ( \12843 , \12842 );
not \U$12501 ( \12844 , \9876 );
not \U$12502 ( \12845 , \11410 );
or \U$12503 ( \12846 , \12844 , \12845 );
not \U$12504 ( \12847 , \8839 );
not \U$12505 ( \12848 , \12847 );
not \U$12506 ( \12849 , \12848 );
and \U$12507 ( \12850 , RI9872130_147, \12849 );
not \U$12508 ( \12851 , RI9872130_147);
and \U$12509 ( \12852 , \12851 , \8575 );
or \U$12510 ( \12853 , \12850 , \12852 );
nand \U$12511 ( \12854 , \12853 , \876 );
nand \U$12512 ( \12855 , \12846 , \12854 );
not \U$12513 ( \12856 , \1518 );
not \U$12514 ( \12857 , \11620 );
or \U$12515 ( \12858 , \12856 , \12857 );
not \U$12516 ( \12859 , \8668 );
xor \U$12517 ( \12860 , RI9871c80_137, \12859 );
nand \U$12518 ( \12861 , \12860 , \1501 );
nand \U$12519 ( \12862 , \12858 , \12861 );
xor \U$12520 ( \12863 , \12855 , \12862 );
xnor \U$12521 ( \12864 , RI98730a8_180, \779 );
not \U$12522 ( \12865 , \12864 );
or \U$12523 ( \12866 , \12865 , \11351 );
buf \U$12524 ( \12867 , \11342 );
buf \U$12525 ( \12868 , \12867 );
nand \U$12526 ( \12869 , \12868 , RI98730a8_180);
nand \U$12527 ( \12870 , \12866 , \12869 );
and \U$12528 ( \12871 , \12863 , \12870 );
and \U$12529 ( \12872 , \12855 , \12862 );
or \U$12530 ( \12873 , \12871 , \12872 );
not \U$12531 ( \12874 , \12873 );
or \U$12532 ( \12875 , \12843 , \12874 );
nand \U$12533 ( \12876 , \12836 , \12601 );
nand \U$12534 ( \12877 , \12875 , \12876 );
and \U$12535 ( \12878 , \12825 , \12877 );
not \U$12536 ( \12879 , \12825 );
not \U$12537 ( \12880 , \12877 );
and \U$12538 ( \12881 , \12879 , \12880 );
nor \U$12539 ( \12882 , \12878 , \12881 );
not \U$12540 ( \12883 , \12882 );
or \U$12541 ( \12884 , \12708 , \12883 );
nand \U$12542 ( \12885 , \12825 , \12877 );
nand \U$12543 ( \12886 , \12884 , \12885 );
not \U$12544 ( \12887 , \12886 );
xor \U$12545 ( \12888 , \11782 , \12887 );
xnor \U$12546 ( \12889 , \12888 , \11813 );
not \U$12547 ( \12890 , \12889 );
or \U$12548 ( \12891 , \12701 , \12890 );
buf \U$12549 ( \12892 , \11813 );
not \U$12550 ( \12893 , \12892 );
nor \U$12551 ( \12894 , \12893 , \11782 );
not \U$12552 ( \12895 , \11782 );
nor \U$12553 ( \12896 , \12895 , \12892 );
or \U$12554 ( \12897 , \12894 , \12896 );
nand \U$12555 ( \12898 , \12897 , \12886 );
nand \U$12556 ( \12899 , \12891 , \12898 );
and \U$12557 ( \12900 , \12653 , \12899 );
and \U$12558 ( \12901 , \12374 , \12652 );
or \U$12559 ( \12902 , \12900 , \12901 );
not \U$12560 ( \12903 , \12902 );
not \U$12561 ( \12904 , \11660 );
and \U$12562 ( \12905 , \11826 , \12904 );
not \U$12563 ( \12906 , \11826 );
and \U$12564 ( \12907 , \12906 , \11660 );
or \U$12565 ( \12908 , \12905 , \12907 );
not \U$12566 ( \12909 , \12908 );
not \U$12567 ( \12910 , \12909 );
or \U$12568 ( \12911 , \12903 , \12910 );
not \U$12569 ( \12912 , \12902 );
nand \U$12570 ( \12913 , \12908 , \12912 );
nand \U$12571 ( \12914 , \12911 , \12913 );
not \U$12572 ( \12915 , \12914 );
not \U$12573 ( \12916 , \11844 );
not \U$12574 ( \12917 , \11873 );
or \U$12575 ( \12918 , \12916 , \12917 );
or \U$12576 ( \12919 , \11873 , \11844 );
nand \U$12577 ( \12920 , \12918 , \12919 );
not \U$12578 ( \12921 , \12920 );
or \U$12579 ( \12922 , \12915 , \12921 );
nand \U$12580 ( \12923 , \12908 , \12902 );
nand \U$12581 ( \12924 , \12922 , \12923 );
not \U$12582 ( \12925 , \12924 );
xor \U$12583 ( \12926 , \12369 , \12925 );
xor \U$12584 ( \12927 , \11841 , \11878 );
xnor \U$12585 ( \12928 , \12926 , \12927 );
not \U$12586 ( \12929 , \12928 );
buf \U$12587 ( \12930 , \12920 );
and \U$12588 ( \12931 , \12930 , \12914 );
not \U$12589 ( \12932 , \12930 );
not \U$12590 ( \12933 , \12914 );
and \U$12591 ( \12934 , \12932 , \12933 );
nor \U$12592 ( \12935 , \12931 , \12934 );
not \U$12593 ( \12936 , \12935 );
xor \U$12594 ( \12937 , \12374 , \12652 );
xor \U$12595 ( \12938 , \12937 , \12899 );
xor \U$12596 ( \12939 , \12639 , \12455 );
xor \U$12597 ( \12940 , \12939 , \12580 );
not \U$12598 ( \12941 , \12940 );
xor \U$12599 ( \12942 , \12536 , \12575 );
not \U$12600 ( \12943 , \12942 );
xor \U$12601 ( \12944 , \12586 , \12629 );
xnor \U$12602 ( \12945 , \12944 , \12627 );
not \U$12603 ( \12946 , \12945 );
or \U$12604 ( \12947 , \12943 , \12946 );
or \U$12605 ( \12948 , \12942 , \12945 );
nand \U$12606 ( \12949 , \12947 , \12948 );
xor \U$12607 ( \12950 , \12505 , \12526 );
xnor \U$12608 ( \12951 , \12950 , \12513 );
xor \U$12609 ( \12952 , \12420 , \12432 );
xnor \U$12610 ( \12953 , \12952 , \12443 );
xor \U$12611 ( \12954 , \12951 , \12953 );
xor \U$12612 ( \12955 , \12559 , \12547 );
xnor \U$12613 ( \12956 , \12955 , \12566 );
and \U$12614 ( \12957 , \12954 , \12956 );
and \U$12615 ( \12958 , \12951 , \12953 );
or \U$12616 ( \12959 , \12957 , \12958 );
nand \U$12617 ( \12960 , \12949 , \12959 );
not \U$12618 ( \12961 , \12945 );
nand \U$12619 ( \12962 , \12961 , \12942 );
and \U$12620 ( \12963 , \12960 , \12962 );
not \U$12621 ( \12964 , \3465 );
and \U$12622 ( \12965 , \4989 , RI98726d0_159);
not \U$12623 ( \12966 , \4989 );
and \U$12624 ( \12967 , \12966 , \4063 );
nor \U$12625 ( \12968 , \12965 , \12967 );
not \U$12626 ( \12969 , \12968 );
or \U$12627 ( \12970 , \12964 , \12969 );
not \U$12628 ( \12971 , \4710 );
and \U$12629 ( \12972 , RI98726d0_159, \12971 );
not \U$12630 ( \12973 , RI98726d0_159);
and \U$12631 ( \12974 , \12973 , \5623 );
or \U$12632 ( \12975 , \12972 , \12974 );
nand \U$12633 ( \12976 , \12975 , \3467 );
nand \U$12634 ( \12977 , \12970 , \12976 );
not \U$12635 ( \12978 , \12977 );
not \U$12636 ( \12979 , \9196 );
not \U$12637 ( \12980 , \11559 );
and \U$12638 ( \12981 , \9198 , \12980 );
not \U$12639 ( \12982 , \9198 );
and \U$12640 ( \12983 , \12982 , \5721 );
nor \U$12641 ( \12984 , \12981 , \12983 );
not \U$12642 ( \12985 , \12984 );
or \U$12643 ( \12986 , \12979 , \12985 );
nand \U$12644 ( \12987 , \12610 , \9214 );
nand \U$12645 ( \12988 , \12986 , \12987 );
not \U$12646 ( \12989 , \12988 );
not \U$12647 ( \12990 , \12475 );
not \U$12648 ( \12991 , \12990 );
not \U$12649 ( \12992 , \932 );
and \U$12650 ( \12993 , \12991 , \12992 );
and \U$12651 ( \12994 , \9750 , \1347 );
not \U$12652 ( \12995 , \9750 );
and \U$12653 ( \12996 , \12995 , RI9871d70_139);
or \U$12654 ( \12997 , \12994 , \12996 );
and \U$12655 ( \12998 , \12997 , \859 );
nor \U$12656 ( \12999 , \12993 , \12998 );
nand \U$12657 ( \13000 , \12989 , \12999 );
not \U$12658 ( \13001 , \13000 );
or \U$12659 ( \13002 , \12978 , \13001 );
not \U$12660 ( \13003 , \12999 );
nand \U$12661 ( \13004 , \13003 , \12988 );
nand \U$12662 ( \13005 , \13002 , \13004 );
xor \U$12663 ( \13006 , \12722 , \12733 );
xor \U$12664 ( \13007 , \13006 , \12744 );
xor \U$12665 ( \13008 , \13005 , \13007 );
not \U$12666 ( \13009 , \8028 );
not \U$12667 ( \13010 , RI9872a18_166);
not \U$12668 ( \13011 , \1366 );
or \U$12669 ( \13012 , \13010 , \13011 );
or \U$12670 ( \13013 , \1369 , RI9872a18_166);
nand \U$12671 ( \13014 , \13012 , \13013 );
not \U$12672 ( \13015 , \13014 );
or \U$12673 ( \13016 , \13009 , \13015 );
buf \U$12674 ( \13017 , \9071 );
nand \U$12675 ( \13018 , \12485 , \13017 );
nand \U$12676 ( \13019 , \13016 , \13018 );
not \U$12677 ( \13020 , \11351 );
not \U$12678 ( \13021 , \13020 );
not \U$12679 ( \13022 , RI98730a8_180);
not \U$12680 ( \13023 , \13022 );
not \U$12681 ( \13024 , \2982 );
or \U$12682 ( \13025 , \13023 , \13024 );
or \U$12683 ( \13026 , \1393 , \13022 );
nand \U$12684 ( \13027 , \13025 , \13026 );
not \U$12685 ( \13028 , \13027 );
or \U$12686 ( \13029 , \13021 , \13028 );
nand \U$12687 ( \13030 , \12864 , \12868 );
nand \U$12688 ( \13031 , \13029 , \13030 );
xor \U$12689 ( \13032 , \13019 , \13031 );
buf \U$12690 ( \13033 , \3163 );
not \U$12691 ( \13034 , \13033 );
and \U$12692 ( \13035 , \7028 , RI9872310_151);
not \U$12693 ( \13036 , \7028 );
and \U$12694 ( \13037 , \13036 , \3154 );
nor \U$12695 ( \13038 , \13035 , \13037 );
not \U$12696 ( \13039 , \13038 );
or \U$12697 ( \13040 , \13034 , \13039 );
nand \U$12698 ( \13041 , \12521 , \12514 );
nand \U$12699 ( \13042 , \13040 , \13041 );
and \U$12700 ( \13043 , \13032 , \13042 );
and \U$12701 ( \13044 , \13019 , \13031 );
nor \U$12702 ( \13045 , \13043 , \13044 );
not \U$12703 ( \13046 , \13045 );
and \U$12704 ( \13047 , \13008 , \13046 );
and \U$12705 ( \13048 , \13005 , \13007 );
or \U$12706 ( \13049 , \13047 , \13048 );
not \U$12707 ( \13050 , \13049 );
xor \U$12708 ( \13051 , \12489 , \12478 );
not \U$12709 ( \13052 , \5847 );
not \U$12710 ( \13053 , \12620 );
or \U$12711 ( \13054 , \13052 , \13053 );
and \U$12712 ( \13055 , RI98725e0_157, \6617 );
not \U$12713 ( \13056 , RI98725e0_157);
buf \U$12714 ( \13057 , \4408 );
not \U$12715 ( \13058 , \13057 );
and \U$12716 ( \13059 , \13056 , \13058 );
or \U$12717 ( \13060 , \13055 , \13059 );
nand \U$12718 ( \13061 , \13060 , \4101 );
nand \U$12719 ( \13062 , \13054 , \13061 );
not \U$12720 ( \13063 , \13062 );
not \U$12721 ( \13064 , \1367 );
buf \U$12722 ( \13065 , \9137 );
not \U$12723 ( \13066 , \13065 );
not \U$12724 ( \13067 , \13066 );
not \U$12725 ( \13068 , \13067 );
or \U$12726 ( \13069 , \13064 , \13068 );
buf \U$12727 ( \13070 , \13065 );
buf \U$12728 ( \13071 , \13070 );
or \U$12729 ( \13072 , \13071 , \1367 );
nand \U$12730 ( \13073 , \13069 , \13072 );
not \U$12731 ( \13074 , \13073 );
not \U$12732 ( \13075 , \13074 );
not \U$12733 ( \13076 , \6194 );
and \U$12734 ( \13077 , \13075 , \13076 );
not \U$12735 ( \13078 , RI9871e60_141);
not \U$12736 ( \13079 , \11371 );
or \U$12737 ( \13080 , \13078 , \13079 );
or \U$12738 ( \13081 , \9722 , RI9871e60_141);
nand \U$12739 ( \13082 , \13080 , \13081 );
and \U$12740 ( \13083 , \13082 , \1352 );
nor \U$12741 ( \13084 , \13077 , \13083 );
nand \U$12742 ( \13085 , \13063 , \13084 );
not \U$12743 ( \13086 , \13085 );
not \U$12744 ( \13087 , \9668 );
not \U$12745 ( \13088 , \12564 );
or \U$12746 ( \13089 , \13087 , \13088 );
not \U$12747 ( \13090 , RI9872bf8_170);
not \U$12748 ( \13091 , \2216 );
or \U$12749 ( \13092 , \13090 , \13091 );
or \U$12750 ( \13093 , \848 , RI9872bf8_170);
nand \U$12751 ( \13094 , \13092 , \13093 );
nand \U$12752 ( \13095 , \13094 , \9670 );
nand \U$12753 ( \13096 , \13089 , \13095 );
not \U$12754 ( \13097 , \13096 );
or \U$12755 ( \13098 , \13086 , \13097 );
not \U$12756 ( \13099 , \13084 );
nand \U$12757 ( \13100 , \13099 , \13062 );
nand \U$12758 ( \13101 , \13098 , \13100 );
xor \U$12759 ( \13102 , \13051 , \13101 );
xor \U$12760 ( \13103 , \12855 , \12862 );
xor \U$12761 ( \13104 , \13103 , \12870 );
and \U$12762 ( \13105 , \13102 , \13104 );
and \U$12763 ( \13106 , \13051 , \13101 );
or \U$12764 ( \13107 , \13105 , \13106 );
not \U$12765 ( \13108 , \13107 );
buf \U$12766 ( \13109 , \12507 );
not \U$12767 ( \13110 , \13109 );
and \U$12768 ( \13111 , RI9873030_179, \1097 );
not \U$12769 ( \13112 , RI9873030_179);
and \U$12770 ( \13113 , \13112 , \1106 );
or \U$12771 ( \13114 , \13111 , \13113 );
not \U$12772 ( \13115 , \13114 );
or \U$12773 ( \13116 , \13110 , \13115 );
nand \U$12774 ( \13117 , \12509 , \9937 );
nand \U$12775 ( \13118 , \13116 , \13117 );
not \U$12776 ( \13119 , \13118 );
not \U$12777 ( \13120 , \5642 );
not \U$12778 ( \13121 , RI9872568_156);
not \U$12779 ( \13122 , \6378 );
or \U$12780 ( \13123 , \13121 , \13122 );
nand \U$12781 ( \13124 , \2110 , \5644 );
nand \U$12782 ( \13125 , \13123 , \13124 );
not \U$12783 ( \13126 , \13125 );
or \U$12784 ( \13127 , \13120 , \13126 );
nand \U$12785 ( \13128 , \5653 , \12441 );
nand \U$12786 ( \13129 , \13127 , \13128 );
not \U$12787 ( \13130 , \13129 );
not \U$12788 ( \13131 , \6284 );
and \U$12789 ( \13132 , \1190 , \5632 );
not \U$12790 ( \13133 , \1190 );
and \U$12791 ( \13134 , \13133 , RI98728b0_163);
nor \U$12792 ( \13135 , \13132 , \13134 );
not \U$12793 ( \13136 , \13135 );
or \U$12794 ( \13137 , \13131 , \13136 );
nand \U$12795 ( \13138 , \12395 , \6611 );
nand \U$12796 ( \13139 , \13137 , \13138 );
xnor \U$12797 ( \13140 , \13130 , \13139 );
not \U$12798 ( \13141 , \13140 );
or \U$12799 ( \13142 , \13119 , \13141 );
nand \U$12800 ( \13143 , \13139 , \13129 );
nand \U$12801 ( \13144 , \13142 , \13143 );
not \U$12802 ( \13145 , \5036 );
not \U$12803 ( \13146 , \12553 );
or \U$12804 ( \13147 , \13145 , \13146 );
and \U$12805 ( \13148 , RI9872478_154, \3860 );
not \U$12806 ( \13149 , RI9872478_154);
and \U$12807 ( \13150 , \13149 , \3859 );
nor \U$12808 ( \13151 , \13148 , \13150 );
nand \U$12809 ( \13152 , \13151 , \5034 );
nand \U$12810 ( \13153 , \13147 , \13152 );
not \U$12811 ( \13154 , \13153 );
not \U$12812 ( \13155 , \4919 );
not \U$12813 ( \13156 , RI9872388_152);
not \U$12814 ( \13157 , \10699 );
or \U$12815 ( \13158 , \13156 , \13157 );
or \U$12816 ( \13159 , \11672 , RI9872388_152);
nand \U$12817 ( \13160 , \13158 , \13159 );
not \U$12818 ( \13161 , \13160 );
or \U$12819 ( \13162 , \13155 , \13161 );
nand \U$12820 ( \13163 , \12545 , \4925 );
nand \U$12821 ( \13164 , \13162 , \13163 );
not \U$12822 ( \13165 , \13164 );
nand \U$12823 ( \13166 , \13154 , \13165 );
not \U$12824 ( \13167 , \13166 );
not \U$12825 ( \13168 , \10251 );
not \U$12826 ( \13169 , \6442 );
and \U$12827 ( \13170 , \13169 , RI9872d60_173);
not \U$12828 ( \13171 , \13169 );
and \U$12829 ( \13172 , \13171 , \8807 );
nor \U$12830 ( \13173 , \13170 , \13172 );
not \U$12831 ( \13174 , \13173 );
or \U$12832 ( \13175 , \13168 , \13174 );
nand \U$12833 ( \13176 , \12429 , \8802 );
nand \U$12834 ( \13177 , \13175 , \13176 );
not \U$12835 ( \13178 , \13177 );
or \U$12836 ( \13179 , \13167 , \13178 );
nand \U$12837 ( \13180 , \13153 , \13164 );
nand \U$12838 ( \13181 , \13179 , \13180 );
not \U$12839 ( \13182 , \13181 );
not \U$12840 ( \13183 , \7325 );
not \U$12841 ( \13184 , RI98729a0_165);
not \U$12842 ( \13185 , \6330 );
or \U$12843 ( \13186 , \13184 , \13185 );
or \U$12844 ( \13187 , \9326 , RI98729a0_165);
nand \U$12845 ( \13188 , \13186 , \13187 );
not \U$12846 ( \13189 , \13188 );
or \U$12847 ( \13190 , \13183 , \13189 );
nand \U$12848 ( \13191 , \7338 , \12384 );
nand \U$12849 ( \13192 , \13190 , \13191 );
not \U$12850 ( \13193 , \13192 );
not \U$12851 ( \13194 , \9273 );
not \U$12852 ( \13195 , \12402 );
or \U$12853 ( \13196 , \13194 , \13195 );
not \U$12854 ( \13197 , RI9872e50_175);
not \U$12855 ( \13198 , \1581 );
or \U$12856 ( \13199 , \13197 , \13198 );
or \U$12857 ( \13200 , \1581 , RI9872e50_175);
nand \U$12858 ( \13201 , \13199 , \13200 );
nand \U$12859 ( \13202 , \13201 , \9686 );
nand \U$12860 ( \13203 , \13196 , \13202 );
not \U$12861 ( \13204 , \13203 );
or \U$12862 ( \13205 , \13193 , \13204 );
or \U$12863 ( \13206 , \13203 , \13192 );
not \U$12864 ( \13207 , \9527 );
and \U$12865 ( \13208 , RI9872f40_177, \2492 );
not \U$12866 ( \13209 , RI9872f40_177);
and \U$12867 ( \13210 , \13209 , \10674 );
or \U$12868 ( \13211 , \13208 , \13210 );
not \U$12869 ( \13212 , \13211 );
or \U$12870 ( \13213 , \13207 , \13212 );
buf \U$12871 ( \13214 , \8752 );
nand \U$12872 ( \13215 , \12416 , \13214 );
nand \U$12873 ( \13216 , \13213 , \13215 );
nand \U$12874 ( \13217 , \13206 , \13216 );
nand \U$12875 ( \13218 , \13205 , \13217 );
not \U$12876 ( \13219 , \13218 );
nand \U$12877 ( \13220 , \13182 , \13219 );
nand \U$12878 ( \13221 , \13144 , \13220 );
not \U$12879 ( \13222 , \13219 );
nand \U$12880 ( \13223 , \13222 , \13181 );
and \U$12881 ( \13224 , \13221 , \13223 );
not \U$12882 ( \13225 , \13224 );
or \U$12883 ( \13226 , \13108 , \13225 );
not \U$12884 ( \13227 , \13223 );
not \U$12885 ( \13228 , \13221 );
or \U$12886 ( \13229 , \13227 , \13228 );
not \U$12887 ( \13230 , \13107 );
nand \U$12888 ( \13231 , \13229 , \13230 );
nand \U$12889 ( \13232 , \13226 , \13231 );
not \U$12890 ( \13233 , \13232 );
or \U$12891 ( \13234 , \13050 , \13233 );
not \U$12892 ( \13235 , \13223 );
not \U$12893 ( \13236 , \13221 );
or \U$12894 ( \13237 , \13235 , \13236 );
nand \U$12895 ( \13238 , \13237 , \13107 );
nand \U$12896 ( \13239 , \13234 , \13238 );
not \U$12897 ( \13240 , \13239 );
and \U$12898 ( \13241 , \12963 , \13240 );
not \U$12899 ( \13242 , \12963 );
and \U$12900 ( \13243 , \13242 , \13239 );
nor \U$12901 ( \13244 , \13241 , \13243 );
not \U$12902 ( \13245 , \13244 );
or \U$12903 ( \13246 , \12941 , \13245 );
not \U$12904 ( \13247 , \12962 );
not \U$12905 ( \13248 , \12960 );
or \U$12906 ( \13249 , \13247 , \13248 );
nand \U$12907 ( \13250 , \13249 , \13239 );
nand \U$12908 ( \13251 , \13246 , \13250 );
not \U$12909 ( \13252 , \13251 );
xor \U$12910 ( \13253 , \12642 , \12647 );
xor \U$12911 ( \13254 , \12707 , \12882 );
not \U$12912 ( \13255 , \13254 );
xnor \U$12913 ( \13256 , \11600 , \11575 );
not \U$12914 ( \13257 , \13256 );
xor \U$12915 ( \13258 , \11680 , \11701 );
xor \U$12916 ( \13259 , \13258 , \11694 );
not \U$12917 ( \13260 , \13259 );
or \U$12918 ( \13261 , \13257 , \13260 );
or \U$12919 ( \13262 , \13259 , \13256 );
nand \U$12920 ( \13263 , \13261 , \13262 );
xor \U$12921 ( \13264 , \12796 , \12811 );
not \U$12922 ( \13265 , \13264 );
not \U$12923 ( \13266 , \1162 );
not \U$12924 ( \13267 , \8678 );
buf \U$12925 ( \13268 , \12772 );
not \U$12926 ( \13269 , \13268 );
or \U$12927 ( \13270 , \13267 , \13269 );
or \U$12928 ( \13271 , \13268 , \8679 );
nand \U$12929 ( \13272 , \13270 , \13271 );
not \U$12930 ( \13273 , \13272 );
or \U$12931 ( \13274 , \13266 , \13273 );
nand \U$12932 ( \13275 , \12790 , \1220 );
nand \U$12933 ( \13276 , \13274 , \13275 );
not \U$12934 ( \13277 , \479 );
nand \U$12935 ( \13278 , \13277 , \488 );
buf \U$12936 ( \13279 , \12761 );
xnor \U$12937 ( \13280 , \13278 , \13279 );
buf \U$12938 ( \13281 , \13280 );
and \U$12939 ( \13282 , \13281 , \5753 );
or \U$12940 ( \13283 , \13276 , \13282 );
not \U$12941 ( \13284 , \13283 );
not \U$12942 ( \13285 , RI9871aa0_133);
not \U$12943 ( \13286 , \5705 );
or \U$12944 ( \13287 , \13285 , \13286 );
or \U$12945 ( \13288 , \8895 , RI9871aa0_133);
nand \U$12946 ( \13289 , \13287 , \13288 );
nand \U$12947 ( \13290 , \13289 , \2072 );
nand \U$12948 ( \13291 , \12503 , \2087 );
nand \U$12949 ( \13292 , \13290 , \13291 );
not \U$12950 ( \13293 , \13292 );
or \U$12951 ( \13294 , \13284 , \13293 );
nand \U$12952 ( \13295 , \13276 , \13282 );
nand \U$12953 ( \13296 , \13294 , \13295 );
not \U$12954 ( \13297 , \876 );
buf \U$12955 ( \13298 , \8554 );
and \U$12956 ( \13299 , \13298 , \919 );
not \U$12957 ( \13300 , \13298 );
and \U$12958 ( \13301 , \13300 , RI9872130_147);
nor \U$12959 ( \13302 , \13299 , \13301 );
not \U$12960 ( \13303 , \13302 );
or \U$12961 ( \13304 , \13297 , \13303 );
nand \U$12962 ( \13305 , \12853 , \9876 );
nand \U$12963 ( \13306 , \13304 , \13305 );
not \U$12964 ( \13307 , \1518 );
not \U$12965 ( \13308 , \12860 );
or \U$12966 ( \13309 , \13307 , \13308 );
and \U$12967 ( \13310 , RI9871c80_137, \8650 );
not \U$12968 ( \13311 , RI9871c80_137);
and \U$12969 ( \13312 , \13311 , \8642 );
or \U$12970 ( \13313 , \13310 , \13312 );
nand \U$12971 ( \13314 , \13313 , \1501 );
nand \U$12972 ( \13315 , \13309 , \13314 );
xor \U$12973 ( \13316 , \13306 , \13315 );
not \U$12974 ( \13317 , \12720 );
not \U$12975 ( \13318 , \1283 );
not \U$12976 ( \13319 , \8597 );
or \U$12977 ( \13320 , \13318 , \13319 );
or \U$12978 ( \13321 , \8597 , \1283 );
nand \U$12979 ( \13322 , \13320 , \13321 );
not \U$12980 ( \13323 , \13322 );
or \U$12981 ( \13324 , \13317 , \13323 );
nand \U$12982 ( \13325 , \12719 , \1323 );
nand \U$12983 ( \13326 , \13324 , \13325 );
and \U$12984 ( \13327 , \13316 , \13326 );
and \U$12985 ( \13328 , \13306 , \13315 );
or \U$12986 ( \13329 , \13327 , \13328 );
xor \U$12987 ( \13330 , \13296 , \13329 );
not \U$12988 ( \13331 , \13330 );
or \U$12989 ( \13332 , \13265 , \13331 );
nand \U$12990 ( \13333 , \13296 , \13329 );
nand \U$12991 ( \13334 , \13332 , \13333 );
nand \U$12992 ( \13335 , \13263 , \13334 );
not \U$12993 ( \13336 , \13256 );
nand \U$12994 ( \13337 , \13336 , \13259 );
nand \U$12995 ( \13338 , \13335 , \13337 );
not \U$12996 ( \13339 , \12841 );
not \U$12997 ( \13340 , \12873 );
or \U$12998 ( \13341 , \13339 , \13340 );
or \U$12999 ( \13342 , \12873 , \12841 );
nand \U$13000 ( \13343 , \13341 , \13342 );
not \U$13001 ( \13344 , \13343 );
not \U$13002 ( \13345 , \11433 );
not \U$13003 ( \13346 , \6568 );
not \U$13004 ( \13347 , \6528 );
or \U$13005 ( \13348 , \13346 , \13347 );
or \U$13006 ( \13349 , \8934 , \1078 );
nand \U$13007 ( \13350 , \13348 , \13349 );
not \U$13008 ( \13351 , \13350 );
or \U$13009 ( \13352 , \13345 , \13351 );
nand \U$13010 ( \13353 , \12809 , \796 );
nand \U$13011 ( \13354 , \13352 , \13353 );
not \U$13012 ( \13355 , \1455 );
and \U$13013 ( \13356 , RI9871c08_136, \9599 );
not \U$13014 ( \13357 , RI9871c08_136);
not \U$13015 ( \13358 , \8074 );
and \U$13016 ( \13359 , \13357 , \13358 );
or \U$13017 ( \13360 , \13356 , \13359 );
not \U$13018 ( \13361 , \13360 );
or \U$13019 ( \13362 , \13355 , \13361 );
nand \U$13020 ( \13363 , \12731 , \1429 );
nand \U$13021 ( \13364 , \13362 , \13363 );
or \U$13022 ( \13365 , \13354 , \13364 );
not \U$13023 ( \13366 , \6672 );
not \U$13024 ( \13367 , \12742 );
or \U$13025 ( \13368 , \13366 , \13367 );
not \U$13026 ( \13369 , \1111 );
not \U$13027 ( \13370 , \9569 );
or \U$13028 ( \13371 , \13369 , \13370 );
nand \U$13029 ( \13372 , \8924 , RI98718c0_129);
nand \U$13030 ( \13373 , \13371 , \13372 );
nand \U$13031 ( \13374 , \13373 , \1083 );
nand \U$13032 ( \13375 , \13368 , \13374 );
nand \U$13033 ( \13376 , \13365 , \13375 );
nand \U$13034 ( \13377 , \13354 , \13364 );
nand \U$13035 ( \13378 , \13376 , \13377 );
not \U$13036 ( \13379 , \13378 );
nand \U$13037 ( \13380 , RI9873288_184, RI9873300_185);
nand \U$13038 ( \13381 , \13380 , RI9873210_183);
not \U$13039 ( \13382 , \1013 );
not \U$13040 ( \13383 , \12599 );
or \U$13041 ( \13384 , \13382 , \13383 );
not \U$13042 ( \13385 , \12592 );
not \U$13043 ( \13386 , \13385 );
not \U$13044 ( \13387 , \10063 );
not \U$13045 ( \13388 , \13387 );
not \U$13046 ( \13389 , \13388 );
or \U$13047 ( \13390 , \13386 , \13389 );
buf \U$13048 ( \13391 , \10063 );
or \U$13049 ( \13392 , \13391 , \8085 );
nand \U$13050 ( \13393 , \13390 , \13392 );
nand \U$13051 ( \13394 , \13393 , \1018 );
nand \U$13052 ( \13395 , \13384 , \13394 );
xor \U$13053 ( \13396 , \13381 , \13395 );
not \U$13054 ( \13397 , \1380 );
not \U$13055 ( \13398 , \13082 );
or \U$13056 ( \13399 , \13397 , \13398 );
nand \U$13057 ( \13400 , \12464 , \1352 );
nand \U$13058 ( \13401 , \13399 , \13400 );
and \U$13059 ( \13402 , \13396 , \13401 );
and \U$13060 ( \13403 , \13381 , \13395 );
nor \U$13061 ( \13404 , \13402 , \13403 );
not \U$13062 ( \13405 , \13404 );
not \U$13063 ( \13406 , \3467 );
not \U$13064 ( \13407 , \12834 );
or \U$13065 ( \13408 , \13406 , \13407 );
buf \U$13066 ( \13409 , \3465 );
nand \U$13067 ( \13410 , \12975 , \13409 );
nand \U$13068 ( \13411 , \13408 , \13410 );
not \U$13069 ( \13412 , \13411 );
or \U$13070 ( \13413 , \13405 , \13412 );
or \U$13071 ( \13414 , \13411 , \13404 );
nand \U$13072 ( \13415 , \13413 , \13414 );
not \U$13073 ( \13416 , \13415 );
or \U$13074 ( \13417 , \13379 , \13416 );
not \U$13075 ( \13418 , \13404 );
nand \U$13076 ( \13419 , \13418 , \13411 );
nand \U$13077 ( \13420 , \13417 , \13419 );
not \U$13078 ( \13421 , \13420 );
or \U$13079 ( \13422 , \13344 , \13421 );
xnor \U$13080 ( \13423 , \12820 , \12747 );
not \U$13081 ( \13424 , \13423 );
xor \U$13082 ( \13425 , \13420 , \13343 );
nand \U$13083 ( \13426 , \13424 , \13425 );
nand \U$13084 ( \13427 , \13422 , \13426 );
xor \U$13085 ( \13428 , \13338 , \13427 );
not \U$13086 ( \13429 , \13428 );
or \U$13087 ( \13430 , \13255 , \13429 );
not \U$13088 ( \13431 , \13337 );
not \U$13089 ( \13432 , \13335 );
or \U$13090 ( \13433 , \13431 , \13432 );
nand \U$13091 ( \13434 , \13433 , \13427 );
nand \U$13092 ( \13435 , \13430 , \13434 );
xor \U$13093 ( \13436 , \13253 , \13435 );
not \U$13094 ( \13437 , \13436 );
or \U$13095 ( \13438 , \13252 , \13437 );
xor \U$13096 ( \13439 , \12642 , \12647 );
nand \U$13097 ( \13440 , \13439 , \13435 );
nand \U$13098 ( \13441 , \13438 , \13440 );
and \U$13099 ( \13442 , \12938 , \13441 );
not \U$13100 ( \13443 , \12938 );
not \U$13101 ( \13444 , \13441 );
and \U$13102 ( \13445 , \13443 , \13444 );
nor \U$13103 ( \13446 , \13442 , \13445 );
not \U$13104 ( \13447 , \13446 );
xnor \U$13105 ( \13448 , \13264 , \13330 );
not \U$13106 ( \13449 , \13448 );
not \U$13107 ( \13450 , \13449 );
not \U$13108 ( \13451 , \9876 );
not \U$13109 ( \13452 , \13302 );
or \U$13110 ( \13453 , \13451 , \13452 );
not \U$13111 ( \13454 , \8722 );
xnor \U$13112 ( \13455 , \13454 , RI9872130_147);
nand \U$13113 ( \13456 , \13455 , \6431 );
nand \U$13114 ( \13457 , \13453 , \13456 );
not \U$13115 ( \13458 , \13457 );
not \U$13116 ( \13459 , \832 );
not \U$13117 ( \13460 , \12997 );
or \U$13118 ( \13461 , \13459 , \13460 );
and \U$13119 ( \13462 , \9850 , \12108 );
not \U$13120 ( \13463 , \9850 );
and \U$13121 ( \13464 , \13463 , RI9871d70_139);
nor \U$13122 ( \13465 , \13462 , \13464 );
nand \U$13123 ( \13466 , \13465 , \859 );
nand \U$13124 ( \13467 , \13461 , \13466 );
not \U$13125 ( \13468 , \13467 );
not \U$13126 ( \13469 , \13468 );
not \U$13127 ( \13470 , \13380 );
nor \U$13128 ( \13471 , RI9873288_184, RI9873300_185);
nor \U$13129 ( \13472 , \13470 , \13471 );
xnor \U$13130 ( \13473 , RI9873300_185, RI9873210_183);
or \U$13131 ( \13474 , \13472 , \13473 );
not \U$13132 ( \13475 , \13474 );
buf \U$13133 ( \13476 , \13475 );
buf \U$13134 ( \13477 , \13476 );
not \U$13135 ( \13478 , \13477 );
xor \U$13136 ( \13479 , RI9873210_183, \1690 );
not \U$13137 ( \13480 , \13479 );
or \U$13138 ( \13481 , \13478 , \13480 );
buf \U$13139 ( \13482 , \13472 );
buf \U$13140 ( \13483 , \13482 );
buf \U$13141 ( \13484 , \13483 );
nand \U$13142 ( \13485 , \13484 , RI9873210_183);
nand \U$13143 ( \13486 , \13481 , \13485 );
not \U$13144 ( \13487 , \13486 );
or \U$13145 ( \13488 , \13469 , \13487 );
or \U$13146 ( \13489 , \13486 , \13468 );
nand \U$13147 ( \13490 , \13488 , \13489 );
not \U$13148 ( \13491 , \13490 );
or \U$13149 ( \13492 , \13458 , \13491 );
not \U$13150 ( \13493 , \13468 );
buf \U$13151 ( \13494 , \13486 );
nand \U$13152 ( \13495 , \13493 , \13494 );
nand \U$13153 ( \13496 , \13492 , \13495 );
xnor \U$13154 ( \13497 , \13396 , \13401 );
not \U$13155 ( \13498 , \13497 );
not \U$13156 ( \13499 , \13282 );
not \U$13157 ( \13500 , \13276 );
or \U$13158 ( \13501 , \13499 , \13500 );
or \U$13159 ( \13502 , \13276 , \13282 );
nand \U$13160 ( \13503 , \13501 , \13502 );
or \U$13161 ( \13504 , \13292 , \13503 );
not \U$13162 ( \13505 , \13291 );
not \U$13163 ( \13506 , \13290 );
or \U$13164 ( \13507 , \13505 , \13506 );
nand \U$13165 ( \13508 , \13507 , \13503 );
nand \U$13166 ( \13509 , \13504 , \13508 );
not \U$13167 ( \13510 , \13509 );
or \U$13168 ( \13511 , \13498 , \13510 );
or \U$13169 ( \13512 , \13509 , \13497 );
nand \U$13170 ( \13513 , \13511 , \13512 );
nand \U$13171 ( \13514 , \13496 , \13513 );
not \U$13172 ( \13515 , \13497 );
nand \U$13173 ( \13516 , \13515 , \13509 );
nand \U$13174 ( \13517 , \13514 , \13516 );
xor \U$13175 ( \13518 , \13415 , \13378 );
xor \U$13176 ( \13519 , \13517 , \13518 );
not \U$13177 ( \13520 , \13519 );
or \U$13178 ( \13521 , \13450 , \13520 );
not \U$13179 ( \13522 , \13516 );
not \U$13180 ( \13523 , \13514 );
or \U$13181 ( \13524 , \13522 , \13523 );
nand \U$13182 ( \13525 , \13524 , \13518 );
nand \U$13183 ( \13526 , \13521 , \13525 );
not \U$13184 ( \13527 , \13526 );
not \U$13185 ( \13528 , \13423 );
not \U$13186 ( \13529 , \13425 );
or \U$13187 ( \13530 , \13528 , \13529 );
or \U$13188 ( \13531 , \13425 , \13423 );
nand \U$13189 ( \13532 , \13530 , \13531 );
not \U$13190 ( \13533 , \13532 );
not \U$13191 ( \13534 , \12691 );
not \U$13192 ( \13535 , \12678 );
and \U$13193 ( \13536 , \13534 , \13535 );
and \U$13194 ( \13537 , \12691 , \12678 );
nor \U$13195 ( \13538 , \13536 , \13537 );
not \U$13196 ( \13539 , \13538 );
or \U$13197 ( \13540 , \13533 , \13539 );
or \U$13198 ( \13541 , \13538 , \13532 );
nand \U$13199 ( \13542 , \13540 , \13541 );
not \U$13200 ( \13543 , \13542 );
or \U$13201 ( \13544 , \13527 , \13543 );
not \U$13202 ( \13545 , \13538 );
nand \U$13203 ( \13546 , \13545 , \13532 );
nand \U$13204 ( \13547 , \13544 , \13546 );
not \U$13205 ( \13548 , \13547 );
xor \U$13206 ( \13549 , \13256 , \13334 );
xnor \U$13207 ( \13550 , \13549 , \13259 );
not \U$13208 ( \13551 , \13550 );
and \U$13209 ( \13552 , \12613 , \12624 );
not \U$13210 ( \13553 , \12613 );
not \U$13211 ( \13554 , \12624 );
and \U$13212 ( \13555 , \13553 , \13554 );
nor \U$13213 ( \13556 , \13552 , \13555 );
xor \U$13214 ( \13557 , \12386 , \12397 );
xor \U$13215 ( \13558 , \13557 , \12406 );
xor \U$13216 ( \13559 , \13556 , \13558 );
not \U$13217 ( \13560 , \1323 );
not \U$13218 ( \13561 , \13322 );
or \U$13219 ( \13562 , \13560 , \13561 );
and \U$13220 ( \13563 , RI9871b18_134, \9885 );
not \U$13221 ( \13564 , RI9871b18_134);
and \U$13222 ( \13565 , \13564 , \8668 );
nor \U$13223 ( \13566 , \13563 , \13565 );
nand \U$13224 ( \13567 , \13566 , \1292 );
nand \U$13225 ( \13568 , \13562 , \13567 );
not \U$13226 ( \13569 , \13568 );
not \U$13227 ( \13570 , \1429 );
not \U$13228 ( \13571 , \13360 );
or \U$13229 ( \13572 , \13570 , \13571 );
not \U$13230 ( \13573 , RI9871c08_136);
not \U$13231 ( \13574 , \12712 );
or \U$13232 ( \13575 , \13573 , \13574 );
nand \U$13233 ( \13576 , \10597 , \1850 );
nand \U$13234 ( \13577 , \13575 , \13576 );
nand \U$13235 ( \13578 , \13577 , \1455 );
nand \U$13236 ( \13579 , \13572 , \13578 );
not \U$13237 ( \13580 , \1518 );
not \U$13238 ( \13581 , \13313 );
or \U$13239 ( \13582 , \13580 , \13581 );
and \U$13240 ( \13583 , RI9871c80_137, \8579 );
not \U$13241 ( \13584 , RI9871c80_137);
and \U$13242 ( \13585 , \13584 , \8845 );
or \U$13243 ( \13586 , \13583 , \13585 );
nand \U$13244 ( \13587 , \1501 , \13586 );
nand \U$13245 ( \13588 , \13582 , \13587 );
xor \U$13246 ( \13589 , \13579 , \13588 );
not \U$13247 ( \13590 , \13589 );
or \U$13248 ( \13591 , \13569 , \13590 );
nand \U$13249 ( \13592 , \13579 , \13588 );
nand \U$13250 ( \13593 , \13591 , \13592 );
not \U$13251 ( \13594 , \13593 );
not \U$13252 ( \13595 , \1013 );
not \U$13253 ( \13596 , \13393 );
or \U$13254 ( \13597 , \13595 , \13596 );
not \U$13255 ( \13598 , \8085 );
not \U$13256 ( \13599 , \12788 );
or \U$13257 ( \13600 , \13598 , \13599 );
not \U$13258 ( \13601 , \12784 );
nand \U$13259 ( \13602 , \13601 , \1043 );
nand \U$13260 ( \13603 , \13600 , \13602 );
not \U$13261 ( \13604 , \13603 );
or \U$13262 ( \13605 , \13604 , \1612 );
nand \U$13263 ( \13606 , \13597 , \13605 );
not \U$13264 ( \13607 , \13606 );
not \U$13265 ( \13608 , \518 );
not \U$13266 ( \13609 , \13608 );
buf \U$13267 ( \13610 , \9093 );
not \U$13268 ( \13611 , \13610 );
or \U$13269 ( \13612 , \13609 , \13611 );
nand \U$13270 ( \13613 , RI986fac0_65, RI986fb38_66);
buf \U$13271 ( \13614 , \13613 );
nand \U$13272 ( \13615 , \13612 , \13614 );
not \U$13273 ( \13616 , \13615 );
not \U$13274 ( \13617 , \516 );
nand \U$13275 ( \13618 , \13617 , \484 );
not \U$13276 ( \13619 , \13618 );
and \U$13277 ( \13620 , \13616 , \13619 );
and \U$13278 ( \13621 , \13615 , \13618 );
nor \U$13279 ( \13622 , \13620 , \13621 );
not \U$13280 ( \13623 , \13622 );
not \U$13281 ( \13624 , \13623 );
not \U$13282 ( \13625 , \13624 );
and \U$13283 ( \13626 , \8679 , \13625 );
not \U$13284 ( \13627 , \6316 );
not \U$13285 ( \13628 , \13272 );
or \U$13286 ( \13629 , \13627 , \13628 );
and \U$13287 ( \13630 , \13281 , \8678 );
not \U$13288 ( \13631 , \13281 );
and \U$13289 ( \13632 , \13631 , \1166 );
nor \U$13290 ( \13633 , \13630 , \13632 );
nand \U$13291 ( \13634 , \9429 , \13633 );
nand \U$13292 ( \13635 , \13629 , \13634 );
xor \U$13293 ( \13636 , \13626 , \13635 );
not \U$13294 ( \13637 , \13636 );
or \U$13295 ( \13638 , \13607 , \13637 );
nand \U$13296 ( \13639 , \13635 , \13626 );
nand \U$13297 ( \13640 , \13638 , \13639 );
not \U$13298 ( \13641 , \13640 );
not \U$13299 ( \13642 , \796 );
not \U$13300 ( \13643 , \13350 );
or \U$13301 ( \13644 , \13642 , \13643 );
not \U$13302 ( \13645 , \8947 );
not \U$13303 ( \13646 , RI98719b0_131);
and \U$13304 ( \13647 , \13645 , \13646 );
not \U$13305 ( \13648 , \13645 );
and \U$13306 ( \13649 , \13648 , RI98719b0_131);
nor \U$13307 ( \13650 , \13647 , \13649 );
nand \U$13308 ( \13651 , \13650 , \793 );
nand \U$13309 ( \13652 , \13644 , \13651 );
not \U$13310 ( \13653 , \13652 );
not \U$13311 ( \13654 , \2085 );
not \U$13312 ( \13655 , \13289 );
or \U$13313 ( \13656 , \13654 , \13655 );
not \U$13314 ( \13657 , RI9871aa0_133);
not \U$13315 ( \13658 , \8904 );
or \U$13316 ( \13659 , \13657 , \13658 );
not \U$13317 ( \13660 , \12806 );
or \U$13318 ( \13661 , \13660 , RI9871aa0_133);
nand \U$13319 ( \13662 , \13659 , \13661 );
nand \U$13320 ( \13663 , \13662 , \2071 );
nand \U$13321 ( \13664 , \13656 , \13663 );
not \U$13322 ( \13665 , \13664 );
or \U$13323 ( \13666 , \13653 , \13665 );
or \U$13324 ( \13667 , \13664 , \13652 );
not \U$13325 ( \13668 , \1083 );
not \U$13326 ( \13669 , \1111 );
not \U$13327 ( \13670 , \8916 );
or \U$13328 ( \13671 , \13669 , \13670 );
nand \U$13329 ( \13672 , \9895 , RI98718c0_129);
nand \U$13330 ( \13673 , \13671 , \13672 );
not \U$13331 ( \13674 , \13673 );
or \U$13332 ( \13675 , \13668 , \13674 );
nand \U$13333 ( \13676 , \13373 , \1136 );
nand \U$13334 ( \13677 , \13675 , \13676 );
nand \U$13335 ( \13678 , \13667 , \13677 );
nand \U$13336 ( \13679 , \13666 , \13678 );
not \U$13337 ( \13680 , \13679 );
not \U$13338 ( \13681 , \13680 );
or \U$13339 ( \13682 , \13641 , \13681 );
not \U$13340 ( \13683 , \13640 );
nand \U$13341 ( \13684 , \13683 , \13679 );
nand \U$13342 ( \13685 , \13682 , \13684 );
not \U$13343 ( \13686 , \13685 );
or \U$13344 ( \13687 , \13594 , \13686 );
nand \U$13345 ( \13688 , \13679 , \13640 );
nand \U$13346 ( \13689 , \13687 , \13688 );
and \U$13347 ( \13690 , \13559 , \13689 );
and \U$13348 ( \13691 , \13556 , \13558 );
nor \U$13349 ( \13692 , \13690 , \13691 );
not \U$13350 ( \13693 , \13692 );
xor \U$13351 ( \13694 , \12410 , \12451 );
not \U$13352 ( \13695 , \13694 );
or \U$13353 ( \13696 , \13693 , \13695 );
or \U$13354 ( \13697 , \13694 , \13692 );
nand \U$13355 ( \13698 , \13696 , \13697 );
not \U$13356 ( \13699 , \13698 );
or \U$13357 ( \13700 , \13551 , \13699 );
not \U$13358 ( \13701 , \13692 );
nand \U$13359 ( \13702 , \13701 , \13694 );
nand \U$13360 ( \13703 , \13700 , \13702 );
not \U$13361 ( \13704 , \13703 );
xor \U$13362 ( \13705 , \12655 , \12663 );
xnor \U$13363 ( \13706 , \13705 , \12695 );
not \U$13364 ( \13707 , \13706 );
or \U$13365 ( \13708 , \13704 , \13707 );
or \U$13366 ( \13709 , \13706 , \13703 );
nand \U$13367 ( \13710 , \13708 , \13709 );
not \U$13368 ( \13711 , \13710 );
or \U$13369 ( \13712 , \13548 , \13711 );
not \U$13370 ( \13713 , \13706 );
nand \U$13371 ( \13714 , \13713 , \13703 );
nand \U$13372 ( \13715 , \13712 , \13714 );
not \U$13373 ( \13716 , \13715 );
xnor \U$13374 ( \13717 , \12889 , \12700 );
nand \U$13375 ( \13718 , \13716 , \13717 );
not \U$13376 ( \13719 , \13718 );
xor \U$13377 ( \13720 , \11481 , \11484 );
xor \U$13378 ( \13721 , \13720 , \11489 );
not \U$13379 ( \13722 , \11535 );
xor \U$13380 ( \13723 , \11650 , \13722 );
xnor \U$13381 ( \13724 , \13723 , \11514 );
xor \U$13382 ( \13725 , \13721 , \13724 );
xor \U$13383 ( \13726 , \11501 , \11505 );
xnor \U$13384 ( \13727 , \13726 , \11508 );
and \U$13385 ( \13728 , \11531 , \11516 );
not \U$13386 ( \13729 , \11531 );
not \U$13387 ( \13730 , \11516 );
and \U$13388 ( \13731 , \13729 , \13730 );
nor \U$13389 ( \13732 , \13728 , \13731 );
xor \U$13390 ( \13733 , \13727 , \13732 );
xor \U$13391 ( \13734 , \11775 , \11779 );
xor \U$13392 ( \13735 , \13734 , \11704 );
not \U$13393 ( \13736 , \13735 );
and \U$13394 ( \13737 , \13733 , \13736 );
and \U$13395 ( \13738 , \13727 , \13732 );
or \U$13396 ( \13739 , \13737 , \13738 );
not \U$13397 ( \13740 , \13739 );
xor \U$13398 ( \13741 , \13725 , \13740 );
not \U$13399 ( \13742 , \13741 );
or \U$13400 ( \13743 , \13719 , \13742 );
not \U$13401 ( \13744 , \13717 );
nand \U$13402 ( \13745 , \13744 , \13715 );
nand \U$13403 ( \13746 , \13743 , \13745 );
not \U$13404 ( \13747 , \13746 );
or \U$13405 ( \13748 , \13447 , \13747 );
nand \U$13406 ( \13749 , \13441 , \12938 );
nand \U$13407 ( \13750 , \13748 , \13749 );
not \U$13408 ( \13751 , \13750 );
xor \U$13409 ( \13752 , \11851 , \11856 );
xor \U$13410 ( \13753 , \13752 , \11860 );
not \U$13411 ( \13754 , \13753 );
not \U$13412 ( \13755 , \13754 );
xnor \U$13413 ( \13756 , \11498 , \11655 );
not \U$13414 ( \13757 , \13756 );
not \U$13415 ( \13758 , \13757 );
or \U$13416 ( \13759 , \13755 , \13758 );
nand \U$13417 ( \13760 , \13756 , \13753 );
nand \U$13418 ( \13761 , \13759 , \13760 );
not \U$13419 ( \13762 , \13761 );
not \U$13420 ( \13763 , \13721 );
not \U$13421 ( \13764 , \13763 );
not \U$13422 ( \13765 , \13724 );
and \U$13423 ( \13766 , \13740 , \13765 );
not \U$13424 ( \13767 , \13740 );
and \U$13425 ( \13768 , \13767 , \13724 );
nor \U$13426 ( \13769 , \13766 , \13768 );
not \U$13427 ( \13770 , \13769 );
or \U$13428 ( \13771 , \13764 , \13770 );
nand \U$13429 ( \13772 , \13739 , \13724 );
nand \U$13430 ( \13773 , \13771 , \13772 );
not \U$13431 ( \13774 , \13773 );
or \U$13432 ( \13775 , \13762 , \13774 );
nand \U$13433 ( \13776 , \13757 , \13753 );
nand \U$13434 ( \13777 , \13775 , \13776 );
not \U$13435 ( \13778 , \13777 );
and \U$13436 ( \13779 , \13751 , \13778 );
not \U$13437 ( \13780 , \13751 );
and \U$13438 ( \13781 , \13780 , \13777 );
nor \U$13439 ( \13782 , \13779 , \13781 );
not \U$13440 ( \13783 , \13782 );
or \U$13441 ( \13784 , \12936 , \13783 );
not \U$13442 ( \13785 , \13751 );
nand \U$13443 ( \13786 , \13785 , \13777 );
nand \U$13444 ( \13787 , \13784 , \13786 );
not \U$13445 ( \13788 , \13787 );
nand \U$13446 ( \13789 , \12929 , \13788 );
buf \U$13447 ( \13790 , \13789 );
xor \U$13448 ( \13791 , \12935 , \13782 );
not \U$13449 ( \13792 , \13791 );
xnor \U$13450 ( \13793 , \13773 , \13761 );
not \U$13451 ( \13794 , \13793 );
not \U$13452 ( \13795 , \13794 );
xor \U$13453 ( \13796 , \13446 , \13746 );
not \U$13454 ( \13797 , \13796 );
or \U$13455 ( \13798 , \13795 , \13797 );
or \U$13456 ( \13799 , \13796 , \13794 );
xor \U$13457 ( \13800 , \13710 , \13547 );
not \U$13458 ( \13801 , \13800 );
not \U$13459 ( \13802 , \12940 );
and \U$13460 ( \13803 , \13244 , \13802 );
not \U$13461 ( \13804 , \13244 );
and \U$13462 ( \13805 , \13804 , \12940 );
nor \U$13463 ( \13806 , \13803 , \13805 );
not \U$13464 ( \13807 , \13806 );
not \U$13465 ( \13808 , \13807 );
xor \U$13466 ( \13809 , \13698 , \13550 );
not \U$13467 ( \13810 , \13809 );
xor \U$13468 ( \13811 , \12999 , \12977 );
xnor \U$13469 ( \13812 , \13811 , \12988 );
xor \U$13470 ( \13813 , \13216 , \13203 );
and \U$13471 ( \13814 , \13813 , \13192 );
not \U$13472 ( \13815 , \13813 );
not \U$13473 ( \13816 , \13192 );
and \U$13474 ( \13817 , \13815 , \13816 );
nor \U$13475 ( \13818 , \13814 , \13817 );
xor \U$13476 ( \13819 , \13812 , \13818 );
not \U$13477 ( \13820 , \793 );
not \U$13478 ( \13821 , \5367 );
not \U$13479 ( \13822 , \7467 );
or \U$13480 ( \13823 , \13821 , \13822 );
buf \U$13481 ( \13824 , \7465 );
nand \U$13482 ( \13825 , \13824 , RI98719b0_131);
nand \U$13483 ( \13826 , \13823 , \13825 );
not \U$13484 ( \13827 , \13826 );
or \U$13485 ( \13828 , \13820 , \13827 );
nand \U$13486 ( \13829 , \13650 , \796 );
nand \U$13487 ( \13830 , \13828 , \13829 );
not \U$13488 ( \13831 , \13830 );
not \U$13489 ( \13832 , \13831 );
not \U$13490 ( \13833 , \1455 );
xor \U$13491 ( \13834 , \8597 , RI9871c08_136);
not \U$13492 ( \13835 , \13834 );
or \U$13493 ( \13836 , \13833 , \13835 );
nand \U$13494 ( \13837 , \13577 , \1429 );
nand \U$13495 ( \13838 , \13836 , \13837 );
not \U$13496 ( \13839 , \13838 );
not \U$13497 ( \13840 , \13839 );
or \U$13498 ( \13841 , \13832 , \13840 );
not \U$13499 ( \13842 , \1083 );
and \U$13500 ( \13843 , RI98718c0_129, \10392 );
not \U$13501 ( \13844 , RI98718c0_129);
and \U$13502 ( \13845 , \13844 , \13358 );
or \U$13503 ( \13846 , \13843 , \13845 );
not \U$13504 ( \13847 , \13846 );
or \U$13505 ( \13848 , \13842 , \13847 );
nand \U$13506 ( \13849 , \13673 , \1136 );
nand \U$13507 ( \13850 , \13848 , \13849 );
nand \U$13508 ( \13851 , \13841 , \13850 );
nand \U$13509 ( \13852 , \13838 , \13830 );
nand \U$13510 ( \13853 , \13851 , \13852 );
not \U$13511 ( \13854 , \13610 );
nand \U$13512 ( \13855 , \13608 , \13613 );
not \U$13513 ( \13856 , \13855 );
and \U$13514 ( \13857 , \13854 , \13856 );
and \U$13515 ( \13858 , \13610 , \13855 );
nor \U$13516 ( \13859 , \13857 , \13858 );
buf \U$13517 ( \13860 , \13859 );
not \U$13518 ( \13861 , \13860 );
and \U$13519 ( \13862 , \13861 , \1165 );
not \U$13520 ( \13863 , \13862 );
nand \U$13521 ( \13864 , RI9873378_186, RI98733f0_187);
and \U$13522 ( \13865 , \13864 , RI9873288_184);
not \U$13523 ( \13866 , \13865 );
and \U$13524 ( \13867 , \13863 , \13866 );
and \U$13525 ( \13868 , \13862 , \13865 );
nor \U$13526 ( \13869 , \13867 , \13868 );
not \U$13527 ( \13870 , \13869 );
not \U$13528 ( \13871 , \13870 );
not \U$13529 ( \13872 , \1353 );
not \U$13530 ( \13873 , \13073 );
or \U$13531 ( \13874 , \13872 , \13873 );
not \U$13532 ( \13875 , \5616 );
not \U$13533 ( \13876 , \13391 );
not \U$13534 ( \13877 , \13876 );
or \U$13535 ( \13878 , \13875 , \13877 );
nand \U$13536 ( \13879 , RI9871e60_141, \10064 );
nand \U$13537 ( \13880 , \13878 , \13879 );
nand \U$13538 ( \13881 , \13880 , \1380 );
nand \U$13539 ( \13882 , \13874 , \13881 );
not \U$13540 ( \13883 , \13882 );
or \U$13541 ( \13884 , \13871 , \13883 );
not \U$13542 ( \13885 , \13865 );
nand \U$13543 ( \13886 , \13885 , \13862 );
nand \U$13544 ( \13887 , \13884 , \13886 );
xor \U$13545 ( \13888 , \13853 , \13887 );
not \U$13546 ( \13889 , \13888 );
not \U$13547 ( \13890 , \2071 );
not \U$13548 ( \13891 , \2076 );
not \U$13549 ( \13892 , \7905 );
or \U$13550 ( \13893 , \13891 , \13892 );
or \U$13551 ( \13894 , \8934 , \2076 );
nand \U$13552 ( \13895 , \13893 , \13894 );
not \U$13553 ( \13896 , \13895 );
or \U$13554 ( \13897 , \13890 , \13896 );
nand \U$13555 ( \13898 , \13662 , \2085 );
nand \U$13556 ( \13899 , \13897 , \13898 );
not \U$13557 ( \13900 , \13899 );
not \U$13558 ( \13901 , \6653 );
and \U$13559 ( \13902 , RI9872310_151, \6308 );
not \U$13560 ( \13903 , RI9872310_151);
and \U$13561 ( \13904 , \13903 , \11438 );
or \U$13562 ( \13905 , \13902 , \13904 );
not \U$13563 ( \13906 , \13905 );
or \U$13564 ( \13907 , \13901 , \13906 );
and \U$13565 ( \13908 , RI9872310_151, \5761 );
not \U$13566 ( \13909 , RI9872310_151);
and \U$13567 ( \13910 , \13909 , \5766 );
or \U$13568 ( \13911 , \13908 , \13910 );
nand \U$13569 ( \13912 , \13911 , \3170 );
nand \U$13570 ( \13913 , \13907 , \13912 );
not \U$13571 ( \13914 , \13913 );
not \U$13572 ( \13915 , \530 );
and \U$13573 ( \13916 , \533 , \528 );
not \U$13574 ( \13917 , \13916 );
not \U$13575 ( \13918 , \515 );
or \U$13576 ( \13919 , \13917 , \13918 );
not \U$13577 ( \13920 , \579 );
nand \U$13578 ( \13921 , \13919 , \13920 );
not \U$13579 ( \13922 , \13921 );
or \U$13580 ( \13923 , \13915 , \13922 );
not \U$13581 ( \13924 , \583 );
nand \U$13582 ( \13925 , \13923 , \13924 );
nor \U$13583 ( \13926 , \573 , \585 );
and \U$13584 ( \13927 , \13925 , \13926 );
not \U$13585 ( \13928 , \13925 );
not \U$13586 ( \13929 , \13926 );
and \U$13587 ( \13930 , \13928 , \13929 );
nor \U$13588 ( \13931 , \13927 , \13930 );
not \U$13589 ( \13932 , \13931 );
not \U$13590 ( \13933 , \13932 );
not \U$13591 ( \13934 , \13933 );
or \U$13592 ( \13935 , \13934 , \9723 );
and \U$13593 ( \13936 , \13914 , \13935 );
not \U$13594 ( \13937 , \13914 );
not \U$13595 ( \13938 , \13935 );
and \U$13596 ( \13939 , \13937 , \13938 );
nor \U$13597 ( \13940 , \13936 , \13939 );
not \U$13598 ( \13941 , \13940 );
or \U$13599 ( \13942 , \13900 , \13941 );
not \U$13600 ( \13943 , \13914 );
nand \U$13601 ( \13944 , \13943 , \13938 );
nand \U$13602 ( \13945 , \13942 , \13944 );
not \U$13603 ( \13946 , \13945 );
or \U$13604 ( \13947 , \13889 , \13946 );
not \U$13605 ( \13948 , \13852 );
not \U$13606 ( \13949 , \13851 );
or \U$13607 ( \13950 , \13948 , \13949 );
nand \U$13608 ( \13951 , \13950 , \13887 );
nand \U$13609 ( \13952 , \13947 , \13951 );
and \U$13610 ( \13953 , \13819 , \13952 );
and \U$13611 ( \13954 , \13812 , \13818 );
or \U$13612 ( \13955 , \13953 , \13954 );
xor \U$13613 ( \13956 , \13181 , \13218 );
xor \U$13614 ( \13957 , \13956 , \13144 );
xor \U$13615 ( \13958 , \13955 , \13957 );
xor \U$13616 ( \13959 , \12951 , \12953 );
xor \U$13617 ( \13960 , \13959 , \12956 );
and \U$13618 ( \13961 , \13958 , \13960 );
and \U$13619 ( \13962 , \13955 , \13957 );
or \U$13620 ( \13963 , \13961 , \13962 );
and \U$13621 ( \13964 , \12949 , \12959 );
not \U$13622 ( \13965 , \12949 );
not \U$13623 ( \13966 , \12959 );
and \U$13624 ( \13967 , \13965 , \13966 );
nor \U$13625 ( \13968 , \13964 , \13967 );
xor \U$13626 ( \13969 , \13963 , \13968 );
not \U$13627 ( \13970 , \13969 );
or \U$13628 ( \13971 , \13810 , \13970 );
nand \U$13629 ( \13972 , \13968 , \13963 );
nand \U$13630 ( \13973 , \13971 , \13972 );
not \U$13631 ( \13974 , \13973 );
not \U$13632 ( \13975 , \13974 );
or \U$13633 ( \13976 , \13808 , \13975 );
nand \U$13634 ( \13977 , \13806 , \13973 );
nand \U$13635 ( \13978 , \13976 , \13977 );
not \U$13636 ( \13979 , \13978 );
or \U$13637 ( \13980 , \13801 , \13979 );
nand \U$13638 ( \13981 , \13807 , \13973 );
nand \U$13639 ( \13982 , \13980 , \13981 );
not \U$13640 ( \13983 , \13982 );
buf \U$13641 ( \13984 , \13436 );
not \U$13642 ( \13985 , \13251 );
and \U$13643 ( \13986 , \13984 , \13985 );
not \U$13644 ( \13987 , \13984 );
and \U$13645 ( \13988 , \13987 , \13251 );
nor \U$13646 ( \13989 , \13986 , \13988 );
xor \U$13647 ( \13990 , \13732 , \13735 );
xor \U$13648 ( \13991 , \13990 , \13727 );
not \U$13649 ( \13992 , \13991 );
xor \U$13650 ( \13993 , \13254 , \13428 );
not \U$13651 ( \13994 , \13993 );
and \U$13652 ( \13995 , \13992 , \13994 );
and \U$13653 ( \13996 , \13991 , \13993 );
nor \U$13654 ( \13997 , \13995 , \13996 );
not \U$13655 ( \13998 , \13997 );
not \U$13656 ( \13999 , \3170 );
not \U$13657 ( \14000 , \13038 );
or \U$13658 ( \14001 , \13999 , \14000 );
nand \U$13659 ( \14002 , \13911 , \13033 );
nand \U$13660 ( \14003 , \14001 , \14002 );
not \U$13661 ( \14004 , \14003 );
not \U$13662 ( \14005 , \3467 );
not \U$13663 ( \14006 , \12968 );
or \U$13664 ( \14007 , \14005 , \14006 );
and \U$13665 ( \14008 , RI98726d0_159, \5736 );
not \U$13666 ( \14009 , RI98726d0_159);
and \U$13667 ( \14010 , \14009 , \5325 );
or \U$13668 ( \14011 , \14008 , \14010 );
nand \U$13669 ( \14012 , \14011 , \3465 );
nand \U$13670 ( \14013 , \14007 , \14012 );
not \U$13671 ( \14014 , \14013 );
or \U$13672 ( \14015 , \14004 , \14014 );
or \U$13673 ( \14016 , \14013 , \14003 );
not \U$13674 ( \14017 , \11692 );
and \U$13675 ( \14018 , \1341 , RI9872b80_169);
not \U$13676 ( \14019 , \1341 );
and \U$13677 ( \14020 , \14019 , \9198 );
nor \U$13678 ( \14021 , \14018 , \14020 );
not \U$13679 ( \14022 , \14021 );
or \U$13680 ( \14023 , \14017 , \14022 );
nand \U$13681 ( \14024 , \12984 , \9214 );
nand \U$13682 ( \14025 , \14023 , \14024 );
nand \U$13683 ( \14026 , \14016 , \14025 );
nand \U$13684 ( \14027 , \14015 , \14026 );
not \U$13685 ( \14028 , \7338 );
not \U$13686 ( \14029 , \13188 );
or \U$13687 ( \14030 , \14028 , \14029 );
not \U$13688 ( \14031 , \7333 );
not \U$13689 ( \14032 , \9263 );
not \U$13690 ( \14033 , \14032 );
or \U$13691 ( \14034 , \14031 , \14033 );
nand \U$13692 ( \14035 , \12393 , RI98729a0_165);
nand \U$13693 ( \14036 , \14034 , \14035 );
nand \U$13694 ( \14037 , \14036 , \7325 );
nand \U$13695 ( \14038 , \14030 , \14037 );
not \U$13696 ( \14039 , \10333 );
not \U$13697 ( \14040 , \13201 );
or \U$13698 ( \14041 , \14039 , \14040 );
not \U$13699 ( \14042 , RI9872e50_175);
not \U$13700 ( \14043 , \6585 );
or \U$13701 ( \14044 , \14042 , \14043 );
or \U$13702 ( \14045 , \6585 , RI9872e50_175);
nand \U$13703 ( \14046 , \14044 , \14045 );
nand \U$13704 ( \14047 , \14046 , \9686 );
nand \U$13705 ( \14048 , \14041 , \14047 );
xor \U$13706 ( \14049 , \14038 , \14048 );
not \U$13707 ( \14050 , \6611 );
not \U$13708 ( \14051 , \13135 );
or \U$13709 ( \14052 , \14050 , \14051 );
and \U$13710 ( \14053 , RI98728b0_163, \10235 );
not \U$13711 ( \14054 , RI98728b0_163);
and \U$13712 ( \14055 , \14054 , \6382 );
or \U$13713 ( \14056 , \14053 , \14055 );
nand \U$13714 ( \14057 , \14056 , \6284 );
nand \U$13715 ( \14058 , \14052 , \14057 );
and \U$13716 ( \14059 , \14049 , \14058 );
and \U$13717 ( \14060 , \14038 , \14048 );
or \U$13718 ( \14061 , \14059 , \14060 );
xor \U$13719 ( \14062 , \14027 , \14061 );
not \U$13720 ( \14063 , \8041 );
not \U$13721 ( \14064 , \13014 );
or \U$13722 ( \14065 , \14063 , \14064 );
xor \U$13723 ( \14066 , RI9872a18_166, \6573 );
nand \U$13724 ( \14067 , \14066 , \8029 );
nand \U$13725 ( \14068 , \14065 , \14067 );
not \U$13726 ( \14069 , \11350 );
and \U$13727 ( \14070 , RI98730a8_180, \1126 );
not \U$13728 ( \14071 , RI98730a8_180);
and \U$13729 ( \14072 , \14071 , \2398 );
nor \U$13730 ( \14073 , \14070 , \14072 );
not \U$13731 ( \14074 , \14073 );
or \U$13732 ( \14075 , \14069 , \14074 );
nand \U$13733 ( \14076 , \13027 , \12868 );
nand \U$13734 ( \14077 , \14075 , \14076 );
xor \U$13735 ( \14078 , \14068 , \14077 );
not \U$13736 ( \14079 , \8743 );
not \U$13737 ( \14080 , RI9872f40_177);
and \U$13738 ( \14081 , \9230 , \14080 );
not \U$13739 ( \14082 , \9230 );
and \U$13740 ( \14083 , \14082 , RI9872f40_177);
nor \U$13741 ( \14084 , \14081 , \14083 );
not \U$13742 ( \14085 , \14084 );
or \U$13743 ( \14086 , \14079 , \14085 );
nand \U$13744 ( \14087 , \13211 , \8752 );
nand \U$13745 ( \14088 , \14086 , \14087 );
and \U$13746 ( \14089 , \14078 , \14088 );
and \U$13747 ( \14090 , \14068 , \14077 );
or \U$13748 ( \14091 , \14089 , \14090 );
and \U$13749 ( \14092 , \14062 , \14091 );
and \U$13750 ( \14093 , \14027 , \14061 );
or \U$13751 ( \14094 , \14092 , \14093 );
xor \U$13752 ( \14095 , \13007 , \13005 );
xnor \U$13753 ( \14096 , \14095 , \13045 );
xor \U$13754 ( \14097 , \14094 , \14096 );
xor \U$13755 ( \14098 , \13306 , \13315 );
xor \U$13756 ( \14099 , \14098 , \13326 );
not \U$13757 ( \14100 , \14099 );
xor \U$13758 ( \14101 , \13364 , \13375 );
buf \U$13759 ( \14102 , \13354 );
xnor \U$13760 ( \14103 , \14101 , \14102 );
nand \U$13761 ( \14104 , \14100 , \14103 );
not \U$13762 ( \14105 , \14104 );
not \U$13763 ( \14106 , \5642 );
and \U$13764 ( \14107 , RI9872568_156, \5885 );
not \U$13765 ( \14108 , RI9872568_156);
and \U$13766 ( \14109 , \14108 , \2948 );
or \U$13767 ( \14110 , \14107 , \14109 );
not \U$13768 ( \14111 , \14110 );
or \U$13769 ( \14112 , \14106 , \14111 );
nand \U$13770 ( \14113 , \13125 , \5653 );
nand \U$13771 ( \14114 , \14112 , \14113 );
not \U$13772 ( \14115 , \14114 );
not \U$13773 ( \14116 , \10242 );
not \U$13774 ( \14117 , \13173 );
or \U$13775 ( \14118 , \14116 , \14117 );
and \U$13776 ( \14119 , RI9872d60_173, \8006 );
not \U$13777 ( \14120 , RI9872d60_173);
and \U$13778 ( \14121 , \14120 , \8005 );
or \U$13779 ( \14122 , \14119 , \14121 );
nand \U$13780 ( \14123 , \14122 , \9312 );
nand \U$13781 ( \14124 , \14118 , \14123 );
not \U$13782 ( \14125 , \14124 );
or \U$13783 ( \14126 , \14115 , \14125 );
xor \U$13784 ( \14127 , \14114 , \14124 );
not \U$13785 ( \14128 , \9952 );
not \U$13786 ( \14129 , RI9873030_179);
not \U$13787 ( \14130 , \1416 );
or \U$13788 ( \14131 , \14129 , \14130 );
not \U$13789 ( \14132 , RI9873030_179);
nand \U$13790 ( \14133 , \10144 , \14132 );
nand \U$13791 ( \14134 , \14131 , \14133 );
not \U$13792 ( \14135 , \14134 );
or \U$13793 ( \14136 , \14128 , \14135 );
nand \U$13794 ( \14137 , \13114 , \9937 );
nand \U$13795 ( \14138 , \14136 , \14137 );
nand \U$13796 ( \14139 , \14127 , \14138 );
nand \U$13797 ( \14140 , \14126 , \14139 );
not \U$13798 ( \14141 , \14140 );
or \U$13799 ( \14142 , \14105 , \14141 );
not \U$13800 ( \14143 , \14103 );
nand \U$13801 ( \14144 , \14143 , \14099 );
nand \U$13802 ( \14145 , \14142 , \14144 );
and \U$13803 ( \14146 , \14097 , \14145 );
and \U$13804 ( \14147 , \14094 , \14096 );
or \U$13805 ( \14148 , \14146 , \14147 );
xor \U$13806 ( \14149 , \13232 , \13049 );
xor \U$13807 ( \14150 , \14148 , \14149 );
xor \U$13808 ( \14151 , \13130 , \13118 );
xnor \U$13809 ( \14152 , \14151 , \13139 );
xor \U$13810 ( \14153 , \13153 , \13165 );
xnor \U$13811 ( \14154 , \14153 , \13177 );
nor \U$13812 ( \14155 , \14152 , \14154 );
xor \U$13813 ( \14156 , \13042 , \13019 );
xnor \U$13814 ( \14157 , \14156 , \13031 );
or \U$13815 ( \14158 , \14155 , \14157 );
nand \U$13816 ( \14159 , \14152 , \14154 );
nand \U$13817 ( \14160 , \14158 , \14159 );
xor \U$13818 ( \14161 , \13051 , \13101 );
xor \U$13819 ( \14162 , \14161 , \13104 );
nor \U$13820 ( \14163 , \14160 , \14162 );
not \U$13821 ( \14164 , \5796 );
not \U$13822 ( \14165 , \13151 );
or \U$13823 ( \14166 , \14164 , \14165 );
xor \U$13824 ( \14167 , RI9872478_154, \3537 );
nand \U$13825 ( \14168 , \14167 , \5034 );
nand \U$13826 ( \14169 , \14166 , \14168 );
xor \U$13827 ( \14170 , \13084 , \14169 );
not \U$13828 ( \14171 , \6553 );
and \U$13829 ( \14172 , RI9872388_152, \5596 );
not \U$13830 ( \14173 , RI9872388_152);
and \U$13831 ( \14174 , \14173 , \11029 );
or \U$13832 ( \14175 , \14172 , \14174 );
not \U$13833 ( \14176 , \14175 );
or \U$13834 ( \14177 , \14171 , \14176 );
nand \U$13835 ( \14178 , \13160 , \4925 );
nand \U$13836 ( \14179 , \14177 , \14178 );
and \U$13837 ( \14180 , \14170 , \14179 );
and \U$13838 ( \14181 , \13084 , \14169 );
or \U$13839 ( \14182 , \14180 , \14181 );
xor \U$13840 ( \14183 , \8679 , \13625 );
not \U$13841 ( \14184 , \14183 );
not \U$13842 ( \14185 , \1162 );
or \U$13843 ( \14186 , \14184 , \14185 );
nand \U$13844 ( \14187 , \1220 , \13633 );
nand \U$13845 ( \14188 , \14186 , \14187 );
not \U$13846 ( \14189 , \1018 );
not \U$13847 ( \14190 , \1042 );
not \U$13848 ( \14191 , \12773 );
or \U$13849 ( \14192 , \14190 , \14191 );
not \U$13850 ( \14193 , \13268 );
nand \U$13851 ( \14194 , \14193 , \3271 );
nand \U$13852 ( \14195 , \14192 , \14194 );
not \U$13853 ( \14196 , \14195 );
or \U$13854 ( \14197 , \14189 , \14196 );
nand \U$13855 ( \14198 , \13603 , \1013 );
nand \U$13856 ( \14199 , \14197 , \14198 );
xor \U$13857 ( \14200 , \14188 , \14199 );
not \U$13858 ( \14201 , \859 );
and \U$13859 ( \14202 , \1347 , \9722 );
not \U$13860 ( \14203 , \1347 );
and \U$13861 ( \14204 , \14203 , \11370 );
nor \U$13862 ( \14205 , \14202 , \14204 );
not \U$13863 ( \14206 , \14205 );
or \U$13864 ( \14207 , \14201 , \14206 );
nand \U$13865 ( \14208 , \13465 , \832 );
nand \U$13866 ( \14209 , \14207 , \14208 );
and \U$13867 ( \14210 , \14200 , \14209 );
and \U$13868 ( \14211 , \14188 , \14199 );
nor \U$13869 ( \14212 , \14210 , \14211 );
not \U$13870 ( \14213 , \14212 );
not \U$13871 ( \14214 , \4085 );
not \U$13872 ( \14215 , \13060 );
or \U$13873 ( \14216 , \14214 , \14215 );
xnor \U$13874 ( \14217 , \12971 , RI98725e0_157);
nand \U$13875 ( \14218 , \14217 , \4101 );
nand \U$13876 ( \14219 , \14216 , \14218 );
not \U$13877 ( \14220 , \14219 );
not \U$13878 ( \14221 , \14220 );
or \U$13879 ( \14222 , \14213 , \14221 );
not \U$13880 ( \14223 , \10487 );
not \U$13881 ( \14224 , \13094 );
or \U$13882 ( \14225 , \14223 , \14224 );
not \U$13883 ( \14226 , \9244 );
not \U$13884 ( \14227 , \944 );
or \U$13885 ( \14228 , \14226 , \14227 );
or \U$13886 ( \14229 , \3836 , \9244 );
nand \U$13887 ( \14230 , \14228 , \14229 );
nand \U$13888 ( \14231 , \14230 , \9670 );
nand \U$13889 ( \14232 , \14225 , \14231 );
nand \U$13890 ( \14233 , \14222 , \14232 );
not \U$13891 ( \14234 , \14212 );
nand \U$13892 ( \14235 , \14234 , \14219 );
nand \U$13893 ( \14236 , \14233 , \14235 );
xor \U$13894 ( \14237 , \14182 , \14236 );
xor \U$13895 ( \14238 , \13084 , \13062 );
xnor \U$13896 ( \14239 , \14238 , \13096 );
and \U$13897 ( \14240 , \14237 , \14239 );
and \U$13898 ( \14241 , \14182 , \14236 );
or \U$13899 ( \14242 , \14240 , \14241 );
not \U$13900 ( \14243 , \14242 );
or \U$13901 ( \14244 , \14163 , \14243 );
nand \U$13902 ( \14245 , \14160 , \14162 );
nand \U$13903 ( \14246 , \14244 , \14245 );
and \U$13904 ( \14247 , \14150 , \14246 );
and \U$13905 ( \14248 , \14148 , \14149 );
or \U$13906 ( \14249 , \14247 , \14248 );
not \U$13907 ( \14250 , \14249 );
not \U$13908 ( \14251 , \14250 );
and \U$13909 ( \14252 , \13998 , \14251 );
not \U$13910 ( \14253 , \13993 );
nor \U$13911 ( \14254 , \14253 , \13991 );
nor \U$13912 ( \14255 , \14252 , \14254 );
nand \U$13913 ( \14256 , \13989 , \14255 );
not \U$13914 ( \14257 , \14256 );
or \U$13915 ( \14258 , \13983 , \14257 );
not \U$13916 ( \14259 , \13989 );
not \U$13917 ( \14260 , \14255 );
nand \U$13918 ( \14261 , \14259 , \14260 );
nand \U$13919 ( \14262 , \14258 , \14261 );
nand \U$13920 ( \14263 , \13799 , \14262 );
nand \U$13921 ( \14264 , \13798 , \14263 );
not \U$13922 ( \14265 , \14264 );
nand \U$13923 ( \14266 , \13792 , \14265 );
nand \U$13924 ( \14267 , \13790 , \14266 );
not \U$13925 ( \14268 , \14267 );
xor \U$13926 ( \14269 , \10364 , \11883 );
xnor \U$13927 ( \14270 , \14269 , \11331 );
not \U$13928 ( \14271 , \12927 );
buf \U$13929 ( \14272 , \12369 );
xnor \U$13930 ( \14273 , \14272 , \12925 );
not \U$13931 ( \14274 , \14273 );
or \U$13932 ( \14275 , \14271 , \14274 );
nand \U$13933 ( \14276 , \12924 , \14272 );
nand \U$13934 ( \14277 , \14275 , \14276 );
nor \U$13935 ( \14278 , \14270 , \14277 );
not \U$13936 ( \14279 , \14278 );
and \U$13937 ( \14280 , \12367 , \14268 , \14279 );
not \U$13938 ( \14281 , \11982 );
not \U$13939 ( \14282 , \11995 );
or \U$13940 ( \14283 , \14281 , \14282 );
nand \U$13941 ( \14284 , \11990 , \11994 );
nand \U$13942 ( \14285 , \14283 , \14284 );
not \U$13943 ( \14286 , \14285 );
not \U$13944 ( \14287 , \11954 );
nand \U$13945 ( \14288 , \14287 , \11904 );
and \U$13946 ( \14289 , \14288 , \11935 );
nor \U$13947 ( \14290 , \14287 , \11904 );
nor \U$13948 ( \14291 , \14289 , \14290 );
not \U$13949 ( \14292 , \11946 );
xnor \U$13950 ( \14293 , \11953 , \11940 );
not \U$13951 ( \14294 , \14293 );
or \U$13952 ( \14295 , \14292 , \14294 );
not \U$13953 ( \14296 , \11940 );
nand \U$13954 ( \14297 , \14296 , \11953 );
nand \U$13955 ( \14298 , \14295 , \14297 );
or \U$13956 ( \14299 , \12290 , \1293 );
and \U$13957 ( \14300 , RI9871b18_134, \4986 );
not \U$13958 ( \14301 , RI9871b18_134);
and \U$13959 ( \14302 , \14301 , \5739 );
nor \U$13960 ( \14303 , \14300 , \14302 );
or \U$13961 ( \14304 , \14303 , \1543 );
nand \U$13962 ( \14305 , \14299 , \14304 );
not \U$13963 ( \14306 , \1455 );
not \U$13964 ( \14307 , \12247 );
or \U$13965 ( \14308 , \14306 , \14307 );
xnor \U$13966 ( \14309 , \4471 , RI9871c08_136);
nand \U$13967 ( \14310 , \14309 , \1430 );
nand \U$13968 ( \14311 , \14308 , \14310 );
xor \U$13969 ( \14312 , \14305 , \14311 );
not \U$13970 ( \14313 , \9670 );
not \U$13971 ( \14314 , \12312 );
or \U$13972 ( \14315 , \14313 , \14314 );
not \U$13973 ( \14316 , \9185 );
not \U$13974 ( \14317 , \1692 );
or \U$13975 ( \14318 , \14316 , \14317 );
or \U$13976 ( \14319 , \7330 , \9244 );
nand \U$13977 ( \14320 , \14318 , \14319 );
nand \U$13978 ( \14321 , \14320 , \10487 );
nand \U$13979 ( \14322 , \14315 , \14321 );
xnor \U$13980 ( \14323 , \14312 , \14322 );
not \U$13981 ( \14324 , \14323 );
not \U$13982 ( \14325 , \3466 );
not \U$13983 ( \14326 , \12277 );
or \U$13984 ( \14327 , \14325 , \14326 );
and \U$13985 ( \14328 , RI98726d0_159, \7604 );
not \U$13986 ( \14329 , RI98726d0_159);
and \U$13987 ( \14330 , \14329 , \1211 );
or \U$13988 ( \14331 , \14328 , \14330 );
nand \U$13989 ( \14332 , \14331 , \3467 );
nand \U$13990 ( \14333 , \14327 , \14332 );
not \U$13991 ( \14334 , \9214 );
not \U$13992 ( \14335 , RI9872b80_169);
not \U$13993 ( \14336 , \1724 );
or \U$13994 ( \14337 , \14335 , \14336 );
or \U$13995 ( \14338 , \9276 , RI9872b80_169);
nand \U$13996 ( \14339 , \14337 , \14338 );
not \U$13997 ( \14340 , \14339 );
or \U$13998 ( \14341 , \14334 , \14340 );
nand \U$13999 ( \14342 , \12269 , \10679 );
nand \U$14000 ( \14343 , \14341 , \14342 );
not \U$14001 ( \14344 , \14343 );
and \U$14002 ( \14345 , \14333 , \14344 );
not \U$14003 ( \14346 , \14333 );
and \U$14004 ( \14347 , \14346 , \14343 );
nor \U$14005 ( \14348 , \14345 , \14347 );
not \U$14006 ( \14349 , \7325 );
not \U$14007 ( \14350 , \12215 );
or \U$14008 ( \14351 , \14349 , \14350 );
and \U$14009 ( \14352 , RI98729a0_165, \1309 );
not \U$14010 ( \14353 , RI98729a0_165);
and \U$14011 ( \14354 , \14353 , \1320 );
nor \U$14012 ( \14355 , \14352 , \14354 );
nand \U$14013 ( \14356 , \14355 , \7338 );
nand \U$14014 ( \14357 , \14351 , \14356 );
not \U$14015 ( \14358 , \14357 );
and \U$14016 ( \14359 , \14348 , \14358 );
not \U$14017 ( \14360 , \14348 );
and \U$14018 ( \14361 , \14360 , \14357 );
nor \U$14019 ( \14362 , \14359 , \14361 );
not \U$14020 ( \14363 , \14362 );
or \U$14021 ( \14364 , \14324 , \14363 );
or \U$14022 ( \14365 , \14362 , \14323 );
nand \U$14023 ( \14366 , \14364 , \14365 );
xor \U$14024 ( \14367 , \14298 , \14366 );
xor \U$14025 ( \14368 , \14291 , \14367 );
xor \U$14026 ( \14369 , \14286 , \14368 );
not \U$14027 ( \14370 , \12009 );
not \U$14028 ( \14371 , \12067 );
or \U$14029 ( \14372 , \14370 , \14371 );
nand \U$14030 ( \14373 , \12008 , \11999 );
nand \U$14031 ( \14374 , \14372 , \14373 );
xor \U$14032 ( \14375 , \14369 , \14374 );
not \U$14033 ( \14376 , \12183 );
not \U$14034 ( \14377 , \12225 );
nand \U$14035 ( \14378 , \14377 , \12189 );
not \U$14036 ( \14379 , \14378 );
or \U$14037 ( \14380 , \14376 , \14379 );
nand \U$14038 ( \14381 , \12225 , \12188 );
nand \U$14039 ( \14382 , \14380 , \14381 );
buf \U$14040 ( \14383 , \12160 );
and \U$14041 ( \14384 , \14383 , \1501 );
xor \U$14042 ( \14385 , \5766 , RI9871c80_137);
and \U$14043 ( \14386 , \14385 , \1518 );
nor \U$14044 ( \14387 , \14384 , \14386 );
not \U$14045 ( \14388 , \876 );
not \U$14046 ( \14389 , \12100 );
or \U$14047 ( \14390 , \14388 , \14389 );
and \U$14048 ( \14391 , RI9872130_147, \12802 );
not \U$14049 ( \14392 , RI9872130_147);
and \U$14050 ( \14393 , \14392 , \8054 );
nor \U$14051 ( \14394 , \14391 , \14393 );
nand \U$14052 ( \14395 , \14394 , \924 );
nand \U$14053 ( \14396 , \14390 , \14395 );
nand \U$14054 ( \14397 , RI9872dd8_174, RI9872e50_175);
and \U$14055 ( \14398 , \14397 , RI9872d60_173);
and \U$14056 ( \14399 , \14396 , \14398 );
not \U$14057 ( \14400 , \14396 );
not \U$14058 ( \14401 , \14398 );
and \U$14059 ( \14402 , \14400 , \14401 );
or \U$14060 ( \14403 , \14399 , \14402 );
xnor \U$14061 ( \14404 , \14387 , \14403 );
not \U$14062 ( \14405 , \12251 );
not \U$14063 ( \14406 , \12242 );
not \U$14064 ( \14407 , \14406 );
or \U$14065 ( \14408 , \14405 , \14407 );
not \U$14066 ( \14409 , \12241 );
nand \U$14067 ( \14410 , \14409 , \12240 );
nand \U$14068 ( \14411 , \14408 , \14410 );
xor \U$14069 ( \14412 , \14404 , \14411 );
xor \U$14070 ( \14413 , \12262 , \12271 );
and \U$14071 ( \14414 , \14413 , \12281 );
and \U$14072 ( \14415 , \12262 , \12271 );
or \U$14073 ( \14416 , \14414 , \14415 );
xor \U$14074 ( \14417 , \14412 , \14416 );
xnor \U$14075 ( \14418 , \14382 , \14417 );
not \U$14076 ( \14419 , \12315 );
not \U$14077 ( \14420 , \12286 );
or \U$14078 ( \14421 , \14419 , \14420 );
not \U$14079 ( \14422 , \12252 );
nand \U$14080 ( \14423 , \14422 , \12282 );
nand \U$14081 ( \14424 , \14421 , \14423 );
and \U$14082 ( \14425 , \14418 , \14424 );
not \U$14083 ( \14426 , \14418 );
not \U$14084 ( \14427 , \14424 );
and \U$14085 ( \14428 , \14426 , \14427 );
nor \U$14086 ( \14429 , \14425 , \14428 );
not \U$14087 ( \14430 , \12133 );
not \U$14088 ( \14431 , \12120 );
or \U$14089 ( \14432 , \14430 , \14431 );
nand \U$14090 ( \14433 , \12104 , \12115 );
nand \U$14091 ( \14434 , \14432 , \14433 );
buf \U$14092 ( \14435 , \12165 );
not \U$14093 ( \14436 , \14435 );
and \U$14094 ( \14437 , \14434 , \14436 );
not \U$14095 ( \14438 , \14434 );
and \U$14096 ( \14439 , \14438 , \14435 );
nor \U$14097 ( \14440 , \14437 , \14439 );
not \U$14098 ( \14441 , \12032 );
or \U$14099 ( \14442 , \12038 , \12022 );
not \U$14100 ( \14443 , \14442 );
or \U$14101 ( \14444 , \14441 , \14443 );
nand \U$14102 ( \14445 , \12038 , \12022 );
nand \U$14103 ( \14446 , \14444 , \14445 );
xnor \U$14104 ( \14447 , \14440 , \14446 );
not \U$14105 ( \14448 , \14447 );
not \U$14106 ( \14449 , \12048 );
not \U$14107 ( \14450 , \12054 );
or \U$14108 ( \14451 , \14449 , \14450 );
not \U$14109 ( \14452 , \12039 );
nand \U$14110 ( \14453 , \14452 , \12044 );
nand \U$14111 ( \14454 , \14451 , \14453 );
not \U$14112 ( \14455 , \14454 );
or \U$14113 ( \14456 , \14448 , \14455 );
or \U$14114 ( \14457 , \14454 , \14447 );
nand \U$14115 ( \14458 , \14456 , \14457 );
not \U$14116 ( \14459 , \12138 );
not \U$14117 ( \14460 , \14459 );
not \U$14118 ( \14461 , \12089 );
or \U$14119 ( \14462 , \14460 , \14461 );
not \U$14120 ( \14463 , \12134 );
nand \U$14121 ( \14464 , \14463 , \12094 );
nand \U$14122 ( \14465 , \14462 , \14464 );
not \U$14123 ( \14466 , \14465 );
and \U$14124 ( \14467 , \14458 , \14466 );
not \U$14125 ( \14468 , \14458 );
and \U$14126 ( \14469 , \14468 , \14465 );
nor \U$14127 ( \14470 , \14467 , \14469 );
not \U$14128 ( \14471 , \14470 );
xor \U$14129 ( \14472 , \14429 , \14471 );
not \U$14130 ( \14473 , \12016 );
xnor \U$14131 ( \14474 , \12065 , \12059 );
not \U$14132 ( \14475 , \14474 );
or \U$14133 ( \14476 , \14473 , \14475 );
not \U$14134 ( \14477 , \12059 );
nand \U$14135 ( \14478 , \14477 , \12066 );
nand \U$14136 ( \14479 , \14476 , \14478 );
xnor \U$14137 ( \14480 , \14472 , \14479 );
xor \U$14138 ( \14481 , \14375 , \14480 );
not \U$14139 ( \14482 , \12322 );
not \U$14140 ( \14483 , \12330 );
or \U$14141 ( \14484 , \14482 , \14483 );
not \U$14142 ( \14485 , \12327 );
not \U$14143 ( \14486 , \12321 );
or \U$14144 ( \14487 , \14485 , \14486 );
nand \U$14145 ( \14488 , \14487 , \12338 );
nand \U$14146 ( \14489 , \14484 , \14488 );
not \U$14147 ( \14490 , \14489 );
not \U$14148 ( \14491 , \4919 );
not \U$14149 ( \14492 , \12299 );
or \U$14150 ( \14493 , \14491 , \14492 );
and \U$14151 ( \14494 , RI9872388_152, \1344 );
not \U$14152 ( \14495 , RI9872388_152);
and \U$14153 ( \14496 , \14495 , \1341 );
or \U$14154 ( \14497 , \14494 , \14496 );
nand \U$14155 ( \14498 , \14497 , \4925 );
nand \U$14156 ( \14499 , \14493 , \14498 );
not \U$14157 ( \14500 , \5530 );
not \U$14158 ( \14501 , \12195 );
or \U$14159 ( \14502 , \14500 , \14501 );
not \U$14160 ( \14503 , \4088 );
not \U$14161 ( \14504 , \1062 );
or \U$14162 ( \14505 , \14503 , \14504 );
or \U$14163 ( \14506 , \10133 , \4088 );
nand \U$14164 ( \14507 , \14505 , \14506 );
nand \U$14165 ( \14508 , \14507 , \5847 );
nand \U$14166 ( \14509 , \14502 , \14508 );
xor \U$14167 ( \14510 , \14499 , \14509 );
not \U$14168 ( \14511 , \8029 );
not \U$14169 ( \14512 , \12205 );
or \U$14170 ( \14513 , \14511 , \14512 );
not \U$14171 ( \14514 , RI9872a18_166);
not \U$14172 ( \14515 , \6174 );
or \U$14173 ( \14516 , \14514 , \14515 );
or \U$14174 ( \14517 , \1416 , RI9872a18_166);
nand \U$14175 ( \14518 , \14516 , \14517 );
nand \U$14176 ( \14519 , \14518 , \9072 );
nand \U$14177 ( \14520 , \14513 , \14519 );
xor \U$14178 ( \14521 , \14510 , \14520 );
not \U$14179 ( \14522 , \2087 );
and \U$14180 ( \14523 , RI9871aa0_133, \2948 );
not \U$14181 ( \14524 , RI9871aa0_133);
and \U$14182 ( \14525 , \14524 , \3691 );
nor \U$14183 ( \14526 , \14523 , \14525 );
not \U$14184 ( \14527 , \14526 );
or \U$14185 ( \14528 , \14522 , \14527 );
or \U$14186 ( \14529 , \11909 , \2073 );
nand \U$14187 ( \14530 , \14528 , \14529 );
not \U$14188 ( \14531 , \3164 );
not \U$14189 ( \14532 , \12258 );
or \U$14190 ( \14533 , \14531 , \14532 );
xor \U$14191 ( \14534 , \6382 , RI9872310_151);
nand \U$14192 ( \14535 , \14534 , \3170 );
nand \U$14193 ( \14536 , \14533 , \14535 );
xor \U$14194 ( \14537 , \14530 , \14536 );
not \U$14195 ( \14538 , \6284 );
not \U$14196 ( \14539 , \11930 );
or \U$14197 ( \14540 , \14538 , \14539 );
not \U$14198 ( \14541 , RI98728b0_163);
not \U$14199 ( \14542 , \916 );
or \U$14200 ( \14543 , \14541 , \14542 );
or \U$14201 ( \14544 , \5480 , RI98728b0_163);
nand \U$14202 ( \14545 , \14543 , \14544 );
nand \U$14203 ( \14546 , \14545 , \6611 );
nand \U$14204 ( \14547 , \14540 , \14546 );
xor \U$14205 ( \14548 , \14537 , \14547 );
xor \U$14206 ( \14549 , \14521 , \14548 );
not \U$14207 ( \14550 , \793 );
not \U$14208 ( \14551 , \12176 );
or \U$14209 ( \14552 , \14550 , \14551 );
not \U$14210 ( \14553 , \1078 );
not \U$14211 ( \14554 , \3537 );
or \U$14212 ( \14555 , \14553 , \14554 );
or \U$14213 ( \14556 , \3543 , \1078 );
nand \U$14214 ( \14557 , \14555 , \14556 );
nand \U$14215 ( \14558 , \14557 , \796 );
nand \U$14216 ( \14559 , \14552 , \14558 );
not \U$14217 ( \14560 , \6673 );
not \U$14218 ( \14561 , RI98718c0_129);
not \U$14219 ( \14562 , \4177 );
not \U$14220 ( \14563 , \14562 );
or \U$14221 ( \14564 , \14561 , \14563 );
or \U$14222 ( \14565 , \12616 , RI98718c0_129);
nand \U$14223 ( \14566 , \14564 , \14565 );
not \U$14224 ( \14567 , \14566 );
or \U$14225 ( \14568 , \14560 , \14567 );
nand \U$14226 ( \14569 , \12146 , \1083 );
nand \U$14227 ( \14570 , \14568 , \14569 );
not \U$14228 ( \14571 , \14570 );
xor \U$14229 ( \14572 , \14559 , \14571 );
not \U$14230 ( \14573 , \7188 );
and \U$14231 ( \14574 , RI9872568_156, \8006 );
not \U$14232 ( \14575 , RI9872568_156);
and \U$14233 ( \14576 , \14575 , \821 );
or \U$14234 ( \14577 , \14574 , \14576 );
not \U$14235 ( \14578 , \14577 );
or \U$14236 ( \14579 , \14573 , \14578 );
nand \U$14237 ( \14580 , \11919 , \5642 );
nand \U$14238 ( \14581 , \14579 , \14580 );
xnor \U$14239 ( \14582 , \14572 , \14581 );
xor \U$14240 ( \14583 , \14549 , \14582 );
not \U$14241 ( \14584 , \14583 );
and \U$14242 ( \14585 , \12028 , \1018 );
xor \U$14243 ( \14586 , \3271 , \8624 );
and \U$14244 ( \14587 , \14586 , \1067 );
nor \U$14245 ( \14588 , \14585 , \14587 );
not \U$14246 ( \14589 , \14588 );
not \U$14247 ( \14590 , \832 );
not \U$14248 ( \14591 , \10583 );
xor \U$14249 ( \14592 , RI9871d70_139, \14591 );
not \U$14250 ( \14593 , \14592 );
or \U$14251 ( \14594 , \14590 , \14593 );
nand \U$14252 ( \14595 , \12113 , \859 );
nand \U$14253 ( \14596 , \14594 , \14595 );
not \U$14254 ( \14597 , \14596 );
not \U$14255 ( \14598 , \1381 );
not \U$14256 ( \14599 , \12128 );
or \U$14257 ( \14600 , \14598 , \14599 );
and \U$14258 ( \14601 , RI9871e60_141, \9895 );
not \U$14259 ( \14602 , RI9871e60_141);
and \U$14260 ( \14603 , \14602 , \8916 );
or \U$14261 ( \14604 , \14601 , \14603 );
nand \U$14262 ( \14605 , \14604 , \1352 );
nand \U$14263 ( \14606 , \14600 , \14605 );
not \U$14264 ( \14607 , \14606 );
not \U$14265 ( \14608 , \14607 );
or \U$14266 ( \14609 , \14597 , \14608 );
or \U$14267 ( \14610 , \14607 , \14596 );
nand \U$14268 ( \14611 , \14609 , \14610 );
not \U$14269 ( \14612 , \14611 );
or \U$14270 ( \14613 , \14589 , \14612 );
or \U$14271 ( \14614 , \14588 , \14611 );
nand \U$14272 ( \14615 , \14613 , \14614 );
and \U$14273 ( \14616 , \1165 , \8575 );
not \U$14274 ( \14617 , \1162 );
not \U$14275 ( \14618 , \12018 );
or \U$14276 ( \14619 , \14617 , \14618 );
xor \U$14277 ( \14620 , \1716 , \8858 );
not \U$14278 ( \14621 , \14620 );
nand \U$14279 ( \14622 , \14621 , \6316 );
nand \U$14280 ( \14623 , \14619 , \14622 );
xor \U$14281 ( \14624 , \14616 , \14623 );
not \U$14282 ( \14625 , \5796 );
xor \U$14283 ( \14626 , RI9872478_154, \944 );
not \U$14284 ( \14627 , \14626 );
or \U$14285 ( \14628 , \14625 , \14627 );
nand \U$14286 ( \14629 , \12238 , \5034 );
nand \U$14287 ( \14630 , \14628 , \14629 );
xor \U$14288 ( \14631 , \14624 , \14630 );
xor \U$14289 ( \14632 , \14615 , \14631 );
xor \U$14290 ( \14633 , \11913 , \11923 );
and \U$14291 ( \14634 , \14633 , \11934 );
and \U$14292 ( \14635 , \11913 , \11923 );
or \U$14293 ( \14636 , \14634 , \14635 );
xor \U$14294 ( \14637 , \14632 , \14636 );
not \U$14295 ( \14638 , \12178 );
not \U$14296 ( \14639 , \12169 );
or \U$14297 ( \14640 , \14638 , \14639 );
nand \U$14298 ( \14641 , \12150 , \14435 );
nand \U$14299 ( \14642 , \14640 , \14641 );
xor \U$14300 ( \14643 , \12293 , \12303 );
and \U$14301 ( \14644 , \14643 , \12314 );
and \U$14302 ( \14645 , \12293 , \12303 );
or \U$14303 ( \14646 , \14644 , \14645 );
xor \U$14304 ( \14647 , \14642 , \14646 );
not \U$14305 ( \14648 , \12199 );
not \U$14306 ( \14649 , \12224 );
or \U$14307 ( \14650 , \14648 , \14649 );
nand \U$14308 ( \14651 , \12209 , \12219 );
nand \U$14309 ( \14652 , \14650 , \14651 );
xor \U$14310 ( \14653 , \14647 , \14652 );
xnor \U$14311 ( \14654 , \14637 , \14653 );
not \U$14312 ( \14655 , \14654 );
or \U$14313 ( \14656 , \14584 , \14655 );
not \U$14314 ( \14657 , \14654 );
not \U$14315 ( \14658 , \14583 );
nand \U$14316 ( \14659 , \14657 , \14658 );
nand \U$14317 ( \14660 , \14656 , \14659 );
or \U$14318 ( \14661 , \11901 , \11955 );
nand \U$14319 ( \14662 , \14661 , \11965 );
nand \U$14320 ( \14663 , \11901 , \11955 );
nand \U$14321 ( \14664 , \14662 , \14663 );
not \U$14322 ( \14665 , \14664 );
xor \U$14323 ( \14666 , \14660 , \14665 );
not \U$14324 ( \14667 , \12316 );
not \U$14325 ( \14668 , \12230 );
or \U$14326 ( \14669 , \14667 , \14668 );
not \U$14327 ( \14670 , \12142 );
nand \U$14328 ( \14671 , \14670 , \12226 );
nand \U$14329 ( \14672 , \14669 , \14671 );
not \U$14330 ( \14673 , \14672 );
xnor \U$14331 ( \14674 , \14666 , \14673 );
not \U$14332 ( \14675 , \14674 );
or \U$14333 ( \14676 , \14490 , \14675 );
or \U$14334 ( \14677 , \14674 , \14489 );
nand \U$14335 ( \14678 , \14676 , \14677 );
xor \U$14336 ( \14679 , \11967 , \11974 );
and \U$14337 ( \14680 , \14679 , \12068 );
and \U$14338 ( \14681 , \11967 , \11974 );
or \U$14339 ( \14682 , \14680 , \14681 );
xor \U$14340 ( \14683 , \14678 , \14682 );
xor \U$14341 ( \14684 , \14481 , \14683 );
not \U$14342 ( \14685 , \12352 );
not \U$14343 ( \14686 , \12078 );
nand \U$14344 ( \14687 , \14686 , \12343 );
not \U$14345 ( \14688 , \14687 );
or \U$14346 ( \14689 , \14685 , \14688 );
not \U$14347 ( \14690 , \12343 );
nand \U$14348 ( \14691 , \14690 , \12078 );
nand \U$14349 ( \14692 , \14689 , \14691 );
and \U$14350 ( \14693 , \14684 , \14692 );
and \U$14351 ( \14694 , \14481 , \14683 );
nor \U$14352 ( \14695 , \14693 , \14694 );
not \U$14353 ( \14696 , \14695 );
or \U$14354 ( \14697 , \14368 , \14286 );
not \U$14355 ( \14698 , \14291 );
nand \U$14356 ( \14699 , \14698 , \14367 );
nand \U$14357 ( \14700 , \14697 , \14699 );
not \U$14358 ( \14701 , \14653 );
not \U$14359 ( \14702 , \14637 );
or \U$14360 ( \14703 , \14701 , \14702 );
or \U$14361 ( \14704 , \14637 , \14653 );
nand \U$14362 ( \14705 , \14704 , \14583 );
nand \U$14363 ( \14706 , \14703 , \14705 );
not \U$14364 ( \14707 , \14706 );
xor \U$14365 ( \14708 , \14615 , \14631 );
and \U$14366 ( \14709 , \14708 , \14636 );
and \U$14367 ( \14710 , \14615 , \14631 );
or \U$14368 ( \14711 , \14709 , \14710 );
not \U$14369 ( \14712 , \14387 );
not \U$14370 ( \14713 , \14712 );
not \U$14371 ( \14714 , \14403 );
or \U$14372 ( \14715 , \14713 , \14714 );
nand \U$14373 ( \14716 , \14396 , \14401 );
nand \U$14374 ( \14717 , \14715 , \14716 );
not \U$14375 ( \14718 , \1430 );
and \U$14376 ( \14719 , \5615 , RI9871c08_136);
not \U$14377 ( \14720 , \5615 );
and \U$14378 ( \14721 , \14720 , \1850 );
nor \U$14379 ( \14722 , \14719 , \14721 );
not \U$14380 ( \14723 , \14722 );
or \U$14381 ( \14724 , \14718 , \14723 );
nand \U$14382 ( \14725 , \14309 , \1455 );
nand \U$14383 ( \14726 , \14724 , \14725 );
not \U$14384 ( \14727 , \924 );
not \U$14385 ( \14728 , RI9872130_147);
not \U$14386 ( \14729 , \5707 );
or \U$14387 ( \14730 , \14728 , \14729 );
or \U$14388 ( \14731 , \5707 , RI9872130_147);
nand \U$14389 ( \14732 , \14730 , \14731 );
not \U$14390 ( \14733 , \14732 );
or \U$14391 ( \14734 , \14727 , \14733 );
nand \U$14392 ( \14735 , \14394 , \876 );
nand \U$14393 ( \14736 , \14734 , \14735 );
not \U$14394 ( \14737 , \14736 );
not \U$14395 ( \14738 , \14737 );
and \U$14396 ( \14739 , \14726 , \14738 );
not \U$14397 ( \14740 , \14726 );
and \U$14398 ( \14741 , \14740 , \14737 );
nor \U$14399 ( \14742 , \14739 , \14741 );
not \U$14400 ( \14743 , \14742 );
and \U$14401 ( \14744 , \14717 , \14743 );
not \U$14402 ( \14745 , \14717 );
and \U$14403 ( \14746 , \14745 , \14742 );
nor \U$14404 ( \14747 , \14744 , \14746 );
and \U$14405 ( \14748 , \14711 , \14747 );
not \U$14406 ( \14749 , \14711 );
not \U$14407 ( \14750 , \14747 );
and \U$14408 ( \14751 , \14749 , \14750 );
or \U$14409 ( \14752 , \14748 , \14751 );
not \U$14410 ( \14753 , \14752 );
xor \U$14411 ( \14754 , \14404 , \14411 );
and \U$14412 ( \14755 , \14754 , \14416 );
and \U$14413 ( \14756 , \14404 , \14411 );
or \U$14414 ( \14757 , \14755 , \14756 );
not \U$14415 ( \14758 , \14757 );
not \U$14416 ( \14759 , \14758 );
or \U$14417 ( \14760 , \14753 , \14759 );
or \U$14418 ( \14761 , \14752 , \14758 );
nand \U$14419 ( \14762 , \14760 , \14761 );
xor \U$14420 ( \14763 , \14707 , \14762 );
not \U$14421 ( \14764 , \14417 );
not \U$14422 ( \14765 , \14424 );
or \U$14423 ( \14766 , \14764 , \14765 );
or \U$14424 ( \14767 , \14424 , \14417 );
nand \U$14425 ( \14768 , \14767 , \14382 );
nand \U$14426 ( \14769 , \14766 , \14768 );
xor \U$14427 ( \14770 , \14763 , \14769 );
xor \U$14428 ( \14771 , \14700 , \14770 );
not \U$14429 ( \14772 , \14479 );
not \U$14430 ( \14773 , \14470 );
and \U$14431 ( \14774 , \14772 , \14773 );
and \U$14432 ( \14775 , \14479 , \14470 );
nor \U$14433 ( \14776 , \14774 , \14775 );
or \U$14434 ( \14777 , \14776 , \14429 );
nand \U$14435 ( \14778 , \14479 , \14471 );
nand \U$14436 ( \14779 , \14777 , \14778 );
xor \U$14437 ( \14780 , \14771 , \14779 );
not \U$14438 ( \14781 , \14780 );
not \U$14439 ( \14782 , \14682 );
not \U$14440 ( \14783 , \14678 );
or \U$14441 ( \14784 , \14782 , \14783 );
not \U$14442 ( \14785 , \14674 );
nand \U$14443 ( \14786 , \14785 , \14489 );
nand \U$14444 ( \14787 , \14784 , \14786 );
not \U$14445 ( \14788 , \14787 );
not \U$14446 ( \14789 , \14788 );
or \U$14447 ( \14790 , \14781 , \14789 );
or \U$14448 ( \14791 , \14780 , \14788 );
nand \U$14449 ( \14792 , \14790 , \14791 );
xor \U$14450 ( \14793 , \14642 , \14646 );
and \U$14451 ( \14794 , \14793 , \14652 );
and \U$14452 ( \14795 , \14642 , \14646 );
or \U$14453 ( \14796 , \14794 , \14795 );
xor \U$14454 ( \14797 , \14499 , \14509 );
and \U$14455 ( \14798 , \14797 , \14520 );
and \U$14456 ( \14799 , \14499 , \14509 );
or \U$14457 ( \14800 , \14798 , \14799 );
not \U$14458 ( \14801 , \14357 );
not \U$14459 ( \14802 , \14333 );
or \U$14460 ( \14803 , \14801 , \14802 );
or \U$14461 ( \14804 , \14333 , \14357 );
nand \U$14462 ( \14805 , \14804 , \14343 );
nand \U$14463 ( \14806 , \14803 , \14805 );
xor \U$14464 ( \14807 , \14800 , \14806 );
not \U$14465 ( \14808 , \14305 );
not \U$14466 ( \14809 , \14311 );
or \U$14467 ( \14810 , \14808 , \14809 );
or \U$14468 ( \14811 , \14311 , \14305 );
nand \U$14469 ( \14812 , \14811 , \14322 );
nand \U$14470 ( \14813 , \14810 , \14812 );
not \U$14471 ( \14814 , \14813 );
and \U$14472 ( \14815 , \14807 , \14814 );
not \U$14473 ( \14816 , \14807 );
and \U$14474 ( \14817 , \14816 , \14813 );
nor \U$14475 ( \14818 , \14815 , \14817 );
xor \U$14476 ( \14819 , \14796 , \14818 );
not \U$14477 ( \14820 , \14559 );
not \U$14478 ( \14821 , \14571 );
not \U$14479 ( \14822 , \14581 );
or \U$14480 ( \14823 , \14821 , \14822 );
or \U$14481 ( \14824 , \14581 , \14571 );
nand \U$14482 ( \14825 , \14823 , \14824 );
not \U$14483 ( \14826 , \14825 );
or \U$14484 ( \14827 , \14820 , \14826 );
nand \U$14485 ( \14828 , \14581 , \14570 );
nand \U$14486 ( \14829 , \14827 , \14828 );
and \U$14487 ( \14830 , \5753 , \8642 );
not \U$14488 ( \14831 , \9670 );
not \U$14489 ( \14832 , \14320 );
or \U$14490 ( \14833 , \14831 , \14832 );
nand \U$14491 ( \14834 , \9227 , RI9872bf8_170);
nand \U$14492 ( \14835 , \14833 , \14834 );
xor \U$14493 ( \14836 , \14830 , \14835 );
not \U$14494 ( \14837 , \14620 );
not \U$14495 ( \14838 , \1809 );
and \U$14496 ( \14839 , \14837 , \14838 );
not \U$14497 ( \14840 , \8679 );
not \U$14498 ( \14841 , \8607 );
or \U$14499 ( \14842 , \14840 , \14841 );
nand \U$14500 ( \14843 , \8597 , \1716 );
nand \U$14501 ( \14844 , \14842 , \14843 );
and \U$14502 ( \14845 , \14844 , \1220 );
nor \U$14503 ( \14846 , \14839 , \14845 );
not \U$14504 ( \14847 , \14846 );
xor \U$14505 ( \14848 , \14836 , \14847 );
not \U$14506 ( \14849 , \14848 );
not \U$14507 ( \14850 , \14588 );
not \U$14508 ( \14851 , \14850 );
not \U$14509 ( \14852 , \14611 );
or \U$14510 ( \14853 , \14851 , \14852 );
nand \U$14511 ( \14854 , \14606 , \14596 );
nand \U$14512 ( \14855 , \14853 , \14854 );
not \U$14513 ( \14856 , \14855 );
nand \U$14514 ( \14857 , \14849 , \14856 );
not \U$14515 ( \14858 , \14856 );
nand \U$14516 ( \14859 , \14858 , \14848 );
nand \U$14517 ( \14860 , \14857 , \14859 );
xor \U$14518 ( \14861 , \14829 , \14860 );
xnor \U$14519 ( \14862 , \14819 , \14861 );
xor \U$14520 ( \14863 , \14521 , \14548 );
and \U$14521 ( \14864 , \14863 , \14582 );
and \U$14522 ( \14865 , \14521 , \14548 );
or \U$14523 ( \14866 , \14864 , \14865 );
not \U$14524 ( \14867 , \14866 );
not \U$14525 ( \14868 , \14867 );
xor \U$14526 ( \14869 , \14616 , \14623 );
and \U$14527 ( \14870 , \14869 , \14630 );
and \U$14528 ( \14871 , \14616 , \14623 );
or \U$14529 ( \14872 , \14870 , \14871 );
not \U$14530 ( \14873 , \1067 );
and \U$14531 ( \14874 , \3271 , \8074 );
not \U$14532 ( \14875 , \3271 );
and \U$14533 ( \14876 , \14875 , \8075 );
nor \U$14534 ( \14877 , \14874 , \14876 );
not \U$14535 ( \14878 , \14877 );
or \U$14536 ( \14879 , \14873 , \14878 );
nand \U$14537 ( \14880 , \14586 , \1018 );
nand \U$14538 ( \14881 , \14879 , \14880 );
not \U$14539 ( \14882 , \1353 );
not \U$14540 ( \14883 , \1367 );
not \U$14541 ( \14884 , \8925 );
or \U$14542 ( \14885 , \14883 , \14884 );
or \U$14543 ( \14886 , \7467 , \1367 );
nand \U$14544 ( \14887 , \14885 , \14886 );
not \U$14545 ( \14888 , \14887 );
or \U$14546 ( \14889 , \14882 , \14888 );
nand \U$14547 ( \14890 , \14604 , \6195 );
nand \U$14548 ( \14891 , \14889 , \14890 );
xor \U$14549 ( \14892 , \14881 , \14891 );
not \U$14550 ( \14893 , \832 );
not \U$14551 ( \14894 , \12108 );
not \U$14552 ( \14895 , \6530 );
or \U$14553 ( \14896 , \14894 , \14895 );
nand \U$14554 ( \14897 , \6529 , RI9871d70_139);
nand \U$14555 ( \14898 , \14896 , \14897 );
not \U$14556 ( \14899 , \14898 );
or \U$14557 ( \14900 , \14893 , \14899 );
nand \U$14558 ( \14901 , \14592 , \6635 );
nand \U$14559 ( \14902 , \14900 , \14901 );
xor \U$14560 ( \14903 , \14892 , \14902 );
xor \U$14561 ( \14904 , \14872 , \14903 );
xor \U$14562 ( \14905 , \14530 , \14536 );
and \U$14563 ( \14906 , \14905 , \14547 );
and \U$14564 ( \14907 , \14530 , \14536 );
or \U$14565 ( \14908 , \14906 , \14907 );
xnor \U$14566 ( \14909 , \14904 , \14908 );
not \U$14567 ( \14910 , \14909 );
not \U$14568 ( \14911 , \14910 );
or \U$14569 ( \14912 , \14868 , \14911 );
nand \U$14570 ( \14913 , \14909 , \14866 );
nand \U$14571 ( \14914 , \14912 , \14913 );
not \U$14572 ( \14915 , \796 );
and \U$14573 ( \14916 , RI98719b0_131, \3861 );
not \U$14574 ( \14917 , RI98719b0_131);
and \U$14575 ( \14918 , \14917 , \3240 );
or \U$14576 ( \14919 , \14916 , \14918 );
not \U$14577 ( \14920 , \14919 );
or \U$14578 ( \14921 , \14915 , \14920 );
nand \U$14579 ( \14922 , \14557 , \793 );
nand \U$14580 ( \14923 , \14921 , \14922 );
not \U$14581 ( \14924 , \1083 );
not \U$14582 ( \14925 , \14566 );
or \U$14583 ( \14926 , \14924 , \14925 );
not \U$14584 ( \14927 , \1111 );
not \U$14585 ( \14928 , \4153 );
or \U$14586 ( \14929 , \14927 , \14928 );
buf \U$14587 ( \14930 , \3567 );
nand \U$14588 ( \14931 , \14930 , RI98718c0_129);
nand \U$14589 ( \14932 , \14929 , \14931 );
nand \U$14590 ( \14933 , \14932 , \6673 );
nand \U$14591 ( \14934 , \14926 , \14933 );
xor \U$14592 ( \14935 , \14923 , \14934 );
not \U$14593 ( \14936 , \5796 );
and \U$14594 ( \14937 , RI9872478_154, \2216 );
not \U$14595 ( \14938 , RI9872478_154);
and \U$14596 ( \14939 , \14938 , \847 );
or \U$14597 ( \14940 , \14937 , \14939 );
not \U$14598 ( \14941 , \14940 );
or \U$14599 ( \14942 , \14936 , \14941 );
nand \U$14600 ( \14943 , \14626 , \5034 );
nand \U$14601 ( \14944 , \14942 , \14943 );
xor \U$14602 ( \14945 , \14935 , \14944 );
not \U$14603 ( \14946 , \4085 );
and \U$14604 ( \14947 , RI98725e0_157, \4455 );
not \U$14605 ( \14948 , RI98725e0_157);
and \U$14606 ( \14949 , \14948 , \1604 );
or \U$14607 ( \14950 , \14947 , \14949 );
not \U$14608 ( \14951 , \14950 );
or \U$14609 ( \14952 , \14946 , \14951 );
nand \U$14610 ( \14953 , \14507 , \8790 );
nand \U$14611 ( \14954 , \14952 , \14953 );
not \U$14612 ( \14955 , \9196 );
not \U$14613 ( \14956 , \14339 );
or \U$14614 ( \14957 , \14955 , \14956 );
not \U$14615 ( \14958 , \9198 );
not \U$14616 ( \14959 , \2982 );
or \U$14617 ( \14960 , \14958 , \14959 );
or \U$14618 ( \14961 , \1393 , \9198 );
nand \U$14619 ( \14962 , \14960 , \14961 );
nand \U$14620 ( \14963 , \14962 , \9214 );
nand \U$14621 ( \14964 , \14957 , \14963 );
xor \U$14622 ( \14965 , \14954 , \14964 );
not \U$14623 ( \14966 , \7338 );
not \U$14624 ( \14967 , RI98729a0_165);
not \U$14625 ( \14968 , \1447 );
or \U$14626 ( \14969 , \14967 , \14968 );
or \U$14627 ( \14970 , \1447 , RI98729a0_165);
nand \U$14628 ( \14971 , \14969 , \14970 );
not \U$14629 ( \14972 , \14971 );
or \U$14630 ( \14973 , \14966 , \14972 );
nand \U$14631 ( \14974 , \14355 , \7325 );
nand \U$14632 ( \14975 , \14973 , \14974 );
xor \U$14633 ( \14976 , \14965 , \14975 );
xor \U$14634 ( \14977 , \14945 , \14976 );
not \U$14635 ( \14978 , \2074 );
not \U$14636 ( \14979 , \14526 );
or \U$14637 ( \14980 , \14978 , \14979 );
xnor \U$14638 ( \14981 , RI9871aa0_133, \2962 );
nand \U$14639 ( \14982 , \14981 , \2087 );
nand \U$14640 ( \14983 , \14980 , \14982 );
not \U$14641 ( \14984 , \9072 );
xnor \U$14642 ( \14985 , RI9872a18_166, \1098 );
not \U$14643 ( \14986 , \14985 );
or \U$14644 ( \14987 , \14984 , \14986 );
nand \U$14645 ( \14988 , \14518 , \9079 );
nand \U$14646 ( \14989 , \14987 , \14988 );
xor \U$14647 ( \14990 , \14983 , \14989 );
not \U$14648 ( \14991 , RI9872568_156);
not \U$14649 ( \14992 , \6443 );
or \U$14650 ( \14993 , \14991 , \14992 );
or \U$14651 ( \14994 , \6443 , RI9872568_156);
nand \U$14652 ( \14995 , \14993 , \14994 );
not \U$14653 ( \14996 , \14995 );
or \U$14654 ( \14997 , \14996 , \7677 );
not \U$14655 ( \14998 , \14577 );
or \U$14656 ( \14999 , \14998 , \7845 );
nand \U$14657 ( \15000 , \14997 , \14999 );
xor \U$14658 ( \15001 , \14990 , \15000 );
xor \U$14659 ( \15002 , \14977 , \15001 );
not \U$14660 ( \15003 , \15002 );
and \U$14661 ( \15004 , \14914 , \15003 );
not \U$14662 ( \15005 , \14914 );
and \U$14663 ( \15006 , \15005 , \15002 );
nor \U$14664 ( \15007 , \15004 , \15006 );
xor \U$14665 ( \15008 , \14862 , \15007 );
not \U$14666 ( \15009 , \14465 );
not \U$14667 ( \15010 , \14458 );
or \U$14668 ( \15011 , \15009 , \15010 );
not \U$14669 ( \15012 , \14447 );
nand \U$14670 ( \15013 , \15012 , \14454 );
nand \U$14671 ( \15014 , \15011 , \15013 );
not \U$14672 ( \15015 , \14366 );
not \U$14673 ( \15016 , \14298 );
or \U$14674 ( \15017 , \15015 , \15016 );
not \U$14675 ( \15018 , \14323 );
nand \U$14676 ( \15019 , \15018 , \14362 );
nand \U$14677 ( \15020 , \15017 , \15019 );
not \U$14678 ( \15021 , \1501 );
not \U$14679 ( \15022 , \14385 );
or \U$14680 ( \15023 , \15021 , \15022 );
and \U$14681 ( \15024 , \5776 , \1800 );
not \U$14682 ( \15025 , \5776 );
and \U$14683 ( \15026 , \15025 , RI9871c80_137);
nor \U$14684 ( \15027 , \15024 , \15026 );
nand \U$14685 ( \15028 , \15027 , \1518 );
nand \U$14686 ( \15029 , \15023 , \15028 );
not \U$14687 ( \15030 , \1323 );
and \U$14688 ( \15031 , \4960 , RI9871b18_134);
not \U$14689 ( \15032 , \4960 );
and \U$14690 ( \15033 , \15032 , \2479 );
nor \U$14691 ( \15034 , \15031 , \15033 );
not \U$14692 ( \15035 , \15034 );
or \U$14693 ( \15036 , \15030 , \15035 );
not \U$14694 ( \15037 , \14303 );
nand \U$14695 ( \15038 , \15037 , \1292 );
nand \U$14696 ( \15039 , \15036 , \15038 );
xor \U$14697 ( \15040 , \15029 , \15039 );
not \U$14698 ( \15041 , \4925 );
and \U$14699 ( \15042 , \1658 , \4902 );
not \U$14700 ( \15043 , \1658 );
and \U$14701 ( \15044 , \15043 , RI9872388_152);
nor \U$14702 ( \15045 , \15042 , \15044 );
not \U$14703 ( \15046 , \15045 );
or \U$14704 ( \15047 , \15041 , \15046 );
nand \U$14705 ( \15048 , \14497 , \6553 );
nand \U$14706 ( \15049 , \15047 , \15048 );
xor \U$14707 ( \15050 , \15040 , \15049 );
not \U$14708 ( \15051 , \3467 );
not \U$14709 ( \15052 , RI98726d0_159);
not \U$14710 ( \15053 , \9323 );
or \U$14711 ( \15054 , \15052 , \15053 );
or \U$14712 ( \15055 , \6330 , RI98726d0_159);
nand \U$14713 ( \15056 , \15054 , \15055 );
not \U$14714 ( \15057 , \15056 );
or \U$14715 ( \15058 , \15051 , \15057 );
nand \U$14716 ( \15059 , \14331 , \3466 );
nand \U$14717 ( \15060 , \15058 , \15059 );
not \U$14718 ( \15061 , \6611 );
not \U$14719 ( \15062 , RI98728b0_163);
not \U$14720 ( \15063 , \7064 );
or \U$14721 ( \15064 , \15062 , \15063 );
or \U$14722 ( \15065 , \7064 , RI98728b0_163);
nand \U$14723 ( \15066 , \15064 , \15065 );
not \U$14724 ( \15067 , \15066 );
or \U$14725 ( \15068 , \15061 , \15067 );
nand \U$14726 ( \15069 , \14545 , \6284 );
nand \U$14727 ( \15070 , \15068 , \15069 );
xor \U$14728 ( \15071 , \15060 , \15070 );
and \U$14729 ( \15072 , RI9872310_151, \5948 );
not \U$14730 ( \15073 , RI9872310_151);
and \U$14731 ( \15074 , \15073 , \3969 );
nor \U$14732 ( \15075 , \15072 , \15074 );
or \U$14733 ( \15076 , \15075 , \4261 );
not \U$14734 ( \15077 , \14534 );
or \U$14735 ( \15078 , \15077 , \3962 );
nand \U$14736 ( \15079 , \15076 , \15078 );
xor \U$14737 ( \15080 , \15071 , \15079 );
xor \U$14738 ( \15081 , \15050 , \15080 );
not \U$14739 ( \15082 , \14446 );
not \U$14740 ( \15083 , \14440 );
or \U$14741 ( \15084 , \15082 , \15083 );
nand \U$14742 ( \15085 , \14434 , \14436 );
nand \U$14743 ( \15086 , \15084 , \15085 );
xor \U$14744 ( \15087 , \15081 , \15086 );
xor \U$14745 ( \15088 , \15020 , \15087 );
xnor \U$14746 ( \15089 , \15014 , \15088 );
not \U$14747 ( \15090 , \15089 );
and \U$14748 ( \15091 , \15008 , \15090 );
not \U$14749 ( \15092 , \15008 );
and \U$14750 ( \15093 , \15092 , \15089 );
nor \U$14751 ( \15094 , \15091 , \15093 );
not \U$14752 ( \15095 , \15094 );
not \U$14753 ( \15096 , \14660 );
not \U$14754 ( \15097 , \14672 );
not \U$14755 ( \15098 , \14665 );
or \U$14756 ( \15099 , \15097 , \15098 );
or \U$14757 ( \15100 , \14665 , \14672 );
nand \U$14758 ( \15101 , \15099 , \15100 );
not \U$14759 ( \15102 , \15101 );
or \U$14760 ( \15103 , \15096 , \15102 );
nand \U$14761 ( \15104 , \14664 , \14672 );
nand \U$14762 ( \15105 , \15103 , \15104 );
not \U$14763 ( \15106 , \15105 );
or \U$14764 ( \15107 , \15095 , \15106 );
or \U$14765 ( \15108 , \15105 , \15094 );
nand \U$14766 ( \15109 , \15107 , \15108 );
not \U$14767 ( \15110 , \15109 );
not \U$14768 ( \15111 , \14480 );
not \U$14769 ( \15112 , \14375 );
or \U$14770 ( \15113 , \15111 , \15112 );
nand \U$14771 ( \15114 , \14374 , \14369 );
nand \U$14772 ( \15115 , \15113 , \15114 );
not \U$14773 ( \15116 , \15115 );
not \U$14774 ( \15117 , \15116 );
or \U$14775 ( \15118 , \15110 , \15117 );
not \U$14776 ( \15119 , \15109 );
nand \U$14777 ( \15120 , \15119 , \15115 );
nand \U$14778 ( \15121 , \15118 , \15120 );
xor \U$14779 ( \15122 , \14792 , \15121 );
not \U$14780 ( \15123 , \15122 );
or \U$14781 ( \15124 , \14696 , \15123 );
not \U$14782 ( \15125 , \15014 );
not \U$14783 ( \15126 , \15088 );
or \U$14784 ( \15127 , \15125 , \15126 );
nand \U$14785 ( \15128 , \15020 , \15087 );
nand \U$14786 ( \15129 , \15127 , \15128 );
not \U$14787 ( \15130 , \15129 );
not \U$14788 ( \15131 , \14706 );
not \U$14789 ( \15132 , \14762 );
not \U$14790 ( \15133 , \15132 );
or \U$14791 ( \15134 , \15131 , \15133 );
not \U$14792 ( \15135 , \14707 );
not \U$14793 ( \15136 , \14762 );
or \U$14794 ( \15137 , \15135 , \15136 );
nand \U$14795 ( \15138 , \15137 , \14769 );
nand \U$14796 ( \15139 , \15134 , \15138 );
and \U$14797 ( \15140 , \15130 , \15139 );
not \U$14798 ( \15141 , \15130 );
not \U$14799 ( \15142 , \15139 );
and \U$14800 ( \15143 , \15141 , \15142 );
nor \U$14801 ( \15144 , \15140 , \15143 );
not \U$14802 ( \15145 , \15144 );
nand \U$14803 ( \15146 , \14861 , \14818 );
and \U$14804 ( \15147 , \15146 , \14796 );
nor \U$14805 ( \15148 , \14861 , \14818 );
nor \U$14806 ( \15149 , \15147 , \15148 );
not \U$14807 ( \15150 , \1162 );
not \U$14808 ( \15151 , \14844 );
or \U$14809 ( \15152 , \15150 , \15151 );
xor \U$14810 ( \15153 , \8679 , \8621 );
nand \U$14811 ( \15154 , \15153 , \1220 );
nand \U$14812 ( \15155 , \15152 , \15154 );
not \U$14813 ( \15156 , \1018 );
not \U$14814 ( \15157 , \14877 );
or \U$14815 ( \15158 , \15156 , \15157 );
not \U$14816 ( \15159 , \8086 );
not \U$14817 ( \15160 , \8335 );
or \U$14818 ( \15161 , \15159 , \15160 );
or \U$14819 ( \15162 , \8335 , \3271 );
nand \U$14820 ( \15163 , \15161 , \15162 );
nand \U$14821 ( \15164 , \15163 , \1013 );
nand \U$14822 ( \15165 , \15158 , \15164 );
xor \U$14823 ( \15166 , \15155 , \15165 );
not \U$14824 ( \15167 , \1381 );
not \U$14825 ( \15168 , \14887 );
or \U$14826 ( \15169 , \15167 , \15168 );
not \U$14827 ( \15170 , \1367 );
not \U$14828 ( \15171 , \10584 );
or \U$14829 ( \15172 , \15170 , \15171 );
not \U$14830 ( \15173 , \7004 );
nand \U$14831 ( \15174 , \15173 , RI9871e60_141);
nand \U$14832 ( \15175 , \15172 , \15174 );
nand \U$14833 ( \15176 , \15175 , \1353 );
nand \U$14834 ( \15177 , \15169 , \15176 );
xor \U$14835 ( \15178 , \15166 , \15177 );
xor \U$14836 ( \15179 , \14881 , \14891 );
and \U$14837 ( \15180 , \15179 , \14902 );
and \U$14838 ( \15181 , \14881 , \14891 );
or \U$14839 ( \15182 , \15180 , \15181 );
xor \U$14840 ( \15183 , \15178 , \15182 );
xor \U$14841 ( \15184 , \14830 , \14835 );
not \U$14842 ( \15185 , \14846 );
and \U$14843 ( \15186 , \15184 , \15185 );
and \U$14844 ( \15187 , \14830 , \14835 );
or \U$14845 ( \15188 , \15186 , \15187 );
xor \U$14846 ( \15189 , \15183 , \15188 );
not \U$14847 ( \15190 , \14813 );
not \U$14848 ( \15191 , \14807 );
or \U$14849 ( \15192 , \15190 , \15191 );
nand \U$14850 ( \15193 , \14806 , \14800 );
nand \U$14851 ( \15194 , \15192 , \15193 );
xor \U$14852 ( \15195 , \15189 , \15194 );
xor \U$14853 ( \15196 , \14945 , \14976 );
and \U$14854 ( \15197 , \15196 , \15001 );
and \U$14855 ( \15198 , \14945 , \14976 );
or \U$14856 ( \15199 , \15197 , \15198 );
xor \U$14857 ( \15200 , \15195 , \15199 );
xor \U$14858 ( \15201 , \15149 , \15200 );
not \U$14859 ( \15202 , \14743 );
not \U$14860 ( \15203 , \14717 );
or \U$14861 ( \15204 , \15202 , \15203 );
nand \U$14862 ( \15205 , \14726 , \14737 );
nand \U$14863 ( \15206 , \15204 , \15205 );
not \U$14864 ( \15207 , \15206 );
or \U$14865 ( \15208 , \14872 , \14903 );
not \U$14866 ( \15209 , \15208 );
not \U$14867 ( \15210 , \14908 );
or \U$14868 ( \15211 , \15209 , \15210 );
nand \U$14869 ( \15212 , \14903 , \14872 );
nand \U$14870 ( \15213 , \15211 , \15212 );
xor \U$14871 ( \15214 , \15207 , \15213 );
not \U$14872 ( \15215 , \14829 );
not \U$14873 ( \15216 , \14857 );
or \U$14874 ( \15217 , \15215 , \15216 );
nand \U$14875 ( \15218 , \15217 , \14859 );
xor \U$14876 ( \15219 , \15214 , \15218 );
xor \U$14877 ( \15220 , \15201 , \15219 );
not \U$14878 ( \15221 , \15220 );
and \U$14879 ( \15222 , \15145 , \15221 );
and \U$14880 ( \15223 , \15220 , \15144 );
nor \U$14881 ( \15224 , \15222 , \15223 );
buf \U$14882 ( \15225 , \14711 );
buf \U$14883 ( \15226 , \14747 );
or \U$14884 ( \15227 , \15225 , \15226 );
nand \U$14885 ( \15228 , \15227 , \14757 );
nand \U$14886 ( \15229 , \15225 , \15226 );
nand \U$14887 ( \15230 , \15228 , \15229 );
not \U$14888 ( \15231 , \15230 );
not \U$14889 ( \15232 , \15231 );
nor \U$14890 ( \15233 , \8857 , \1716 );
not \U$14891 ( \15234 , \1292 );
not \U$14892 ( \15235 , \15034 );
or \U$14893 ( \15236 , \15234 , \15235 );
and \U$14894 ( \15237 , \4471 , \1283 );
not \U$14895 ( \15238 , \4471 );
and \U$14896 ( \15239 , \15238 , RI9871b18_134);
nor \U$14897 ( \15240 , \15237 , \15239 );
nand \U$14898 ( \15241 , \15240 , \1323 );
nand \U$14899 ( \15242 , \15236 , \15241 );
xor \U$14900 ( \15243 , \15233 , \15242 );
not \U$14901 ( \15244 , \5937 );
not \U$14902 ( \15245 , \4902 );
not \U$14903 ( \15246 , \944 );
or \U$14904 ( \15247 , \15245 , \15246 );
or \U$14905 ( \15248 , \944 , \4902 );
nand \U$14906 ( \15249 , \15247 , \15248 );
not \U$14907 ( \15250 , \15249 );
or \U$14908 ( \15251 , \15244 , \15250 );
nand \U$14909 ( \15252 , \15045 , \4920 );
nand \U$14910 ( \15253 , \15251 , \15252 );
xor \U$14911 ( \15254 , \15243 , \15253 );
not \U$14912 ( \15255 , \1430 );
and \U$14913 ( \15256 , \14562 , \3487 );
not \U$14914 ( \15257 , \14562 );
and \U$14915 ( \15258 , \15257 , RI9871c08_136);
nor \U$14916 ( \15259 , \15256 , \15258 );
not \U$14917 ( \15260 , \15259 );
or \U$14918 ( \15261 , \15255 , \15260 );
nand \U$14919 ( \15262 , \14722 , \1455 );
nand \U$14920 ( \15263 , \15261 , \15262 );
not \U$14921 ( \15264 , \15263 );
not \U$14922 ( \15265 , \15264 );
not \U$14923 ( \15266 , \1083 );
not \U$14924 ( \15267 , \14932 );
or \U$14925 ( \15268 , \15266 , \15267 );
and \U$14926 ( \15269 , RI98718c0_129, \3537 );
not \U$14927 ( \15270 , RI98718c0_129);
and \U$14928 ( \15271 , \15270 , \3542 );
nor \U$14929 ( \15272 , \15269 , \15271 );
nand \U$14930 ( \15273 , \15272 , \6672 );
nand \U$14931 ( \15274 , \15268 , \15273 );
not \U$14932 ( \15275 , \15274 );
not \U$14933 ( \15276 , \15275 );
not \U$14934 ( \15277 , \14736 );
or \U$14935 ( \15278 , \15276 , \15277 );
or \U$14936 ( \15279 , \15275 , \14736 );
nand \U$14937 ( \15280 , \15278 , \15279 );
not \U$14938 ( \15281 , \15280 );
or \U$14939 ( \15282 , \15265 , \15281 );
or \U$14940 ( \15283 , \15264 , \15280 );
nand \U$14941 ( \15284 , \15282 , \15283 );
xor \U$14942 ( \15285 , \15254 , \15284 );
not \U$14943 ( \15286 , \7326 );
not \U$14944 ( \15287 , \14971 );
or \U$14945 ( \15288 , \15286 , \15287 );
not \U$14946 ( \15289 , RI98729a0_165);
not \U$14947 ( \15290 , \6692 );
or \U$14948 ( \15291 , \15289 , \15290 );
or \U$14949 ( \15292 , \10145 , RI98729a0_165);
nand \U$14950 ( \15293 , \15291 , \15292 );
nand \U$14951 ( \15294 , \15293 , \7338 );
nand \U$14952 ( \15295 , \15288 , \15294 );
not \U$14953 ( \15296 , \6611 );
not \U$14954 ( \15297 , RI98728b0_163);
not \U$14955 ( \15298 , \1320 );
or \U$14956 ( \15299 , \15297 , \15298 );
or \U$14957 ( \15300 , \1320 , RI98728b0_163);
nand \U$14958 ( \15301 , \15299 , \15300 );
not \U$14959 ( \15302 , \15301 );
or \U$14960 ( \15303 , \15296 , \15302 );
nand \U$14961 ( \15304 , \15066 , \6284 );
nand \U$14962 ( \15305 , \15303 , \15304 );
and \U$14963 ( \15306 , \15295 , \15305 );
not \U$14964 ( \15307 , \15295 );
not \U$14965 ( \15308 , \15305 );
and \U$14966 ( \15309 , \15307 , \15308 );
nor \U$14967 ( \15310 , \15306 , \15309 );
not \U$14968 ( \15311 , \3600 );
not \U$14969 ( \15312 , \15056 );
or \U$14970 ( \15313 , \15311 , \15312 );
xor \U$14971 ( \15314 , RI98726d0_159, \10133 );
nand \U$14972 ( \15315 , \15314 , \3467 );
nand \U$14973 ( \15316 , \15313 , \15315 );
not \U$14974 ( \15317 , \15316 );
and \U$14975 ( \15318 , \15310 , \15317 );
not \U$14976 ( \15319 , \15310 );
and \U$14977 ( \15320 , \15319 , \15316 );
nor \U$14978 ( \15321 , \15318 , \15320 );
not \U$14979 ( \15322 , \15321 );
and \U$14980 ( \15323 , \15285 , \15322 );
not \U$14981 ( \15324 , \15285 );
and \U$14982 ( \15325 , \15324 , \15321 );
nor \U$14983 ( \15326 , \15323 , \15325 );
not \U$14984 ( \15327 , \793 );
not \U$14985 ( \15328 , \14919 );
or \U$14986 ( \15329 , \15327 , \15328 );
and \U$14987 ( \15330 , RI98719b0_131, \3691 );
not \U$14988 ( \15331 , RI98719b0_131);
and \U$14989 ( \15332 , \15331 , \10942 );
or \U$14990 ( \15333 , \15330 , \15332 );
nand \U$14991 ( \15334 , \15333 , \6145 );
nand \U$14992 ( \15335 , \15329 , \15334 );
not \U$14993 ( \15336 , \2074 );
not \U$14994 ( \15337 , \14981 );
or \U$14995 ( \15338 , \15336 , \15337 );
and \U$14996 ( \15339 , RI9871aa0_133, \2116 );
not \U$14997 ( \15340 , RI9871aa0_133);
and \U$14998 ( \15341 , \15340 , \3275 );
or \U$14999 ( \15342 , \15339 , \15341 );
nand \U$15000 ( \15343 , \15342 , \2087 );
nand \U$15001 ( \15344 , \15338 , \15343 );
xor \U$15002 ( \15345 , \15335 , \15344 );
not \U$15003 ( \15346 , \5796 );
and \U$15004 ( \15347 , RI9872478_154, \8006 );
not \U$15005 ( \15348 , RI9872478_154);
and \U$15006 ( \15349 , \15348 , \7691 );
or \U$15007 ( \15350 , \15347 , \15349 );
not \U$15008 ( \15351 , \15350 );
or \U$15009 ( \15352 , \15346 , \15351 );
nand \U$15010 ( \15353 , \14940 , \5034 );
nand \U$15011 ( \15354 , \15352 , \15353 );
xor \U$15012 ( \15355 , \15345 , \15354 );
and \U$15013 ( \15356 , \1800 , \5739 );
not \U$15014 ( \15357 , \1800 );
and \U$15015 ( \15358 , \15357 , \10873 );
nor \U$15016 ( \15359 , \15356 , \15358 );
or \U$15017 ( \15360 , \15359 , \1746 );
not \U$15018 ( \15361 , \15027 );
or \U$15019 ( \15362 , \15361 , \1591 );
nand \U$15020 ( \15363 , \15360 , \15362 );
not \U$15021 ( \15364 , \10679 );
not \U$15022 ( \15365 , \14962 );
or \U$15023 ( \15366 , \15364 , \15365 );
and \U$15024 ( \15367 , RI9872b80_169, \1690 );
not \U$15025 ( \15368 , RI9872b80_169);
and \U$15026 ( \15369 , \15368 , \779 );
nor \U$15027 ( \15370 , \15367 , \15369 );
nand \U$15028 ( \15371 , \15370 , \9214 );
nand \U$15029 ( \15372 , \15366 , \15371 );
xor \U$15030 ( \15373 , \15363 , \15372 );
not \U$15031 ( \15374 , \4101 );
not \U$15032 ( \15375 , \14950 );
or \U$15033 ( \15376 , \15374 , \15375 );
not \U$15034 ( \15377 , RI98725e0_157);
not \U$15035 ( \15378 , \1340 );
or \U$15036 ( \15379 , \15377 , \15378 );
or \U$15037 ( \15380 , \1344 , RI98725e0_157);
nand \U$15038 ( \15381 , \15379 , \15380 );
nand \U$15039 ( \15382 , \15381 , \5847 );
nand \U$15040 ( \15383 , \15376 , \15382 );
xor \U$15041 ( \15384 , \15373 , \15383 );
xor \U$15042 ( \15385 , \15355 , \15384 );
not \U$15043 ( \15386 , \9079 );
not \U$15044 ( \15387 , \14985 );
or \U$15045 ( \15388 , \15386 , \15387 );
not \U$15046 ( \15389 , RI9872a18_166);
and \U$15047 ( \15390 , \1725 , \15389 );
not \U$15048 ( \15391 , \1725 );
and \U$15049 ( \15392 , \15391 , RI9872a18_166);
nor \U$15050 ( \15393 , \15390 , \15392 );
nand \U$15051 ( \15394 , \15393 , \9072 );
nand \U$15052 ( \15395 , \15388 , \15394 );
not \U$15053 ( \15396 , \6653 );
not \U$15054 ( \15397 , \15075 );
not \U$15055 ( \15398 , \15397 );
or \U$15056 ( \15399 , \15396 , \15398 );
and \U$15057 ( \15400 , \7605 , RI9872310_151);
not \U$15058 ( \15401 , \7605 );
and \U$15059 ( \15402 , \15401 , \3154 );
nor \U$15060 ( \15403 , \15400 , \15402 );
nand \U$15061 ( \15404 , \15403 , \3170 );
nand \U$15062 ( \15405 , \15399 , \15404 );
xor \U$15063 ( \15406 , \15395 , \15405 );
not \U$15064 ( \15407 , \5642 );
not \U$15065 ( \15408 , \14995 );
or \U$15066 ( \15409 , \15407 , \15408 );
not \U$15067 ( \15410 , RI9872568_156);
not \U$15068 ( \15411 , \5480 );
or \U$15069 ( \15412 , \15410 , \15411 );
or \U$15070 ( \15413 , \918 , RI9872568_156);
nand \U$15071 ( \15414 , \15412 , \15413 );
nand \U$15072 ( \15415 , \15414 , \7188 );
nand \U$15073 ( \15416 , \15409 , \15415 );
xor \U$15074 ( \15417 , \15406 , \15416 );
not \U$15075 ( \15418 , \15417 );
xnor \U$15076 ( \15419 , \15385 , \15418 );
xor \U$15077 ( \15420 , \15326 , \15419 );
not \U$15078 ( \15421 , \15420 );
or \U$15079 ( \15422 , \15232 , \15421 );
or \U$15080 ( \15423 , \15420 , \15231 );
nand \U$15081 ( \15424 , \15422 , \15423 );
not \U$15082 ( \15425 , RI9872d60_173);
not \U$15083 ( \15426 , RI9872ce8_172);
or \U$15084 ( \15427 , \15425 , \15426 );
nand \U$15085 ( \15428 , \15427 , RI9872bf8_170);
not \U$15086 ( \15429 , \6635 );
not \U$15087 ( \15430 , \14898 );
or \U$15088 ( \15431 , \15429 , \15430 );
not \U$15089 ( \15432 , \1347 );
not \U$15090 ( \15433 , \12802 );
or \U$15091 ( \15434 , \15432 , \15433 );
nand \U$15092 ( \15435 , \8054 , RI9871d70_139);
nand \U$15093 ( \15436 , \15434 , \15435 );
nand \U$15094 ( \15437 , \15436 , \832 );
nand \U$15095 ( \15438 , \15431 , \15437 );
xor \U$15096 ( \15439 , \15428 , \15438 );
not \U$15097 ( \15440 , \876 );
not \U$15098 ( \15441 , \14732 );
or \U$15099 ( \15442 , \15440 , \15441 );
and \U$15100 ( \15443 , \10795 , RI9872130_147);
and \U$15101 ( \15444 , \6060 , \919 );
nor \U$15102 ( \15445 , \15443 , \15444 );
or \U$15103 ( \15446 , \15445 , \1470 );
nand \U$15104 ( \15447 , \15442 , \15446 );
xor \U$15105 ( \15448 , \15439 , \15447 );
xor \U$15106 ( \15449 , \14923 , \14934 );
and \U$15107 ( \15450 , \15449 , \14944 );
and \U$15108 ( \15451 , \14923 , \14934 );
or \U$15109 ( \15452 , \15450 , \15451 );
xor \U$15110 ( \15453 , \15448 , \15452 );
not \U$15111 ( \15454 , \15039 );
xor \U$15112 ( \15455 , \15049 , \15029 );
not \U$15113 ( \15456 , \15455 );
or \U$15114 ( \15457 , \15454 , \15456 );
nand \U$15115 ( \15458 , \15049 , \15029 );
nand \U$15116 ( \15459 , \15457 , \15458 );
xor \U$15117 ( \15460 , \15453 , \15459 );
xor \U$15118 ( \15461 , \14954 , \14964 );
and \U$15119 ( \15462 , \15461 , \14975 );
and \U$15120 ( \15463 , \14954 , \14964 );
or \U$15121 ( \15464 , \15462 , \15463 );
xor \U$15122 ( \15465 , \15060 , \15070 );
and \U$15123 ( \15466 , \15465 , \15079 );
and \U$15124 ( \15467 , \15060 , \15070 );
or \U$15125 ( \15468 , \15466 , \15467 );
xor \U$15126 ( \15469 , \15464 , \15468 );
xor \U$15127 ( \15470 , \14983 , \14989 );
and \U$15128 ( \15471 , \15470 , \15000 );
and \U$15129 ( \15472 , \14983 , \14989 );
or \U$15130 ( \15473 , \15471 , \15472 );
xor \U$15131 ( \15474 , \15469 , \15473 );
xor \U$15132 ( \15475 , \15460 , \15474 );
xor \U$15133 ( \15476 , \15050 , \15080 );
and \U$15134 ( \15477 , \15476 , \15086 );
and \U$15135 ( \15478 , \15050 , \15080 );
or \U$15136 ( \15479 , \15477 , \15478 );
xor \U$15137 ( \15480 , \15475 , \15479 );
not \U$15138 ( \15481 , \15480 );
not \U$15139 ( \15482 , \15002 );
nand \U$15140 ( \15483 , \14909 , \14867 );
not \U$15141 ( \15484 , \15483 );
or \U$15142 ( \15485 , \15482 , \15484 );
nand \U$15143 ( \15486 , \14910 , \14866 );
nand \U$15144 ( \15487 , \15485 , \15486 );
not \U$15145 ( \15488 , \15487 );
not \U$15146 ( \15489 , \15488 );
or \U$15147 ( \15490 , \15481 , \15489 );
or \U$15148 ( \15491 , \15488 , \15480 );
nand \U$15149 ( \15492 , \15490 , \15491 );
xor \U$15150 ( \15493 , \15424 , \15492 );
and \U$15151 ( \15494 , \14862 , \15007 );
or \U$15152 ( \15495 , \15089 , \15494 );
or \U$15153 ( \15496 , \15007 , \14862 );
nand \U$15154 ( \15497 , \15495 , \15496 );
nand \U$15155 ( \15498 , \15493 , \15497 );
not \U$15156 ( \15499 , \15497 );
not \U$15157 ( \15500 , \15493 );
nand \U$15158 ( \15501 , \15499 , \15500 );
nand \U$15159 ( \15502 , \15498 , \15501 );
xor \U$15160 ( \15503 , \15224 , \15502 );
xor \U$15161 ( \15504 , \14700 , \14770 );
and \U$15162 ( \15505 , \15504 , \14779 );
and \U$15163 ( \15506 , \14700 , \14770 );
or \U$15164 ( \15507 , \15505 , \15506 );
xnor \U$15165 ( \15508 , \15503 , \15507 );
or \U$15166 ( \15509 , \15105 , \15094 );
not \U$15167 ( \15510 , \15509 );
not \U$15168 ( \15511 , \15115 );
or \U$15169 ( \15512 , \15510 , \15511 );
nand \U$15170 ( \15513 , \15105 , \15094 );
nand \U$15171 ( \15514 , \15512 , \15513 );
and \U$15172 ( \15515 , \15508 , \15514 );
not \U$15173 ( \15516 , \15508 );
not \U$15174 ( \15517 , \15514 );
and \U$15175 ( \15518 , \15516 , \15517 );
nor \U$15176 ( \15519 , \15515 , \15518 );
not \U$15177 ( \15520 , \15121 );
not \U$15178 ( \15521 , \14792 );
or \U$15179 ( \15522 , \15520 , \15521 );
not \U$15180 ( \15523 , \14780 );
nand \U$15181 ( \15524 , \15523 , \14788 );
nand \U$15182 ( \15525 , \15522 , \15524 );
nand \U$15183 ( \15526 , \15519 , \15525 );
nand \U$15184 ( \15527 , \15124 , \15526 );
buf \U$15185 ( \15528 , \15527 );
xor \U$15186 ( \15529 , \15502 , \15507 );
buf \U$15187 ( \15530 , \15224 );
nand \U$15188 ( \15531 , \15529 , \15530 );
not \U$15189 ( \15532 , \15531 );
not \U$15190 ( \15533 , \15514 );
or \U$15191 ( \15534 , \15532 , \15533 );
or \U$15192 ( \15535 , \15529 , \15530 );
nand \U$15193 ( \15536 , \15534 , \15535 );
not \U$15194 ( \15537 , \15263 );
not \U$15195 ( \15538 , \15280 );
or \U$15196 ( \15539 , \15537 , \15538 );
nand \U$15197 ( \15540 , \14738 , \15274 );
nand \U$15198 ( \15541 , \15539 , \15540 );
not \U$15199 ( \15542 , \5796 );
not \U$15200 ( \15543 , RI9872478_154);
not \U$15201 ( \15544 , \893 );
or \U$15202 ( \15545 , \15543 , \15544 );
or \U$15203 ( \15546 , \893 , RI9872478_154);
nand \U$15204 ( \15547 , \15545 , \15546 );
not \U$15205 ( \15548 , \15547 );
or \U$15206 ( \15549 , \15542 , \15548 );
nand \U$15207 ( \15550 , \15350 , \5034 );
nand \U$15208 ( \15551 , \15549 , \15550 );
not \U$15209 ( \15552 , \793 );
not \U$15210 ( \15553 , \15333 );
or \U$15211 ( \15554 , \15552 , \15553 );
and \U$15212 ( \15555 , RI98719b0_131, \7164 );
not \U$15213 ( \15556 , RI98719b0_131);
and \U$15214 ( \15557 , \15556 , \2111 );
or \U$15215 ( \15558 , \15555 , \15557 );
nand \U$15216 ( \15559 , \15558 , \796 );
nand \U$15217 ( \15560 , \15554 , \15559 );
not \U$15218 ( \15561 , \15560 );
not \U$15219 ( \15562 , \1136 );
and \U$15220 ( \15563 , RI98718c0_129, \3860 );
not \U$15221 ( \15564 , RI98718c0_129);
and \U$15222 ( \15565 , \15564 , \3861 );
nor \U$15223 ( \15566 , \15563 , \15565 );
not \U$15224 ( \15567 , \15566 );
or \U$15225 ( \15568 , \15562 , \15567 );
nand \U$15226 ( \15569 , \15272 , \1083 );
nand \U$15227 ( \15570 , \15568 , \15569 );
not \U$15228 ( \15571 , \15570 );
xor \U$15229 ( \15572 , \15561 , \15571 );
xor \U$15230 ( \15573 , \15551 , \15572 );
xor \U$15231 ( \15574 , \15541 , \15573 );
not \U$15232 ( \15575 , \3170 );
and \U$15233 ( \15576 , \1040 , \3154 );
not \U$15234 ( \15577 , \1040 );
and \U$15235 ( \15578 , \15577 , RI9872310_151);
nor \U$15236 ( \15579 , \15576 , \15578 );
not \U$15237 ( \15580 , \15579 );
or \U$15238 ( \15581 , \15575 , \15580 );
nand \U$15239 ( \15582 , \15403 , \3163 );
nand \U$15240 ( \15583 , \15581 , \15582 );
not \U$15241 ( \15584 , \6284 );
not \U$15242 ( \15585 , \15301 );
or \U$15243 ( \15586 , \15584 , \15585 );
and \U$15244 ( \15587 , RI98728b0_163, \1447 );
not \U$15245 ( \15588 , RI98728b0_163);
and \U$15246 ( \15589 , \15588 , \10674 );
or \U$15247 ( \15590 , \15587 , \15589 );
nand \U$15248 ( \15591 , \15590 , \6611 );
nand \U$15249 ( \15592 , \15586 , \15591 );
xor \U$15250 ( \15593 , \15583 , \15592 );
not \U$15251 ( \15594 , \3467 );
and \U$15252 ( \15595 , RI98726d0_159, \1605 );
not \U$15253 ( \15596 , RI98726d0_159);
and \U$15254 ( \15597 , \15596 , \1606 );
nor \U$15255 ( \15598 , \15595 , \15597 );
not \U$15256 ( \15599 , \15598 );
or \U$15257 ( \15600 , \15594 , \15599 );
nand \U$15258 ( \15601 , \15314 , \3600 );
nand \U$15259 ( \15602 , \15600 , \15601 );
xor \U$15260 ( \15603 , \15593 , \15602 );
xor \U$15261 ( \15604 , \15574 , \15603 );
xor \U$15262 ( \15605 , \15335 , \15344 );
and \U$15263 ( \15606 , \15605 , \15354 );
and \U$15264 ( \15607 , \15335 , \15344 );
or \U$15265 ( \15608 , \15606 , \15607 );
and \U$15266 ( \15609 , \919 , \7028 );
not \U$15267 ( \15610 , \919 );
and \U$15268 ( \15611 , \15610 , \5776 );
nor \U$15269 ( \15612 , \15609 , \15611 );
or \U$15270 ( \15613 , \15612 , \1470 );
or \U$15271 ( \15614 , \15445 , \7927 );
nand \U$15272 ( \15615 , \15613 , \15614 );
not \U$15273 ( \15616 , \8029 );
not \U$15274 ( \15617 , \15393 );
or \U$15275 ( \15618 , \15616 , \15617 );
not \U$15276 ( \15619 , \8031 );
not \U$15277 ( \15620 , \2982 );
or \U$15278 ( \15621 , \15619 , \15620 );
or \U$15279 ( \15622 , \2982 , \8031 );
nand \U$15280 ( \15623 , \15621 , \15622 );
nand \U$15281 ( \15624 , \15623 , \9072 );
nand \U$15282 ( \15625 , \15618 , \15624 );
xor \U$15283 ( \15626 , \15615 , \15625 );
not \U$15284 ( \15627 , \1518 );
and \U$15285 ( \15628 , \10639 , RI9871c80_137);
not \U$15286 ( \15629 , \10639 );
and \U$15287 ( \15630 , \15629 , \1584 );
nor \U$15288 ( \15631 , \15628 , \15630 );
not \U$15289 ( \15632 , \15631 );
or \U$15290 ( \15633 , \15627 , \15632 );
or \U$15291 ( \15634 , \15359 , \1591 );
nand \U$15292 ( \15635 , \15633 , \15634 );
xor \U$15293 ( \15636 , \15626 , \15635 );
xor \U$15294 ( \15637 , \15608 , \15636 );
not \U$15295 ( \15638 , \7188 );
xnor \U$15296 ( \15639 , RI9872568_156, \1583 );
not \U$15297 ( \15640 , \15639 );
or \U$15298 ( \15641 , \15638 , \15640 );
nand \U$15299 ( \15642 , \15414 , \5642 );
nand \U$15300 ( \15643 , \15641 , \15642 );
not \U$15301 ( \15644 , \7338 );
not \U$15302 ( \15645 , RI98729a0_165);
not \U$15303 ( \15646 , \1097 );
or \U$15304 ( \15647 , \15645 , \15646 );
or \U$15305 ( \15648 , \1098 , RI98729a0_165);
nand \U$15306 ( \15649 , \15647 , \15648 );
not \U$15307 ( \15650 , \15649 );
or \U$15308 ( \15651 , \15644 , \15650 );
nand \U$15309 ( \15652 , \15293 , \7326 );
nand \U$15310 ( \15653 , \15651 , \15652 );
xor \U$15311 ( \15654 , \15643 , \15653 );
and \U$15312 ( \15655 , RI9871aa0_133, \5948 );
not \U$15313 ( \15656 , RI9871aa0_133);
and \U$15314 ( \15657 , \15656 , \1194 );
or \U$15315 ( \15658 , \15655 , \15657 );
not \U$15316 ( \15659 , \15658 );
or \U$15317 ( \15660 , \15659 , \2086 );
not \U$15318 ( \15661 , \15342 );
or \U$15319 ( \15662 , \15661 , \2073 );
nand \U$15320 ( \15663 , \15660 , \15662 );
xor \U$15321 ( \15664 , \15654 , \15663 );
xor \U$15322 ( \15665 , \15637 , \15664 );
xor \U$15323 ( \15666 , \15604 , \15665 );
not \U$15324 ( \15667 , \15213 );
not \U$15325 ( \15668 , \15207 );
not \U$15326 ( \15669 , \15218 );
or \U$15327 ( \15670 , \15668 , \15669 );
or \U$15328 ( \15671 , \15218 , \15207 );
nand \U$15329 ( \15672 , \15670 , \15671 );
not \U$15330 ( \15673 , \15672 );
or \U$15331 ( \15674 , \15667 , \15673 );
not \U$15332 ( \15675 , \15207 );
nand \U$15333 ( \15676 , \15675 , \15218 );
nand \U$15334 ( \15677 , \15674 , \15676 );
xor \U$15335 ( \15678 , \15666 , \15677 );
xor \U$15336 ( \15679 , \15448 , \15452 );
and \U$15337 ( \15680 , \15679 , \15459 );
and \U$15338 ( \15681 , \15448 , \15452 );
or \U$15339 ( \15682 , \15680 , \15681 );
not \U$15340 ( \15683 , \1323 );
not \U$15341 ( \15684 , \1283 );
not \U$15342 ( \15685 , \5614 );
not \U$15343 ( \15686 , \15685 );
or \U$15344 ( \15687 , \15684 , \15686 );
or \U$15345 ( \15688 , \5611 , \1283 );
nand \U$15346 ( \15689 , \15687 , \15688 );
not \U$15347 ( \15690 , \15689 );
or \U$15348 ( \15691 , \15683 , \15690 );
nand \U$15349 ( \15692 , \15240 , \1292 );
nand \U$15350 ( \15693 , \15691 , \15692 );
not \U$15351 ( \15694 , \1456 );
not \U$15352 ( \15695 , \15259 );
or \U$15353 ( \15696 , \15694 , \15695 );
and \U$15354 ( \15697 , \10699 , \3487 );
not \U$15355 ( \15698 , \10699 );
and \U$15356 ( \15699 , \15698 , RI9871c08_136);
nor \U$15357 ( \15700 , \15697 , \15699 );
nand \U$15358 ( \15701 , \15700 , \1430 );
nand \U$15359 ( \15702 , \15696 , \15701 );
xor \U$15360 ( \15703 , \15693 , \15702 );
not \U$15361 ( \15704 , \4925 );
xor \U$15362 ( \15705 , RI9872388_152, \847 );
not \U$15363 ( \15706 , \15705 );
or \U$15364 ( \15707 , \15704 , \15706 );
nand \U$15365 ( \15708 , \4920 , \15249 );
nand \U$15366 ( \15709 , \15707 , \15708 );
xor \U$15367 ( \15710 , \15703 , \15709 );
xor \U$15368 ( \15711 , \15155 , \15165 );
and \U$15369 ( \15712 , \15711 , \15177 );
and \U$15370 ( \15713 , \15155 , \15165 );
or \U$15371 ( \15714 , \15712 , \15713 );
not \U$15372 ( \15715 , \10679 );
not \U$15373 ( \15716 , \15370 );
or \U$15374 ( \15717 , \15715 , \15716 );
nand \U$15375 ( \15718 , \9214 , RI9872b80_169);
nand \U$15376 ( \15719 , \15717 , \15718 );
and \U$15377 ( \15720 , \15714 , \15719 );
not \U$15378 ( \15721 , \15714 );
not \U$15379 ( \15722 , \15719 );
and \U$15380 ( \15723 , \15721 , \15722 );
or \U$15381 ( \15724 , \15720 , \15723 );
not \U$15382 ( \15725 , \15724 );
xor \U$15383 ( \15726 , \15428 , \15438 );
and \U$15384 ( \15727 , \15726 , \15447 );
and \U$15385 ( \15728 , \15428 , \15438 );
nor \U$15386 ( \15729 , \15727 , \15728 );
not \U$15387 ( \15730 , \15729 );
or \U$15388 ( \15731 , \15725 , \15730 );
or \U$15389 ( \15732 , \15729 , \15724 );
nand \U$15390 ( \15733 , \15731 , \15732 );
xor \U$15391 ( \15734 , \15710 , \15733 );
xor \U$15392 ( \15735 , \15682 , \15734 );
xor \U$15393 ( \15736 , \15189 , \15194 );
and \U$15394 ( \15737 , \15736 , \15199 );
and \U$15395 ( \15738 , \15189 , \15194 );
or \U$15396 ( \15739 , \15737 , \15738 );
xor \U$15397 ( \15740 , \15735 , \15739 );
xor \U$15398 ( \15741 , \15178 , \15182 );
and \U$15399 ( \15742 , \15741 , \15188 );
and \U$15400 ( \15743 , \15178 , \15182 );
or \U$15401 ( \15744 , \15742 , \15743 );
xor \U$15402 ( \15745 , \15464 , \15468 );
and \U$15403 ( \15746 , \15745 , \15473 );
and \U$15404 ( \15747 , \15464 , \15468 );
or \U$15405 ( \15748 , \15746 , \15747 );
xor \U$15406 ( \15749 , \15744 , \15748 );
xor \U$15407 ( \15750 , \15363 , \15372 );
and \U$15408 ( \15751 , \15750 , \15383 );
and \U$15409 ( \15752 , \15363 , \15372 );
or \U$15410 ( \15753 , \15751 , \15752 );
not \U$15411 ( \15754 , \15317 );
not \U$15412 ( \15755 , \15308 );
or \U$15413 ( \15756 , \15754 , \15755 );
nand \U$15414 ( \15757 , \15756 , \15295 );
nand \U$15415 ( \15758 , \15305 , \15316 );
nand \U$15416 ( \15759 , \15757 , \15758 );
xor \U$15417 ( \15760 , \15753 , \15759 );
xor \U$15418 ( \15761 , \15395 , \15405 );
and \U$15419 ( \15762 , \15761 , \15416 );
and \U$15420 ( \15763 , \15395 , \15405 );
or \U$15421 ( \15764 , \15762 , \15763 );
xor \U$15422 ( \15765 , \15760 , \15764 );
and \U$15423 ( \15766 , \15749 , \15765 );
not \U$15424 ( \15767 , \15749 );
not \U$15425 ( \15768 , \15765 );
and \U$15426 ( \15769 , \15767 , \15768 );
nor \U$15427 ( \15770 , \15766 , \15769 );
xor \U$15428 ( \15771 , \15740 , \15770 );
xor \U$15429 ( \15772 , \15678 , \15771 );
not \U$15430 ( \15773 , \15149 );
not \U$15431 ( \15774 , \15773 );
not \U$15432 ( \15775 , \15200 );
nand \U$15433 ( \15776 , \15775 , \15219 );
not \U$15434 ( \15777 , \15776 );
or \U$15435 ( \15778 , \15774 , \15777 );
not \U$15436 ( \15779 , \15219 );
nand \U$15437 ( \15780 , \15779 , \15200 );
nand \U$15438 ( \15781 , \15778 , \15780 );
xor \U$15439 ( \15782 , \15772 , \15781 );
not \U$15440 ( \15783 , \15220 );
nand \U$15441 ( \15784 , \15130 , \15142 );
not \U$15442 ( \15785 , \15784 );
or \U$15443 ( \15786 , \15783 , \15785 );
nand \U$15444 ( \15787 , \15129 , \15139 );
nand \U$15445 ( \15788 , \15786 , \15787 );
not \U$15446 ( \15789 , \15480 );
nand \U$15447 ( \15790 , \15789 , \15488 );
not \U$15448 ( \15791 , \15790 );
not \U$15449 ( \15792 , \15424 );
or \U$15450 ( \15793 , \15791 , \15792 );
nand \U$15451 ( \15794 , \15487 , \15480 );
nand \U$15452 ( \15795 , \15793 , \15794 );
not \U$15453 ( \15796 , \15230 );
not \U$15454 ( \15797 , \15420 );
or \U$15455 ( \15798 , \15796 , \15797 );
nand \U$15456 ( \15799 , \15419 , \15326 );
nand \U$15457 ( \15800 , \15798 , \15799 );
not \U$15458 ( \15801 , \15800 );
xor \U$15459 ( \15802 , \15460 , \15474 );
and \U$15460 ( \15803 , \15802 , \15479 );
and \U$15461 ( \15804 , \15460 , \15474 );
or \U$15462 ( \15805 , \15803 , \15804 );
not \U$15463 ( \15806 , \15805 );
not \U$15464 ( \15807 , \15806 );
not \U$15465 ( \15808 , \15384 );
nand \U$15466 ( \15809 , \15808 , \15418 );
not \U$15467 ( \15810 , \15809 );
not \U$15468 ( \15811 , \15355 );
or \U$15469 ( \15812 , \15810 , \15811 );
nand \U$15470 ( \15813 , \15417 , \15384 );
nand \U$15471 ( \15814 , \15812 , \15813 );
not \U$15472 ( \15815 , \15814 );
not \U$15473 ( \15816 , \15284 );
nand \U$15474 ( \15817 , \15816 , \15321 );
not \U$15475 ( \15818 , \15817 );
not \U$15476 ( \15819 , \15254 );
or \U$15477 ( \15820 , \15818 , \15819 );
nand \U$15478 ( \15821 , \15322 , \15284 );
nand \U$15479 ( \15822 , \15820 , \15821 );
not \U$15480 ( \15823 , \15822 );
not \U$15481 ( \15824 , \1013 );
not \U$15482 ( \15825 , \8086 );
not \U$15483 ( \15826 , \7467 );
or \U$15484 ( \15827 , \15825 , \15826 );
or \U$15485 ( \15828 , \8925 , \1043 );
nand \U$15486 ( \15829 , \15827 , \15828 );
not \U$15487 ( \15830 , \15829 );
or \U$15488 ( \15831 , \15824 , \15830 );
nand \U$15489 ( \15832 , \15163 , \1018 );
nand \U$15490 ( \15833 , \15831 , \15832 );
not \U$15491 ( \15834 , \15833 );
nand \U$15492 ( \15835 , \8597 , \1165 );
not \U$15493 ( \15836 , \15835 );
and \U$15494 ( \15837 , \15834 , \15836 );
and \U$15495 ( \15838 , \15833 , \15835 );
nor \U$15496 ( \15839 , \15837 , \15838 );
not \U$15497 ( \15840 , \15839 );
not \U$15498 ( \15841 , \4101 );
not \U$15499 ( \15842 , \15381 );
or \U$15500 ( \15843 , \15841 , \15842 );
and \U$15501 ( \15844 , RI98725e0_157, \5721 );
not \U$15502 ( \15845 , RI98725e0_157);
and \U$15503 ( \15846 , \15845 , \7019 );
nor \U$15504 ( \15847 , \15844 , \15846 );
nand \U$15505 ( \15848 , \15847 , \4085 );
nand \U$15506 ( \15849 , \15843 , \15848 );
not \U$15507 ( \15850 , \15849 );
and \U$15508 ( \15851 , \15840 , \15850 );
and \U$15509 ( \15852 , \15839 , \15849 );
nor \U$15510 ( \15853 , \15851 , \15852 );
not \U$15511 ( \15854 , \15853 );
not \U$15512 ( \15855 , \1220 );
and \U$15513 ( \15856 , \9599 , \1716 );
not \U$15514 ( \15857 , \9599 );
and \U$15515 ( \15858 , \15857 , \8679 );
nor \U$15516 ( \15859 , \15856 , \15858 );
not \U$15517 ( \15860 , \15859 );
or \U$15518 ( \15861 , \15855 , \15860 );
nand \U$15519 ( \15862 , \15153 , \1162 );
nand \U$15520 ( \15863 , \15861 , \15862 );
not \U$15521 ( \15864 , \832 );
and \U$15522 ( \15865 , \6304 , RI9871d70_139);
not \U$15523 ( \15866 , \6304 );
and \U$15524 ( \15867 , \15866 , \12108 );
nor \U$15525 ( \15868 , \15865 , \15867 );
not \U$15526 ( \15869 , \15868 );
or \U$15527 ( \15870 , \15864 , \15869 );
nand \U$15528 ( \15871 , \15436 , \5350 );
nand \U$15529 ( \15872 , \15870 , \15871 );
xor \U$15530 ( \15873 , \15863 , \15872 );
not \U$15531 ( \15874 , \1353 );
not \U$15532 ( \15875 , \7905 );
and \U$15533 ( \15876 , RI9871e60_141, \15875 );
not \U$15534 ( \15877 , RI9871e60_141);
and \U$15535 ( \15878 , \15877 , \6530 );
or \U$15536 ( \15879 , \15876 , \15878 );
not \U$15537 ( \15880 , \15879 );
or \U$15538 ( \15881 , \15874 , \15880 );
nand \U$15539 ( \15882 , \15175 , \1381 );
nand \U$15540 ( \15883 , \15881 , \15882 );
not \U$15541 ( \15884 , \15883 );
xnor \U$15542 ( \15885 , \15873 , \15884 );
not \U$15543 ( \15886 , \15885 );
or \U$15544 ( \15887 , \15854 , \15886 );
or \U$15545 ( \15888 , \15853 , \15885 );
nand \U$15546 ( \15889 , \15887 , \15888 );
xor \U$15547 ( \15890 , \15233 , \15242 );
and \U$15548 ( \15891 , \15890 , \15253 );
and \U$15549 ( \15892 , \15233 , \15242 );
or \U$15550 ( \15893 , \15891 , \15892 );
xnor \U$15551 ( \15894 , \15889 , \15893 );
not \U$15552 ( \15895 , \15894 );
and \U$15553 ( \15896 , \15823 , \15895 );
and \U$15554 ( \15897 , \15822 , \15894 );
nor \U$15555 ( \15898 , \15896 , \15897 );
not \U$15556 ( \15899 , \15898 );
or \U$15557 ( \15900 , \15815 , \15899 );
or \U$15558 ( \15901 , \15814 , \15898 );
nand \U$15559 ( \15902 , \15900 , \15901 );
not \U$15560 ( \15903 , \15902 );
or \U$15561 ( \15904 , \15807 , \15903 );
or \U$15562 ( \15905 , \15902 , \15806 );
nand \U$15563 ( \15906 , \15904 , \15905 );
not \U$15564 ( \15907 , \15906 );
and \U$15565 ( \15908 , \15801 , \15907 );
and \U$15566 ( \15909 , \15800 , \15906 );
nor \U$15567 ( \15910 , \15908 , \15909 );
xor \U$15568 ( \15911 , \15795 , \15910 );
xor \U$15569 ( \15912 , \15788 , \15911 );
xor \U$15570 ( \15913 , \15782 , \15912 );
not \U$15571 ( \15914 , \15501 );
not \U$15572 ( \15915 , \15507 );
or \U$15573 ( \15916 , \15914 , \15915 );
nand \U$15574 ( \15917 , \15916 , \15498 );
xor \U$15575 ( \15918 , \15913 , \15917 );
nor \U$15576 ( \15919 , \15536 , \15918 );
not \U$15577 ( \15920 , \14692 );
and \U$15578 ( \15921 , \14684 , \15920 );
not \U$15579 ( \15922 , \14684 );
and \U$15580 ( \15923 , \15922 , \14692 );
nor \U$15581 ( \15924 , \15921 , \15923 );
not \U$15582 ( \15925 , \15924 );
not \U$15583 ( \15926 , \12358 );
not \U$15584 ( \15927 , \12069 );
or \U$15585 ( \15928 , \15926 , \15927 );
not \U$15586 ( \15929 , \12070 );
not \U$15587 ( \15930 , \12357 );
or \U$15588 ( \15931 , \15929 , \15930 );
nand \U$15589 ( \15932 , \15931 , \11894 );
nand \U$15590 ( \15933 , \15928 , \15932 );
nor \U$15591 ( \15934 , \15925 , \15933 );
nor \U$15592 ( \15935 , \15528 , \15919 , \15934 );
buf \U$15593 ( \15936 , \15935 );
nand \U$15594 ( \15937 , \14280 , \15936 );
not \U$15595 ( \15938 , \924 );
not \U$15596 ( \15939 , \7795 );
or \U$15597 ( \15940 , \15938 , \15939 );
and \U$15598 ( \15941 , RI9872130_147, \10873 );
not \U$15599 ( \15942 , RI9872130_147);
and \U$15600 ( \15943 , \15942 , \5325 );
nor \U$15601 ( \15944 , \15941 , \15943 );
not \U$15602 ( \15945 , \15944 );
nand \U$15603 ( \15946 , \15945 , \6431 );
nand \U$15604 ( \15947 , \15940 , \15946 );
not \U$15605 ( \15948 , \1162 );
and \U$15606 ( \15949 , \8334 , \1199 );
not \U$15607 ( \15950 , \8334 );
and \U$15608 ( \15951 , \15950 , \4708 );
nor \U$15609 ( \15952 , \15949 , \15951 );
not \U$15610 ( \15953 , \15952 );
or \U$15611 ( \15954 , \15948 , \15953 );
nand \U$15612 ( \15955 , \8339 , \1220 );
nand \U$15613 ( \15956 , \15954 , \15955 );
xor \U$15614 ( \15957 , \15947 , \15956 );
or \U$15615 ( \15958 , \8351 , \3591 );
xnor \U$15616 ( \15959 , RI98726d0_159, \1949 );
not \U$15617 ( \15960 , \3466 );
or \U$15618 ( \15961 , \15959 , \15960 );
nand \U$15619 ( \15962 , \15958 , \15961 );
xor \U$15620 ( \15963 , \15957 , \15962 );
xor \U$15621 ( \15964 , \8215 , \8190 );
xor \U$15622 ( \15965 , \15963 , \15964 );
xor \U$15623 ( \15966 , \7981 , \7991 );
xor \U$15624 ( \15967 , \15966 , \8012 );
xor \U$15625 ( \15968 , \15965 , \15967 );
not \U$15626 ( \15969 , \15853 );
not \U$15627 ( \15970 , \15885 );
not \U$15628 ( \15971 , \15970 );
or \U$15629 ( \15972 , \15969 , \15971 );
nand \U$15630 ( \15973 , \15972 , \15893 );
not \U$15631 ( \15974 , \15853 );
nand \U$15632 ( \15975 , \15974 , \15885 );
nand \U$15633 ( \15976 , \15973 , \15975 );
xor \U$15634 ( \15977 , \15541 , \15573 );
and \U$15635 ( \15978 , \15977 , \15603 );
and \U$15636 ( \15979 , \15541 , \15573 );
or \U$15637 ( \15980 , \15978 , \15979 );
xor \U$15638 ( \15981 , \15976 , \15980 );
xor \U$15639 ( \15982 , \15753 , \15759 );
and \U$15640 ( \15983 , \15982 , \15764 );
and \U$15641 ( \15984 , \15753 , \15759 );
or \U$15642 ( \15985 , \15983 , \15984 );
and \U$15643 ( \15986 , \15981 , \15985 );
and \U$15644 ( \15987 , \15976 , \15980 );
or \U$15645 ( \15988 , \15986 , \15987 );
xor \U$15646 ( \15989 , \15968 , \15988 );
xor \U$15647 ( \15990 , \15615 , \15625 );
and \U$15648 ( \15991 , \15990 , \15635 );
and \U$15649 ( \15992 , \15615 , \15625 );
nor \U$15650 ( \15993 , \15991 , \15992 );
not \U$15651 ( \15994 , \15993 );
not \U$15652 ( \15995 , \15994 );
xor \U$15653 ( \15996 , \15643 , \15653 );
and \U$15654 ( \15997 , \15996 , \15663 );
and \U$15655 ( \15998 , \15643 , \15653 );
or \U$15656 ( \15999 , \15997 , \15998 );
not \U$15657 ( \16000 , \15999 );
and \U$15658 ( \16001 , \15593 , \15602 );
and \U$15659 ( \16002 , \15583 , \15592 );
nor \U$15660 ( \16003 , \16001 , \16002 );
not \U$15661 ( \16004 , \16003 );
or \U$15662 ( \16005 , \16000 , \16004 );
or \U$15663 ( \16006 , \16003 , \15999 );
nand \U$15664 ( \16007 , \16005 , \16006 );
not \U$15665 ( \16008 , \16007 );
or \U$15666 ( \16009 , \15995 , \16008 );
not \U$15667 ( \16010 , \16003 );
nand \U$15668 ( \16011 , \16010 , \15999 );
nand \U$15669 ( \16012 , \16009 , \16011 );
not \U$15670 ( \16013 , \16012 );
nand \U$15671 ( \16014 , \9188 , RI9872b80_169);
not \U$15672 ( \16015 , \16014 );
not \U$15673 ( \16016 , \859 );
not \U$15674 ( \16017 , \15868 );
or \U$15675 ( \16018 , \16016 , \16017 );
or \U$15676 ( \16019 , \8116 , \932 );
nand \U$15677 ( \16020 , \16018 , \16019 );
not \U$15678 ( \16021 , \16020 );
or \U$15679 ( \16022 , \16015 , \16021 );
or \U$15680 ( \16023 , \16020 , \16014 );
not \U$15681 ( \16024 , \1381 );
not \U$15682 ( \16025 , \15879 );
or \U$15683 ( \16026 , \16024 , \16025 );
nand \U$15684 ( \16027 , \8058 , \1353 );
nand \U$15685 ( \16028 , \16026 , \16027 );
nand \U$15686 ( \16029 , \16023 , \16028 );
nand \U$15687 ( \16030 , \16022 , \16029 );
not \U$15688 ( \16031 , \16030 );
and \U$15689 ( \16032 , \8679 , \8621 );
not \U$15690 ( \16033 , \1162 );
not \U$15691 ( \16034 , \15859 );
or \U$15692 ( \16035 , \16033 , \16034 );
nand \U$15693 ( \16036 , \15952 , \1220 );
nand \U$15694 ( \16037 , \16035 , \16036 );
xor \U$15695 ( \16038 , \16032 , \16037 );
not \U$15696 ( \16039 , \15829 );
or \U$15697 ( \16040 , \16039 , \1612 );
not \U$15698 ( \16041 , \8088 );
or \U$15699 ( \16042 , \16041 , \1014 );
nand \U$15700 ( \16043 , \16040 , \16042 );
and \U$15701 ( \16044 , \16038 , \16043 );
and \U$15702 ( \16045 , \16032 , \16037 );
nor \U$15703 ( \16046 , \16044 , \16045 );
not \U$15704 ( \16047 , \16046 );
or \U$15705 ( \16048 , \16031 , \16047 );
or \U$15706 ( \16049 , \16030 , \16046 );
nand \U$15707 ( \16050 , \16048 , \16049 );
not \U$15708 ( \16051 , \8060 );
and \U$15709 ( \16052 , \8094 , \16051 );
not \U$15710 ( \16053 , \8094 );
and \U$15711 ( \16054 , \16053 , \8060 );
nor \U$15712 ( \16055 , \16052 , \16054 );
and \U$15713 ( \16056 , \16050 , \16055 );
not \U$15714 ( \16057 , \16050 );
and \U$15715 ( \16058 , \8094 , \16051 );
not \U$15716 ( \16059 , \8094 );
and \U$15717 ( \16060 , \16059 , \8060 );
or \U$15718 ( \16061 , \16058 , \16060 );
and \U$15719 ( \16062 , \16057 , \16061 );
or \U$15720 ( \16063 , \16056 , \16062 );
not \U$15721 ( \16064 , \16063 );
xor \U$15722 ( \16065 , \16014 , \16020 );
xnor \U$15723 ( \16066 , \16065 , \16028 );
not \U$15724 ( \16067 , \15839 );
and \U$15725 ( \16068 , \16067 , \15849 );
not \U$15726 ( \16069 , \15833 );
nor \U$15727 ( \16070 , \16069 , \15835 );
nor \U$15728 ( \16071 , \16068 , \16070 );
nand \U$15729 ( \16072 , \16066 , \16071 );
xor \U$15730 ( \16073 , \16032 , \16037 );
xor \U$15731 ( \16074 , \16073 , \16043 );
nand \U$15732 ( \16075 , \16072 , \16074 );
or \U$15733 ( \16076 , \16066 , \16071 );
and \U$15734 ( \16077 , \16075 , \16076 );
not \U$15735 ( \16078 , \16077 );
and \U$15736 ( \16079 , \16064 , \16078 );
and \U$15737 ( \16080 , \16063 , \16077 );
nor \U$15738 ( \16081 , \16079 , \16080 );
not \U$15739 ( \16082 , \16081 );
and \U$15740 ( \16083 , \16013 , \16082 );
and \U$15741 ( \16084 , \16012 , \16081 );
nor \U$15742 ( \16085 , \16083 , \16084 );
and \U$15743 ( \16086 , \15989 , \16085 );
not \U$15744 ( \16087 , \15989 );
not \U$15745 ( \16088 , \16085 );
and \U$15746 ( \16089 , \16087 , \16088 );
nor \U$15747 ( \16090 , \16086 , \16089 );
xor \U$15748 ( \16091 , \15976 , \15980 );
xor \U$15749 ( \16092 , \16091 , \15985 );
not \U$15750 ( \16093 , \16092 );
or \U$15751 ( \16094 , \15872 , \15863 );
and \U$15752 ( \16095 , \16094 , \15883 );
and \U$15753 ( \16096 , \15872 , \15863 );
nor \U$15754 ( \16097 , \16095 , \16096 );
not \U$15755 ( \16098 , \16097 );
not \U$15756 ( \16099 , \15722 );
not \U$15757 ( \16100 , \1323 );
and \U$15758 ( \16101 , RI9871b18_134, \5596 );
not \U$15759 ( \16102 , RI9871b18_134);
and \U$15760 ( \16103 , \16102 , \5599 );
or \U$15761 ( \16104 , \16101 , \16103 );
not \U$15762 ( \16105 , \16104 );
or \U$15763 ( \16106 , \16100 , \16105 );
nand \U$15764 ( \16107 , \1292 , \15689 );
nand \U$15765 ( \16108 , \16106 , \16107 );
not \U$15766 ( \16109 , \16108 );
or \U$15767 ( \16110 , \16099 , \16109 );
or \U$15768 ( \16111 , \16108 , \15722 );
nand \U$15769 ( \16112 , \16110 , \16111 );
not \U$15770 ( \16113 , \16112 );
and \U$15771 ( \16114 , \16098 , \16113 );
and \U$15772 ( \16115 , \16097 , \16112 );
nor \U$15773 ( \16116 , \16114 , \16115 );
not \U$15774 ( \16117 , \16116 );
not \U$15775 ( \16118 , \1455 );
not \U$15776 ( \16119 , \15700 );
or \U$15777 ( \16120 , \16118 , \16119 );
nand \U$15778 ( \16121 , \8147 , \1430 );
nand \U$15779 ( \16122 , \16120 , \16121 );
and \U$15780 ( \16123 , \8158 , \6673 );
and \U$15781 ( \16124 , \15566 , \1083 );
nor \U$15782 ( \16125 , \16123 , \16124 );
xor \U$15783 ( \16126 , \16122 , \16125 );
not \U$15784 ( \16127 , \5937 );
not \U$15785 ( \16128 , \8008 );
or \U$15786 ( \16129 , \16127 , \16128 );
nand \U$15787 ( \16130 , \15705 , \5942 );
nand \U$15788 ( \16131 , \16129 , \16130 );
xnor \U$15789 ( \16132 , \16126 , \16131 );
not \U$15790 ( \16133 , \16132 );
or \U$15791 ( \16134 , \16117 , \16133 );
or \U$15792 ( \16135 , \16132 , \16116 );
nand \U$15793 ( \16136 , \16134 , \16135 );
not \U$15794 ( \16137 , \15724 );
not \U$15795 ( \16138 , \15729 );
not \U$15796 ( \16139 , \16138 );
or \U$15797 ( \16140 , \16137 , \16139 );
nand \U$15798 ( \16141 , \15714 , \15722 );
nand \U$15799 ( \16142 , \16140 , \16141 );
not \U$15800 ( \16143 , \16142 );
and \U$15801 ( \16144 , \16136 , \16143 );
not \U$15802 ( \16145 , \16136 );
and \U$15803 ( \16146 , \16145 , \16142 );
nor \U$15804 ( \16147 , \16144 , \16146 );
nand \U$15805 ( \16148 , \16093 , \16147 );
not \U$15806 ( \16149 , \15765 );
not \U$15807 ( \16150 , \15749 );
or \U$15808 ( \16151 , \16149 , \16150 );
nand \U$15809 ( \16152 , \15748 , \15744 );
nand \U$15810 ( \16153 , \16151 , \16152 );
buf \U$15811 ( \16154 , \16153 );
and \U$15812 ( \16155 , \16148 , \16154 );
nor \U$15813 ( \16156 , \16093 , \16147 );
nor \U$15814 ( \16157 , \16155 , \16156 );
xor \U$15815 ( \16158 , \16090 , \16157 );
not \U$15816 ( \16159 , \3600 );
not \U$15817 ( \16160 , \15598 );
or \U$15818 ( \16161 , \16159 , \16160 );
not \U$15819 ( \16162 , \15959 );
nand \U$15820 ( \16163 , \16162 , \3467 );
nand \U$15821 ( \16164 , \16161 , \16163 );
not \U$15822 ( \16165 , \8029 );
not \U$15823 ( \16166 , \15623 );
or \U$15824 ( \16167 , \16165 , \16166 );
nand \U$15825 ( \16168 , \8036 , \8041 );
nand \U$15826 ( \16169 , \16167 , \16168 );
not \U$15827 ( \16170 , \6284 );
not \U$15828 ( \16171 , \15590 );
or \U$15829 ( \16172 , \16170 , \16171 );
nand \U$15830 ( \16173 , \7979 , \6611 );
nand \U$15831 ( \16174 , \16172 , \16173 );
xor \U$15832 ( \16175 , \16169 , \16174 );
xor \U$15833 ( \16176 , \16164 , \16175 );
not \U$15834 ( \16177 , \3164 );
not \U$15835 ( \16178 , \15579 );
or \U$15836 ( \16179 , \16177 , \16178 );
nand \U$15837 ( \16180 , \8122 , \3170 );
nand \U$15838 ( \16181 , \16179 , \16180 );
not \U$15839 ( \16182 , \2074 );
not \U$15840 ( \16183 , \15658 );
or \U$15841 ( \16184 , \16182 , \16183 );
nand \U$15842 ( \16185 , \8187 , \2087 );
nand \U$15843 ( \16186 , \16184 , \16185 );
xor \U$15844 ( \16187 , \16181 , \16186 );
not \U$15845 ( \16188 , \5642 );
not \U$15846 ( \16189 , \15639 );
or \U$15847 ( \16190 , \16188 , \16189 );
nand \U$15848 ( \16191 , \8206 , \7188 );
nand \U$15849 ( \16192 , \16190 , \16191 );
xnor \U$15850 ( \16193 , \16187 , \16192 );
not \U$15851 ( \16194 , \16193 );
xor \U$15852 ( \16195 , \16176 , \16194 );
not \U$15853 ( \16196 , \7988 );
not \U$15854 ( \16197 , \6145 );
not \U$15855 ( \16198 , \16197 );
and \U$15856 ( \16199 , \16196 , \16198 );
and \U$15857 ( \16200 , \15558 , \793 );
nor \U$15858 ( \16201 , \16199 , \16200 );
nand \U$15859 ( \16202 , \8131 , \7338 );
nand \U$15860 ( \16203 , \15649 , \7325 );
and \U$15861 ( \16204 , \16202 , \16203 );
xor \U$15862 ( \16205 , \16201 , \16204 );
not \U$15863 ( \16206 , \5034 );
not \U$15864 ( \16207 , \15547 );
or \U$15865 ( \16208 , \16206 , \16207 );
nand \U$15866 ( \16209 , \8199 , \5796 );
nand \U$15867 ( \16210 , \16208 , \16209 );
xnor \U$15868 ( \16211 , \16205 , \16210 );
xor \U$15869 ( \16212 , \16195 , \16211 );
not \U$15870 ( \16213 , \16212 );
nand \U$15871 ( \16214 , \16076 , \16072 );
and \U$15872 ( \16215 , \16214 , \16074 );
not \U$15873 ( \16216 , \16214 );
not \U$15874 ( \16217 , \16074 );
and \U$15875 ( \16218 , \16216 , \16217 );
nor \U$15876 ( \16219 , \16215 , \16218 );
not \U$15877 ( \16220 , \16219 );
and \U$15878 ( \16221 , \16213 , \16220 );
xor \U$15879 ( \16222 , \16176 , \16219 );
not \U$15880 ( \16223 , \16211 );
and \U$15881 ( \16224 , \16194 , \16223 );
not \U$15882 ( \16225 , \16194 );
and \U$15883 ( \16226 , \16225 , \16211 );
nor \U$15884 ( \16227 , \16224 , \16226 );
not \U$15885 ( \16228 , \16227 );
xor \U$15886 ( \16229 , \16222 , \16228 );
and \U$15887 ( \16230 , \15734 , \15682 );
and \U$15888 ( \16231 , \15710 , \15733 );
nor \U$15889 ( \16232 , \16230 , \16231 );
not \U$15890 ( \16233 , \16232 );
and \U$15891 ( \16234 , \16229 , \16233 );
nor \U$15892 ( \16235 , \16221 , \16234 );
and \U$15893 ( \16236 , \16158 , \16235 );
and \U$15894 ( \16237 , \16090 , \16157 );
or \U$15895 ( \16238 , \16236 , \16237 );
not \U$15896 ( \16239 , \15814 );
not \U$15897 ( \16240 , \15898 );
not \U$15898 ( \16241 , \16240 );
or \U$15899 ( \16242 , \16239 , \16241 );
not \U$15900 ( \16243 , \15894 );
nand \U$15901 ( \16244 , \16243 , \15822 );
nand \U$15902 ( \16245 , \16242 , \16244 );
xor \U$15903 ( \16246 , \15608 , \15636 );
and \U$15904 ( \16247 , \16246 , \15664 );
and \U$15905 ( \16248 , \15608 , \15636 );
or \U$15906 ( \16249 , \16247 , \16248 );
xor \U$15907 ( \16250 , \15693 , \15702 );
and \U$15908 ( \16251 , \16250 , \15709 );
and \U$15909 ( \16252 , \15693 , \15702 );
or \U$15910 ( \16253 , \16251 , \16252 );
not \U$15911 ( \16254 , \15551 );
not \U$15912 ( \16255 , \15570 );
and \U$15913 ( \16256 , \15561 , \16255 );
not \U$15914 ( \16257 , \16256 );
not \U$15915 ( \16258 , \16257 );
or \U$15916 ( \16259 , \16254 , \16258 );
nand \U$15917 ( \16260 , \15560 , \15570 );
nand \U$15918 ( \16261 , \16259 , \16260 );
xor \U$15919 ( \16262 , \16253 , \16261 );
not \U$15920 ( \16263 , \1501 );
not \U$15921 ( \16264 , \15631 );
or \U$15922 ( \16265 , \16263 , \16264 );
xnor \U$15923 ( \16266 , \4712 , RI9871c80_137);
or \U$15924 ( \16267 , \16266 , \1746 );
nand \U$15925 ( \16268 , \16265 , \16267 );
or \U$15926 ( \16269 , \8171 , \6048 );
not \U$15927 ( \16270 , \15847 );
or \U$15928 ( \16271 , \16270 , \4102 );
nand \U$15929 ( \16272 , \16269 , \16271 );
xor \U$15930 ( \16273 , \16268 , \16272 );
or \U$15931 ( \16274 , \15944 , \1470 );
not \U$15932 ( \16275 , \6431 );
or \U$15933 ( \16276 , \15612 , \16275 );
nand \U$15934 ( \16277 , \16274 , \16276 );
xor \U$15935 ( \16278 , \16273 , \16277 );
xor \U$15936 ( \16279 , \16262 , \16278 );
xor \U$15937 ( \16280 , \16249 , \16279 );
not \U$15938 ( \16281 , \15993 );
not \U$15939 ( \16282 , \16007 );
or \U$15940 ( \16283 , \16281 , \16282 );
or \U$15941 ( \16284 , \16007 , \15993 );
nand \U$15942 ( \16285 , \16283 , \16284 );
xor \U$15943 ( \16286 , \16280 , \16285 );
xor \U$15944 ( \16287 , \16245 , \16286 );
xor \U$15945 ( \16288 , \16219 , \16232 );
xnor \U$15946 ( \16289 , \16288 , \16212 );
and \U$15947 ( \16290 , \16287 , \16289 );
and \U$15948 ( \16291 , \16245 , \16286 );
or \U$15949 ( \16292 , \16290 , \16291 );
xor \U$15950 ( \16293 , \16249 , \16279 );
and \U$15951 ( \16294 , \16293 , \16285 );
and \U$15952 ( \16295 , \16249 , \16279 );
or \U$15953 ( \16296 , \16294 , \16295 );
not \U$15954 ( \16297 , \1518 );
not \U$15955 ( \16298 , \8300 );
or \U$15956 ( \16299 , \16297 , \16298 );
or \U$15957 ( \16300 , \16266 , \1591 );
nand \U$15958 ( \16301 , \16299 , \16300 );
not \U$15959 ( \16302 , \16301 );
not \U$15960 ( \16303 , \8043 );
or \U$15961 ( \16304 , \16302 , \16303 );
or \U$15962 ( \16305 , \8043 , \16301 );
nand \U$15963 ( \16306 , \16304 , \16305 );
not \U$15964 ( \16307 , \8288 );
or \U$15965 ( \16308 , \16307 , \1543 );
not \U$15966 ( \16309 , \16104 );
or \U$15967 ( \16310 , \16309 , \1293 );
nand \U$15968 ( \16311 , \16308 , \16310 );
xnor \U$15969 ( \16312 , \16306 , \16311 );
not \U$15970 ( \16313 , \16312 );
not \U$15971 ( \16314 , \16122 );
not \U$15972 ( \16315 , \16314 );
not \U$15973 ( \16316 , \16131 );
or \U$15974 ( \16317 , \16315 , \16316 );
or \U$15975 ( \16318 , \16131 , \16314 );
nand \U$15976 ( \16319 , \16317 , \16318 );
not \U$15977 ( \16320 , \16319 );
not \U$15978 ( \16321 , \16125 );
not \U$15979 ( \16322 , \16321 );
or \U$15980 ( \16323 , \16320 , \16322 );
nand \U$15981 ( \16324 , \16131 , \16122 );
nand \U$15982 ( \16325 , \16323 , \16324 );
not \U$15983 ( \16326 , \16325 );
not \U$15984 ( \16327 , \16201 );
xor \U$15985 ( \16328 , \16327 , \16210 );
not \U$15986 ( \16329 , \16204 );
and \U$15987 ( \16330 , \16328 , \16329 );
and \U$15988 ( \16331 , \16327 , \16210 );
nor \U$15989 ( \16332 , \16330 , \16331 );
not \U$15990 ( \16333 , \16332 );
or \U$15991 ( \16334 , \16326 , \16333 );
or \U$15992 ( \16335 , \16332 , \16325 );
nand \U$15993 ( \16336 , \16334 , \16335 );
not \U$15994 ( \16337 , \16336 );
or \U$15995 ( \16338 , \16313 , \16337 );
or \U$15996 ( \16339 , \16336 , \16312 );
nand \U$15997 ( \16340 , \16338 , \16339 );
not \U$15998 ( \16341 , \16340 );
nand \U$15999 ( \16342 , \16223 , \16194 );
not \U$16000 ( \16343 , \16193 );
not \U$16001 ( \16344 , \16211 );
or \U$16002 ( \16345 , \16343 , \16344 );
nand \U$16003 ( \16346 , \16345 , \16176 );
nand \U$16004 ( \16347 , \16342 , \16346 );
xor \U$16005 ( \16348 , \16253 , \16261 );
and \U$16006 ( \16349 , \16348 , \16278 );
and \U$16007 ( \16350 , \16253 , \16261 );
or \U$16008 ( \16351 , \16349 , \16350 );
not \U$16009 ( \16352 , \16351 );
and \U$16010 ( \16353 , \16347 , \16352 );
not \U$16011 ( \16354 , \16347 );
and \U$16012 ( \16355 , \16354 , \16351 );
or \U$16013 ( \16356 , \16353 , \16355 );
not \U$16014 ( \16357 , \16356 );
not \U$16015 ( \16358 , \16357 );
or \U$16016 ( \16359 , \16341 , \16358 );
not \U$16017 ( \16360 , \16340 );
nand \U$16018 ( \16361 , \16360 , \16356 );
nand \U$16019 ( \16362 , \16359 , \16361 );
xor \U$16020 ( \16363 , \16296 , \16362 );
xor \U$16021 ( \16364 , \8118 , \8124 );
xor \U$16022 ( \16365 , \16364 , \8135 );
not \U$16023 ( \16366 , \16108 );
not \U$16024 ( \16367 , \15719 );
or \U$16025 ( \16368 , \16366 , \16367 );
not \U$16026 ( \16369 , \16097 );
nand \U$16027 ( \16370 , \16369 , \16112 );
nand \U$16028 ( \16371 , \16368 , \16370 );
xor \U$16029 ( \16372 , \16365 , \16371 );
xor \U$16030 ( \16373 , \8160 , \8149 );
xor \U$16031 ( \16374 , \16373 , \8174 );
xor \U$16032 ( \16375 , \16372 , \16374 );
not \U$16033 ( \16376 , \16142 );
not \U$16034 ( \16377 , \16136 );
or \U$16035 ( \16378 , \16376 , \16377 );
not \U$16036 ( \16379 , \16116 );
nand \U$16037 ( \16380 , \16379 , \16132 );
nand \U$16038 ( \16381 , \16378 , \16380 );
not \U$16039 ( \16382 , \16381 );
xor \U$16040 ( \16383 , \16375 , \16382 );
xor \U$16041 ( \16384 , \16268 , \16272 );
and \U$16042 ( \16385 , \16384 , \16277 );
and \U$16043 ( \16386 , \16268 , \16272 );
nor \U$16044 ( \16387 , \16385 , \16386 );
not \U$16045 ( \16388 , \16387 );
or \U$16046 ( \16389 , \16186 , \16181 );
nand \U$16047 ( \16390 , \16389 , \16192 );
nand \U$16048 ( \16391 , \16186 , \16181 );
nand \U$16049 ( \16392 , \16390 , \16391 );
not \U$16050 ( \16393 , \16164 );
not \U$16051 ( \16394 , \16175 );
or \U$16052 ( \16395 , \16393 , \16394 );
nand \U$16053 ( \16396 , \16174 , \16169 );
nand \U$16054 ( \16397 , \16395 , \16396 );
xor \U$16055 ( \16398 , \16392 , \16397 );
not \U$16056 ( \16399 , \16398 );
or \U$16057 ( \16400 , \16388 , \16399 );
or \U$16058 ( \16401 , \16398 , \16387 );
nand \U$16059 ( \16402 , \16400 , \16401 );
xnor \U$16060 ( \16403 , \16383 , \16402 );
xor \U$16061 ( \16404 , \16363 , \16403 );
xor \U$16062 ( \16405 , \16292 , \16404 );
xor \U$16063 ( \16406 , \15604 , \15665 );
and \U$16064 ( \16407 , \16406 , \15677 );
and \U$16065 ( \16408 , \15604 , \15665 );
or \U$16066 ( \16409 , \16407 , \16408 );
xor \U$16067 ( \16410 , \15735 , \15739 );
and \U$16068 ( \16411 , \16410 , \15770 );
and \U$16069 ( \16412 , \15735 , \15739 );
or \U$16070 ( \16413 , \16411 , \16412 );
xor \U$16071 ( \16414 , \16409 , \16413 );
xor \U$16072 ( \16415 , \16147 , \16153 );
xnor \U$16073 ( \16416 , \16415 , \16092 );
and \U$16074 ( \16417 , \16414 , \16416 );
and \U$16075 ( \16418 , \16409 , \16413 );
or \U$16076 ( \16419 , \16417 , \16418 );
and \U$16077 ( \16420 , \16405 , \16419 );
and \U$16078 ( \16421 , \16292 , \16404 );
or \U$16079 ( \16422 , \16420 , \16421 );
not \U$16080 ( \16423 , \16422 );
xor \U$16081 ( \16424 , \16238 , \16423 );
xor \U$16082 ( \16425 , \16296 , \16362 );
and \U$16083 ( \16426 , \16425 , \16403 );
and \U$16084 ( \16427 , \16296 , \16362 );
or \U$16085 ( \16428 , \16426 , \16427 );
not \U$16086 ( \16429 , \16428 );
not \U$16087 ( \16430 , \16429 );
not \U$16088 ( \16431 , \16356 );
not \U$16089 ( \16432 , \16340 );
or \U$16090 ( \16433 , \16431 , \16432 );
not \U$16091 ( \16434 , \16342 );
not \U$16092 ( \16435 , \16346 );
or \U$16093 ( \16436 , \16434 , \16435 );
nand \U$16094 ( \16437 , \16436 , \16351 );
nand \U$16095 ( \16438 , \16433 , \16437 );
not \U$16096 ( \16439 , \16375 );
xnor \U$16097 ( \16440 , \16382 , \16402 );
not \U$16098 ( \16441 , \16440 );
or \U$16099 ( \16442 , \16439 , \16441 );
nand \U$16100 ( \16443 , \16402 , \16381 );
nand \U$16101 ( \16444 , \16442 , \16443 );
not \U$16102 ( \16445 , \16444 );
xor \U$16103 ( \16446 , \16438 , \16445 );
not \U$16104 ( \16447 , \15962 );
not \U$16105 ( \16448 , \15957 );
or \U$16106 ( \16449 , \16447 , \16448 );
nand \U$16107 ( \16450 , \15947 , \15956 );
nand \U$16108 ( \16451 , \16449 , \16450 );
xor \U$16109 ( \16452 , \8347 , \8354 );
xor \U$16110 ( \16453 , \16451 , \16452 );
not \U$16111 ( \16454 , \7898 );
not \U$16112 ( \16455 , \16454 );
buf \U$16113 ( \16456 , \7917 );
not \U$16114 ( \16457 , \16456 );
or \U$16115 ( \16458 , \16455 , \16457 );
or \U$16116 ( \16459 , \16456 , \16454 );
nand \U$16117 ( \16460 , \16458 , \16459 );
xnor \U$16118 ( \16461 , \16453 , \16460 );
xor \U$16119 ( \16462 , \8138 , \8220 );
xnor \U$16120 ( \16463 , \16462 , \8179 );
xor \U$16121 ( \16464 , \16461 , \16463 );
not \U$16122 ( \16465 , \16312 );
not \U$16123 ( \16466 , \16465 );
not \U$16124 ( \16467 , \16336 );
or \U$16125 ( \16468 , \16466 , \16467 );
not \U$16126 ( \16469 , \16332 );
nand \U$16127 ( \16470 , \16469 , \16325 );
nand \U$16128 ( \16471 , \16468 , \16470 );
not \U$16129 ( \16472 , \16471 );
xnor \U$16130 ( \16473 , \16464 , \16472 );
xor \U$16131 ( \16474 , \16446 , \16473 );
not \U$16132 ( \16475 , \16474 );
or \U$16133 ( \16476 , \16430 , \16475 );
or \U$16134 ( \16477 , \16429 , \16474 );
nand \U$16135 ( \16478 , \16476 , \16477 );
not \U$16136 ( \16479 , \16478 );
xor \U$16137 ( \16480 , \8015 , \8103 );
not \U$16138 ( \16481 , \16061 );
not \U$16139 ( \16482 , \16050 );
or \U$16140 ( \16483 , \16481 , \16482 );
not \U$16141 ( \16484 , \16046 );
nand \U$16142 ( \16485 , \16484 , \16030 );
nand \U$16143 ( \16486 , \16483 , \16485 );
not \U$16144 ( \16487 , \16486 );
xnor \U$16145 ( \16488 , \16480 , \16487 );
not \U$16146 ( \16489 , \16387 );
not \U$16147 ( \16490 , \16489 );
not \U$16148 ( \16491 , \16398 );
or \U$16149 ( \16492 , \16490 , \16491 );
nand \U$16150 ( \16493 , \16397 , \16392 );
nand \U$16151 ( \16494 , \16492 , \16493 );
xor \U$16152 ( \16495 , \16488 , \16494 );
xor \U$16153 ( \16496 , \8293 , \8302 );
xor \U$16154 ( \16497 , \16496 , \8308 );
xor \U$16155 ( \16498 , \7827 , \7836 );
xor \U$16156 ( \16499 , \16498 , \7847 );
xor \U$16157 ( \16500 , \16497 , \16499 );
xor \U$16158 ( \16501 , \7861 , \7872 );
xor \U$16159 ( \16502 , \16501 , \7882 );
xor \U$16160 ( \16503 , \16500 , \16502 );
not \U$16161 ( \16504 , \16081 );
not \U$16162 ( \16505 , \16504 );
not \U$16163 ( \16506 , \16012 );
or \U$16164 ( \16507 , \16505 , \16506 );
not \U$16165 ( \16508 , \16077 );
nand \U$16166 ( \16509 , \16508 , \16063 );
nand \U$16167 ( \16510 , \16507 , \16509 );
xor \U$16168 ( \16511 , \16503 , \16510 );
xor \U$16169 ( \16512 , \16495 , \16511 );
and \U$16170 ( \16513 , \15989 , \16088 );
and \U$16171 ( \16514 , \15968 , \15988 );
nor \U$16172 ( \16515 , \16513 , \16514 );
xor \U$16173 ( \16516 , \16365 , \16371 );
and \U$16174 ( \16517 , \16516 , \16374 );
and \U$16175 ( \16518 , \16365 , \16371 );
or \U$16176 ( \16519 , \16517 , \16518 );
xor \U$16177 ( \16520 , \15963 , \15964 );
and \U$16178 ( \16521 , \16520 , \15967 );
and \U$16179 ( \16522 , \15963 , \15964 );
or \U$16180 ( \16523 , \16521 , \16522 );
xor \U$16181 ( \16524 , \16519 , \16523 );
xor \U$16182 ( \16525 , \7788 , \7803 );
xor \U$16183 ( \16526 , \16525 , \7814 );
and \U$16184 ( \16527 , \16311 , \16306 );
and \U$16185 ( \16528 , \8044 , \16301 );
nor \U$16186 ( \16529 , \16527 , \16528 );
xor \U$16187 ( \16530 , \16526 , \16529 );
xor \U$16188 ( \16531 , \8369 , \8379 );
xnor \U$16189 ( \16532 , \16531 , \8375 );
xnor \U$16190 ( \16533 , \16530 , \16532 );
xnor \U$16191 ( \16534 , \16524 , \16533 );
and \U$16192 ( \16535 , \16515 , \16534 );
not \U$16193 ( \16536 , \16515 );
not \U$16194 ( \16537 , \16534 );
and \U$16195 ( \16538 , \16536 , \16537 );
nor \U$16196 ( \16539 , \16535 , \16538 );
xnor \U$16197 ( \16540 , \16512 , \16539 );
not \U$16198 ( \16541 , \16540 );
and \U$16199 ( \16542 , \16479 , \16541 );
and \U$16200 ( \16543 , \16478 , \16540 );
nor \U$16201 ( \16544 , \16542 , \16543 );
xor \U$16202 ( \16545 , \16424 , \16544 );
xor \U$16203 ( \16546 , \16409 , \16413 );
xor \U$16204 ( \16547 , \16546 , \16416 );
not \U$16205 ( \16548 , \16547 );
not \U$16206 ( \16549 , \16548 );
buf \U$16207 ( \16550 , \15902 );
nand \U$16208 ( \16551 , \16550 , \15805 );
not \U$16209 ( \16552 , \16551 );
not \U$16210 ( \16553 , \15800 );
not \U$16211 ( \16554 , \16553 );
or \U$16212 ( \16555 , \16552 , \16554 );
not \U$16213 ( \16556 , \16550 );
nand \U$16214 ( \16557 , \16556 , \15806 );
nand \U$16215 ( \16558 , \16555 , \16557 );
xor \U$16216 ( \16559 , \16245 , \16286 );
xor \U$16217 ( \16560 , \16559 , \16289 );
and \U$16218 ( \16561 , \16558 , \16560 );
not \U$16219 ( \16562 , \16558 );
not \U$16220 ( \16563 , \16560 );
and \U$16221 ( \16564 , \16562 , \16563 );
or \U$16222 ( \16565 , \16561 , \16564 );
not \U$16223 ( \16566 , \16565 );
or \U$16224 ( \16567 , \16549 , \16566 );
nand \U$16225 ( \16568 , \16558 , \16563 );
nand \U$16226 ( \16569 , \16567 , \16568 );
not \U$16227 ( \16570 , \16569 );
xor \U$16228 ( \16571 , \16090 , \16157 );
xor \U$16229 ( \16572 , \16571 , \16235 );
not \U$16230 ( \16573 , \16572 );
xor \U$16231 ( \16574 , \16292 , \16404 );
xor \U$16232 ( \16575 , \16574 , \16419 );
buf \U$16233 ( \16576 , \16575 );
not \U$16234 ( \16577 , \16576 );
or \U$16235 ( \16578 , \16573 , \16577 );
or \U$16236 ( \16579 , \16576 , \16572 );
nand \U$16237 ( \16580 , \16578 , \16579 );
not \U$16238 ( \16581 , \16580 );
or \U$16239 ( \16582 , \16570 , \16581 );
not \U$16240 ( \16583 , \16576 );
nand \U$16241 ( \16584 , \16583 , \16572 );
nand \U$16242 ( \16585 , \16582 , \16584 );
nand \U$16243 ( \16586 , \16545 , \16585 );
buf \U$16244 ( \16587 , \16586 );
xor \U$16245 ( \16588 , \16451 , \16460 );
and \U$16246 ( \16589 , \16588 , \16452 );
and \U$16247 ( \16590 , \16451 , \16460 );
nor \U$16248 ( \16591 , \16589 , \16590 );
xor \U$16249 ( \16592 , \16499 , \16502 );
and \U$16250 ( \16593 , \16592 , \16497 );
and \U$16251 ( \16594 , \16499 , \16502 );
nor \U$16252 ( \16595 , \16593 , \16594 );
xor \U$16253 ( \16596 , \16591 , \16595 );
not \U$16254 ( \16597 , \16526 );
xor \U$16255 ( \16598 , \8369 , \16529 );
xnor \U$16256 ( \16599 , \16598 , \8383 );
not \U$16257 ( \16600 , \16599 );
or \U$16258 ( \16601 , \16597 , \16600 );
not \U$16259 ( \16602 , \16529 );
nand \U$16260 ( \16603 , \16602 , \16532 );
nand \U$16261 ( \16604 , \16601 , \16603 );
xnor \U$16262 ( \16605 , \16596 , \16604 );
and \U$16263 ( \16606 , \16511 , \16495 );
and \U$16264 ( \16607 , \16503 , \16510 );
nor \U$16265 ( \16608 , \16606 , \16607 );
xor \U$16266 ( \16609 , \16605 , \16608 );
xor \U$16267 ( \16610 , \8281 , \8312 );
not \U$16268 ( \16611 , \16610 );
not \U$16269 ( \16612 , \8109 );
not \U$16270 ( \16613 , \8228 );
or \U$16271 ( \16614 , \16612 , \16613 );
or \U$16272 ( \16615 , \8228 , \8109 );
nand \U$16273 ( \16616 , \16614 , \16615 );
not \U$16274 ( \16617 , \16616 );
not \U$16275 ( \16618 , \16617 );
or \U$16276 ( \16619 , \16611 , \16618 );
not \U$16277 ( \16620 , \16610 );
nand \U$16278 ( \16621 , \16620 , \16616 );
nand \U$16279 ( \16622 , \16619 , \16621 );
not \U$16280 ( \16623 , \16488 );
not \U$16281 ( \16624 , \16494 );
or \U$16282 ( \16625 , \16623 , \16624 );
not \U$16283 ( \16626 , \16487 );
nand \U$16284 ( \16627 , \16626 , \16480 );
nand \U$16285 ( \16628 , \16625 , \16627 );
xnor \U$16286 ( \16629 , \16622 , \16628 );
xor \U$16287 ( \16630 , \16609 , \16629 );
not \U$16288 ( \16631 , \16630 );
not \U$16289 ( \16632 , \16631 );
not \U$16290 ( \16633 , \16478 );
not \U$16291 ( \16634 , \16540 );
not \U$16292 ( \16635 , \16634 );
or \U$16293 ( \16636 , \16633 , \16635 );
nand \U$16294 ( \16637 , \16474 , \16428 );
nand \U$16295 ( \16638 , \16636 , \16637 );
not \U$16296 ( \16639 , \16638 );
not \U$16297 ( \16640 , \16639 );
or \U$16298 ( \16641 , \16632 , \16640 );
nand \U$16299 ( \16642 , \16638 , \16630 );
nand \U$16300 ( \16643 , \16641 , \16642 );
not \U$16301 ( \16644 , \16512 );
not \U$16302 ( \16645 , \16539 );
or \U$16303 ( \16646 , \16644 , \16645 );
not \U$16304 ( \16647 , \16515 );
nand \U$16305 ( \16648 , \16647 , \16537 );
nand \U$16306 ( \16649 , \16646 , \16648 );
xor \U$16307 ( \16650 , \7817 , \7850 );
xor \U$16308 ( \16651 , \16650 , \7885 );
not \U$16309 ( \16652 , \8388 );
not \U$16310 ( \16653 , \8362 );
and \U$16311 ( \16654 , \16652 , \16653 );
and \U$16312 ( \16655 , \8388 , \8362 );
nor \U$16313 ( \16656 , \16654 , \16655 );
xnor \U$16314 ( \16657 , \16651 , \16656 );
not \U$16315 ( \16658 , \16657 );
xor \U$16316 ( \16659 , \8269 , \8271 );
xor \U$16317 ( \16660 , \16659 , \8274 );
not \U$16318 ( \16661 , \16660 );
and \U$16319 ( \16662 , \16658 , \16661 );
and \U$16320 ( \16663 , \16657 , \16660 );
nor \U$16321 ( \16664 , \16662 , \16663 );
and \U$16322 ( \16665 , \16533 , \16524 );
and \U$16323 ( \16666 , \16519 , \16523 );
nor \U$16324 ( \16667 , \16665 , \16666 );
xor \U$16325 ( \16668 , \16664 , \16667 );
not \U$16326 ( \16669 , \16472 );
not \U$16327 ( \16670 , \16461 );
and \U$16328 ( \16671 , \16669 , \16670 );
not \U$16329 ( \16672 , \16461 );
not \U$16330 ( \16673 , \16471 );
or \U$16331 ( \16674 , \16672 , \16673 );
or \U$16332 ( \16675 , \16471 , \16461 );
nand \U$16333 ( \16676 , \16674 , \16675 );
and \U$16334 ( \16677 , \16676 , \16463 );
nor \U$16335 ( \16678 , \16671 , \16677 );
xor \U$16336 ( \16679 , \16668 , \16678 );
not \U$16337 ( \16680 , \16679 );
not \U$16338 ( \16681 , \16473 );
and \U$16339 ( \16682 , \16681 , \16438 );
not \U$16340 ( \16683 , \16681 );
not \U$16341 ( \16684 , \16438 );
and \U$16342 ( \16685 , \16683 , \16684 );
nor \U$16343 ( \16686 , \16682 , \16685 );
not \U$16344 ( \16687 , \16686 );
not \U$16345 ( \16688 , \16444 );
or \U$16346 ( \16689 , \16687 , \16688 );
nand \U$16347 ( \16690 , \16681 , \16438 );
nand \U$16348 ( \16691 , \16689 , \16690 );
not \U$16349 ( \16692 , \16691 );
or \U$16350 ( \16693 , \16680 , \16692 );
or \U$16351 ( \16694 , \16691 , \16679 );
nand \U$16352 ( \16695 , \16693 , \16694 );
xor \U$16353 ( \16696 , \16649 , \16695 );
not \U$16354 ( \16697 , \16696 );
and \U$16355 ( \16698 , \16643 , \16697 );
not \U$16356 ( \16699 , \16643 );
and \U$16357 ( \16700 , \16699 , \16696 );
nor \U$16358 ( \16701 , \16698 , \16700 );
xor \U$16359 ( \16702 , \16238 , \16423 );
and \U$16360 ( \16703 , \16702 , \16544 );
and \U$16361 ( \16704 , \16238 , \16423 );
or \U$16362 ( \16705 , \16703 , \16704 );
nand \U$16363 ( \16706 , \16701 , \16705 );
xor \U$16364 ( \16707 , \16572 , \16575 );
xnor \U$16365 ( \16708 , \16707 , \16569 );
xor \U$16366 ( \16709 , \16547 , \16565 );
not \U$16367 ( \16710 , \16709 );
not \U$16368 ( \16711 , \16710 );
and \U$16369 ( \16712 , \15795 , \15910 );
or \U$16370 ( \16713 , \16712 , \15788 );
or \U$16371 ( \16714 , \15910 , \15795 );
nand \U$16372 ( \16715 , \16713 , \16714 );
not \U$16373 ( \16716 , \16715 );
xor \U$16374 ( \16717 , \15678 , \15771 );
and \U$16375 ( \16718 , \16717 , \15781 );
and \U$16376 ( \16719 , \15678 , \15771 );
nor \U$16377 ( \16720 , \16718 , \16719 );
xnor \U$16378 ( \16721 , \16716 , \16720 );
not \U$16379 ( \16722 , \16721 );
or \U$16380 ( \16723 , \16711 , \16722 );
not \U$16381 ( \16724 , \16716 );
nand \U$16382 ( \16725 , \16724 , \16720 );
nand \U$16383 ( \16726 , \16723 , \16725 );
nand \U$16384 ( \16727 , \16708 , \16726 );
xor \U$16385 ( \16728 , \15782 , \15912 );
and \U$16386 ( \16729 , \16728 , \15917 );
and \U$16387 ( \16730 , \15782 , \15912 );
or \U$16388 ( \16731 , \16729 , \16730 );
not \U$16389 ( \16732 , \16731 );
not \U$16390 ( \16733 , \16710 );
not \U$16391 ( \16734 , \16721 );
not \U$16392 ( \16735 , \16734 );
or \U$16393 ( \16736 , \16733 , \16735 );
nand \U$16394 ( \16737 , \16721 , \16709 );
nand \U$16395 ( \16738 , \16736 , \16737 );
nand \U$16396 ( \16739 , \16732 , \16738 );
and \U$16397 ( \16740 , \16727 , \16739 );
and \U$16398 ( \16741 , \16587 , \16706 , \16740 );
nand \U$16399 ( \16742 , \16643 , \16696 );
xor \U$16400 ( \16743 , \8243 , \8245 );
xor \U$16401 ( \16744 , \16743 , \8248 );
not \U$16402 ( \16745 , \16744 );
not \U$16403 ( \16746 , \7958 );
not \U$16404 ( \16747 , \7965 );
or \U$16405 ( \16748 , \16746 , \16747 );
nand \U$16406 ( \16749 , \7966 , \7957 );
nand \U$16407 ( \16750 , \16748 , \16749 );
not \U$16408 ( \16751 , \8233 );
and \U$16409 ( \16752 , \16750 , \16751 );
not \U$16410 ( \16753 , \16750 );
and \U$16411 ( \16754 , \16753 , \8233 );
nor \U$16412 ( \16755 , \16752 , \16754 );
not \U$16413 ( \16756 , \16755 );
or \U$16414 ( \16757 , \16745 , \16756 );
or \U$16415 ( \16758 , \16755 , \16744 );
nand \U$16416 ( \16759 , \16757 , \16758 );
not \U$16417 ( \16760 , \16628 );
not \U$16418 ( \16761 , \16622 );
or \U$16419 ( \16762 , \16760 , \16761 );
nand \U$16420 ( \16763 , \16616 , \16610 );
nand \U$16421 ( \16764 , \16762 , \16763 );
xor \U$16422 ( \16765 , \16759 , \16764 );
xor \U$16423 ( \16766 , \16664 , \16667 );
and \U$16424 ( \16767 , \16766 , \16678 );
and \U$16425 ( \16768 , \16664 , \16667 );
or \U$16426 ( \16769 , \16767 , \16768 );
not \U$16427 ( \16770 , \8398 );
not \U$16428 ( \16771 , \8277 );
and \U$16429 ( \16772 , \16770 , \16771 );
and \U$16430 ( \16773 , \8398 , \8277 );
nor \U$16431 ( \16774 , \16772 , \16773 );
not \U$16432 ( \16775 , \16774 );
not \U$16433 ( \16776 , \16775 );
not \U$16434 ( \16777 , \16591 );
nor \U$16435 ( \16778 , \16604 , \16777 );
or \U$16436 ( \16779 , \16778 , \16595 );
nand \U$16437 ( \16780 , \16604 , \16777 );
nand \U$16438 ( \16781 , \16779 , \16780 );
not \U$16439 ( \16782 , \16781 );
not \U$16440 ( \16783 , \16782 );
or \U$16441 ( \16784 , \16776 , \16783 );
nand \U$16442 ( \16785 , \16781 , \16774 );
nand \U$16443 ( \16786 , \16784 , \16785 );
not \U$16444 ( \16787 , \16786 );
not \U$16445 ( \16788 , \16660 );
not \U$16446 ( \16789 , \16788 );
not \U$16447 ( \16790 , \16657 );
or \U$16448 ( \16791 , \16789 , \16790 );
not \U$16449 ( \16792 , \16656 );
nand \U$16450 ( \16793 , \16792 , \16651 );
nand \U$16451 ( \16794 , \16791 , \16793 );
not \U$16452 ( \16795 , \16794 );
not \U$16453 ( \16796 , \16795 );
and \U$16454 ( \16797 , \16787 , \16796 );
and \U$16455 ( \16798 , \16786 , \16795 );
nor \U$16456 ( \16799 , \16797 , \16798 );
xor \U$16457 ( \16800 , \16769 , \16799 );
xor \U$16458 ( \16801 , \16605 , \16608 );
and \U$16459 ( \16802 , \16801 , \16629 );
and \U$16460 ( \16803 , \16605 , \16608 );
or \U$16461 ( \16804 , \16802 , \16803 );
xor \U$16462 ( \16805 , \16800 , \16804 );
xor \U$16463 ( \16806 , \16765 , \16805 );
not \U$16464 ( \16807 , \16649 );
not \U$16465 ( \16808 , \16695 );
or \U$16466 ( \16809 , \16807 , \16808 );
not \U$16467 ( \16810 , \16679 );
nand \U$16468 ( \16811 , \16810 , \16691 );
nand \U$16469 ( \16812 , \16809 , \16811 );
xor \U$16470 ( \16813 , \16806 , \16812 );
nand \U$16471 ( \16814 , \16638 , \16631 );
nand \U$16472 ( \16815 , \16742 , \16813 , \16814 );
not \U$16473 ( \16816 , \16765 );
nand \U$16474 ( \16817 , \16816 , \16805 );
not \U$16475 ( \16818 , \16817 );
not \U$16476 ( \16819 , \16812 );
or \U$16477 ( \16820 , \16818 , \16819 );
not \U$16478 ( \16821 , \16805 );
nand \U$16479 ( \16822 , \16821 , \16765 );
nand \U$16480 ( \16823 , \16820 , \16822 );
not \U$16481 ( \16824 , \16823 );
not \U$16482 ( \16825 , \16755 );
not \U$16483 ( \16826 , \16744 );
not \U$16484 ( \16827 , \16826 );
and \U$16485 ( \16828 , \16825 , \16827 );
and \U$16486 ( \16829 , \16759 , \16764 );
nor \U$16487 ( \16830 , \16828 , \16829 );
xor \U$16488 ( \16831 , \16769 , \16799 );
and \U$16489 ( \16832 , \16831 , \16804 );
and \U$16490 ( \16833 , \16769 , \16799 );
or \U$16491 ( \16834 , \16832 , \16833 );
xor \U$16492 ( \16835 , \16830 , \16834 );
and \U$16493 ( \16836 , \8262 , \8403 );
not \U$16494 ( \16837 , \8262 );
and \U$16495 ( \16838 , \16837 , \8402 );
or \U$16496 ( \16839 , \16836 , \16838 );
xor \U$16497 ( \16840 , \7948 , \7950 );
xor \U$16498 ( \16841 , \16840 , \8235 );
xor \U$16499 ( \16842 , \16839 , \16841 );
not \U$16500 ( \16843 , \16794 );
not \U$16501 ( \16844 , \16786 );
or \U$16502 ( \16845 , \16843 , \16844 );
nand \U$16503 ( \16846 , \16781 , \16775 );
nand \U$16504 ( \16847 , \16845 , \16846 );
xnor \U$16505 ( \16848 , \16842 , \16847 );
xor \U$16506 ( \16849 , \16835 , \16848 );
nand \U$16507 ( \16850 , \16824 , \16849 );
xor \U$16508 ( \16851 , \16830 , \16834 );
and \U$16509 ( \16852 , \16851 , \16848 );
and \U$16510 ( \16853 , \16830 , \16834 );
or \U$16511 ( \16854 , \16852 , \16853 );
xor \U$16512 ( \16855 , \8422 , \8417 );
xor \U$16513 ( \16856 , \16855 , \8420 );
xor \U$16514 ( \16857 , \8238 , \8240 );
xor \U$16515 ( \16858 , \16857 , \8405 );
xor \U$16516 ( \16859 , \16856 , \16858 );
not \U$16517 ( \16860 , \16839 );
not \U$16518 ( \16861 , \16847 );
or \U$16519 ( \16862 , \16860 , \16861 );
or \U$16520 ( \16863 , \16847 , \16839 );
nand \U$16521 ( \16864 , \16863 , \16841 );
nand \U$16522 ( \16865 , \16862 , \16864 );
xnor \U$16523 ( \16866 , \16859 , \16865 );
nand \U$16524 ( \16867 , \16854 , \16866 );
and \U$16525 ( \16868 , \16815 , \16850 , \16867 );
or \U$16526 ( \16869 , \16856 , \16858 );
nand \U$16527 ( \16870 , \16869 , \16865 );
not \U$16528 ( \16871 , \8427 );
not \U$16529 ( \16872 , \7768 );
xor \U$16530 ( \16873 , \16871 , \16872 );
xnor \U$16531 ( \16874 , \16873 , \8408 );
nand \U$16532 ( \16875 , \16858 , \16856 );
nand \U$16533 ( \16876 , \16870 , \16874 , \16875 );
nand \U$16534 ( \16877 , \16741 , \16868 , \16876 );
nor \U$16535 ( \16878 , \15937 , \16877 );
not \U$16536 ( \16879 , \16878 );
not \U$16537 ( \16880 , \7338 );
not \U$16538 ( \16881 , RI98729a0_165);
not \U$16539 ( \16882 , \4370 );
or \U$16540 ( \16883 , \16881 , \16882 );
or \U$16541 ( \16884 , \3859 , RI98729a0_165);
nand \U$16542 ( \16885 , \16883 , \16884 );
not \U$16543 ( \16886 , \16885 );
or \U$16544 ( \16887 , \16880 , \16886 );
not \U$16545 ( \16888 , \3536 );
not \U$16546 ( \16889 , \7333 );
and \U$16547 ( \16890 , \16888 , \16889 );
not \U$16548 ( \16891 , \12543 );
not \U$16549 ( \16892 , RI98729a0_165);
and \U$16550 ( \16893 , \16891 , \16892 );
nor \U$16551 ( \16894 , \16890 , \16893 );
not \U$16552 ( \16895 , \16894 );
nand \U$16553 ( \16896 , \16895 , \7325 );
nand \U$16554 ( \16897 , \16887 , \16896 );
not \U$16555 ( \16898 , \6284 );
not \U$16556 ( \16899 , RI98728b0_163);
not \U$16557 ( \16900 , \4176 );
or \U$16558 ( \16901 , \16899 , \16900 );
or \U$16559 ( \16902 , \11028 , RI98728b0_163);
nand \U$16560 ( \16903 , \16901 , \16902 );
not \U$16561 ( \16904 , \16903 );
or \U$16562 ( \16905 , \16898 , \16904 );
not \U$16563 ( \16906 , \14930 );
not \U$16564 ( \16907 , \16906 );
not \U$16565 ( \16908 , RI98728b0_163);
and \U$16566 ( \16909 , \16907 , \16908 );
and \U$16567 ( \16910 , \10698 , RI98728b0_163);
nor \U$16568 ( \16911 , \16909 , \16910 );
nand \U$16569 ( \16912 , \16911 , \6610 );
nand \U$16570 ( \16913 , \16905 , \16912 );
xor \U$16571 ( \16914 , \16897 , \16913 );
not \U$16572 ( \16915 , \9527 );
not \U$16573 ( \16916 , \8732 );
not \U$16574 ( \16917 , \943 );
or \U$16575 ( \16918 , \16916 , \16917 );
or \U$16576 ( \16919 , \8732 , \1550 );
nand \U$16577 ( \16920 , \16918 , \16919 );
not \U$16578 ( \16921 , \16920 );
or \U$16579 ( \16922 , \16915 , \16921 );
not \U$16580 ( \16923 , \845 );
buf \U$16581 ( \16924 , \16923 );
not \U$16582 ( \16925 , \16924 );
not \U$16583 ( \16926 , \16925 );
xor \U$16584 ( \16927 , RI9872f40_177, \16926 );
not \U$16585 ( \16928 , \11199 );
or \U$16586 ( \16929 , \16927 , \16928 );
nand \U$16587 ( \16930 , \16922 , \16929 );
and \U$16588 ( \16931 , \16914 , \16930 );
and \U$16589 ( \16932 , \16897 , \16913 );
or \U$16590 ( \16933 , \16931 , \16932 );
not \U$16591 ( \16934 , \11433 );
and \U$16592 ( \16935 , RI98719b0_131, \8606 );
not \U$16593 ( \16936 , RI98719b0_131);
and \U$16594 ( \16937 , \16936 , \10308 );
nor \U$16595 ( \16938 , \16935 , \16937 );
not \U$16596 ( \16939 , \16938 );
or \U$16597 ( \16940 , \16934 , \16939 );
not \U$16598 ( \16941 , RI98719b0_131);
not \U$16599 ( \16942 , \8877 );
not \U$16600 ( \16943 , \16942 );
or \U$16601 ( \16944 , \16941 , \16943 );
buf \U$16602 ( \16945 , \8873 );
not \U$16603 ( \16946 , \16945 );
or \U$16604 ( \16947 , \16946 , RI98719b0_131);
nand \U$16605 ( \16948 , \16944 , \16947 );
nand \U$16606 ( \16949 , \16948 , \796 );
nand \U$16607 ( \16950 , \16940 , \16949 );
not \U$16608 ( \16951 , \16950 );
not \U$16609 ( \16952 , \6672 );
xnor \U$16610 ( \16953 , \8857 , RI98718c0_129);
not \U$16611 ( \16954 , \16953 );
or \U$16612 ( \16955 , \16952 , \16954 );
and \U$16613 ( \16956 , RI98718c0_129, \8650 );
not \U$16614 ( \16957 , RI98718c0_129);
and \U$16615 ( \16958 , \16957 , \8642 );
or \U$16616 ( \16959 , \16956 , \16958 );
nand \U$16617 ( \16960 , \16959 , \1083 );
nand \U$16618 ( \16961 , \16955 , \16960 );
not \U$16619 ( \16962 , \16961 );
not \U$16620 ( \16963 , \16962 );
or \U$16621 ( \16964 , \16951 , \16963 );
or \U$16622 ( \16965 , \16962 , \16950 );
nand \U$16623 ( \16966 , \16964 , \16965 );
not \U$16624 ( \16967 , \2087 );
and \U$16625 ( \16968 , RI9871aa0_133, \12727 );
not \U$16626 ( \16969 , RI9871aa0_133);
and \U$16627 ( \16970 , \16969 , \8333 );
nor \U$16628 ( \16971 , \16968 , \16970 );
not \U$16629 ( \16972 , \16971 );
or \U$16630 ( \16973 , \16967 , \16972 );
not \U$16631 ( \16974 , RI9871aa0_133);
not \U$16632 ( \16975 , \8074 );
or \U$16633 ( \16976 , \16974 , \16975 );
or \U$16634 ( \16977 , \11628 , RI9871aa0_133);
nand \U$16635 ( \16978 , \16976 , \16977 );
nand \U$16636 ( \16979 , \16978 , \2071 );
nand \U$16637 ( \16980 , \16973 , \16979 );
not \U$16638 ( \16981 , \16980 );
and \U$16639 ( \16982 , \16966 , \16981 );
not \U$16640 ( \16983 , \16966 );
and \U$16641 ( \16984 , \16983 , \16980 );
nor \U$16642 ( \16985 , \16982 , \16984 );
buf \U$16643 ( \16986 , \515 );
buf \U$16644 ( \16987 , \533 );
buf \U$16645 ( \16988 , \576 );
nand \U$16646 ( \16989 , \16987 , \16988 );
not \U$16647 ( \16990 , \16989 );
and \U$16648 ( \16991 , \16986 , \16990 );
not \U$16649 ( \16992 , \16986 );
and \U$16650 ( \16993 , \16992 , \16989 );
nor \U$16651 ( \16994 , \16991 , \16993 );
buf \U$16652 ( \16995 , \16994 );
not \U$16653 ( \16996 , \16995 );
or \U$16654 ( \16997 , \1164 , \16996 );
and \U$16655 ( \16998 , RI9873558_190, RI98735d0_191);
not \U$16656 ( \16999 , RI98734e0_189);
nor \U$16657 ( \17000 , \16998 , \16999 );
xor \U$16658 ( \17001 , \16997 , \17000 );
not \U$16659 ( \17002 , \1017 );
buf \U$16660 ( \17003 , \13931 );
not \U$16661 ( \17004 , \17003 );
not \U$16662 ( \17005 , \17004 );
and \U$16663 ( \17006 , \17005 , \1157 );
not \U$16664 ( \17007 , \17005 );
and \U$16665 ( \17008 , \17007 , \12592 );
nor \U$16666 ( \17009 , \17006 , \17008 );
not \U$16667 ( \17010 , \17009 );
or \U$16668 ( \17011 , \17002 , \17010 );
not \U$16669 ( \17012 , \1157 );
buf \U$16670 ( \17013 , \13859 );
not \U$16671 ( \17014 , \17013 );
not \U$16672 ( \17015 , \17014 );
not \U$16673 ( \17016 , \17015 );
or \U$16674 ( \17017 , \17012 , \17016 );
nand \U$16675 ( \17018 , \13861 , \1043 );
nand \U$16676 ( \17019 , \17017 , \17018 );
nand \U$16677 ( \17020 , \17019 , \1013 );
nand \U$16678 ( \17021 , \17011 , \17020 );
xnor \U$16679 ( \17022 , \17001 , \17021 );
not \U$16680 ( \17023 , \1323 );
and \U$16681 ( \17024 , RI9871b18_134, \12471 );
not \U$16682 ( \17025 , RI9871b18_134);
and \U$16683 ( \17026 , \17025 , \12470 );
or \U$16684 ( \17027 , \17024 , \17026 );
not \U$16685 ( \17028 , \17027 );
or \U$16686 ( \17029 , \17023 , \17028 );
not \U$16687 ( \17030 , \4044 );
not \U$16688 ( \17031 , \9750 );
or \U$16689 ( \17032 , \17030 , \17031 );
not \U$16690 ( \17033 , \8697 );
nand \U$16691 ( \17034 , \17033 , RI9871b18_134);
nand \U$16692 ( \17035 , \17032 , \17034 );
nand \U$16693 ( \17036 , \17035 , \12720 );
nand \U$16694 ( \17037 , \17029 , \17036 );
xor \U$16695 ( \17038 , \17022 , \17037 );
not \U$16696 ( \17039 , \1455 );
and \U$16697 ( \17040 , \10369 , \1619 );
not \U$16698 ( \17041 , \10369 );
and \U$16699 ( \17042 , \17041 , RI9871c08_136);
nor \U$16700 ( \17043 , \17040 , \17042 );
not \U$16701 ( \17044 , \17043 );
or \U$16702 ( \17045 , \17039 , \17044 );
and \U$16703 ( \17046 , \8580 , RI9871c08_136);
not \U$16704 ( \17047 , \8580 );
and \U$16705 ( \17048 , \17047 , \3487 );
nor \U$16706 ( \17049 , \17046 , \17048 );
nand \U$16707 ( \17050 , \17049 , \1429 );
nand \U$16708 ( \17051 , \17045 , \17050 );
xor \U$16709 ( \17052 , \17038 , \17051 );
not \U$16710 ( \17053 , \17052 );
and \U$16711 ( \17054 , \16985 , \17053 );
not \U$16712 ( \17055 , \16985 );
and \U$16713 ( \17056 , \17055 , \17052 );
nor \U$16714 ( \17057 , \17054 , \17056 );
not \U$16715 ( \17058 , \17057 );
xor \U$16716 ( \17059 , \16933 , \17058 );
xor \U$16717 ( \17060 , \16897 , \16913 );
xor \U$16718 ( \17061 , \17060 , \16930 );
not \U$16719 ( \17062 , \17061 );
not \U$16720 ( \17063 , \3467 );
not \U$16721 ( \17064 , \3593 );
not \U$16722 ( \17065 , \6530 );
or \U$16723 ( \17066 , \17064 , \17065 );
or \U$16724 ( \17067 , \8934 , \4063 );
nand \U$16725 ( \17068 , \17066 , \17067 );
not \U$16726 ( \17069 , \17068 );
or \U$16727 ( \17070 , \17063 , \17069 );
not \U$16728 ( \17071 , RI98726d0_159);
xor \U$16729 ( \17072 , \6995 , \6997 );
not \U$16730 ( \17073 , \17072 );
or \U$16731 ( \17074 , \17071 , \17073 );
or \U$16732 ( \17075 , \7002 , RI98726d0_159);
nand \U$16733 ( \17076 , \17074 , \17075 );
nand \U$16734 ( \17077 , \17076 , \3465 );
nand \U$16735 ( \17078 , \17070 , \17077 );
not \U$16736 ( \17079 , \17078 );
not \U$16737 ( \17080 , \17079 );
not \U$16738 ( \17081 , \12772 );
and \U$16739 ( \17082 , RI9871d70_139, \17081 );
not \U$16740 ( \17083 , RI9871d70_139);
and \U$16741 ( \17084 , \17083 , \13268 );
nor \U$16742 ( \17085 , \17082 , \17084 );
not \U$16743 ( \17086 , \17085 );
not \U$16744 ( \17087 , \17086 );
not \U$16745 ( \17088 , \932 );
and \U$16746 ( \17089 , \17087 , \17088 );
not \U$16747 ( \17090 , \13281 );
and \U$16748 ( \17091 , \1347 , \17090 );
not \U$16749 ( \17092 , \1347 );
and \U$16750 ( \17093 , \17092 , \13281 );
nor \U$16751 ( \17094 , \17091 , \17093 );
and \U$16752 ( \17095 , \17094 , \859 );
nor \U$16753 ( \17096 , \17089 , \17095 );
not \U$16754 ( \17097 , \17096 );
buf \U$16755 ( \17098 , \5847 );
not \U$16756 ( \17099 , \17098 );
not \U$16757 ( \17100 , \4088 );
not \U$16758 ( \17101 , \11438 );
or \U$16759 ( \17102 , \17100 , \17101 );
or \U$16760 ( \17103 , \7112 , \6042 );
nand \U$16761 ( \17104 , \17102 , \17103 );
not \U$16762 ( \17105 , \17104 );
or \U$16763 ( \17106 , \17099 , \17105 );
not \U$16764 ( \17107 , \4088 );
not \U$16765 ( \17108 , \12802 );
or \U$16766 ( \17109 , \17107 , \17108 );
nand \U$16767 ( \17110 , \8904 , RI98725e0_157);
nand \U$16768 ( \17111 , \17109 , \17110 );
nand \U$16769 ( \17112 , \17111 , \8790 );
nand \U$16770 ( \17113 , \17106 , \17112 );
not \U$16771 ( \17114 , \17113 );
or \U$16772 ( \17115 , \17097 , \17114 );
or \U$16773 ( \17116 , \17113 , \17096 );
nand \U$16774 ( \17117 , \17115 , \17116 );
buf \U$16775 ( \17118 , \17117 );
not \U$16776 ( \17119 , \17118 );
or \U$16777 ( \17120 , \17080 , \17119 );
or \U$16778 ( \17121 , \17118 , \17079 );
nand \U$16779 ( \17122 , \17120 , \17121 );
buf \U$16780 ( \17123 , \13483 );
not \U$16781 ( \17124 , \17123 );
not \U$16782 ( \17125 , RI9873210_183);
not \U$16783 ( \17126 , \1318 );
or \U$16784 ( \17127 , \17125 , \17126 );
or \U$16785 ( \17128 , \1319 , RI9873210_183);
nand \U$16786 ( \17129 , \17127 , \17128 );
not \U$16787 ( \17130 , \17129 );
or \U$16788 ( \17131 , \17124 , \17130 );
and \U$16789 ( \17132 , RI9873210_183, \1273 );
not \U$16790 ( \17133 , RI9873210_183);
and \U$16791 ( \17134 , \17133 , \1581 );
nor \U$16792 ( \17135 , \17132 , \17134 );
nand \U$16793 ( \17136 , \17135 , \13476 );
nand \U$16794 ( \17137 , \17131 , \17136 );
not \U$16795 ( \17138 , \9312 );
not \U$16796 ( \17139 , RI9872d60_173);
not \U$16797 ( \17140 , \1037 );
not \U$16798 ( \17141 , \17140 );
or \U$16799 ( \17142 , \17139 , \17141 );
buf \U$16800 ( \17143 , \17140 );
or \U$16801 ( \17144 , \17143 , RI9872d60_173);
nand \U$16802 ( \17145 , \17142 , \17144 );
not \U$16803 ( \17146 , \17145 );
or \U$16804 ( \17147 , \17138 , \17146 );
not \U$16805 ( \17148 , \8807 );
not \U$16806 ( \17149 , \1062 );
or \U$16807 ( \17150 , \17148 , \17149 );
or \U$16808 ( \17151 , \6573 , \8811 );
nand \U$16809 ( \17152 , \17150 , \17151 );
nand \U$16810 ( \17153 , \17152 , \8802 );
nand \U$16811 ( \17154 , \17147 , \17153 );
xor \U$16812 ( \17155 , \17137 , \17154 );
not \U$16813 ( \17156 , \9670 );
not \U$16814 ( \17157 , RI9872bf8_170);
not \U$16815 ( \17158 , \5946 );
or \U$16816 ( \17159 , \17157 , \17158 );
or \U$16817 ( \17160 , \1190 , RI9872bf8_170);
nand \U$16818 ( \17161 , \17159 , \17160 );
not \U$16819 ( \17162 , \17161 );
or \U$16820 ( \17163 , \17156 , \17162 );
not \U$16821 ( \17164 , RI9872bf8_170);
not \U$16822 ( \17165 , \17164 );
not \U$16823 ( \17166 , \6020 );
or \U$16824 ( \17167 , \17165 , \17166 );
nand \U$16825 ( \17168 , \1210 , RI9872bf8_170);
nand \U$16826 ( \17169 , \17167 , \17168 );
nand \U$16827 ( \17170 , \17169 , \9668 );
nand \U$16828 ( \17171 , \17163 , \17170 );
and \U$16829 ( \17172 , \17155 , \17171 );
and \U$16830 ( \17173 , \17137 , \17154 );
or \U$16831 ( \17174 , \17172 , \17173 );
xor \U$16832 ( \17175 , \17122 , \17174 );
not \U$16833 ( \17176 , \17175 );
or \U$16834 ( \17177 , \17062 , \17176 );
nand \U$16835 ( \17178 , \17174 , \17122 );
nand \U$16836 ( \17179 , \17177 , \17178 );
xor \U$16837 ( \17180 , \17059 , \17179 );
not \U$16838 ( \17181 , \4925 );
not \U$16839 ( \17182 , RI9872388_152);
not \U$16840 ( \17183 , \5775 );
or \U$16841 ( \17184 , \17182 , \17183 );
nand \U$16842 ( \17185 , \5393 , \4902 );
nand \U$16843 ( \17186 , \17184 , \17185 );
not \U$16844 ( \17187 , \17186 );
or \U$16845 ( \17188 , \17181 , \17187 );
xor \U$16846 ( \17189 , \5766 , RI9872388_152);
nand \U$16847 ( \17190 , \17189 , \4919 );
nand \U$16848 ( \17191 , \17188 , \17190 );
not \U$16849 ( \17192 , \6698 );
not \U$16850 ( \17193 , \4960 );
not \U$16851 ( \17194 , RI9872478_154);
and \U$16852 ( \17195 , \17193 , \17194 );
and \U$16853 ( \17196 , \4960 , RI9872478_154);
nor \U$16854 ( \17197 , \17195 , \17196 );
not \U$16855 ( \17198 , \17197 );
or \U$16856 ( \17199 , \17192 , \17198 );
and \U$16857 ( \17200 , RI9872478_154, \5739 );
not \U$16858 ( \17201 , RI9872478_154);
and \U$16859 ( \17202 , \17201 , \5736 );
nor \U$16860 ( \17203 , \17200 , \17202 );
nand \U$16861 ( \17204 , \17203 , \5034 );
nand \U$16862 ( \17205 , \17199 , \17204 );
xor \U$16863 ( \17206 , \17191 , \17205 );
not \U$16864 ( \17207 , \10333 );
and \U$16865 ( \17208 , RI9872e50_175, \11559 );
not \U$16866 ( \17209 , RI9872e50_175);
and \U$16867 ( \17210 , \17209 , \7019 );
nor \U$16868 ( \17211 , \17208 , \17210 );
not \U$16869 ( \17212 , \17211 );
or \U$16870 ( \17213 , \17207 , \17212 );
not \U$16871 ( \17214 , \9690 );
not \U$16872 ( \17215 , \5712 );
or \U$16873 ( \17216 , \17214 , \17215 );
nand \U$16874 ( \17217 , \1340 , RI9872e50_175);
nand \U$16875 ( \17218 , \17216 , \17217 );
nand \U$16876 ( \17219 , \17218 , \9294 );
nand \U$16877 ( \17220 , \17213 , \17219 );
and \U$16878 ( \17221 , \17206 , \17220 );
and \U$16879 ( \17222 , \17191 , \17205 );
or \U$16880 ( \17223 , \17221 , \17222 );
not \U$16881 ( \17224 , \10624 );
and \U$16882 ( \17225 , RI9872d60_173, \1603 );
not \U$16883 ( \17226 , RI9872d60_173);
and \U$16884 ( \17227 , \17226 , \4454 );
or \U$16885 ( \17228 , \17225 , \17227 );
not \U$16886 ( \17229 , \17228 );
or \U$16887 ( \17230 , \17224 , \17229 );
nand \U$16888 ( \17231 , \17152 , \9312 );
nand \U$16889 ( \17232 , \17230 , \17231 );
not \U$16890 ( \17233 , \17232 );
buf \U$16891 ( \17234 , \13484 );
not \U$16892 ( \17235 , \17234 );
not \U$16893 ( \17236 , RI9873210_183);
not \U$16894 ( \17237 , \1447 );
or \U$16895 ( \17238 , \17236 , \17237 );
or \U$16896 ( \17239 , \2492 , RI9873210_183);
nand \U$16897 ( \17240 , \17238 , \17239 );
not \U$16898 ( \17241 , \17240 );
or \U$16899 ( \17242 , \17235 , \17241 );
not \U$16900 ( \17243 , \13474 );
nand \U$16901 ( \17244 , \17243 , \17129 );
nand \U$16902 ( \17245 , \17242 , \17244 );
or \U$16903 ( \17246 , RI98733f0_187, RI98734e0_189);
not \U$16904 ( \17247 , RI9873468_188);
nand \U$16905 ( \17248 , \17247 , RI98734e0_189);
nand \U$16906 ( \17249 , RI98733f0_187, RI9873468_188);
nand \U$16907 ( \17250 , \17246 , \17248 , \17249 );
not \U$16908 ( \17251 , \17250 );
buf \U$16909 ( \17252 , \17251 );
not \U$16910 ( \17253 , \17252 );
and \U$16911 ( \17254 , RI98733f0_187, \1125 );
not \U$16912 ( \17255 , RI98733f0_187);
and \U$16913 ( \17256 , \17255 , \2398 );
nor \U$16914 ( \17257 , \17254 , \17256 );
not \U$16915 ( \17258 , \17257 );
or \U$16916 ( \17259 , \17253 , \17258 );
xor \U$16917 ( \17260 , RI98733f0_187, \2982 );
nand \U$16918 ( \17261 , \16999 , RI9873468_188);
and \U$16919 ( \17262 , \17261 , \17248 );
not \U$16920 ( \17263 , \17262 );
nand \U$16921 ( \17264 , \17260 , \17263 );
nand \U$16922 ( \17265 , \17259 , \17264 );
and \U$16923 ( \17266 , \17245 , \17265 );
not \U$16924 ( \17267 , \17245 );
not \U$16925 ( \17268 , \17265 );
and \U$16926 ( \17269 , \17267 , \17268 );
nor \U$16927 ( \17270 , \17266 , \17269 );
not \U$16928 ( \17271 , \17270 );
or \U$16929 ( \17272 , \17233 , \17271 );
nand \U$16930 ( \17273 , \17245 , \17265 );
nand \U$16931 ( \17274 , \17272 , \17273 );
xor \U$16932 ( \17275 , \17223 , \17274 );
not \U$16933 ( \17276 , \9214 );
and \U$16934 ( \17277 , \5946 , \11688 );
not \U$16935 ( \17278 , \5946 );
and \U$16936 ( \17279 , \17278 , RI9872b80_169);
nor \U$16937 ( \17280 , \17277 , \17279 );
not \U$16938 ( \17281 , \17280 );
or \U$16939 ( \17282 , \17276 , \17281 );
and \U$16940 ( \17283 , RI9872b80_169, \1485 );
not \U$16941 ( \17284 , RI9872b80_169);
and \U$16942 ( \17285 , \17284 , \3275 );
or \U$16943 ( \17286 , \17283 , \17285 );
nand \U$16944 ( \17287 , \17286 , \10679 );
nand \U$16945 ( \17288 , \17282 , \17287 );
not \U$16946 ( \17289 , \17288 );
not \U$16947 ( \17290 , \12868 );
and \U$16948 ( \17291 , RI98730a8_180, \1581 );
not \U$16949 ( \17292 , RI98730a8_180);
and \U$16950 ( \17293 , \17292 , \1273 );
or \U$16951 ( \17294 , \17291 , \17293 );
not \U$16952 ( \17295 , \17294 );
or \U$16953 ( \17296 , \17290 , \17295 );
not \U$16954 ( \17297 , RI98730a8_180);
not \U$16955 ( \17298 , \915 );
or \U$16956 ( \17299 , \17297 , \17298 );
or \U$16957 ( \17300 , \5480 , RI98730a8_180);
nand \U$16958 ( \17301 , \17299 , \17300 );
nand \U$16959 ( \17302 , \17301 , \13020 );
nand \U$16960 ( \17303 , \17296 , \17302 );
not \U$16961 ( \17304 , \9227 );
xor \U$16962 ( \17305 , \1038 , RI9872bf8_170);
not \U$16963 ( \17306 , \17305 );
or \U$16964 ( \17307 , \17304 , \17306 );
nand \U$16965 ( \17308 , \17169 , \9249 );
nand \U$16966 ( \17309 , \17307 , \17308 );
and \U$16967 ( \17310 , \17303 , \17309 );
not \U$16968 ( \17311 , \17303 );
not \U$16969 ( \17312 , \17309 );
and \U$16970 ( \17313 , \17311 , \17312 );
nor \U$16971 ( \17314 , \17310 , \17313 );
not \U$16972 ( \17315 , \17314 );
or \U$16973 ( \17316 , \17289 , \17315 );
nand \U$16974 ( \17317 , \17309 , \17303 );
nand \U$16975 ( \17318 , \17316 , \17317 );
xor \U$16976 ( \17319 , \17275 , \17318 );
and \U$16977 ( \17320 , \17180 , \17319 );
and \U$16978 ( \17321 , \17059 , \17179 );
or \U$16979 ( \17322 , \17320 , \17321 );
not \U$16980 ( \17323 , \9670 );
not \U$16981 ( \17324 , \17305 );
or \U$16982 ( \17325 , \17323 , \17324 );
not \U$16983 ( \17326 , \9244 );
not \U$16984 ( \17327 , \6573 );
or \U$16985 ( \17328 , \17326 , \17327 );
or \U$16986 ( \17329 , \1062 , \9244 );
nand \U$16987 ( \17330 , \17328 , \17329 );
nand \U$16988 ( \17331 , \17330 , \9668 );
nand \U$16989 ( \17332 , \17325 , \17331 );
not \U$16990 ( \17333 , \17332 );
not \U$16991 ( \17334 , \17333 );
not \U$16992 ( \17335 , \9196 );
not \U$16993 ( \17336 , \17280 );
or \U$16994 ( \17337 , \17335 , \17336 );
and \U$16995 ( \17338 , RI9872b80_169, \6678 );
not \U$16996 ( \17339 , RI9872b80_169);
and \U$16997 ( \17340 , \17339 , \1211 );
or \U$16998 ( \17341 , \17338 , \17340 );
nand \U$16999 ( \17342 , \17341 , \9214 );
nand \U$17000 ( \17343 , \17337 , \17342 );
not \U$17001 ( \17344 , \17343 );
not \U$17002 ( \17345 , \17344 );
or \U$17003 ( \17346 , \17334 , \17345 );
buf \U$17004 ( \17347 , \11342 );
not \U$17005 ( \17348 , \17347 );
xnor \U$17006 ( \17349 , \1308 , RI98730a8_180);
not \U$17007 ( \17350 , \17349 );
or \U$17008 ( \17351 , \17348 , \17350 );
nand \U$17009 ( \17352 , \17294 , \11350 );
nand \U$17010 ( \17353 , \17351 , \17352 );
nand \U$17011 ( \17354 , \17346 , \17353 );
nand \U$17012 ( \17355 , \17343 , \17332 );
nand \U$17013 ( \17356 , \17354 , \17355 );
not \U$17014 ( \17357 , \17356 );
not \U$17015 ( \17358 , \8819 );
not \U$17016 ( \17359 , \17228 );
or \U$17017 ( \17360 , \17358 , \17359 );
not \U$17018 ( \17361 , RI9872d60_173);
not \U$17019 ( \17362 , \1339 );
not \U$17020 ( \17363 , \17362 );
not \U$17021 ( \17364 , \17363 );
or \U$17022 ( \17365 , \17361 , \17364 );
or \U$17023 ( \17366 , \17363 , RI9872d60_173);
nand \U$17024 ( \17367 , \17365 , \17366 );
nand \U$17025 ( \17368 , \17367 , \8802 );
nand \U$17026 ( \17369 , \17360 , \17368 );
not \U$17027 ( \17370 , \17369 );
buf \U$17028 ( \17371 , \17251 );
not \U$17029 ( \17372 , \17371 );
not \U$17030 ( \17373 , \17260 );
or \U$17031 ( \17374 , \17372 , \17373 );
and \U$17032 ( \17375 , RI98733f0_187, \1691 );
not \U$17033 ( \17376 , RI98733f0_187);
and \U$17034 ( \17377 , \17376 , \1690 );
or \U$17035 ( \17378 , \17375 , \17377 );
nand \U$17036 ( \17379 , \17378 , \17263 );
nand \U$17037 ( \17380 , \17374 , \17379 );
buf \U$17038 ( \17381 , \17380 );
not \U$17039 ( \17382 , \17381 );
or \U$17040 ( \17383 , \17370 , \17382 );
not \U$17041 ( \17384 , \17380 );
not \U$17042 ( \17385 , \17369 );
nand \U$17043 ( \17386 , \17384 , \17385 );
not \U$17044 ( \17387 , \17234 );
not \U$17045 ( \17388 , RI9873210_183);
not \U$17046 ( \17389 , \6692 );
or \U$17047 ( \17390 , \17388 , \17389 );
or \U$17048 ( \17391 , \10145 , RI9873210_183);
nand \U$17049 ( \17392 , \17390 , \17391 );
not \U$17050 ( \17393 , \17392 );
or \U$17051 ( \17394 , \17387 , \17393 );
nand \U$17052 ( \17395 , \17240 , \17243 );
nand \U$17053 ( \17396 , \17394 , \17395 );
nand \U$17054 ( \17397 , \17386 , \17396 );
nand \U$17055 ( \17398 , \17383 , \17397 );
not \U$17056 ( \17399 , \17398 );
not \U$17057 ( \17400 , \4919 );
not \U$17058 ( \17401 , \17186 );
or \U$17059 ( \17402 , \17400 , \17401 );
xor \U$17060 ( \17403 , RI9872388_152, \9374 );
nand \U$17061 ( \17404 , \17403 , \5047 );
nand \U$17062 ( \17405 , \17402 , \17404 );
not \U$17063 ( \17406 , \5034 );
not \U$17064 ( \17407 , \17197 );
or \U$17065 ( \17408 , \17406 , \17407 );
and \U$17066 ( \17409 , \4470 , \5025 );
not \U$17067 ( \17410 , \4470 );
and \U$17068 ( \17411 , \17410 , RI9872478_154);
nor \U$17069 ( \17412 , \17409 , \17411 );
nand \U$17070 ( \17413 , \17412 , \5796 );
nand \U$17071 ( \17414 , \17408 , \17413 );
xor \U$17072 ( \17415 , \17405 , \17414 );
not \U$17073 ( \17416 , \10332 );
not \U$17074 ( \17417 , \9690 );
not \U$17075 ( \17418 , \6651 );
or \U$17076 ( \17419 , \17417 , \17418 );
or \U$17077 ( \17420 , \943 , \9690 );
nand \U$17078 ( \17421 , \17419 , \17420 );
not \U$17079 ( \17422 , \17421 );
or \U$17080 ( \17423 , \17416 , \17422 );
nand \U$17081 ( \17424 , \17211 , \9294 );
nand \U$17082 ( \17425 , \17423 , \17424 );
and \U$17083 ( \17426 , \17415 , \17425 );
and \U$17084 ( \17427 , \17405 , \17414 );
or \U$17085 ( \17428 , \17426 , \17427 );
not \U$17086 ( \17429 , \17428 );
not \U$17087 ( \17430 , \17429 );
and \U$17088 ( \17431 , \17399 , \17430 );
and \U$17089 ( \17432 , \17398 , \17429 );
nor \U$17090 ( \17433 , \17431 , \17432 );
not \U$17091 ( \17434 , \17433 );
or \U$17092 ( \17435 , \17357 , \17434 );
or \U$17093 ( \17436 , \17356 , \17433 );
nand \U$17094 ( \17437 , \17435 , \17436 );
not \U$17095 ( \17438 , \3163 );
not \U$17096 ( \17439 , \3154 );
not \U$17097 ( \17440 , \9569 );
not \U$17098 ( \17441 , \17440 );
not \U$17099 ( \17442 , \17441 );
or \U$17100 ( \17443 , \17439 , \17442 );
nand \U$17101 ( \17444 , \8924 , RI9872310_151);
nand \U$17102 ( \17445 , \17443 , \17444 );
not \U$17103 ( \17446 , \17445 );
or \U$17104 ( \17447 , \17438 , \17446 );
not \U$17105 ( \17448 , \3154 );
not \U$17106 ( \17449 , \10582 );
not \U$17107 ( \17450 , \17449 );
or \U$17108 ( \17451 , \17448 , \17450 );
nand \U$17109 ( \17452 , \8948 , RI9872310_151);
nand \U$17110 ( \17453 , \17451 , \17452 );
nand \U$17111 ( \17454 , \17453 , \12514 );
nand \U$17112 ( \17455 , \17447 , \17454 );
not \U$17113 ( \17456 , \3465 );
not \U$17114 ( \17457 , \17068 );
or \U$17115 ( \17458 , \17456 , \17457 );
not \U$17116 ( \17459 , RI98726d0_159);
not \U$17117 ( \17460 , \8904 );
or \U$17118 ( \17461 , \17459 , \17460 );
or \U$17119 ( \17462 , \13660 , RI98726d0_159);
nand \U$17120 ( \17463 , \17461 , \17462 );
nand \U$17121 ( \17464 , \17463 , \3467 );
nand \U$17122 ( \17465 , \17458 , \17464 );
xor \U$17123 ( \17466 , \17455 , \17465 );
not \U$17124 ( \17467 , \8790 );
not \U$17125 ( \17468 , \17104 );
or \U$17126 ( \17469 , \17467 , \17468 );
and \U$17127 ( \17470 , \5761 , RI98725e0_157);
and \U$17128 ( \17471 , \5762 , \4088 );
nor \U$17129 ( \17472 , \17470 , \17471 );
not \U$17130 ( \17473 , \17472 );
nand \U$17131 ( \17474 , \17473 , \5847 );
nand \U$17132 ( \17475 , \17469 , \17474 );
xor \U$17133 ( \17476 , \17466 , \17475 );
not \U$17134 ( \17477 , \6284 );
not \U$17135 ( \17478 , \16911 );
or \U$17136 ( \17479 , \17477 , \17478 );
not \U$17137 ( \17480 , \5632 );
not \U$17138 ( \17481 , \6718 );
or \U$17139 ( \17482 , \17480 , \17481 );
or \U$17140 ( \17483 , \6718 , \7049 );
nand \U$17141 ( \17484 , \17482 , \17483 );
nand \U$17142 ( \17485 , \17484 , \6286 );
nand \U$17143 ( \17486 , \17479 , \17485 );
not \U$17144 ( \17487 , \7326 );
not \U$17145 ( \17488 , \16885 );
or \U$17146 ( \17489 , \17487 , \17488 );
not \U$17147 ( \17490 , RI98729a0_165);
not \U$17148 ( \17491 , \3691 );
or \U$17149 ( \17492 , \17490 , \17491 );
or \U$17150 ( \17493 , \4287 , RI98729a0_165);
nand \U$17151 ( \17494 , \17492 , \17493 );
nand \U$17152 ( \17495 , \17494 , \7338 );
nand \U$17153 ( \17496 , \17489 , \17495 );
xor \U$17154 ( \17497 , \17486 , \17496 );
not \U$17155 ( \17498 , \11199 );
and \U$17156 ( \17499 , RI9872f40_177, \7691 );
not \U$17157 ( \17500 , RI9872f40_177);
and \U$17158 ( \17501 , \17500 , \820 );
nor \U$17159 ( \17502 , \17499 , \17501 );
not \U$17160 ( \17503 , \17502 );
or \U$17161 ( \17504 , \17498 , \17503 );
not \U$17162 ( \17505 , \16927 );
nand \U$17163 ( \17506 , \17505 , \8743 );
nand \U$17164 ( \17507 , \17504 , \17506 );
xor \U$17165 ( \17508 , \17497 , \17507 );
xor \U$17166 ( \17509 , \17476 , \17508 );
not \U$17167 ( \17510 , \8041 );
xnor \U$17168 ( \17511 , \7164 , RI9872a18_166);
not \U$17169 ( \17512 , \17511 );
or \U$17170 ( \17513 , \17510 , \17512 );
not \U$17171 ( \17514 , RI9872a18_166);
not \U$17172 ( \17515 , \2947 );
or \U$17173 ( \17516 , \17514 , \17515 );
or \U$17174 ( \17517 , \2947 , RI9872a18_166);
nand \U$17175 ( \17518 , \17516 , \17517 );
nand \U$17176 ( \17519 , \17518 , \8029 );
nand \U$17177 ( \17520 , \17513 , \17519 );
not \U$17178 ( \17521 , RI9873378_186);
not \U$17179 ( \17522 , RI98733f0_187);
not \U$17180 ( \17523 , \17522 );
or \U$17181 ( \17524 , \17521 , \17523 );
not \U$17182 ( \17525 , RI9873378_186);
nand \U$17183 ( \17526 , \17525 , RI98733f0_187);
nand \U$17184 ( \17527 , \17524 , \17526 );
buf \U$17185 ( \17528 , \17527 );
not \U$17186 ( \17529 , \17528 );
xor \U$17187 ( \17530 , \1106 , RI9873288_184);
not \U$17188 ( \17531 , \17530 );
or \U$17189 ( \17532 , \17529 , \17531 );
not \U$17190 ( \17533 , RI9873288_184);
not \U$17191 ( \17534 , \6692 );
or \U$17192 ( \17535 , \17533 , \17534 );
or \U$17193 ( \17536 , \6692 , RI9873288_184);
nand \U$17194 ( \17537 , \17535 , \17536 );
not \U$17195 ( \17538 , RI9873288_184);
not \U$17196 ( \17539 , RI98733f0_187);
nand \U$17197 ( \17540 , \17538 , \17539 );
nand \U$17198 ( \17541 , RI9873288_184, RI9873378_186);
and \U$17199 ( \17542 , \17540 , \17526 , \17541 );
buf \U$17200 ( \17543 , \17542 );
buf \U$17201 ( \17544 , \17543 );
buf \U$17202 ( \17545 , \17544 );
nand \U$17203 ( \17546 , \17537 , \17545 );
nand \U$17204 ( \17547 , \17532 , \17546 );
xor \U$17205 ( \17548 , \17520 , \17547 );
not \U$17206 ( \17549 , \9937 );
not \U$17207 ( \17550 , RI9873030_179);
not \U$17208 ( \17551 , \893 );
or \U$17209 ( \17552 , \17550 , \17551 );
or \U$17210 ( \17553 , \1506 , RI9873030_179);
nand \U$17211 ( \17554 , \17552 , \17553 );
not \U$17212 ( \17555 , \17554 );
or \U$17213 ( \17556 , \17549 , \17555 );
not \U$17214 ( \17557 , \14132 );
not \U$17215 ( \17558 , \8004 );
or \U$17216 ( \17559 , \17557 , \17558 );
not \U$17217 ( \17560 , RI9873030_179);
or \U$17218 ( \17561 , \8004 , \17560 );
nand \U$17219 ( \17562 , \17559 , \17561 );
nand \U$17220 ( \17563 , \17562 , \9952 );
nand \U$17221 ( \17564 , \17556 , \17563 );
and \U$17222 ( \17565 , \17548 , \17564 );
and \U$17223 ( \17566 , \17520 , \17547 );
or \U$17224 ( \17567 , \17565 , \17566 );
and \U$17225 ( \17568 , \17509 , \17567 );
and \U$17226 ( \17569 , \17476 , \17508 );
or \U$17227 ( \17570 , \17568 , \17569 );
xor \U$17228 ( \17571 , \17437 , \17570 );
not \U$17229 ( \17572 , \6144 );
not \U$17230 ( \17573 , RI98719b0_131);
not \U$17231 ( \17574 , \10392 );
or \U$17232 ( \17575 , \17573 , \17574 );
or \U$17233 ( \17576 , \8074 , RI98719b0_131);
nand \U$17234 ( \17577 , \17575 , \17576 );
not \U$17235 ( \17578 , \17577 );
or \U$17236 ( \17579 , \17572 , \17578 );
nand \U$17237 ( \17580 , \16948 , \793 );
nand \U$17238 ( \17581 , \17579 , \17580 );
not \U$17239 ( \17582 , \2087 );
not \U$17240 ( \17583 , \2076 );
not \U$17241 ( \17584 , \9569 );
or \U$17242 ( \17585 , \17583 , \17584 );
nand \U$17243 ( \17586 , \7466 , RI9871aa0_133);
nand \U$17244 ( \17587 , \17585 , \17586 );
not \U$17245 ( \17588 , \17587 );
or \U$17246 ( \17589 , \17582 , \17588 );
nand \U$17247 ( \17590 , \16971 , \2071 );
nand \U$17248 ( \17591 , \17589 , \17590 );
and \U$17249 ( \17592 , \17581 , \17591 );
not \U$17250 ( \17593 , \17581 );
not \U$17251 ( \17594 , \17591 );
and \U$17252 ( \17595 , \17593 , \17594 );
nor \U$17253 ( \17596 , \17592 , \17595 );
not \U$17254 ( \17597 , \1083 );
not \U$17255 ( \17598 , \16953 );
or \U$17256 ( \17599 , \17597 , \17598 );
not \U$17257 ( \17600 , RI98718c0_129);
not \U$17258 ( \17601 , \8607 );
or \U$17259 ( \17602 , \17600 , \17601 );
or \U$17260 ( \17603 , \10309 , RI98718c0_129);
nand \U$17261 ( \17604 , \17602 , \17603 );
nand \U$17262 ( \17605 , \1136 , \17604 );
nand \U$17263 ( \17606 , \17599 , \17605 );
xor \U$17264 ( \17607 , \17596 , \17606 );
not \U$17265 ( \17608 , \1323 );
and \U$17266 ( \17609 , RI9871b18_134, \8555 );
not \U$17267 ( \17610 , RI9871b18_134);
and \U$17268 ( \17611 , \17610 , \10372 );
or \U$17269 ( \17612 , \17609 , \17611 );
not \U$17270 ( \17613 , \17612 );
or \U$17271 ( \17614 , \17608 , \17613 );
nand \U$17272 ( \17615 , \17027 , \12720 );
nand \U$17273 ( \17616 , \17614 , \17615 );
not \U$17274 ( \17617 , \17371 );
not \U$17275 ( \17618 , \17378 );
or \U$17276 ( \17619 , \17617 , \17618 );
not \U$17277 ( \17620 , \17263 );
not \U$17278 ( \17621 , \17620 );
nand \U$17279 ( \17622 , \17621 , RI98733f0_187);
nand \U$17280 ( \17623 , \17619 , \17622 );
xor \U$17281 ( \17624 , \17616 , \17623 );
not \U$17282 ( \17625 , \1430 );
not \U$17283 ( \17626 , RI9871c08_136);
not \U$17284 ( \17627 , \8650 );
or \U$17285 ( \17628 , \17626 , \17627 );
or \U$17286 ( \17629 , \11406 , RI9871c08_136);
nand \U$17287 ( \17630 , \17628 , \17629 );
not \U$17288 ( \17631 , \17630 );
or \U$17289 ( \17632 , \17625 , \17631 );
nand \U$17290 ( \17633 , \17049 , \1455 );
nand \U$17291 ( \17634 , \17632 , \17633 );
xor \U$17292 ( \17635 , \17624 , \17634 );
xor \U$17293 ( \17636 , \17607 , \17635 );
not \U$17294 ( \17637 , \9952 );
not \U$17295 ( \17638 , \17554 );
or \U$17296 ( \17639 , \17637 , \17638 );
not \U$17297 ( \17640 , RI9873030_179);
not \U$17298 ( \17641 , \916 );
or \U$17299 ( \17642 , \17640 , \17641 );
or \U$17300 ( \17643 , \916 , RI9873030_179);
nand \U$17301 ( \17644 , \17642 , \17643 );
nand \U$17302 ( \17645 , \17644 , \9937 );
nand \U$17303 ( \17646 , \17639 , \17645 );
not \U$17304 ( \17647 , \17646 );
not \U$17305 ( \17648 , \17545 );
not \U$17306 ( \17649 , \17530 );
or \U$17307 ( \17650 , \17648 , \17649 );
not \U$17308 ( \17651 , RI9873288_184);
not \U$17309 ( \17652 , \9276 );
or \U$17310 ( \17653 , \17651 , \17652 );
or \U$17311 ( \17654 , \1127 , RI9873288_184);
nand \U$17312 ( \17655 , \17653 , \17654 );
nand \U$17313 ( \17656 , \17655 , \17528 );
nand \U$17314 ( \17657 , \17650 , \17656 );
not \U$17315 ( \17658 , \17657 );
or \U$17316 ( \17659 , \17647 , \17658 );
and \U$17317 ( \17660 , \17511 , \9079 );
and \U$17318 ( \17661 , RI9872a18_166, \1485 );
not \U$17319 ( \17662 , RI9872a18_166);
and \U$17320 ( \17663 , \17662 , \1486 );
or \U$17321 ( \17664 , \17661 , \17663 );
and \U$17322 ( \17665 , \17664 , \9072 );
nor \U$17323 ( \17666 , \17660 , \17665 );
not \U$17324 ( \17667 , \17666 );
not \U$17325 ( \17668 , \17657 );
not \U$17326 ( \17669 , \17668 );
not \U$17327 ( \17670 , \17646 );
or \U$17328 ( \17671 , \17669 , \17670 );
or \U$17329 ( \17672 , \17646 , \17668 );
nand \U$17330 ( \17673 , \17671 , \17672 );
nand \U$17331 ( \17674 , \17667 , \17673 );
nand \U$17332 ( \17675 , \17659 , \17674 );
xor \U$17333 ( \17676 , \17636 , \17675 );
xor \U$17334 ( \17677 , \17571 , \17676 );
xor \U$17335 ( \17678 , \17322 , \17677 );
xor \U$17336 ( \17679 , \17476 , \17508 );
xor \U$17337 ( \17680 , \17679 , \17567 );
not \U$17338 ( \17681 , \17680 );
not \U$17339 ( \17682 , \1154 );
not \U$17340 ( \17683 , \17682 );
not \U$17341 ( \17684 , \497 );
not \U$17342 ( \17685 , \17684 );
buf \U$17343 ( \17686 , \504 );
not \U$17344 ( \17687 , \17686 );
or \U$17345 ( \17688 , \17685 , \17687 );
buf \U$17346 ( \17689 , \511 );
not \U$17347 ( \17690 , \17689 );
nand \U$17348 ( \17691 , \17688 , \17690 );
not \U$17349 ( \17692 , \17691 );
and \U$17350 ( \17693 , RI9870240_81, \508 );
not \U$17351 ( \17694 , RI9870240_81);
and \U$17352 ( \17695 , \17694 , RI98702b8_82);
nor \U$17353 ( \17696 , \17693 , \17695 );
not \U$17354 ( \17697 , \17696 );
and \U$17355 ( \17698 , \17692 , \17697 );
and \U$17356 ( \17699 , \17691 , \17696 );
nor \U$17357 ( \17700 , \17698 , \17699 );
not \U$17358 ( \17701 , \17700 );
buf \U$17359 ( \17702 , \17701 );
buf \U$17360 ( \17703 , \17702 );
not \U$17361 ( \17704 , \17703 );
nor \U$17362 ( \17705 , \17683 , \17704 );
not \U$17363 ( \17706 , \16995 );
not \U$17364 ( \17707 , \12780 );
or \U$17365 ( \17708 , \17706 , \17707 );
nand \U$17366 ( \17709 , \8678 , \16996 );
nand \U$17367 ( \17710 , \17708 , \17709 );
not \U$17368 ( \17711 , \17710 );
not \U$17369 ( \17712 , \1161 );
or \U$17370 ( \17713 , \17711 , \17712 );
not \U$17371 ( \17714 , \16987 );
not \U$17372 ( \17715 , \515 );
or \U$17373 ( \17716 , \17714 , \17715 );
nand \U$17374 ( \17717 , \17716 , \16988 );
xor \U$17375 ( \17718 , RI9870600_89, RI9870678_90);
and \U$17376 ( \17719 , \17717 , \17718 );
not \U$17377 ( \17720 , \17717 );
not \U$17378 ( \17721 , \17718 );
and \U$17379 ( \17722 , \17720 , \17721 );
nor \U$17380 ( \17723 , \17719 , \17722 );
not \U$17381 ( \17724 , \17723 );
not \U$17382 ( \17725 , \17724 );
not \U$17383 ( \17726 , \17725 );
not \U$17384 ( \17727 , \17726 );
xor \U$17385 ( \17728 , \17682 , \17727 );
nand \U$17386 ( \17729 , \6315 , \17728 );
nand \U$17387 ( \17730 , \17713 , \17729 );
xor \U$17388 ( \17731 , \17705 , \17730 );
not \U$17389 ( \17732 , \1013 );
not \U$17390 ( \17733 , \17009 );
or \U$17391 ( \17734 , \17732 , \17733 );
not \U$17392 ( \17735 , \13921 );
nand \U$17393 ( \17736 , \530 , \13924 );
not \U$17394 ( \17737 , \17736 );
and \U$17395 ( \17738 , \17735 , \17737 );
and \U$17396 ( \17739 , \13921 , \17736 );
nor \U$17397 ( \17740 , \17738 , \17739 );
buf \U$17398 ( \17741 , \17740 );
and \U$17399 ( \17742 , \1042 , \17741 );
not \U$17400 ( \17743 , \1042 );
not \U$17401 ( \17744 , \17741 );
and \U$17402 ( \17745 , \17743 , \17744 );
or \U$17403 ( \17746 , \17742 , \17745 );
nand \U$17404 ( \17747 , \1016 , \17746 );
nand \U$17405 ( \17748 , \17734 , \17747 );
and \U$17406 ( \17749 , \17731 , \17748 );
not \U$17407 ( \17750 , \17731 );
not \U$17408 ( \17751 , \17748 );
and \U$17409 ( \17752 , \17750 , \17751 );
nor \U$17410 ( \17753 , \17749 , \17752 );
not \U$17411 ( \17754 , \17753 );
not \U$17412 ( \17755 , \1518 );
not \U$17413 ( \17756 , \9137 );
buf \U$17414 ( \17757 , \17756 );
not \U$17415 ( \17758 , \17757 );
not \U$17416 ( \17759 , \17758 );
not \U$17417 ( \17760 , RI9871c80_137);
and \U$17418 ( \17761 , \17759 , \17760 );
and \U$17419 ( \17762 , \13070 , RI9871c80_137);
nor \U$17420 ( \17763 , \17761 , \17762 );
not \U$17421 ( \17764 , \17763 );
or \U$17422 ( \17765 , \17755 , \17764 );
not \U$17423 ( \17766 , RI9871c80_137);
not \U$17424 ( \17767 , \11358 );
not \U$17425 ( \17768 , \17767 );
or \U$17426 ( \17769 , \17766 , \17768 );
not \U$17427 ( \17770 , \10064 );
nand \U$17428 ( \17771 , \17770 , \1800 );
nand \U$17429 ( \17772 , \17769 , \17771 );
nand \U$17430 ( \17773 , \17772 , \1501 );
nand \U$17431 ( \17774 , \17765 , \17773 );
not \U$17432 ( \17775 , \832 );
not \U$17433 ( \17776 , \17094 );
or \U$17434 ( \17777 , \17775 , \17776 );
not \U$17435 ( \17778 , \13615 );
not \U$17436 ( \17779 , \13618 );
and \U$17437 ( \17780 , \17778 , \17779 );
and \U$17438 ( \17781 , \13615 , \13618 );
nor \U$17439 ( \17782 , \17780 , \17781 );
buf \U$17440 ( \17783 , \17782 );
and \U$17441 ( \17784 , \17783 , \2243 );
not \U$17442 ( \17785 , \17783 );
and \U$17443 ( \17786 , \17785 , RI9871d70_139);
nor \U$17444 ( \17787 , \17784 , \17786 );
nand \U$17445 ( \17788 , \17787 , \859 );
nand \U$17446 ( \17789 , \17777 , \17788 );
and \U$17447 ( \17790 , \17774 , \17789 );
not \U$17448 ( \17791 , \17790 );
or \U$17449 ( \17792 , \17754 , \17791 );
or \U$17450 ( \17793 , \17790 , \17753 );
nand \U$17451 ( \17794 , \17792 , \17793 );
not \U$17452 ( \17795 , \17794 );
not \U$17453 ( \17796 , \17795 );
not \U$17454 ( \17797 , \5653 );
not \U$17455 ( \17798 , \5648 );
not \U$17456 ( \17799 , \4410 );
not \U$17457 ( \17800 , \17799 );
or \U$17458 ( \17801 , \17798 , \17800 );
nand \U$17459 ( \17802 , \5206 , RI9872568_156);
nand \U$17460 ( \17803 , \17801 , \17802 );
not \U$17461 ( \17804 , \17803 );
or \U$17462 ( \17805 , \17797 , \17804 );
and \U$17463 ( \17806 , RI9872568_156, \5623 );
not \U$17464 ( \17807 , RI9872568_156);
and \U$17465 ( \17808 , \17807 , \4470 );
nor \U$17466 ( \17809 , \17806 , \17808 );
nand \U$17467 ( \17810 , \17809 , \9320 );
nand \U$17468 ( \17811 , \17805 , \17810 );
not \U$17469 ( \17812 , \17811 );
or \U$17470 ( \17813 , \17796 , \17812 );
or \U$17471 ( \17814 , \17811 , \17795 );
nand \U$17472 ( \17815 , \17813 , \17814 );
not \U$17473 ( \17816 , \17288 );
not \U$17474 ( \17817 , \17816 );
not \U$17475 ( \17818 , \17314 );
or \U$17476 ( \17819 , \17817 , \17818 );
or \U$17477 ( \17820 , \17314 , \17816 );
nand \U$17478 ( \17821 , \17819 , \17820 );
xor \U$17479 ( \17822 , \17815 , \17821 );
xor \U$17480 ( \17823 , \17520 , \17547 );
xor \U$17481 ( \17824 , \17823 , \17564 );
and \U$17482 ( \17825 , \17822 , \17824 );
and \U$17483 ( \17826 , \17815 , \17821 );
or \U$17484 ( \17827 , \17825 , \17826 );
not \U$17485 ( \17828 , \17827 );
xor \U$17486 ( \17829 , \17191 , \17205 );
xor \U$17487 ( \17830 , \17829 , \17220 );
not \U$17488 ( \17831 , \17830 );
not \U$17489 ( \17832 , \6286 );
not \U$17490 ( \17833 , \16903 );
or \U$17491 ( \17834 , \17832 , \17833 );
not \U$17492 ( \17835 , \7049 );
not \U$17493 ( \17836 , \5208 );
or \U$17494 ( \17837 , \17835 , \17836 );
nand \U$17495 ( \17838 , \13057 , RI98728b0_163);
nand \U$17496 ( \17839 , \17837 , \17838 );
nand \U$17497 ( \17840 , \17839 , \6284 );
nand \U$17498 ( \17841 , \17834 , \17840 );
not \U$17499 ( \17842 , \17841 );
not \U$17500 ( \17843 , \1380 );
not \U$17501 ( \17844 , RI9871e60_141);
and \U$17502 ( \17845 , \13934 , \17844 );
not \U$17503 ( \17846 , \13934 );
and \U$17504 ( \17847 , \17846 , RI9871e60_141);
nor \U$17505 ( \17848 , \17845 , \17847 );
not \U$17506 ( \17849 , \17848 );
or \U$17507 ( \17850 , \17843 , \17849 );
xnor \U$17508 ( \17851 , RI9871e60_141, \13860 );
nand \U$17509 ( \17852 , \17851 , \1352 );
nand \U$17510 ( \17853 , \17850 , \17852 );
not \U$17511 ( \17854 , \17686 );
not \U$17512 ( \17855 , \17689 );
nand \U$17513 ( \17856 , \17855 , \17684 );
and \U$17514 ( \17857 , \17854 , \17856 );
not \U$17515 ( \17858 , \17854 );
not \U$17516 ( \17859 , \17856 );
and \U$17517 ( \17860 , \17858 , \17859 );
nor \U$17518 ( \17861 , \17857 , \17860 );
buf \U$17519 ( \17862 , \17861 );
buf \U$17520 ( \17863 , \17862 );
and \U$17521 ( \17864 , \17682 , \17863 );
not \U$17522 ( \17865 , \1013 );
not \U$17523 ( \17866 , \17746 );
or \U$17524 ( \17867 , \17865 , \17866 );
buf \U$17525 ( \17868 , \17724 );
not \U$17526 ( \17869 , \17868 );
and \U$17527 ( \17870 , \17869 , \1042 );
not \U$17528 ( \17871 , \17869 );
and \U$17529 ( \17872 , \17871 , \12592 );
nor \U$17530 ( \17873 , \17870 , \17872 );
nand \U$17531 ( \17874 , \17873 , \1016 );
nand \U$17532 ( \17875 , \17867 , \17874 );
xor \U$17533 ( \17876 , \17864 , \17875 );
xor \U$17534 ( \17877 , \17853 , \17876 );
not \U$17535 ( \17878 , \832 );
not \U$17536 ( \17879 , \17787 );
or \U$17537 ( \17880 , \17878 , \17879 );
and \U$17538 ( \17881 , RI9871d70_139, \13860 );
not \U$17539 ( \17882 , RI9871d70_139);
not \U$17540 ( \17883 , \17013 );
and \U$17541 ( \17884 , \17882 , \17883 );
or \U$17542 ( \17885 , \17881 , \17884 );
nand \U$17543 ( \17886 , \17885 , \859 );
nand \U$17544 ( \17887 , \17880 , \17886 );
not \U$17545 ( \17888 , \17887 );
not \U$17546 ( \17889 , \1292 );
and \U$17547 ( \17890 , RI9871b18_134, \13065 );
not \U$17548 ( \17891 , RI9871b18_134);
and \U$17549 ( \17892 , \17891 , \17757 );
nor \U$17550 ( \17893 , \17890 , \17892 );
not \U$17551 ( \17894 , \17893 );
or \U$17552 ( \17895 , \17889 , \17894 );
not \U$17553 ( \17896 , \1283 );
not \U$17554 ( \17897 , \9113 );
not \U$17555 ( \17898 , \17897 );
or \U$17556 ( \17899 , \17896 , \17898 );
or \U$17557 ( \17900 , \9119 , \1283 );
nand \U$17558 ( \17901 , \17899 , \17900 );
nand \U$17559 ( \17902 , \17901 , \1323 );
nand \U$17560 ( \17903 , \17895 , \17902 );
not \U$17561 ( \17904 , \17903 );
not \U$17562 ( \17905 , \1352 );
not \U$17563 ( \17906 , \17848 );
or \U$17564 ( \17907 , \17905 , \17906 );
buf \U$17565 ( \17908 , \17740 );
and \U$17566 ( \17909 , RI9871e60_141, \17908 );
not \U$17567 ( \17910 , RI9871e60_141);
buf \U$17568 ( \17911 , \17740 );
not \U$17569 ( \17912 , \17911 );
and \U$17570 ( \17913 , \17910 , \17912 );
or \U$17571 ( \17914 , \17909 , \17913 );
nand \U$17572 ( \17915 , \17914 , \1379 );
nand \U$17573 ( \17916 , \17907 , \17915 );
not \U$17574 ( \17917 , \17916 );
nand \U$17575 ( \17918 , \17904 , \17917 );
not \U$17576 ( \17919 , \17918 );
or \U$17577 ( \17920 , \17888 , \17919 );
nand \U$17578 ( \17921 , \17903 , \17916 );
nand \U$17579 ( \17922 , \17920 , \17921 );
xor \U$17580 ( \17923 , \17877 , \17922 );
not \U$17581 ( \17924 , \17923 );
or \U$17582 ( \17925 , \17842 , \17924 );
nand \U$17583 ( \17926 , \17922 , \17877 );
nand \U$17584 ( \17927 , \17925 , \17926 );
xor \U$17585 ( \17928 , \17232 , \17265 );
xor \U$17586 ( \17929 , \17928 , \17245 );
xor \U$17587 ( \17930 , \17927 , \17929 );
not \U$17588 ( \17931 , \17930 );
or \U$17589 ( \17932 , \17831 , \17931 );
nand \U$17590 ( \17933 , \17929 , \17927 );
nand \U$17591 ( \17934 , \17932 , \17933 );
not \U$17592 ( \17935 , \17934 );
not \U$17593 ( \17936 , \17935 );
or \U$17594 ( \17937 , \17828 , \17936 );
or \U$17595 ( \17938 , \17827 , \17935 );
nand \U$17596 ( \17939 , \17937 , \17938 );
not \U$17597 ( \17940 , \17939 );
or \U$17598 ( \17941 , \17681 , \17940 );
nand \U$17599 ( \17942 , \17827 , \17934 );
nand \U$17600 ( \17943 , \17941 , \17942 );
not \U$17601 ( \17944 , \17943 );
xnor \U$17602 ( \17945 , \17678 , \17944 );
not \U$17603 ( \17946 , \11199 );
not \U$17604 ( \17947 , \1253 );
not \U$17605 ( \17948 , RI9872f40_177);
and \U$17606 ( \17949 , \17947 , \17948 );
and \U$17607 ( \17950 , \5720 , RI9872f40_177);
nor \U$17608 ( \17951 , \17949 , \17950 );
not \U$17609 ( \17952 , \17951 );
not \U$17610 ( \17953 , \17952 );
or \U$17611 ( \17954 , \17946 , \17953 );
not \U$17612 ( \17955 , RI9872f40_177);
not \U$17613 ( \17956 , \1339 );
or \U$17614 ( \17957 , \17955 , \17956 );
or \U$17615 ( \17958 , \17363 , RI9872f40_177);
nand \U$17616 ( \17959 , \17957 , \17958 );
nand \U$17617 ( \17960 , \17959 , \8743 );
nand \U$17618 ( \17961 , \17954 , \17960 );
not \U$17619 ( \17962 , \17961 );
not \U$17620 ( \17963 , \5036 );
not \U$17621 ( \17964 , RI9872478_154);
not \U$17622 ( \17965 , \5776 );
or \U$17623 ( \17966 , \17964 , \17965 );
or \U$17624 ( \17967 , \5776 , RI9872478_154);
nand \U$17625 ( \17968 , \17966 , \17967 );
not \U$17626 ( \17969 , \17968 );
or \U$17627 ( \17970 , \17963 , \17969 );
and \U$17628 ( \17971 , \5762 , RI9872478_154);
not \U$17629 ( \17972 , \5762 );
and \U$17630 ( \17973 , \17972 , \5025 );
nor \U$17631 ( \17974 , \17971 , \17973 );
nand \U$17632 ( \17975 , \17974 , \5034 );
nand \U$17633 ( \17976 , \17970 , \17975 );
not \U$17634 ( \17977 , \7188 );
not \U$17635 ( \17978 , \5648 );
not \U$17636 ( \17979 , \10639 );
or \U$17637 ( \17980 , \17978 , \17979 );
nand \U$17638 ( \17981 , \7007 , RI9872568_156);
nand \U$17639 ( \17982 , \17980 , \17981 );
not \U$17640 ( \17983 , \17982 );
or \U$17641 ( \17984 , \17977 , \17983 );
not \U$17642 ( \17985 , \5648 );
not \U$17643 ( \17986 , \9374 );
or \U$17644 ( \17987 , \17985 , \17986 );
nand \U$17645 ( \17988 , \4986 , RI9872568_156);
nand \U$17646 ( \17989 , \17987 , \17988 );
nand \U$17647 ( \17990 , \17989 , \9320 );
nand \U$17648 ( \17991 , \17984 , \17990 );
xor \U$17649 ( \17992 , \17976 , \17991 );
not \U$17650 ( \17993 , \17992 );
or \U$17651 ( \17994 , \17962 , \17993 );
nand \U$17652 ( \17995 , \17991 , \17976 );
nand \U$17653 ( \17996 , \17994 , \17995 );
not \U$17654 ( \17997 , \10487 );
not \U$17655 ( \17998 , \17161 );
or \U$17656 ( \17999 , \17997 , \17998 );
and \U$17657 ( \18000 , \1478 , \1480 );
not \U$17658 ( \18001 , \1478 );
not \U$17659 ( \18002 , \1480 );
and \U$17660 ( \18003 , \18001 , \18002 );
nor \U$17661 ( \18004 , \18000 , \18003 );
xnor \U$17662 ( \18005 , RI9872bf8_170, \18004 );
nand \U$17663 ( \18006 , \18005 , \9670 );
nand \U$17664 ( \18007 , \17999 , \18006 );
not \U$17665 ( \18008 , \18007 );
not \U$17666 ( \18009 , \13484 );
not \U$17667 ( \18010 , \17135 );
or \U$17668 ( \18011 , \18009 , \18010 );
not \U$17669 ( \18012 , RI9873210_183);
and \U$17670 ( \18013 , \18012 , \915 );
not \U$17671 ( \18014 , \18012 );
and \U$17672 ( \18015 , \18014 , \5479 );
nor \U$17673 ( \18016 , \18013 , \18015 );
nand \U$17674 ( \18017 , \18016 , \13476 );
nand \U$17675 ( \18018 , \18011 , \18017 );
not \U$17676 ( \18019 , \18018 );
not \U$17677 ( \18020 , \18019 );
not \U$17678 ( \18021 , \8802 );
not \U$17679 ( \18022 , \17145 );
or \U$17680 ( \18023 , \18021 , \18022 );
not \U$17681 ( \18024 , \8807 );
not \U$17682 ( \18025 , \3126 );
or \U$17683 ( \18026 , \18024 , \18025 );
nand \U$17684 ( \18027 , \12393 , RI9872d60_173);
nand \U$17685 ( \18028 , \18026 , \18027 );
nand \U$17686 ( \18029 , \18028 , \9312 );
nand \U$17687 ( \18030 , \18023 , \18029 );
not \U$17688 ( \18031 , \18030 );
or \U$17689 ( \18032 , \18020 , \18031 );
or \U$17690 ( \18033 , \18030 , \18019 );
nand \U$17691 ( \18034 , \18032 , \18033 );
not \U$17692 ( \18035 , \18034 );
or \U$17693 ( \18036 , \18008 , \18035 );
nand \U$17694 ( \18037 , \18030 , \18018 );
nand \U$17695 ( \18038 , \18036 , \18037 );
xor \U$17696 ( \18039 , \17996 , \18038 );
not \U$17697 ( \18040 , \17347 );
and \U$17698 ( \18041 , RI98730a8_180, \1505 );
not \U$17699 ( \18042 , RI98730a8_180);
and \U$17700 ( \18043 , \18042 , \13169 );
or \U$17701 ( \18044 , \18041 , \18043 );
not \U$17702 ( \18045 , \18044 );
or \U$17703 ( \18046 , \18040 , \18045 );
not \U$17704 ( \18047 , \13022 );
not \U$17705 ( \18048 , \8004 );
or \U$17706 ( \18049 , \18047 , \18048 );
or \U$17707 ( \18050 , \8004 , \13022 );
nand \U$17708 ( \18051 , \18049 , \18050 );
nand \U$17709 ( \18052 , \18051 , \13020 );
nand \U$17710 ( \18053 , \18046 , \18052 );
not \U$17711 ( \18054 , \10679 );
not \U$17712 ( \18055 , RI9872b80_169);
not \U$17713 ( \18056 , \2947 );
or \U$17714 ( \18057 , \18055 , \18056 );
or \U$17715 ( \18058 , \2947 , RI9872b80_169);
nand \U$17716 ( \18059 , \18057 , \18058 );
not \U$17717 ( \18060 , \18059 );
or \U$17718 ( \18061 , \18054 , \18060 );
and \U$17719 ( \18062 , RI9872b80_169, \9162 );
not \U$17720 ( \18063 , RI9872b80_169);
and \U$17721 ( \18064 , \18063 , \2110 );
nor \U$17722 ( \18065 , \18062 , \18064 );
not \U$17723 ( \18066 , \18065 );
nand \U$17724 ( \18067 , \18066 , \9214 );
nand \U$17725 ( \18068 , \18061 , \18067 );
nand \U$17726 ( \18069 , \18053 , \18068 );
xnor \U$17727 ( \18070 , \1096 , RI98733f0_187);
not \U$17728 ( \18071 , \18070 );
nor \U$17729 ( \18072 , \18071 , \17620 );
not \U$17730 ( \18073 , RI98733f0_187);
not \U$17731 ( \18074 , \6174 );
or \U$17732 ( \18075 , \18073 , \18074 );
or \U$17733 ( \18076 , \1416 , RI98733f0_187);
nand \U$17734 ( \18077 , \18075 , \18076 );
not \U$17735 ( \18078 , \18077 );
not \U$17736 ( \18079 , \17371 );
nor \U$17737 ( \18080 , \18078 , \18079 );
nor \U$17738 ( \18081 , \18072 , \18080 );
and \U$17739 ( \18082 , \18069 , \18081 );
nor \U$17740 ( \18083 , \18053 , \18068 );
nor \U$17741 ( \18084 , \18082 , \18083 );
and \U$17742 ( \18085 , \18039 , \18084 );
and \U$17743 ( \18086 , \17996 , \18038 );
or \U$17744 ( \18087 , \18085 , \18086 );
not \U$17745 ( \18088 , \18087 );
not \U$17746 ( \18089 , \3170 );
and \U$17747 ( \18090 , RI9872310_151, \8333 );
not \U$17748 ( \18091 , RI9872310_151);
and \U$17749 ( \18092 , \18091 , \8916 );
or \U$17750 ( \18093 , \18090 , \18092 );
not \U$17751 ( \18094 , \18093 );
or \U$17752 ( \18095 , \18089 , \18094 );
not \U$17753 ( \18096 , \3154 );
not \U$17754 ( \18097 , \13358 );
or \U$17755 ( \18098 , \18096 , \18097 );
nand \U$17756 ( \18099 , \8074 , RI9872310_151);
nand \U$17757 ( \18100 , \18098 , \18099 );
nand \U$17758 ( \18101 , \18100 , \6653 );
nand \U$17759 ( \18102 , \18095 , \18101 );
not \U$17760 ( \18103 , \18102 );
not \U$17761 ( \18104 , \18103 );
not \U$17762 ( \18105 , \2071 );
not \U$17763 ( \18106 , RI9871aa0_133);
not \U$17764 ( \18107 , \8606 );
not \U$17765 ( \18108 , \18107 );
or \U$17766 ( \18109 , \18106 , \18108 );
not \U$17767 ( \18110 , \8605 );
buf \U$17768 ( \18111 , \18110 );
or \U$17769 ( \18112 , \18111 , RI9871aa0_133);
nand \U$17770 ( \18113 , \18109 , \18112 );
not \U$17771 ( \18114 , \18113 );
or \U$17772 ( \18115 , \18105 , \18114 );
not \U$17773 ( \18116 , RI9871aa0_133);
not \U$17774 ( \18117 , \8878 );
or \U$17775 ( \18118 , \18116 , \18117 );
or \U$17776 ( \18119 , \12712 , RI9871aa0_133);
nand \U$17777 ( \18120 , \18118 , \18119 );
nand \U$17778 ( \18121 , \18120 , \2087 );
nand \U$17779 ( \18122 , \18115 , \18121 );
not \U$17780 ( \18123 , \18122 );
not \U$17781 ( \18124 , \18123 );
or \U$17782 ( \18125 , \18104 , \18124 );
not \U$17783 ( \18126 , \3465 );
not \U$17784 ( \18127 , RI98726d0_159);
not \U$17785 ( \18128 , \9569 );
not \U$17786 ( \18129 , \18128 );
or \U$17787 ( \18130 , \18127 , \18129 );
or \U$17788 ( \18131 , \7466 , RI98726d0_159);
nand \U$17789 ( \18132 , \18130 , \18131 );
not \U$17790 ( \18133 , \18132 );
or \U$17791 ( \18134 , \18126 , \18133 );
nand \U$17792 ( \18135 , \17076 , \3467 );
nand \U$17793 ( \18136 , \18134 , \18135 );
nand \U$17794 ( \18137 , \18125 , \18136 );
nand \U$17795 ( \18138 , \18102 , \18122 );
nand \U$17796 ( \18139 , \18137 , \18138 );
not \U$17797 ( \18140 , \18139 );
not \U$17798 ( \18141 , \18140 );
not \U$17799 ( \18142 , \875 );
not \U$17800 ( \18143 , RI9872130_147);
not \U$17801 ( \18144 , \13268 );
or \U$17802 ( \18145 , \18143 , \18144 );
or \U$17803 ( \18146 , \13268 , RI9872130_147);
nand \U$17804 ( \18147 , \18145 , \18146 );
not \U$17805 ( \18148 , \18147 );
or \U$17806 ( \18149 , \18142 , \18148 );
not \U$17807 ( \18150 , \919 );
buf \U$17808 ( \18151 , \11453 );
not \U$17809 ( \18152 , \18151 );
not \U$17810 ( \18153 , \18152 );
or \U$17811 ( \18154 , \18150 , \18153 );
not \U$17812 ( \18155 , \12783 );
nand \U$17813 ( \18156 , \18155 , RI9872130_147);
nand \U$17814 ( \18157 , \18154 , \18156 );
nand \U$17815 ( \18158 , \18157 , \924 );
nand \U$17816 ( \18159 , \18149 , \18158 );
not \U$17817 ( \18160 , \1292 );
not \U$17818 ( \18161 , \17901 );
or \U$17819 ( \18162 , \18160 , \18161 );
and \U$17820 ( \18163 , \12460 , \4044 );
not \U$17821 ( \18164 , \12460 );
and \U$17822 ( \18165 , \18164 , RI9871b18_134);
nor \U$17823 ( \18166 , \18163 , \18165 );
nand \U$17824 ( \18167 , \18166 , \1323 );
nand \U$17825 ( \18168 , \18162 , \18167 );
xor \U$17826 ( \18169 , \18159 , \18168 );
not \U$17827 ( \18170 , \18169 );
buf \U$17828 ( \18171 , \4101 );
not \U$17829 ( \18172 , \18171 );
not \U$17830 ( \18173 , \4088 );
not \U$17831 ( \18174 , \7905 );
or \U$17832 ( \18175 , \18173 , \18174 );
nand \U$17833 ( \18176 , \6529 , RI98725e0_157);
nand \U$17834 ( \18177 , \18175 , \18176 );
not \U$17835 ( \18178 , \18177 );
or \U$17836 ( \18179 , \18172 , \18178 );
nand \U$17837 ( \18180 , \17111 , \5847 );
nand \U$17838 ( \18181 , \18179 , \18180 );
not \U$17839 ( \18182 , \18181 );
or \U$17840 ( \18183 , \18170 , \18182 );
nand \U$17841 ( \18184 , \18159 , \18168 );
nand \U$17842 ( \18185 , \18183 , \18184 );
xor \U$17843 ( \18186 , RI9870510_87, RI9870588_88);
buf \U$17844 ( \18187 , \500 );
and \U$17845 ( \18188 , \18186 , \18187 );
not \U$17846 ( \18189 , \18186 );
not \U$17847 ( \18190 , \18187 );
and \U$17848 ( \18191 , \18189 , \18190 );
nor \U$17849 ( \18192 , \18188 , \18191 );
buf \U$17850 ( \18193 , \18192 );
buf \U$17851 ( \18194 , \18193 );
not \U$17852 ( \18195 , \18194 );
nand \U$17853 ( \18196 , \12781 , \18195 );
not \U$17854 ( \18197 , \17863 );
not \U$17855 ( \18198 , \1154 );
or \U$17856 ( \18199 , \18197 , \18198 );
or \U$17857 ( \18200 , \12780 , \17863 );
nand \U$17858 ( \18201 , \18199 , \18200 );
not \U$17859 ( \18202 , \18201 );
not \U$17860 ( \18203 , \1160 );
or \U$17861 ( \18204 , \18202 , \18203 );
not \U$17862 ( \18205 , \1218 );
not \U$17863 ( \18206 , \17702 );
not \U$17864 ( \18207 , \1154 );
or \U$17865 ( \18208 , \18206 , \18207 );
not \U$17866 ( \18209 , \17702 );
not \U$17867 ( \18210 , \18209 );
or \U$17868 ( \18211 , \1154 , \18210 );
nand \U$17869 ( \18212 , \18208 , \18211 );
nand \U$17870 ( \18213 , \18205 , \18212 );
nand \U$17871 ( \18214 , \18204 , \18213 );
xnor \U$17872 ( \18215 , \18196 , \18214 );
not \U$17873 ( \18216 , \16995 );
not \U$17874 ( \18217 , \18216 );
not \U$17875 ( \18218 , \1157 );
not \U$17876 ( \18219 , \18218 );
not \U$17877 ( \18220 , \18219 );
or \U$17878 ( \18221 , \18217 , \18220 );
or \U$17879 ( \18222 , \18219 , \18216 );
nand \U$17880 ( \18223 , \18221 , \18222 );
not \U$17881 ( \18224 , \18223 );
not \U$17882 ( \18225 , \1016 );
or \U$17883 ( \18226 , \18224 , \18225 );
nand \U$17884 ( \18227 , \17873 , \1013 );
nand \U$17885 ( \18228 , \18226 , \18227 );
nand \U$17886 ( \18229 , \18215 , \18228 );
buf \U$17887 ( \18230 , \18214 );
not \U$17888 ( \18231 , \18196 );
nand \U$17889 ( \18232 , \18230 , \18231 );
nand \U$17890 ( \18233 , \18229 , \18232 );
not \U$17891 ( \18234 , \18212 );
not \U$17892 ( \18235 , \1161 );
or \U$17893 ( \18236 , \18234 , \18235 );
nand \U$17894 ( \18237 , \6315 , \17710 );
nand \U$17895 ( \18238 , \18236 , \18237 );
not \U$17896 ( \18239 , RI9873558_190);
nor \U$17897 ( \18240 , \18238 , \18239 );
not \U$17898 ( \18241 , \18240 );
nand \U$17899 ( \18242 , \18238 , \18239 );
nand \U$17900 ( \18243 , \18241 , \18242 );
xor \U$17901 ( \18244 , \18233 , \18243 );
not \U$17902 ( \18245 , \18244 );
not \U$17903 ( \18246 , \4919 );
not \U$17904 ( \18247 , RI9872388_152);
not \U$17905 ( \18248 , \7112 );
not \U$17906 ( \18249 , \18248 );
or \U$17907 ( \18250 , \18247 , \18249 );
not \U$17908 ( \18251 , RI9872388_152);
nand \U$17909 ( \18252 , \5706 , \18251 );
nand \U$17910 ( \18253 , \18250 , \18252 );
not \U$17911 ( \18254 , \18253 );
or \U$17912 ( \18255 , \18246 , \18254 );
nand \U$17913 ( \18256 , \17189 , \5047 );
nand \U$17914 ( \18257 , \18255 , \18256 );
not \U$17915 ( \18258 , \18257 );
or \U$17916 ( \18259 , \18245 , \18258 );
not \U$17917 ( \18260 , \18232 );
not \U$17918 ( \18261 , \18229 );
or \U$17919 ( \18262 , \18260 , \18261 );
nand \U$17920 ( \18263 , \18262 , \18243 );
nand \U$17921 ( \18264 , \18259 , \18263 );
xor \U$17922 ( \18265 , \18185 , \18264 );
not \U$17923 ( \18266 , \18265 );
or \U$17924 ( \18267 , \18141 , \18266 );
or \U$17925 ( \18268 , \18265 , \18140 );
nand \U$17926 ( \18269 , \18267 , \18268 );
not \U$17927 ( \18270 , \5034 );
not \U$17928 ( \18271 , \17968 );
or \U$17929 ( \18272 , \18270 , \18271 );
nand \U$17930 ( \18273 , \17203 , \5796 );
nand \U$17931 ( \18274 , \18272 , \18273 );
not \U$17932 ( \18275 , \5642 );
not \U$17933 ( \18276 , \17982 );
or \U$17934 ( \18277 , \18275 , \18276 );
nand \U$17935 ( \18278 , \17809 , \5653 );
nand \U$17936 ( \18279 , \18277 , \18278 );
xor \U$17937 ( \18280 , \18274 , \18279 );
not \U$17938 ( \18281 , \16920 );
not \U$17939 ( \18282 , \8752 );
or \U$17940 ( \18283 , \18281 , \18282 );
not \U$17941 ( \18284 , \8743 );
or \U$17942 ( \18285 , \17951 , \18284 );
nand \U$17943 ( \18286 , \18283 , \18285 );
and \U$17944 ( \18287 , \18280 , \18286 );
and \U$17945 ( \18288 , \18274 , \18279 );
or \U$17946 ( \18289 , \18287 , \18288 );
not \U$17947 ( \18290 , \793 );
and \U$17948 ( \18291 , \8650 , \7075 );
not \U$17949 ( \18292 , \8650 );
and \U$17950 ( \18293 , \18292 , RI98719b0_131);
nor \U$17951 ( \18294 , \18291 , \18293 );
not \U$17952 ( \18295 , \18294 );
or \U$17953 ( \18296 , \18290 , \18295 );
xnor \U$17954 ( \18297 , \9880 , RI98719b0_131);
nand \U$17955 ( \18298 , \6145 , \18297 );
nand \U$17956 ( \18299 , \18296 , \18298 );
not \U$17957 ( \18300 , \1083 );
and \U$17958 ( \18301 , RI98718c0_129, \8555 );
not \U$17959 ( \18302 , RI98718c0_129);
and \U$17960 ( \18303 , \18302 , \9760 );
or \U$17961 ( \18304 , \18301 , \18303 );
not \U$17962 ( \18305 , \18304 );
or \U$17963 ( \18306 , \18300 , \18305 );
not \U$17964 ( \18307 , RI98718c0_129);
not \U$17965 ( \18308 , \8840 );
not \U$17966 ( \18309 , \18308 );
not \U$17967 ( \18310 , \18309 );
or \U$17968 ( \18311 , \18307 , \18310 );
not \U$17969 ( \18312 , \12847 );
nand \U$17970 ( \18313 , \18312 , \1111 );
nand \U$17971 ( \18314 , \18311 , \18313 );
nand \U$17972 ( \18315 , \18314 , \6672 );
nand \U$17973 ( \18316 , \18306 , \18315 );
or \U$17974 ( \18317 , \18299 , \18316 );
not \U$17975 ( \18318 , \1429 );
and \U$17976 ( \18319 , RI9871c08_136, \8723 );
not \U$17977 ( \18320 , RI9871c08_136);
and \U$17978 ( \18321 , \18320 , \8722 );
or \U$17979 ( \18322 , \18319 , \18321 );
not \U$17980 ( \18323 , \18322 );
or \U$17981 ( \18324 , \18318 , \18323 );
not \U$17982 ( \18325 , \3487 );
not \U$17983 ( \18326 , \8695 );
or \U$17984 ( \18327 , \18325 , \18326 );
buf \U$17985 ( \18328 , \8693 );
not \U$17986 ( \18329 , \18328 );
not \U$17987 ( \18330 , \18329 );
nand \U$17988 ( \18331 , \18330 , RI9871c08_136);
nand \U$17989 ( \18332 , \18327 , \18331 );
nand \U$17990 ( \18333 , \18332 , \1455 );
nand \U$17991 ( \18334 , \18324 , \18333 );
nand \U$17992 ( \18335 , \18317 , \18334 );
nand \U$17993 ( \18336 , \18299 , \18316 );
nand \U$17994 ( \18337 , \18335 , \18336 );
not \U$17995 ( \18338 , \1500 );
not \U$17996 ( \18339 , \17763 );
or \U$17997 ( \18340 , \18338 , \18339 );
not \U$17998 ( \18341 , \17897 );
not \U$17999 ( \18342 , RI9871c80_137);
and \U$18000 ( \18343 , \18341 , \18342 );
not \U$18001 ( \18344 , \9113 );
and \U$18002 ( \18345 , \18344 , RI9871c80_137);
nor \U$18003 ( \18346 , \18343 , \18345 );
nand \U$18004 ( \18347 , \18346 , \1517 );
nand \U$18005 ( \18348 , \18340 , \18347 );
not \U$18006 ( \18349 , \1352 );
buf \U$18007 ( \18350 , \13622 );
and \U$18008 ( \18351 , \18350 , \5621 );
not \U$18009 ( \18352 , \18350 );
and \U$18010 ( \18353 , \18352 , RI9871e60_141);
nor \U$18011 ( \18354 , \18351 , \18353 );
not \U$18012 ( \18355 , \18354 );
or \U$18013 ( \18356 , \18349 , \18355 );
nand \U$18014 ( \18357 , \17851 , \1379 );
nand \U$18015 ( \18358 , \18356 , \18357 );
xor \U$18016 ( \18359 , \18348 , \18358 );
not \U$18017 ( \18360 , \9876 );
and \U$18018 ( \18361 , RI9872130_147, \10064 );
not \U$18019 ( \18362 , RI9872130_147);
and \U$18020 ( \18363 , \18362 , \13876 );
or \U$18021 ( \18364 , \18361 , \18363 );
not \U$18022 ( \18365 , \18364 );
or \U$18023 ( \18366 , \18360 , \18365 );
nand \U$18024 ( \18367 , \18157 , \875 );
nand \U$18025 ( \18368 , \18366 , \18367 );
xor \U$18026 ( \18369 , \18359 , \18368 );
xor \U$18027 ( \18370 , \18337 , \18369 );
xor \U$18028 ( \18371 , \18289 , \18370 );
xor \U$18029 ( \18372 , \18269 , \18371 );
not \U$18030 ( \18373 , \18372 );
or \U$18031 ( \18374 , \18088 , \18373 );
nand \U$18032 ( \18375 , \18269 , \18371 );
nand \U$18033 ( \18376 , \18374 , \18375 );
not \U$18034 ( \18377 , \17794 );
not \U$18035 ( \18378 , \17811 );
or \U$18036 ( \18379 , \18377 , \18378 );
not \U$18037 ( \18380 , \17753 );
nand \U$18038 ( \18381 , \18380 , \17790 );
nand \U$18039 ( \18382 , \18379 , \18381 );
xor \U$18040 ( \18383 , \17381 , \18382 );
not \U$18041 ( \18384 , \17385 );
not \U$18042 ( \18385 , \17396 );
or \U$18043 ( \18386 , \18384 , \18385 );
or \U$18044 ( \18387 , \17396 , \17385 );
nand \U$18045 ( \18388 , \18386 , \18387 );
xor \U$18046 ( \18389 , \18383 , \18388 );
xor \U$18047 ( \18390 , \17332 , \17353 );
xor \U$18048 ( \18391 , \18390 , \17344 );
xor \U$18049 ( \18392 , \18389 , \18391 );
not \U$18050 ( \18393 , \18392 );
not \U$18051 ( \18394 , \5653 );
and \U$18052 ( \18395 , \5595 , \5648 );
not \U$18053 ( \18396 , \5595 );
and \U$18054 ( \18397 , \18396 , RI9872568_156);
nor \U$18055 ( \18398 , \18395 , \18397 );
not \U$18056 ( \18399 , \18398 );
or \U$18057 ( \18400 , \18394 , \18399 );
nand \U$18058 ( \18401 , \17803 , \5642 );
nand \U$18059 ( \18402 , \18400 , \18401 );
or \U$18060 ( \18403 , \18348 , \18358 );
nand \U$18061 ( \18404 , \18403 , \18368 );
nand \U$18062 ( \18405 , \18348 , \18358 );
and \U$18063 ( \18406 , \18404 , \18405 );
not \U$18064 ( \18407 , \18406 );
not \U$18065 ( \18408 , \17751 );
not \U$18066 ( \18409 , \17731 );
or \U$18067 ( \18410 , \18408 , \18409 );
nand \U$18068 ( \18411 , \17730 , \17705 );
nand \U$18069 ( \18412 , \18410 , \18411 );
not \U$18070 ( \18413 , \18412 );
and \U$18071 ( \18414 , \18407 , \18413 );
and \U$18072 ( \18415 , \18406 , \18412 );
nor \U$18073 ( \18416 , \18414 , \18415 );
and \U$18074 ( \18417 , \18402 , \18416 );
not \U$18075 ( \18418 , \18402 );
not \U$18076 ( \18419 , \18416 );
and \U$18077 ( \18420 , \18418 , \18419 );
nor \U$18078 ( \18421 , \18417 , \18420 );
not \U$18079 ( \18422 , \18421 );
not \U$18080 ( \18423 , \18422 );
xor \U$18081 ( \18424 , \17405 , \17414 );
xor \U$18082 ( \18425 , \18424 , \17425 );
not \U$18083 ( \18426 , \18425 );
not \U$18084 ( \18427 , \18426 );
or \U$18085 ( \18428 , \18423 , \18427 );
nand \U$18086 ( \18429 , \18425 , \18421 );
nand \U$18087 ( \18430 , \18428 , \18429 );
xor \U$18088 ( \18431 , \17666 , \18430 );
xnor \U$18089 ( \18432 , \18431 , \17673 );
not \U$18090 ( \18433 , \18432 );
or \U$18091 ( \18434 , \18393 , \18433 );
or \U$18092 ( \18435 , \18432 , \18392 );
nand \U$18093 ( \18436 , \18434 , \18435 );
xor \U$18094 ( \18437 , \18376 , \18436 );
not \U$18095 ( \18438 , \18437 );
xor \U$18096 ( \18439 , \17815 , \17821 );
xor \U$18097 ( \18440 , \18439 , \17824 );
not \U$18098 ( \18441 , \18440 );
xor \U$18099 ( \18442 , \17927 , \17830 );
xnor \U$18100 ( \18443 , \18442 , \17929 );
nand \U$18101 ( \18444 , \18441 , \18443 );
not \U$18102 ( \18445 , \18444 );
not \U$18103 ( \18446 , \9668 );
not \U$18104 ( \18447 , \18005 );
or \U$18105 ( \18448 , \18446 , \18447 );
not \U$18106 ( \18449 , \2098 );
and \U$18107 ( \18450 , \2105 , \18449 );
not \U$18108 ( \18451 , \2105 );
and \U$18109 ( \18452 , \18451 , \2098 );
nor \U$18110 ( \18453 , \18450 , \18452 );
and \U$18111 ( \18454 , RI9872bf8_170, \18453 );
not \U$18112 ( \18455 , RI9872bf8_170);
and \U$18113 ( \18456 , \18455 , \9162 );
nor \U$18114 ( \18457 , \18454 , \18456 );
nand \U$18115 ( \18458 , \18457 , \9670 );
nand \U$18116 ( \18459 , \18448 , \18458 );
not \U$18117 ( \18460 , \9214 );
not \U$18118 ( \18461 , \18059 );
or \U$18119 ( \18462 , \18460 , \18461 );
not \U$18120 ( \18463 , RI9872b80_169);
not \U$18121 ( \18464 , \3859 );
or \U$18122 ( \18465 , \18463 , \18464 );
or \U$18123 ( \18466 , \3859 , RI9872b80_169);
nand \U$18124 ( \18467 , \18465 , \18466 );
nand \U$18125 ( \18468 , \18467 , \9196 );
nand \U$18126 ( \18469 , \18462 , \18468 );
xor \U$18127 ( \18470 , \18459 , \18469 );
not \U$18128 ( \18471 , \17263 );
not \U$18129 ( \18472 , \18077 );
or \U$18130 ( \18473 , \18471 , \18472 );
and \U$18131 ( \18474 , RI98733f0_187, \1445 );
not \U$18132 ( \18475 , RI98733f0_187);
and \U$18133 ( \18476 , \18475 , \10673 );
or \U$18134 ( \18477 , \18474 , \18476 );
nand \U$18135 ( \18478 , \18477 , \17251 );
nand \U$18136 ( \18479 , \18473 , \18478 );
and \U$18137 ( \18480 , \18470 , \18479 );
and \U$18138 ( \18481 , \18459 , \18469 );
or \U$18139 ( \18482 , \18480 , \18481 );
not \U$18140 ( \18483 , \18482 );
not \U$18141 ( \18484 , \18483 );
not \U$18142 ( \18485 , \5653 );
not \U$18143 ( \18486 , \17989 );
or \U$18144 ( \18487 , \18485 , \18486 );
not \U$18145 ( \18488 , \5648 );
not \U$18146 ( \18489 , \5393 );
or \U$18147 ( \18490 , \18488 , \18489 );
nand \U$18148 ( \18491 , \5775 , RI9872568_156);
nand \U$18149 ( \18492 , \18490 , \18491 );
nand \U$18150 ( \18493 , \18492 , \5642 );
nand \U$18151 ( \18494 , \18487 , \18493 );
not \U$18152 ( \18495 , \6672 );
and \U$18153 ( \18496 , RI98718c0_129, \12470 );
not \U$18154 ( \18497 , RI98718c0_129);
not \U$18155 ( \18498 , \8722 );
and \U$18156 ( \18499 , \18497 , \18498 );
nor \U$18157 ( \18500 , \18496 , \18499 );
not \U$18158 ( \18501 , \18500 );
or \U$18159 ( \18502 , \18495 , \18501 );
xor \U$18160 ( \18503 , RI98718c0_129, \8695 );
nand \U$18161 ( \18504 , \18503 , \1083 );
nand \U$18162 ( \18505 , \18502 , \18504 );
or \U$18163 ( \18506 , \18494 , \18505 );
not \U$18164 ( \18507 , \18506 );
buf \U$18165 ( \18508 , \17543 );
not \U$18166 ( \18509 , \18508 );
not \U$18167 ( \18510 , RI9873288_184);
not \U$18168 ( \18511 , \1581 );
or \U$18169 ( \18512 , \18510 , \18511 );
or \U$18170 ( \18513 , \1581 , RI9873288_184);
nand \U$18171 ( \18514 , \18512 , \18513 );
not \U$18172 ( \18515 , \18514 );
or \U$18173 ( \18516 , \18509 , \18515 );
not \U$18174 ( \18517 , RI9873288_184);
not \U$18175 ( \18518 , \1319 );
or \U$18176 ( \18519 , \18517 , \18518 );
or \U$18177 ( \18520 , \9230 , RI9873288_184);
nand \U$18178 ( \18521 , \18519 , \18520 );
buf \U$18179 ( \18522 , \17528 );
nand \U$18180 ( \18523 , \18521 , \18522 );
nand \U$18181 ( \18524 , \18516 , \18523 );
not \U$18182 ( \18525 , \18524 );
or \U$18183 ( \18526 , \18507 , \18525 );
nand \U$18184 ( \18527 , \18494 , \18505 );
nand \U$18185 ( \18528 , \18526 , \18527 );
not \U$18186 ( \18529 , \18528 );
not \U$18187 ( \18530 , \18529 );
or \U$18188 ( \18531 , \18484 , \18530 );
not \U$18189 ( \18532 , \9526 );
and \U$18190 ( \18533 , RI9872f40_177, \1365 );
not \U$18191 ( \18534 , RI9872f40_177);
and \U$18192 ( \18535 , \18534 , \1603 );
nor \U$18193 ( \18536 , \18533 , \18535 );
not \U$18194 ( \18537 , \18536 );
or \U$18195 ( \18538 , \18532 , \18537 );
nand \U$18196 ( \18539 , \17959 , \11198 );
nand \U$18197 ( \18540 , \18538 , \18539 );
not \U$18198 ( \18541 , \18540 );
not \U$18199 ( \18542 , RI9873648_192);
and \U$18200 ( \18543 , \18542 , RI9873558_190);
buf \U$18201 ( \18544 , \18543 );
buf \U$18202 ( \18545 , \18544 );
not \U$18203 ( \18546 , \18545 );
xor \U$18204 ( \18547 , RI9873558_190, \1393 );
not \U$18205 ( \18548 , \18547 );
or \U$18206 ( \18549 , \18546 , \18548 );
and \U$18207 ( \18550 , RI9873558_190, \779 );
not \U$18208 ( \18551 , RI9873558_190);
and \U$18209 ( \18552 , \18551 , \1690 );
or \U$18210 ( \18553 , \18550 , \18552 );
nand \U$18211 ( \18554 , \18553 , RI9873648_192);
nand \U$18212 ( \18555 , \18549 , \18554 );
not \U$18213 ( \18556 , \18555 );
not \U$18214 ( \18557 , \18556 );
or \U$18215 ( \18558 , \18541 , \18557 );
or \U$18216 ( \18559 , \18556 , \18540 );
nand \U$18217 ( \18560 , \18558 , \18559 );
not \U$18218 ( \18561 , \18560 );
buf \U$18219 ( \18562 , \9293 );
buf \U$18220 ( \18563 , \18562 );
not \U$18221 ( \18564 , \18563 );
not \U$18222 ( \18565 , RI9872e50_175);
not \U$18223 ( \18566 , \17140 );
or \U$18224 ( \18567 , \18565 , \18566 );
and \U$18225 ( \18568 , \1031 , \1033 );
not \U$18226 ( \18569 , \1031 );
and \U$18227 ( \18570 , \18569 , \1032 );
nor \U$18228 ( \18571 , \18568 , \18570 );
not \U$18229 ( \18572 , \18571 );
or \U$18230 ( \18573 , \18572 , RI9872e50_175);
nand \U$18231 ( \18574 , \18567 , \18573 );
not \U$18232 ( \18575 , \18574 );
or \U$18233 ( \18576 , \18564 , \18575 );
not \U$18234 ( \18577 , \9690 );
not \U$18235 ( \18578 , \1713 );
or \U$18236 ( \18579 , \18577 , \18578 );
or \U$18237 ( \18580 , \1061 , \9694 );
nand \U$18238 ( \18581 , \18579 , \18580 );
nand \U$18239 ( \18582 , \18581 , \9273 );
nand \U$18240 ( \18583 , \18576 , \18582 );
not \U$18241 ( \18584 , \18583 );
or \U$18242 ( \18585 , \18561 , \18584 );
nand \U$18243 ( \18586 , \18555 , \18540 );
nand \U$18244 ( \18587 , \18585 , \18586 );
nand \U$18245 ( \18588 , \18531 , \18587 );
nand \U$18246 ( \18589 , \18528 , \18482 );
nand \U$18247 ( \18590 , \18588 , \18589 );
not \U$18248 ( \18591 , \18590 );
xor \U$18249 ( \18592 , \17789 , \17774 );
and \U$18250 ( \18593 , \18181 , \18169 );
not \U$18251 ( \18594 , \18181 );
not \U$18252 ( \18595 , \18169 );
and \U$18253 ( \18596 , \18594 , \18595 );
nor \U$18254 ( \18597 , \18593 , \18596 );
xor \U$18255 ( \18598 , \18592 , \18597 );
not \U$18256 ( \18599 , \18332 );
not \U$18257 ( \18600 , \1429 );
or \U$18258 ( \18601 , \18599 , \18600 );
and \U$18259 ( \18602 , RI9871c08_136, \12460 );
not \U$18260 ( \18603 , RI9871c08_136);
and \U$18261 ( \18604 , \18603 , \8708 );
or \U$18262 ( \18605 , \18602 , \18604 );
not \U$18263 ( \18606 , \18605 );
or \U$18264 ( \18607 , \18606 , \5411 );
nand \U$18265 ( \18608 , \18601 , \18607 );
not \U$18266 ( \18609 , \1136 );
not \U$18267 ( \18610 , \18304 );
or \U$18268 ( \18611 , \18609 , \18610 );
nand \U$18269 ( \18612 , \18500 , \1083 );
nand \U$18270 ( \18613 , \18611 , \18612 );
xor \U$18271 ( \18614 , \18608 , \18613 );
buf \U$18272 ( \18615 , \18544 );
not \U$18273 ( \18616 , \18615 );
not \U$18274 ( \18617 , \18553 );
or \U$18275 ( \18618 , \18616 , \18617 );
nand \U$18276 ( \18619 , RI9873558_190, RI9873648_192);
nand \U$18277 ( \18620 , \18618 , \18619 );
and \U$18278 ( \18621 , \18614 , \18620 );
and \U$18279 ( \18622 , \18608 , \18613 );
or \U$18280 ( \18623 , \18621 , \18622 );
xnor \U$18281 ( \18624 , \18598 , \18623 );
not \U$18282 ( \18625 , \18624 );
and \U$18283 ( \18626 , \18591 , \18625 );
and \U$18284 ( \18627 , \18590 , \18624 );
nor \U$18285 ( \18628 , \18626 , \18627 );
not \U$18286 ( \18629 , \18628 );
not \U$18287 ( \18630 , \18629 );
xor \U$18288 ( \18631 , \18608 , \18613 );
xor \U$18289 ( \18632 , \18631 , \18620 );
not \U$18290 ( \18633 , \18632 );
not \U$18291 ( \18634 , \6284 );
xor \U$18292 ( \18635 , \4960 , RI98728b0_163);
not \U$18293 ( \18636 , \18635 );
or \U$18294 ( \18637 , \18634 , \18636 );
and \U$18295 ( \18638 , RI98728b0_163, \4711 );
not \U$18296 ( \18639 , RI98728b0_163);
and \U$18297 ( \18640 , \18639 , \4712 );
or \U$18298 ( \18641 , \18638 , \18640 );
nand \U$18299 ( \18642 , \18641 , \6286 );
nand \U$18300 ( \18643 , \18637 , \18642 );
not \U$18301 ( \18644 , \18643 );
not \U$18302 ( \18645 , \7338 );
not \U$18303 ( \18646 , RI98729a0_165);
buf \U$18304 ( \18647 , \4175 );
not \U$18305 ( \18648 , \18647 );
or \U$18306 ( \18649 , \18646 , \18648 );
or \U$18307 ( \18650 , \11028 , RI98729a0_165);
nand \U$18308 ( \18651 , \18649 , \18650 );
not \U$18309 ( \18652 , \18651 );
or \U$18310 ( \18653 , \18645 , \18652 );
not \U$18311 ( \18654 , RI98729a0_165);
not \U$18312 ( \18655 , \5205 );
or \U$18313 ( \18656 , \18654 , \18655 );
or \U$18314 ( \18657 , \5614 , RI98729a0_165);
nand \U$18315 ( \18658 , \18656 , \18657 );
nand \U$18316 ( \18659 , \18658 , \7325 );
nand \U$18317 ( \18660 , \18653 , \18659 );
not \U$18318 ( \18661 , \9937 );
xor \U$18319 ( \18662 , RI9873030_179, \942 );
not \U$18320 ( \18663 , \18662 );
or \U$18321 ( \18664 , \18661 , \18663 );
and \U$18322 ( \18665 , \1246 , \1247 );
not \U$18323 ( \18666 , \1246 );
and \U$18324 ( \18667 , \18666 , \1250 );
nor \U$18325 ( \18668 , \18665 , \18667 );
or \U$18326 ( \18669 , RI9873030_179, \18668 );
or \U$18327 ( \18670 , \5719 , \14132 );
nand \U$18328 ( \18671 , \18669 , \18670 );
buf \U$18329 ( \18672 , \12507 );
nand \U$18330 ( \18673 , \18671 , \18672 );
nand \U$18331 ( \18674 , \18664 , \18673 );
xor \U$18332 ( \18675 , \18660 , \18674 );
not \U$18333 ( \18676 , \18675 );
or \U$18334 ( \18677 , \18644 , \18676 );
nand \U$18335 ( \18678 , \18660 , \18674 );
nand \U$18336 ( \18679 , \18677 , \18678 );
not \U$18337 ( \18680 , \18679 );
not \U$18338 ( \18681 , \9072 );
not \U$18339 ( \18682 , \8031 );
not \U$18340 ( \18683 , \3536 );
or \U$18341 ( \18684 , \18682 , \18683 );
not \U$18342 ( \18685 , \12543 );
or \U$18343 ( \18686 , \18685 , \8031 );
nand \U$18344 ( \18687 , \18684 , \18686 );
not \U$18345 ( \18688 , \18687 );
or \U$18346 ( \18689 , \18681 , \18688 );
not \U$18347 ( \18690 , RI9872a18_166);
not \U$18348 ( \18691 , \3567 );
or \U$18349 ( \18692 , \18690 , \18691 );
or \U$18350 ( \18693 , \3567 , RI9872a18_166);
nand \U$18351 ( \18694 , \18692 , \18693 );
nand \U$18352 ( \18695 , \18694 , \8028 );
nand \U$18353 ( \18696 , \18689 , \18695 );
not \U$18354 ( \18697 , \18696 );
not \U$18355 ( \18698 , \8678 );
and \U$18356 ( \18699 , RI9870498_86, RI9870420_85);
not \U$18357 ( \18700 , RI9870498_86);
not \U$18358 ( \18701 , RI9870420_85);
and \U$18359 ( \18702 , \18700 , \18701 );
nor \U$18360 ( \18703 , \18699 , \18702 );
buf \U$18361 ( \18704 , \18703 );
buf \U$18362 ( \18705 , \18704 );
not \U$18363 ( \18706 , \18705 );
nor \U$18364 ( \18707 , \18698 , \18706 );
not \U$18365 ( \18708 , \859 );
buf \U$18366 ( \18709 , \17003 );
not \U$18367 ( \18710 , \18709 );
and \U$18368 ( \18711 , RI9871d70_139, \18710 );
not \U$18369 ( \18712 , RI9871d70_139);
not \U$18370 ( \18713 , \13934 );
and \U$18371 ( \18714 , \18712 , \18713 );
or \U$18372 ( \18715 , \18711 , \18714 );
not \U$18373 ( \18716 , \18715 );
or \U$18374 ( \18717 , \18708 , \18716 );
nand \U$18375 ( \18718 , \17885 , \832 );
nand \U$18376 ( \18719 , \18717 , \18718 );
xor \U$18377 ( \18720 , \18707 , \18719 );
not \U$18378 ( \18721 , \18196 );
and \U$18379 ( \18722 , \1164 , \18194 );
nor \U$18380 ( \18723 , \18721 , \18722 );
not \U$18381 ( \18724 , \18723 );
not \U$18382 ( \18725 , \1161 );
or \U$18383 ( \18726 , \18724 , \18725 );
nand \U$18384 ( \18727 , \6315 , \18201 );
nand \U$18385 ( \18728 , \18726 , \18727 );
xor \U$18386 ( \18729 , \18720 , \18728 );
not \U$18387 ( \18730 , \18729 );
not \U$18388 ( \18731 , \18730 );
not \U$18389 ( \18732 , \17347 );
not \U$18390 ( \18733 , \18051 );
or \U$18391 ( \18734 , \18732 , \18733 );
and \U$18392 ( \18735 , RI98730a8_180, \846 );
not \U$18393 ( \18736 , RI98730a8_180);
not \U$18394 ( \18737 , \846 );
and \U$18395 ( \18738 , \18736 , \18737 );
nor \U$18396 ( \18739 , \18735 , \18738 );
nand \U$18397 ( \18740 , \18739 , \13020 );
nand \U$18398 ( \18741 , \18734 , \18740 );
not \U$18399 ( \18742 , \18741 );
or \U$18400 ( \18743 , \18731 , \18742 );
or \U$18401 ( \18744 , \18741 , \18730 );
nand \U$18402 ( \18745 , \18743 , \18744 );
not \U$18403 ( \18746 , \18745 );
or \U$18404 ( \18747 , \18697 , \18746 );
nand \U$18405 ( \18748 , \18741 , \18729 );
nand \U$18406 ( \18749 , \18747 , \18748 );
xnor \U$18407 ( \18750 , \18680 , \18749 );
not \U$18408 ( \18751 , \18750 );
or \U$18409 ( \18752 , \18633 , \18751 );
nand \U$18410 ( \18753 , \18749 , \18679 );
nand \U$18411 ( \18754 , \18752 , \18753 );
not \U$18412 ( \18755 , \18754 );
or \U$18413 ( \18756 , \18630 , \18755 );
not \U$18414 ( \18757 , \18624 );
nand \U$18415 ( \18758 , \18757 , \18590 );
nand \U$18416 ( \18759 , \18756 , \18758 );
not \U$18417 ( \18760 , \18759 );
or \U$18418 ( \18761 , \18445 , \18760 );
not \U$18419 ( \18762 , \18443 );
nand \U$18420 ( \18763 , \18762 , \18440 );
nand \U$18421 ( \18764 , \18761 , \18763 );
not \U$18422 ( \18765 , \18764 );
not \U$18423 ( \18766 , \17680 );
and \U$18424 ( \18767 , \17939 , \18766 );
not \U$18425 ( \18768 , \17939 );
and \U$18426 ( \18769 , \18768 , \17680 );
nor \U$18427 ( \18770 , \18767 , \18769 );
buf \U$18428 ( \18771 , \18770 );
and \U$18429 ( \18772 , \18765 , \18771 );
not \U$18430 ( \18773 , \18765 );
not \U$18431 ( \18774 , \18771 );
and \U$18432 ( \18775 , \18773 , \18774 );
nor \U$18433 ( \18776 , \18772 , \18775 );
not \U$18434 ( \18777 , \18776 );
or \U$18435 ( \18778 , \18438 , \18777 );
nand \U$18436 ( \18779 , \18764 , \18774 );
nand \U$18437 ( \18780 , \18778 , \18779 );
xor \U$18438 ( \18781 , \17945 , \18780 );
not \U$18439 ( \18782 , \16997 );
not \U$18440 ( \18783 , \17000 );
and \U$18441 ( \18784 , \18782 , \18783 );
xor \U$18442 ( \18785 , \16997 , \17000 );
and \U$18443 ( \18786 , \17021 , \18785 );
nor \U$18444 ( \18787 , \18784 , \18786 );
not \U$18445 ( \18788 , \18787 );
not \U$18446 ( \18789 , \12514 );
not \U$18447 ( \18790 , \3154 );
not \U$18448 ( \18791 , \7905 );
or \U$18449 ( \18792 , \18790 , \18791 );
buf \U$18450 ( \18793 , \10411 );
not \U$18451 ( \18794 , \18793 );
nand \U$18452 ( \18795 , \18794 , RI9872310_151);
nand \U$18453 ( \18796 , \18792 , \18795 );
not \U$18454 ( \18797 , \18796 );
or \U$18455 ( \18798 , \18789 , \18797 );
nand \U$18456 ( \18799 , \17453 , \13033 );
nand \U$18457 ( \18800 , \18798 , \18799 );
not \U$18458 ( \18801 , \18800 );
or \U$18459 ( \18802 , \18788 , \18801 );
or \U$18460 ( \18803 , \18800 , \18787 );
nand \U$18461 ( \18804 , \18802 , \18803 );
buf \U$18462 ( \18805 , \18804 );
not \U$18463 ( \18806 , \3467 );
not \U$18464 ( \18807 , \4063 );
not \U$18465 ( \18808 , \5704 );
buf \U$18466 ( \18809 , \18808 );
not \U$18467 ( \18810 , \18809 );
or \U$18468 ( \18811 , \18807 , \18810 );
nand \U$18469 ( \18812 , \6308 , RI98726d0_159);
nand \U$18470 ( \18813 , \18811 , \18812 );
not \U$18471 ( \18814 , \18813 );
or \U$18472 ( \18815 , \18806 , \18814 );
nand \U$18473 ( \18816 , \17463 , \3600 );
nand \U$18474 ( \18817 , \18815 , \18816 );
and \U$18475 ( \18818 , \18805 , \18817 );
not \U$18476 ( \18819 , \18805 );
not \U$18477 ( \18820 , \18817 );
and \U$18478 ( \18821 , \18819 , \18820 );
nor \U$18479 ( \18822 , \18818 , \18821 );
xor \U$18480 ( \18823 , \17486 , \17496 );
and \U$18481 ( \18824 , \18823 , \17507 );
and \U$18482 ( \18825 , \17486 , \17496 );
or \U$18483 ( \18826 , \18824 , \18825 );
xor \U$18484 ( \18827 , \18822 , \18826 );
not \U$18485 ( \18828 , \9876 );
and \U$18486 ( \18829 , \9139 , RI9872130_147);
not \U$18487 ( \18830 , \9139 );
and \U$18488 ( \18831 , \18830 , \919 );
nor \U$18489 ( \18832 , \18829 , \18831 );
not \U$18490 ( \18833 , \18832 );
or \U$18491 ( \18834 , \18828 , \18833 );
nand \U$18492 ( \18835 , \18364 , \875 );
nand \U$18493 ( \18836 , \18834 , \18835 );
not \U$18494 ( \18837 , \18836 );
not \U$18495 ( \18838 , \17728 );
not \U$18496 ( \18839 , \9429 );
or \U$18497 ( \18840 , \18838 , \18839 );
not \U$18498 ( \18841 , \17908 );
xnor \U$18499 ( \18842 , \1164 , \18841 );
nand \U$18500 ( \18843 , \6315 , \18842 );
nand \U$18501 ( \18844 , \18840 , \18843 );
xor \U$18502 ( \18845 , \18844 , \17751 );
not \U$18503 ( \18846 , \18845 );
not \U$18504 ( \18847 , \18846 );
or \U$18505 ( \18848 , \18837 , \18847 );
nand \U$18506 ( \18849 , \18844 , \17748 );
nand \U$18507 ( \18850 , \18848 , \18849 );
not \U$18508 ( \18851 , \5796 );
xor \U$18509 ( \18852 , \7355 , RI9872478_154);
not \U$18510 ( \18853 , \18852 );
or \U$18511 ( \18854 , \18851 , \18853 );
nand \U$18512 ( \18855 , \17412 , \5034 );
nand \U$18513 ( \18856 , \18854 , \18855 );
xor \U$18514 ( \18857 , \18850 , \18856 );
not \U$18515 ( \18858 , \10333 );
not \U$18516 ( \18859 , RI9872e50_175);
not \U$18517 ( \18860 , \6224 );
or \U$18518 ( \18861 , \18859 , \18860 );
not \U$18519 ( \18862 , RI9872e50_175);
nand \U$18520 ( \18863 , \16925 , \18862 );
nand \U$18521 ( \18864 , \18861 , \18863 );
not \U$18522 ( \18865 , \18864 );
or \U$18523 ( \18866 , \18858 , \18865 );
nand \U$18524 ( \18867 , \17421 , \9294 );
nand \U$18525 ( \18868 , \18866 , \18867 );
xor \U$18526 ( \18869 , \18857 , \18868 );
xor \U$18527 ( \18870 , \18827 , \18869 );
not \U$18528 ( \18871 , \18391 );
not \U$18529 ( \18872 , \18871 );
not \U$18530 ( \18873 , \18389 );
or \U$18531 ( \18874 , \18872 , \18873 );
xor \U$18532 ( \18875 , \17369 , \17381 );
xor \U$18533 ( \18876 , \18875 , \17396 );
nand \U$18534 ( \18877 , \18876 , \18382 );
nand \U$18535 ( \18878 , \18874 , \18877 );
xor \U$18536 ( \18879 , \18870 , \18878 );
not \U$18537 ( \18880 , \18422 );
not \U$18538 ( \18881 , \18425 );
or \U$18539 ( \18882 , \18880 , \18881 );
xor \U$18540 ( \18883 , \17666 , \17657 );
xnor \U$18541 ( \18884 , \18883 , \17646 );
nand \U$18542 ( \18885 , \18426 , \18421 );
nand \U$18543 ( \18886 , \18884 , \18885 );
nand \U$18544 ( \18887 , \18882 , \18886 );
xor \U$18545 ( \18888 , \18879 , \18887 );
not \U$18546 ( \18889 , \18376 );
not \U$18547 ( \18890 , \18436 );
or \U$18548 ( \18891 , \18889 , \18890 );
not \U$18549 ( \18892 , \18392 );
nand \U$18550 ( \18893 , \18892 , \18432 );
nand \U$18551 ( \18894 , \18891 , \18893 );
xor \U$18552 ( \18895 , \18888 , \18894 );
and \U$18553 ( \18896 , \18402 , \18419 );
not \U$18554 ( \18897 , \18412 );
nor \U$18555 ( \18898 , \18897 , \18406 );
nor \U$18556 ( \18899 , \18896 , \18898 );
not \U$18557 ( \18900 , \9214 );
not \U$18558 ( \18901 , RI9872b80_169);
not \U$18559 ( \18902 , \9323 );
or \U$18560 ( \18903 , \18901 , \18902 );
buf \U$18561 ( \18904 , \6333 );
or \U$18562 ( \18905 , \18904 , RI9872b80_169);
nand \U$18563 ( \18906 , \18903 , \18905 );
not \U$18564 ( \18907 , \18906 );
or \U$18565 ( \18908 , \18900 , \18907 );
nand \U$18566 ( \18909 , \17341 , \9196 );
nand \U$18567 ( \18910 , \18908 , \18909 );
not \U$18568 ( \18911 , \9937 );
not \U$18569 ( \18912 , RI9873030_179);
not \U$18570 ( \18913 , \1581 );
or \U$18571 ( \18914 , \18912 , \18913 );
or \U$18572 ( \18915 , \7064 , RI9873030_179);
nand \U$18573 ( \18916 , \18914 , \18915 );
not \U$18574 ( \18917 , \18916 );
or \U$18575 ( \18918 , \18911 , \18917 );
nand \U$18576 ( \18919 , \17644 , \13109 );
nand \U$18577 ( \18920 , \18918 , \18919 );
xor \U$18578 ( \18921 , \18910 , \18920 );
not \U$18579 ( \18922 , \11350 );
not \U$18580 ( \18923 , \17349 );
or \U$18581 ( \18924 , \18922 , \18923 );
and \U$18582 ( \18925 , RI98730a8_180, \1447 );
not \U$18583 ( \18926 , RI98730a8_180);
and \U$18584 ( \18927 , \18926 , \6165 );
or \U$18585 ( \18928 , \18925 , \18927 );
nand \U$18586 ( \18929 , \18928 , \12868 );
nand \U$18587 ( \18930 , \18924 , \18929 );
xor \U$18588 ( \18931 , \18921 , \18930 );
xor \U$18589 ( \18932 , \18899 , \18931 );
not \U$18590 ( \18933 , \9072 );
not \U$18591 ( \18934 , \11755 );
not \U$18592 ( \18935 , RI9872a18_166);
and \U$18593 ( \18936 , \18934 , \18935 );
not \U$18594 ( \18937 , \9255 );
and \U$18595 ( \18938 , \18937 , RI9872a18_166);
nor \U$18596 ( \18939 , \18936 , \18938 );
not \U$18597 ( \18940 , \18939 );
or \U$18598 ( \18941 , \18933 , \18940 );
nand \U$18599 ( \18942 , \17664 , \8029 );
nand \U$18600 ( \18943 , \18941 , \18942 );
not \U$18601 ( \18944 , \7326 );
not \U$18602 ( \18945 , \17494 );
or \U$18603 ( \18946 , \18944 , \18945 );
and \U$18604 ( \18947 , RI98729a0_165, \6378 );
not \U$18605 ( \18948 , RI98729a0_165);
and \U$18606 ( \18949 , \18948 , \2111 );
or \U$18607 ( \18950 , \18947 , \18949 );
nand \U$18608 ( \18951 , \18950 , \7338 );
nand \U$18609 ( \18952 , \18946 , \18951 );
nor \U$18610 ( \18953 , \18943 , \18952 );
not \U$18611 ( \18954 , \18953 );
nand \U$18612 ( \18955 , \18943 , \18952 );
nand \U$18613 ( \18956 , \18954 , \18955 );
buf \U$18614 ( \18957 , \13476 );
not \U$18615 ( \18958 , \18957 );
not \U$18616 ( \18959 , \17392 );
or \U$18617 ( \18960 , \18958 , \18959 );
not \U$18618 ( \18961 , RI9873210_183);
not \U$18619 ( \18962 , \1097 );
or \U$18620 ( \18963 , \18961 , \18962 );
or \U$18621 ( \18964 , \1097 , RI9873210_183);
nand \U$18622 ( \18965 , \18963 , \18964 );
nand \U$18623 ( \18966 , \18965 , \17234 );
nand \U$18624 ( \18967 , \18960 , \18966 );
not \U$18625 ( \18968 , \18967 );
and \U$18626 ( \18969 , \18956 , \18968 );
not \U$18627 ( \18970 , \18956 );
and \U$18628 ( \18971 , \18970 , \18967 );
nor \U$18629 ( \18972 , \18969 , \18971 );
xnor \U$18630 ( \18973 , \18932 , \18972 );
and \U$18631 ( \18974 , RI9871c80_137, \12460 );
not \U$18632 ( \18975 , RI9871c80_137);
and \U$18633 ( \18976 , \18975 , \8708 );
nor \U$18634 ( \18977 , \18974 , \18976 );
not \U$18635 ( \18978 , \18977 );
not \U$18636 ( \18979 , \1746 );
and \U$18637 ( \18980 , \18978 , \18979 );
and \U$18638 ( \18981 , \18346 , \1501 );
nor \U$18639 ( \18982 , \18980 , \18981 );
not \U$18640 ( \18983 , \18982 );
not \U$18641 ( \18984 , \859 );
not \U$18642 ( \18985 , \17085 );
or \U$18643 ( \18986 , \18984 , \18985 );
not \U$18644 ( \18987 , RI9871d70_139);
not \U$18645 ( \18988 , \11455 );
or \U$18646 ( \18989 , \18987 , \18988 );
or \U$18647 ( \18990 , \18151 , RI9871d70_139);
nand \U$18648 ( \18991 , \18989 , \18990 );
nand \U$18649 ( \18992 , \18991 , \832 );
nand \U$18650 ( \18993 , \18986 , \18992 );
not \U$18651 ( \18994 , \1352 );
not \U$18652 ( \18995 , RI9871e60_141);
not \U$18653 ( \18996 , \17090 );
or \U$18654 ( \18997 , \18995 , \18996 );
nand \U$18655 ( \18998 , \13281 , \5621 );
nand \U$18656 ( \18999 , \18997 , \18998 );
not \U$18657 ( \19000 , \18999 );
or \U$18658 ( \19001 , \18994 , \19000 );
nand \U$18659 ( \19002 , \18354 , \1380 );
nand \U$18660 ( \19003 , \19001 , \19002 );
and \U$18661 ( \19004 , \18993 , \19003 );
not \U$18662 ( \19005 , \18993 );
not \U$18663 ( \19006 , \19003 );
and \U$18664 ( \19007 , \19005 , \19006 );
nor \U$18665 ( \19008 , \19004 , \19007 );
not \U$18666 ( \19009 , \19008 );
or \U$18667 ( \19010 , \18983 , \19009 );
or \U$18668 ( \19011 , \19008 , \18982 );
nand \U$18669 ( \19012 , \19010 , \19011 );
not \U$18670 ( \19013 , \19012 );
xor \U$18671 ( \19014 , \18845 , \18836 );
not \U$18672 ( \19015 , \19014 );
and \U$18673 ( \19016 , \19013 , \19015 );
and \U$18674 ( \19017 , \19012 , \19014 );
nor \U$18675 ( \19018 , \19016 , \19017 );
not \U$18676 ( \19019 , \19018 );
not \U$18677 ( \19020 , \19019 );
not \U$18678 ( \19021 , \1430 );
not \U$18679 ( \19022 , \17043 );
or \U$18680 ( \19023 , \19021 , \19022 );
nand \U$18681 ( \19024 , \18322 , \1455 );
nand \U$18682 ( \19025 , \19023 , \19024 );
not \U$18683 ( \19026 , \19025 );
not \U$18684 ( \19027 , \1323 );
not \U$18685 ( \19028 , \17035 );
or \U$18686 ( \19029 , \19027 , \19028 );
nand \U$18687 ( \19030 , \18166 , \1292 );
nand \U$18688 ( \19031 , \19029 , \19030 );
xnor \U$18689 ( \19032 , RI98735d0_191, RI9873558_190);
xor \U$18690 ( \19033 , RI98734e0_189, RI98735d0_191);
and \U$18691 ( \19034 , \19032 , \19033 );
buf \U$18692 ( \19035 , \19034 );
buf \U$18693 ( \19036 , \19035 );
not \U$18694 ( \19037 , \19036 );
and \U$18695 ( \19038 , RI98734e0_189, \778 );
not \U$18696 ( \19039 , RI98734e0_189);
and \U$18697 ( \19040 , \19039 , \779 );
nor \U$18698 ( \19041 , \19038 , \19040 );
not \U$18699 ( \19042 , \19041 );
or \U$18700 ( \19043 , \19037 , \19042 );
not \U$18701 ( \19044 , \19032 );
buf \U$18702 ( \19045 , \19044 );
buf \U$18703 ( \19046 , \19045 );
nand \U$18704 ( \19047 , \19046 , RI98734e0_189);
nand \U$18705 ( \19048 , \19043 , \19047 );
xor \U$18706 ( \19049 , \19031 , \19048 );
not \U$18707 ( \19050 , \19049 );
or \U$18708 ( \19051 , \19026 , \19050 );
nand \U$18709 ( \19052 , \19048 , \19031 );
nand \U$18710 ( \19053 , \19051 , \19052 );
not \U$18711 ( \19054 , \19053 );
or \U$18712 ( \19055 , \19020 , \19054 );
not \U$18713 ( \19056 , \19014 );
nand \U$18714 ( \19057 , \19056 , \19012 );
nand \U$18715 ( \19058 , \19055 , \19057 );
not \U$18716 ( \19059 , \19058 );
not \U$18717 ( \19060 , \17853 );
not \U$18718 ( \19061 , \17876 );
or \U$18719 ( \19062 , \19060 , \19061 );
nand \U$18720 ( \19063 , \17875 , \17864 );
nand \U$18721 ( \19064 , \19062 , \19063 );
not \U$18722 ( \19065 , \19064 );
buf \U$18723 ( \19066 , \18240 );
nand \U$18724 ( \19067 , \19065 , \19066 );
not \U$18725 ( \19068 , \19067 );
not \U$18726 ( \19069 , \13033 );
not \U$18727 ( \19070 , \18093 );
or \U$18728 ( \19071 , \19069 , \19070 );
nand \U$18729 ( \19072 , \17445 , \3170 );
nand \U$18730 ( \19073 , \19071 , \19072 );
not \U$18731 ( \19074 , \19073 );
or \U$18732 ( \19075 , \19068 , \19074 );
not \U$18733 ( \19076 , \19066 );
nand \U$18734 ( \19077 , \19076 , \19064 );
nand \U$18735 ( \19078 , \19075 , \19077 );
not \U$18736 ( \19079 , \19078 );
not \U$18737 ( \19080 , \19079 );
not \U$18738 ( \19081 , \17078 );
not \U$18739 ( \19082 , \17117 );
or \U$18740 ( \19083 , \19081 , \19082 );
not \U$18741 ( \19084 , \17096 );
nand \U$18742 ( \19085 , \19084 , \17113 );
nand \U$18743 ( \19086 , \19083 , \19085 );
not \U$18744 ( \19087 , \19086 );
not \U$18745 ( \19088 , \19087 );
or \U$18746 ( \19089 , \19080 , \19088 );
not \U$18747 ( \19090 , \6144 );
not \U$18748 ( \19091 , \16938 );
or \U$18749 ( \19092 , \19090 , \19091 );
nand \U$18750 ( \19093 , \18297 , \11433 );
nand \U$18751 ( \19094 , \19092 , \19093 );
not \U$18752 ( \19095 , \2087 );
not \U$18753 ( \19096 , \16978 );
or \U$18754 ( \19097 , \19095 , \19096 );
nand \U$18755 ( \19098 , \18120 , \2071 );
nand \U$18756 ( \19099 , \19097 , \19098 );
or \U$18757 ( \19100 , \19094 , \19099 );
not \U$18758 ( \19101 , \6672 );
not \U$18759 ( \19102 , \16959 );
or \U$18760 ( \19103 , \19101 , \19102 );
nand \U$18761 ( \19104 , \18314 , \1083 );
nand \U$18762 ( \19105 , \19103 , \19104 );
nand \U$18763 ( \19106 , \19100 , \19105 );
nand \U$18764 ( \19107 , \19094 , \19099 );
and \U$18765 ( \19108 , \19106 , \19107 );
not \U$18766 ( \19109 , \19108 );
nand \U$18767 ( \19110 , \19089 , \19109 );
not \U$18768 ( \19111 , \19079 );
nand \U$18769 ( \19112 , \19111 , \19086 );
nand \U$18770 ( \19113 , \19110 , \19112 );
not \U$18771 ( \19114 , \19113 );
not \U$18772 ( \19115 , \19114 );
or \U$18773 ( \19116 , \19059 , \19115 );
or \U$18774 ( \19117 , \19114 , \19058 );
nand \U$18775 ( \19118 , \19116 , \19117 );
xor \U$18776 ( \19119 , \17223 , \17274 );
and \U$18777 ( \19120 , \19119 , \17318 );
and \U$18778 ( \19121 , \17223 , \17274 );
or \U$18779 ( \19122 , \19120 , \19121 );
not \U$18780 ( \19123 , \19122 );
and \U$18781 ( \19124 , \19118 , \19123 );
not \U$18782 ( \19125 , \19118 );
and \U$18783 ( \19126 , \19125 , \19122 );
or \U$18784 ( \19127 , \19124 , \19126 );
xor \U$18785 ( \19128 , \18973 , \19127 );
and \U$18786 ( \19129 , \8695 , RI9871c80_137);
not \U$18787 ( \19130 , \8695 );
and \U$18788 ( \19131 , \19130 , \1800 );
nor \U$18789 ( \19132 , \19129 , \19131 );
not \U$18790 ( \19133 , \19132 );
or \U$18791 ( \19134 , \19133 , \1746 );
or \U$18792 ( \19135 , \18977 , \1591 );
nand \U$18793 ( \19136 , \19134 , \19135 );
not \U$18794 ( \19137 , \4925 );
not \U$18795 ( \19138 , RI9872388_152);
not \U$18796 ( \19139 , \7791 );
or \U$18797 ( \19140 , \19138 , \19139 );
or \U$18798 ( \19141 , \7791 , RI9872388_152);
nand \U$18799 ( \19142 , \19140 , \19141 );
not \U$18800 ( \19143 , \19142 );
or \U$18801 ( \19144 , \19137 , \19143 );
nand \U$18802 ( \19145 , \17403 , \4918 );
nand \U$18803 ( \19146 , \19144 , \19145 );
xor \U$18804 ( \19147 , \19136 , \19146 );
not \U$18805 ( \19148 , \10251 );
not \U$18806 ( \19149 , \17367 );
or \U$18807 ( \19150 , \19148 , \19149 );
not \U$18808 ( \19151 , RI9872d60_173);
not \U$18809 ( \19152 , \5720 );
or \U$18810 ( \19153 , \19151 , \19152 );
or \U$18811 ( \19154 , \1658 , RI9872d60_173);
nand \U$18812 ( \19155 , \19153 , \19154 );
nand \U$18813 ( \19156 , \19155 , \8802 );
nand \U$18814 ( \19157 , \19150 , \19156 );
xnor \U$18815 ( \19158 , \19147 , \19157 );
and \U$18816 ( \19159 , \7028 , RI98725e0_157);
not \U$18817 ( \19160 , \7028 );
and \U$18818 ( \19161 , \19160 , \6042 );
nor \U$18819 ( \19162 , \19159 , \19161 );
not \U$18820 ( \19163 , \19162 );
or \U$18821 ( \19164 , \19163 , \6048 );
not \U$18822 ( \19165 , \8790 );
or \U$18823 ( \19166 , \17472 , \19165 );
nand \U$18824 ( \19167 , \19164 , \19166 );
not \U$18825 ( \19168 , \17330 );
not \U$18826 ( \19169 , \9670 );
or \U$18827 ( \19170 , \19168 , \19169 );
not \U$18828 ( \19171 , \10486 );
not \U$18829 ( \19172 , RI9872bf8_170);
not \U$18830 ( \19173 , \12295 );
or \U$18831 ( \19174 , \19172 , \19173 );
nand \U$18832 ( \19175 , \1370 , \9185 );
nand \U$18833 ( \19176 , \19174 , \19175 );
nand \U$18834 ( \19177 , \19171 , \19176 );
nand \U$18835 ( \19178 , \19170 , \19177 );
xor \U$18836 ( \19179 , \19167 , \19178 );
and \U$18837 ( \19180 , RI9873288_184, \2982 );
not \U$18838 ( \19181 , RI9873288_184);
not \U$18839 ( \19182 , \1393 );
and \U$18840 ( \19183 , \19181 , \19182 );
nor \U$18841 ( \19184 , \19180 , \19183 );
not \U$18842 ( \19185 , \19184 );
not \U$18843 ( \19186 , \17528 );
or \U$18844 ( \19187 , \19185 , \19186 );
not \U$18845 ( \19188 , \17655 );
not \U$18846 ( \19189 , \17545 );
or \U$18847 ( \19190 , \19188 , \19189 );
nand \U$18848 ( \19191 , \19187 , \19190 );
xor \U$18849 ( \19192 , \19179 , \19191 );
xor \U$18850 ( \19193 , \19158 , \19192 );
not \U$18851 ( \19194 , \5642 );
not \U$18852 ( \19195 , \18398 );
or \U$18853 ( \19196 , \19194 , \19195 );
and \U$18854 ( \19197 , RI9872568_156, \3569 );
not \U$18855 ( \19198 , RI9872568_156);
and \U$18856 ( \19199 , \19198 , \10699 );
nor \U$18857 ( \19200 , \19197 , \19199 );
nand \U$18858 ( \19201 , \19200 , \7188 );
nand \U$18859 ( \19202 , \19196 , \19201 );
not \U$18860 ( \19203 , \19202 );
not \U$18861 ( \19204 , \6611 );
and \U$18862 ( \19205 , RI98728b0_163, \3860 );
not \U$18863 ( \19206 , RI98728b0_163);
and \U$18864 ( \19207 , \19206 , \9461 );
nor \U$18865 ( \19208 , \19205 , \19207 );
not \U$18866 ( \19209 , \19208 );
or \U$18867 ( \19210 , \19204 , \19209 );
nand \U$18868 ( \19211 , \17484 , \6284 );
nand \U$18869 ( \19212 , \19210 , \19211 );
xor \U$18870 ( \19213 , \19203 , \19212 );
not \U$18871 ( \19214 , \11199 );
not \U$18872 ( \19215 , RI9872f40_177);
not \U$18873 ( \19216 , \6443 );
or \U$18874 ( \19217 , \19215 , \19216 );
not \U$18875 ( \19218 , \6400 );
or \U$18876 ( \19219 , RI9872f40_177, \19218 );
nand \U$18877 ( \19220 , \19217 , \19219 );
not \U$18878 ( \19221 , \19220 );
or \U$18879 ( \19222 , \19214 , \19221 );
nand \U$18880 ( \19223 , \17502 , \9527 );
nand \U$18881 ( \19224 , \19222 , \19223 );
xnor \U$18882 ( \19225 , \19213 , \19224 );
xnor \U$18883 ( \19226 , \19193 , \19225 );
xor \U$18884 ( \19227 , \19128 , \19226 );
xor \U$18885 ( \19228 , \18895 , \19227 );
xnor \U$18886 ( \19229 , \18781 , \19228 );
not \U$18887 ( \19230 , \18563 );
and \U$18888 ( \19231 , \9690 , \1365 );
not \U$18889 ( \19232 , \9690 );
and \U$18890 ( \19233 , \19232 , \1369 );
or \U$18891 ( \19234 , \19231 , \19233 );
not \U$18892 ( \19235 , \19234 );
or \U$18893 ( \19236 , \19230 , \19235 );
nand \U$18894 ( \19237 , \17218 , \10332 );
nand \U$18895 ( \19238 , \19236 , \19237 );
not \U$18896 ( \19239 , \19046 );
not \U$18897 ( \19240 , \19041 );
or \U$18898 ( \19241 , \19239 , \19240 );
xor \U$18899 ( \19242 , RI98734e0_189, \1393 );
buf \U$18900 ( \19243 , \19035 );
buf \U$18901 ( \19244 , \19243 );
nand \U$18902 ( \19245 , \19242 , \19244 );
nand \U$18903 ( \19246 , \19241 , \19245 );
xor \U$18904 ( \19247 , \19238 , \19246 );
not \U$18905 ( \19248 , \19247 );
not \U$18906 ( \19249 , \17545 );
not \U$18907 ( \19250 , RI9873288_184);
not \U$18908 ( \19251 , \2492 );
or \U$18909 ( \19252 , \19250 , \19251 );
or \U$18910 ( \19253 , \2492 , RI9873288_184);
nand \U$18911 ( \19254 , \19252 , \19253 );
not \U$18912 ( \19255 , \19254 );
or \U$18913 ( \19256 , \19249 , \19255 );
nand \U$18914 ( \19257 , \17537 , \17528 );
nand \U$18915 ( \19258 , \19256 , \19257 );
not \U$18916 ( \19259 , \19258 );
or \U$18917 ( \19260 , \19248 , \19259 );
nand \U$18918 ( \19261 , \19246 , \19238 );
nand \U$18919 ( \19262 , \19260 , \19261 );
not \U$18920 ( \19263 , \19262 );
not \U$18921 ( \19264 , \18065 );
not \U$18922 ( \19265 , \11691 );
and \U$18923 ( \19266 , \19264 , \19265 );
and \U$18924 ( \19267 , \17286 , \9214 );
nor \U$18925 ( \19268 , \19266 , \19267 );
not \U$18926 ( \19269 , \19268 );
not \U$18927 ( \19270 , \19269 );
not \U$18928 ( \19271 , \13020 );
not \U$18929 ( \19272 , \18044 );
or \U$18930 ( \19273 , \19271 , \19272 );
nand \U$18931 ( \19274 , \17301 , \17347 );
nand \U$18932 ( \19275 , \19273 , \19274 );
not \U$18933 ( \19276 , \19275 );
or \U$18934 ( \19277 , \19270 , \19276 );
or \U$18935 ( \19278 , \19275 , \19269 );
not \U$18936 ( \19279 , \17371 );
not \U$18937 ( \19280 , \18070 );
or \U$18938 ( \19281 , \19279 , \19280 );
buf \U$18939 ( \19282 , \17263 );
nand \U$18940 ( \19283 , \17257 , \19282 );
nand \U$18941 ( \19284 , \19281 , \19283 );
nand \U$18942 ( \19285 , \19278 , \19284 );
nand \U$18943 ( \19286 , \19277 , \19285 );
xor \U$18944 ( \19287 , \19263 , \19286 );
not \U$18945 ( \19288 , \16894 );
not \U$18946 ( \19289 , \7338 );
not \U$18947 ( \19290 , \19289 );
and \U$18948 ( \19291 , \19288 , \19290 );
not \U$18949 ( \19292 , RI98729a0_165);
not \U$18950 ( \19293 , \11672 );
or \U$18951 ( \19294 , \19292 , \19293 );
or \U$18952 ( \19295 , \14930 , RI98729a0_165);
nand \U$18953 ( \19296 , \19294 , \19295 );
and \U$18954 ( \19297 , \19296 , \7325 );
nor \U$18955 ( \19298 , \19291 , \19297 );
not \U$18956 ( \19299 , \19298 );
not \U$18957 ( \19300 , \19299 );
not \U$18958 ( \19301 , \8028 );
and \U$18959 ( \19302 , RI9872a18_166, \3859 );
not \U$18960 ( \19303 , RI9872a18_166);
not \U$18961 ( \19304 , \3858 );
and \U$18962 ( \19305 , \19303 , \19304 );
or \U$18963 ( \19306 , \19302 , \19305 );
not \U$18964 ( \19307 , \19306 );
or \U$18965 ( \19308 , \19301 , \19307 );
nand \U$18966 ( \19309 , \17518 , \8041 );
nand \U$18967 ( \19310 , \19308 , \19309 );
not \U$18968 ( \19311 , \19310 );
not \U$18969 ( \19312 , \19311 );
not \U$18970 ( \19313 , \9937 );
not \U$18971 ( \19314 , \17562 );
or \U$18972 ( \19315 , \19313 , \19314 );
and \U$18973 ( \19316 , RI9873030_179, \846 );
not \U$18974 ( \19317 , RI9873030_179);
and \U$18975 ( \19318 , \19317 , \16924 );
nor \U$18976 ( \19319 , \19316 , \19318 );
not \U$18977 ( \19320 , \9952 );
not \U$18978 ( \19321 , \19320 );
nand \U$18979 ( \19322 , \19319 , \19321 );
nand \U$18980 ( \19323 , \19315 , \19322 );
not \U$18981 ( \19324 , \19323 );
or \U$18982 ( \19325 , \19312 , \19324 );
or \U$18983 ( \19326 , \19323 , \19311 );
nand \U$18984 ( \19327 , \19325 , \19326 );
not \U$18985 ( \19328 , \19327 );
or \U$18986 ( \19329 , \19300 , \19328 );
nand \U$18987 ( \19330 , \19323 , \19310 );
nand \U$18988 ( \19331 , \19329 , \19330 );
xnor \U$18989 ( \19332 , \19287 , \19331 );
not \U$18990 ( \19333 , \19332 );
not \U$18991 ( \19334 , \19064 );
not \U$18992 ( \19335 , \19066 );
and \U$18993 ( \19336 , \19334 , \19335 );
and \U$18994 ( \19337 , \19064 , \19066 );
nor \U$18995 ( \19338 , \19336 , \19337 );
xor \U$18996 ( \19339 , \19073 , \19338 );
not \U$18997 ( \19340 , \19099 );
not \U$18998 ( \19341 , \19094 );
or \U$18999 ( \19342 , \19340 , \19341 );
or \U$19000 ( \19343 , \19094 , \19099 );
nand \U$19001 ( \19344 , \19342 , \19343 );
not \U$19002 ( \19345 , \19344 );
not \U$19003 ( \19346 , \19105 );
and \U$19004 ( \19347 , \19345 , \19346 );
and \U$19005 ( \19348 , \19344 , \19105 );
nor \U$19006 ( \19349 , \19347 , \19348 );
not \U$19007 ( \19350 , \19349 );
xor \U$19008 ( \19351 , \19339 , \19350 );
xor \U$19009 ( \19352 , \19025 , \19031 );
xor \U$19010 ( \19353 , \19352 , \19048 );
xor \U$19011 ( \19354 , \19351 , \19353 );
not \U$19012 ( \19355 , \19354 );
not \U$19013 ( \19356 , \19243 );
not \U$19014 ( \19357 , \16999 );
not \U$19015 ( \19358 , \1125 );
or \U$19016 ( \19359 , \19357 , \19358 );
not \U$19017 ( \19360 , \2398 );
not \U$19018 ( \19361 , RI98734e0_189);
or \U$19019 ( \19362 , \19360 , \19361 );
nand \U$19020 ( \19363 , \19359 , \19362 );
not \U$19021 ( \19364 , \19363 );
or \U$19022 ( \19365 , \19356 , \19364 );
nand \U$19023 ( \19366 , \19242 , \19046 );
nand \U$19024 ( \19367 , \19365 , \19366 );
not \U$19025 ( \19368 , \9273 );
not \U$19026 ( \19369 , \19234 );
or \U$19027 ( \19370 , \19368 , \19369 );
nand \U$19028 ( \19371 , \18581 , \9686 );
nand \U$19029 ( \19372 , \19370 , \19371 );
or \U$19030 ( \19373 , \19367 , \19372 );
not \U$19031 ( \19374 , \17528 );
not \U$19032 ( \19375 , \19254 );
or \U$19033 ( \19376 , \19374 , \19375 );
nand \U$19034 ( \19377 , \18521 , \17545 );
nand \U$19035 ( \19378 , \19376 , \19377 );
nand \U$19036 ( \19379 , \19373 , \19378 );
nand \U$19037 ( \19380 , \19367 , \19372 );
nand \U$19038 ( \19381 , \19379 , \19380 );
not \U$19039 ( \19382 , \19381 );
buf \U$19040 ( \19383 , \18704 );
nand \U$19041 ( \19384 , \1147 , \19383 );
nand \U$19042 ( \19385 , \13385 , \1158 );
and \U$19043 ( \19386 , \19384 , \19385 , \8679 );
not \U$19044 ( \19387 , \832 );
not \U$19045 ( \19388 , \18715 );
or \U$19046 ( \19389 , \19387 , \19388 );
and \U$19047 ( \19390 , \13921 , \17736 );
not \U$19048 ( \19391 , \13921 );
not \U$19049 ( \19392 , \17736 );
and \U$19050 ( \19393 , \19391 , \19392 );
nor \U$19051 ( \19394 , \19390 , \19393 );
xnor \U$19052 ( \19395 , RI9871d70_139, \19394 );
nand \U$19053 ( \19396 , \19395 , \859 );
nand \U$19054 ( \19397 , \19389 , \19396 );
and \U$19055 ( \19398 , \19386 , \19397 );
not \U$19056 ( \19399 , \19398 );
not \U$19057 ( \19400 , \17704 );
not \U$19058 ( \19401 , \18219 );
or \U$19059 ( \19402 , \19400 , \19401 );
or \U$19060 ( \19403 , \18219 , \17704 );
nand \U$19061 ( \19404 , \19402 , \19403 );
not \U$19062 ( \19405 , \19404 );
not \U$19063 ( \19406 , \1016 );
or \U$19064 ( \19407 , \19405 , \19406 );
nand \U$19065 ( \19408 , \18223 , \1013 );
nand \U$19066 ( \19409 , \19407 , \19408 );
not \U$19067 ( \19410 , \1379 );
not \U$19068 ( \19411 , \17723 );
not \U$19069 ( \19412 , \19411 );
xor \U$19070 ( \19413 , \19412 , RI9871e60_141);
not \U$19071 ( \19414 , \19413 );
or \U$19072 ( \19415 , \19410 , \19414 );
nand \U$19073 ( \19416 , \17914 , \1352 );
nand \U$19074 ( \19417 , \19415 , \19416 );
and \U$19075 ( \19418 , \19409 , \19417 );
not \U$19076 ( \19419 , \19409 );
not \U$19077 ( \19420 , \19417 );
and \U$19078 ( \19421 , \19419 , \19420 );
nor \U$19079 ( \19422 , \19418 , \19421 );
not \U$19080 ( \19423 , \19422 );
or \U$19081 ( \19424 , \19399 , \19423 );
nand \U$19082 ( \19425 , \19417 , \19409 );
nand \U$19083 ( \19426 , \19424 , \19425 );
not \U$19084 ( \19427 , \19426 );
xor \U$19085 ( \19428 , \18231 , \18228 );
xnor \U$19086 ( \19429 , \19428 , \18230 );
nand \U$19087 ( \19430 , \19427 , \19429 );
not \U$19088 ( \19431 , \19430 );
not \U$19089 ( \19432 , \6610 );
not \U$19090 ( \19433 , \17839 );
or \U$19091 ( \19434 , \19432 , \19433 );
nand \U$19092 ( \19435 , \18641 , \6284 );
nand \U$19093 ( \19436 , \19434 , \19435 );
not \U$19094 ( \19437 , \19436 );
or \U$19095 ( \19438 , \19431 , \19437 );
not \U$19096 ( \19439 , \19429 );
nand \U$19097 ( \19440 , \19439 , \19426 );
nand \U$19098 ( \19441 , \19438 , \19440 );
not \U$19099 ( \19442 , \19441 );
xor \U$19100 ( \19443 , \18244 , \18257 );
not \U$19101 ( \19444 , \19443 );
not \U$19102 ( \19445 , \19444 );
or \U$19103 ( \19446 , \19442 , \19445 );
not \U$19104 ( \19447 , \19441 );
nand \U$19105 ( \19448 , \19447 , \19443 );
nand \U$19106 ( \19449 , \19446 , \19448 );
not \U$19107 ( \19450 , \19449 );
or \U$19108 ( \19451 , \19382 , \19450 );
nand \U$19109 ( \19452 , \19443 , \19441 );
nand \U$19110 ( \19453 , \19451 , \19452 );
not \U$19111 ( \19454 , \19453 );
and \U$19112 ( \19455 , \19355 , \19454 );
and \U$19113 ( \19456 , \19354 , \19453 );
nor \U$19114 ( \19457 , \19455 , \19456 );
not \U$19115 ( \19458 , \19457 );
and \U$19116 ( \19459 , \19333 , \19458 );
and \U$19117 ( \19460 , \19332 , \19457 );
nor \U$19118 ( \19461 , \19459 , \19460 );
not \U$19119 ( \19462 , \19461 );
xor \U$19120 ( \19463 , \17841 , \17923 );
not \U$19121 ( \19464 , \19258 );
not \U$19122 ( \19465 , \19247 );
not \U$19123 ( \19466 , \19465 );
or \U$19124 ( \19467 , \19464 , \19466 );
not \U$19125 ( \19468 , \19258 );
nand \U$19126 ( \19469 , \19468 , \19247 );
nand \U$19127 ( \19470 , \19467 , \19469 );
xor \U$19128 ( \19471 , \19463 , \19470 );
xor \U$19129 ( \19472 , \18274 , \18279 );
xor \U$19130 ( \19473 , \19472 , \18286 );
xnor \U$19131 ( \19474 , \19471 , \19473 );
not \U$19132 ( \19475 , \19474 );
not \U$19133 ( \19476 , \19475 );
xor \U$19134 ( \19477 , \19298 , \19311 );
xnor \U$19135 ( \19478 , \19477 , \19323 );
xor \U$19136 ( \19479 , \17137 , \17154 );
xor \U$19137 ( \19480 , \19479 , \17171 );
and \U$19138 ( \19481 , \19478 , \19480 );
not \U$19139 ( \19482 , \19478 );
not \U$19140 ( \19483 , \19480 );
and \U$19141 ( \19484 , \19482 , \19483 );
or \U$19142 ( \19485 , \19481 , \19484 );
xor \U$19143 ( \19486 , \19268 , \19284 );
xor \U$19144 ( \19487 , \19486 , \19275 );
and \U$19145 ( \19488 , \19485 , \19487 );
not \U$19146 ( \19489 , \19485 );
not \U$19147 ( \19490 , \19487 );
and \U$19148 ( \19491 , \19489 , \19490 );
nor \U$19149 ( \19492 , \19488 , \19491 );
not \U$19150 ( \19493 , \19492 );
not \U$19151 ( \19494 , \19493 );
or \U$19152 ( \19495 , \19476 , \19494 );
not \U$19153 ( \19496 , \19474 );
not \U$19154 ( \19497 , \19492 );
or \U$19155 ( \19498 , \19496 , \19497 );
not \U$19156 ( \19499 , \6653 );
not \U$19157 ( \19500 , RI9872310_151);
not \U$19158 ( \19501 , \18110 );
or \U$19159 ( \19502 , \19500 , \19501 );
or \U$19160 ( \19503 , \18110 , RI9872310_151);
nand \U$19161 ( \19504 , \19502 , \19503 );
not \U$19162 ( \19505 , \19504 );
or \U$19163 ( \19506 , \19499 , \19505 );
and \U$19164 ( \19507 , RI9872310_151, \12713 );
not \U$19165 ( \19508 , RI9872310_151);
and \U$19166 ( \19509 , \19508 , \10598 );
nor \U$19167 ( \19510 , \19507 , \19509 );
nand \U$19168 ( \19511 , \19510 , \3170 );
nand \U$19169 ( \19512 , \19506 , \19511 );
not \U$19170 ( \19513 , \1352 );
not \U$19171 ( \19514 , \19413 );
or \U$19172 ( \19515 , \19513 , \19514 );
and \U$19173 ( \19516 , RI9871e60_141, \18216 );
not \U$19174 ( \19517 , RI9871e60_141);
buf \U$19175 ( \19518 , \16994 );
buf \U$19176 ( \19519 , \19518 );
and \U$19177 ( \19520 , \19517 , \19519 );
or \U$19178 ( \19521 , \19516 , \19520 );
not \U$19179 ( \19522 , \19521 );
or \U$19180 ( \19523 , \19522 , \9922 );
nand \U$19181 ( \19524 , \19515 , \19523 );
not \U$19182 ( \19525 , \19524 );
not \U$19183 ( \19526 , \8678 );
not \U$19184 ( \19527 , \18705 );
and \U$19185 ( \19528 , \19526 , \19527 );
nor \U$19186 ( \19529 , \19528 , \18707 );
not \U$19187 ( \19530 , \19529 );
not \U$19188 ( \19531 , \9429 );
or \U$19189 ( \19532 , \19530 , \19531 );
not \U$19190 ( \19533 , \1219 );
nand \U$19191 ( \19534 , \19533 , \18723 );
nand \U$19192 ( \19535 , \19532 , \19534 );
not \U$19193 ( \19536 , \17686 );
not \U$19194 ( \19537 , \17856 );
and \U$19195 ( \19538 , \19536 , \19537 );
not \U$19196 ( \19539 , \17854 );
and \U$19197 ( \19540 , \19539 , \17856 );
nor \U$19198 ( \19541 , \19538 , \19540 );
buf \U$19199 ( \19542 , \19541 );
not \U$19200 ( \19543 , \19542 );
not \U$19201 ( \19544 , \19543 );
not \U$19202 ( \19545 , \19544 );
not \U$19203 ( \19546 , \1157 );
or \U$19204 ( \19547 , \19545 , \19546 );
or \U$19205 ( \19548 , \1042 , \19544 );
nand \U$19206 ( \19549 , \19547 , \19548 );
not \U$19207 ( \19550 , \19549 );
not \U$19208 ( \19551 , \1017 );
or \U$19209 ( \19552 , \19550 , \19551 );
nand \U$19210 ( \19553 , \1013 , \19404 );
nand \U$19211 ( \19554 , \19552 , \19553 );
or \U$19212 ( \19555 , \19535 , \19554 );
not \U$19213 ( \19556 , \19555 );
or \U$19214 ( \19557 , \19525 , \19556 );
nand \U$19215 ( \19558 , \19535 , \19554 );
nand \U$19216 ( \19559 , \19557 , \19558 );
xnor \U$19217 ( \19560 , \19512 , \19559 );
not \U$19218 ( \19561 , \3467 );
not \U$19219 ( \19562 , RI98726d0_159);
not \U$19220 ( \19563 , \8334 );
or \U$19221 ( \19564 , \19562 , \19563 );
or \U$19222 ( \19565 , \9895 , RI98726d0_159);
nand \U$19223 ( \19566 , \19564 , \19565 );
not \U$19224 ( \19567 , \19566 );
or \U$19225 ( \19568 , \19561 , \19567 );
not \U$19226 ( \19569 , RI98726d0_159);
not \U$19227 ( \19570 , \8074 );
or \U$19228 ( \19571 , \19569 , \19570 );
or \U$19229 ( \19572 , \8074 , RI98726d0_159);
nand \U$19230 ( \19573 , \19571 , \19572 );
nand \U$19231 ( \19574 , \19573 , \13409 );
nand \U$19232 ( \19575 , \19568 , \19574 );
or \U$19233 ( \19576 , \19560 , \19575 );
nand \U$19234 ( \19577 , \19560 , \19575 );
not \U$19235 ( \19578 , \875 );
and \U$19236 ( \19579 , \17783 , \919 );
not \U$19237 ( \19580 , \17783 );
and \U$19238 ( \19581 , \19580 , RI9872130_147);
nor \U$19239 ( \19582 , \19579 , \19581 );
not \U$19240 ( \19583 , \19582 );
or \U$19241 ( \19584 , \19578 , \19583 );
not \U$19242 ( \19585 , RI9872130_147);
not \U$19243 ( \19586 , \13279 );
not \U$19244 ( \19587 , \13278 );
and \U$19245 ( \19588 , \19586 , \19587 );
and \U$19246 ( \19589 , \13279 , \13278 );
nor \U$19247 ( \19590 , \19588 , \19589 );
buf \U$19248 ( \19591 , \19590 );
not \U$19249 ( \19592 , \19591 );
or \U$19250 ( \19593 , \19585 , \19592 );
not \U$19251 ( \19594 , \19590 );
not \U$19252 ( \19595 , \19594 );
or \U$19253 ( \19596 , \19595 , RI9872130_147);
nand \U$19254 ( \19597 , \19593 , \19596 );
nand \U$19255 ( \19598 , \19597 , \924 );
nand \U$19256 ( \19599 , \19584 , \19598 );
not \U$19257 ( \19600 , \1500 );
and \U$19258 ( \19601 , RI9871c80_137, \13268 );
not \U$19259 ( \19602 , RI9871c80_137);
and \U$19260 ( \19603 , \19602 , \17081 );
or \U$19261 ( \19604 , \19601 , \19603 );
not \U$19262 ( \19605 , \19604 );
or \U$19263 ( \19606 , \19600 , \19605 );
not \U$19264 ( \19607 , \18151 );
xor \U$19265 ( \19608 , RI9871c80_137, \19607 );
nand \U$19266 ( \19609 , \19608 , \1518 );
nand \U$19267 ( \19610 , \19606 , \19609 );
xor \U$19268 ( \19611 , \19599 , \19610 );
not \U$19269 ( \19612 , \1455 );
not \U$19270 ( \19613 , RI9871c08_136);
not \U$19271 ( \19614 , \9113 );
or \U$19272 ( \19615 , \19613 , \19614 );
or \U$19273 ( \19616 , \9113 , RI9871c08_136);
nand \U$19274 ( \19617 , \19615 , \19616 );
not \U$19275 ( \19618 , \19617 );
or \U$19276 ( \19619 , \19612 , \19618 );
nand \U$19277 ( \19620 , \18605 , \1429 );
nand \U$19278 ( \19621 , \19619 , \19620 );
xor \U$19279 ( \19622 , \19611 , \19621 );
not \U$19280 ( \19623 , \19622 );
nand \U$19281 ( \19624 , \19576 , \19577 , \19623 );
not \U$19282 ( \19625 , \19624 );
not \U$19283 ( \19626 , \5653 );
not \U$19284 ( \19627 , \18492 );
or \U$19285 ( \19628 , \19626 , \19627 );
and \U$19286 ( \19629 , RI9872568_156, \6059 );
not \U$19287 ( \19630 , RI9872568_156);
and \U$19288 ( \19631 , \19630 , \5766 );
or \U$19289 ( \19632 , \19629 , \19631 );
nand \U$19290 ( \19633 , \19632 , \6063 );
nand \U$19291 ( \19634 , \19628 , \19633 );
not \U$19292 ( \19635 , \19634 );
not \U$19293 ( \19636 , \17528 );
not \U$19294 ( \19637 , \18514 );
or \U$19295 ( \19638 , \19636 , \19637 );
not \U$19296 ( \19639 , \6585 );
xor \U$19297 ( \19640 , RI9873288_184, \19639 );
buf \U$19298 ( \19641 , \17543 );
nand \U$19299 ( \19642 , \19640 , \19641 );
nand \U$19300 ( \19643 , \19638 , \19642 );
not \U$19301 ( \19644 , \19643 );
or \U$19302 ( \19645 , \19635 , \19644 );
not \U$19303 ( \19646 , \13214 );
not \U$19304 ( \19647 , \18536 );
or \U$19305 ( \19648 , \19646 , \19647 );
not \U$19306 ( \19649 , \9529 );
not \U$19307 ( \19650 , \1061 );
or \U$19308 ( \19651 , \19649 , \19650 );
or \U$19309 ( \19652 , \1061 , \8732 );
nand \U$19310 ( \19653 , \19651 , \19652 );
nand \U$19311 ( \19654 , \19653 , \9526 );
nand \U$19312 ( \19655 , \19648 , \19654 );
not \U$19313 ( \19656 , \19655 );
nand \U$19314 ( \19657 , \19645 , \19656 );
not \U$19315 ( \19658 , \19643 );
not \U$19316 ( \19659 , \19634 );
nand \U$19317 ( \19660 , \19658 , \19659 );
and \U$19318 ( \19661 , \19657 , \19660 );
not \U$19319 ( \19662 , \19661 );
or \U$19320 ( \19663 , \19625 , \19662 );
xnor \U$19321 ( \19664 , \19575 , \19560 );
nand \U$19322 ( \19665 , \19664 , \19622 );
nand \U$19323 ( \19666 , \19663 , \19665 );
not \U$19324 ( \19667 , \19666 );
not \U$19325 ( \19668 , \924 );
not \U$19326 ( \19669 , \18147 );
or \U$19327 ( \19670 , \19668 , \19669 );
nand \U$19328 ( \19671 , \19597 , \876 );
nand \U$19329 ( \19672 , \19670 , \19671 );
not \U$19330 ( \19673 , \1518 );
not \U$19331 ( \19674 , \17772 );
or \U$19332 ( \19675 , \19673 , \19674 );
nand \U$19333 ( \19676 , \19608 , \1500 );
nand \U$19334 ( \19677 , \19675 , \19676 );
xor \U$19335 ( \19678 , \19672 , \19677 );
xor \U$19336 ( \19679 , \17887 , \17917 );
xor \U$19337 ( \19680 , \19679 , \17903 );
xor \U$19338 ( \19681 , \19678 , \19680 );
not \U$19339 ( \19682 , \4084 );
not \U$19340 ( \19683 , \18177 );
or \U$19341 ( \19684 , \19682 , \19683 );
not \U$19342 ( \19685 , RI98725e0_157);
not \U$19343 ( \19686 , \10582 );
or \U$19344 ( \19687 , \19685 , \19686 );
or \U$19345 ( \19688 , \8081 , RI98725e0_157);
nand \U$19346 ( \19689 , \19687 , \19688 );
nand \U$19347 ( \19690 , \19689 , \18171 );
nand \U$19348 ( \19691 , \19684 , \19690 );
xnor \U$19349 ( \19692 , \19681 , \19691 );
not \U$19350 ( \19693 , \793 );
not \U$19351 ( \19694 , RI98719b0_131);
not \U$19352 ( \19695 , \8554 );
or \U$19353 ( \19696 , \19694 , \19695 );
or \U$19354 ( \19697 , \8555 , RI98719b0_131);
nand \U$19355 ( \19698 , \19696 , \19697 );
not \U$19356 ( \19699 , \19698 );
or \U$19357 ( \19700 , \19693 , \19699 );
not \U$19358 ( \19701 , \8575 );
and \U$19359 ( \19702 , RI98719b0_131, \19701 );
not \U$19360 ( \19703 , RI98719b0_131);
and \U$19361 ( \19704 , \19703 , \8580 );
or \U$19362 ( \19705 , \19702 , \19704 );
nand \U$19363 ( \19706 , \19705 , \796 );
nand \U$19364 ( \19707 , \19700 , \19706 );
not \U$19365 ( \19708 , \2087 );
and \U$19366 ( \19709 , RI9871aa0_133, \8668 );
not \U$19367 ( \19710 , RI9871aa0_133);
and \U$19368 ( \19711 , \19710 , \9881 );
or \U$19369 ( \19712 , \19709 , \19711 );
not \U$19370 ( \19713 , \19712 );
or \U$19371 ( \19714 , \19708 , \19713 );
not \U$19372 ( \19715 , \11406 );
and \U$19373 ( \19716 , RI9871aa0_133, \19715 );
not \U$19374 ( \19717 , RI9871aa0_133);
and \U$19375 ( \19718 , \19717 , \8650 );
nor \U$19376 ( \19719 , \19716 , \19718 );
nand \U$19377 ( \19720 , \19719 , \2072 );
nand \U$19378 ( \19721 , \19714 , \19720 );
xor \U$19379 ( \19722 , \19707 , \19721 );
not \U$19380 ( \19723 , \5034 );
and \U$19381 ( \19724 , RI9872478_154, \11435 );
not \U$19382 ( \19725 , RI9872478_154);
and \U$19383 ( \19726 , \19725 , \6303 );
or \U$19384 ( \19727 , \19724 , \19726 );
not \U$19385 ( \19728 , \19727 );
or \U$19386 ( \19729 , \19723 , \19728 );
nand \U$19387 ( \19730 , \17974 , \5796 );
nand \U$19388 ( \19731 , \19729 , \19730 );
and \U$19389 ( \19732 , \19722 , \19731 );
and \U$19390 ( \19733 , \19707 , \19721 );
or \U$19391 ( \19734 , \19732 , \19733 );
xnor \U$19392 ( \19735 , \19692 , \19734 );
not \U$19393 ( \19736 , \19735 );
xor \U$19394 ( \19737 , \19707 , \19721 );
xor \U$19395 ( \19738 , \19737 , \19731 );
not \U$19396 ( \19739 , \1292 );
not \U$19397 ( \19740 , RI9871b18_134);
not \U$19398 ( \19741 , \13388 );
or \U$19399 ( \19742 , \19740 , \19741 );
nand \U$19400 ( \19743 , \13387 , \1283 );
nand \U$19401 ( \19744 , \19742 , \19743 );
not \U$19402 ( \19745 , \19744 );
or \U$19403 ( \19746 , \19739 , \19745 );
nand \U$19404 ( \19747 , \17893 , \1323 );
nand \U$19405 ( \19748 , \19746 , \19747 );
not \U$19406 ( \19749 , \4101 );
and \U$19407 ( \19750 , RI98725e0_157, \7466 );
not \U$19408 ( \19751 , RI98725e0_157);
not \U$19409 ( \19752 , \13824 );
and \U$19410 ( \19753 , \19751 , \19752 );
or \U$19411 ( \19754 , \19750 , \19753 );
not \U$19412 ( \19755 , \19754 );
or \U$19413 ( \19756 , \19749 , \19755 );
nand \U$19414 ( \19757 , \19689 , \4084 );
nand \U$19415 ( \19758 , \19756 , \19757 );
xor \U$19416 ( \19759 , \19748 , \19758 );
not \U$19417 ( \19760 , \4919 );
xor \U$19418 ( \19761 , RI9872388_152, \6528 );
not \U$19419 ( \19762 , \19761 );
or \U$19420 ( \19763 , \19760 , \19762 );
not \U$19421 ( \19764 , RI9872388_152);
not \U$19422 ( \19765 , \12805 );
or \U$19423 ( \19766 , \19764 , \19765 );
or \U$19424 ( \19767 , \8053 , RI9872388_152);
nand \U$19425 ( \19768 , \19766 , \19767 );
nand \U$19426 ( \19769 , \19768 , \4923 );
nand \U$19427 ( \19770 , \19763 , \19769 );
buf \U$19428 ( \19771 , \19770 );
xor \U$19429 ( \19772 , \19759 , \19771 );
xor \U$19430 ( \19773 , \19738 , \19772 );
not \U$19431 ( \19774 , \9249 );
not \U$19432 ( \19775 , RI9872bf8_170);
and \U$19433 ( \19776 , \2947 , \19775 );
not \U$19434 ( \19777 , \2947 );
and \U$19435 ( \19778 , \19777 , RI9872bf8_170);
nor \U$19436 ( \19779 , \19776 , \19778 );
not \U$19437 ( \19780 , \19779 );
or \U$19438 ( \19781 , \19774 , \19780 );
nand \U$19439 ( \19782 , \18457 , \9668 );
nand \U$19440 ( \19783 , \19781 , \19782 );
not \U$19441 ( \19784 , \19783 );
and \U$19442 ( \19785 , RI9872d60_173, \1190 );
not \U$19443 ( \19786 , RI9872d60_173);
and \U$19444 ( \19787 , \19786 , \3395 );
or \U$19445 ( \19788 , \19785 , \19787 );
not \U$19446 ( \19789 , \19788 );
not \U$19447 ( \19790 , \10624 );
or \U$19448 ( \19791 , \19789 , \19790 );
and \U$19449 ( \19792 , RI9872d60_173, \6382 );
not \U$19450 ( \19793 , RI9872d60_173);
and \U$19451 ( \19794 , \19793 , \1485 );
nor \U$19452 ( \19795 , \19792 , \19794 );
nand \U$19453 ( \19796 , \19795 , \10251 );
nand \U$19454 ( \19797 , \19791 , \19796 );
not \U$19455 ( \19798 , \19797 );
or \U$19456 ( \19799 , \19784 , \19798 );
and \U$19457 ( \19800 , \19788 , \10624 );
and \U$19458 ( \19801 , \19795 , \9312 );
nor \U$19459 ( \19802 , \19800 , \19801 , \19783 );
not \U$19460 ( \19803 , \19802 );
not \U$19461 ( \19804 , \17234 );
and \U$19462 ( \19805 , RI9873210_183, \892 );
not \U$19463 ( \19806 , RI9873210_183);
and \U$19464 ( \19807 , \19806 , \13169 );
or \U$19465 ( \19808 , \19805 , \19807 );
not \U$19466 ( \19809 , \19808 );
or \U$19467 ( \19810 , \19804 , \19809 );
not \U$19468 ( \19811 , RI9873210_183);
not \U$19469 ( \19812 , \820 );
or \U$19470 ( \19813 , \19811 , \19812 );
or \U$19471 ( \19814 , \820 , RI9873210_183);
nand \U$19472 ( \19815 , \19813 , \19814 );
nand \U$19473 ( \19816 , \19815 , \13476 );
nand \U$19474 ( \19817 , \19810 , \19816 );
nand \U$19475 ( \19818 , \19803 , \19817 );
nand \U$19476 ( \19819 , \19799 , \19818 );
and \U$19477 ( \19820 , \19773 , \19819 );
and \U$19478 ( \19821 , \19738 , \19772 );
or \U$19479 ( \19822 , \19820 , \19821 );
not \U$19480 ( \19823 , \19822 );
or \U$19481 ( \19824 , \19736 , \19823 );
or \U$19482 ( \19825 , \19822 , \19735 );
nand \U$19483 ( \19826 , \19824 , \19825 );
not \U$19484 ( \19827 , \19826 );
or \U$19485 ( \19828 , \19667 , \19827 );
not \U$19486 ( \19829 , \19735 );
nand \U$19487 ( \19830 , \19829 , \19822 );
nand \U$19488 ( \19831 , \19828 , \19830 );
nand \U$19489 ( \19832 , \19498 , \19831 );
nand \U$19490 ( \19833 , \19495 , \19832 );
not \U$19491 ( \19834 , \19833 );
or \U$19492 ( \19835 , \19462 , \19834 );
or \U$19493 ( \19836 , \19833 , \19461 );
nand \U$19494 ( \19837 , \19835 , \19836 );
and \U$19495 ( \19838 , \18443 , \18440 );
not \U$19496 ( \19839 , \18443 );
and \U$19497 ( \19840 , \19839 , \18441 );
nor \U$19498 ( \19841 , \19838 , \19840 );
xnor \U$19499 ( \19842 , \18759 , \19841 );
nand \U$19500 ( \19843 , \19837 , \19842 );
not \U$19501 ( \19844 , \19461 );
nand \U$19502 ( \19845 , \19844 , \19833 );
and \U$19503 ( \19846 , \19843 , \19845 );
not \U$19504 ( \19847 , \19463 );
not \U$19505 ( \19848 , \19470 );
or \U$19506 ( \19849 , \19847 , \19848 );
or \U$19507 ( \19850 , \19470 , \19463 );
nand \U$19508 ( \19851 , \19850 , \19473 );
nand \U$19509 ( \19852 , \19849 , \19851 );
buf \U$19510 ( \19853 , \19480 );
not \U$19511 ( \19854 , \19853 );
not \U$19512 ( \19855 , \19490 );
or \U$19513 ( \19856 , \19854 , \19855 );
not \U$19514 ( \19857 , \19483 );
not \U$19515 ( \19858 , \19487 );
or \U$19516 ( \19859 , \19857 , \19858 );
not \U$19517 ( \19860 , \19478 );
nand \U$19518 ( \19861 , \19859 , \19860 );
nand \U$19519 ( \19862 , \19856 , \19861 );
xor \U$19520 ( \19863 , \19852 , \19862 );
xor \U$19521 ( \19864 , \17061 , \17175 );
xor \U$19522 ( \19865 , \19863 , \19864 );
not \U$19523 ( \19866 , \19865 );
xor \U$19524 ( \19867 , \18087 , \18372 );
not \U$19525 ( \19868 , \19867 );
xor \U$19526 ( \19869 , \18068 , \18053 );
xor \U$19527 ( \19870 , \19869 , \18081 );
not \U$19528 ( \19871 , \19870 );
not \U$19529 ( \19872 , \18034 );
not \U$19530 ( \19873 , \18007 );
not \U$19531 ( \19874 , \19873 );
and \U$19532 ( \19875 , \19872 , \19874 );
and \U$19533 ( \19876 , \18034 , \19873 );
nor \U$19534 ( \19877 , \19875 , \19876 );
not \U$19535 ( \19878 , \19877 );
or \U$19536 ( \19879 , \19871 , \19878 );
not \U$19537 ( \19880 , \9072 );
not \U$19538 ( \19881 , \19306 );
or \U$19539 ( \19882 , \19880 , \19881 );
nand \U$19540 ( \19883 , \18687 , \8028 );
nand \U$19541 ( \19884 , \19882 , \19883 );
not \U$19542 ( \19885 , \7325 );
not \U$19543 ( \19886 , \18651 );
or \U$19544 ( \19887 , \19885 , \19886 );
nand \U$19545 ( \19888 , \19296 , \7338 );
nand \U$19546 ( \19889 , \19887 , \19888 );
xor \U$19547 ( \19890 , \19884 , \19889 );
nand \U$19548 ( \19891 , \19319 , \9937 );
nand \U$19549 ( \19892 , \18662 , \9952 );
nand \U$19550 ( \19893 , \19891 , \19892 );
xor \U$19551 ( \19894 , \19890 , \19893 );
nand \U$19552 ( \19895 , \19879 , \19894 );
not \U$19553 ( \19896 , \19870 );
not \U$19554 ( \19897 , \19877 );
nand \U$19555 ( \19898 , \19896 , \19897 );
and \U$19556 ( \19899 , \19449 , \19381 );
not \U$19557 ( \19900 , \19449 );
not \U$19558 ( \19901 , \19381 );
and \U$19559 ( \19902 , \19900 , \19901 );
or \U$19560 ( \19903 , \19899 , \19902 );
nand \U$19561 ( \19904 , \19895 , \19898 , \19903 );
xor \U$19562 ( \19905 , \19429 , \19426 );
xnor \U$19563 ( \19906 , \19436 , \19905 );
not \U$19564 ( \19907 , \17961 );
not \U$19565 ( \19908 , \19907 );
not \U$19566 ( \19909 , \17992 );
or \U$19567 ( \19910 , \19908 , \19909 );
or \U$19568 ( \19911 , \17992 , \19907 );
nand \U$19569 ( \19912 , \19910 , \19911 );
xor \U$19570 ( \19913 , \19906 , \19912 );
xor \U$19571 ( \19914 , \19372 , \19367 );
xor \U$19572 ( \19915 , \19914 , \19378 );
and \U$19573 ( \19916 , \19913 , \19915 );
and \U$19574 ( \19917 , \19906 , \19912 );
or \U$19575 ( \19918 , \19916 , \19917 );
nand \U$19576 ( \19919 , \19904 , \19918 );
not \U$19577 ( \19920 , \19903 );
nand \U$19578 ( \19921 , \19895 , \19898 );
nand \U$19579 ( \19922 , \19920 , \19921 );
and \U$19580 ( \19923 , \19919 , \19922 );
not \U$19581 ( \19924 , \19923 );
or \U$19582 ( \19925 , \19868 , \19924 );
or \U$19583 ( \19926 , \19923 , \19867 );
nand \U$19584 ( \19927 , \19925 , \19926 );
not \U$19585 ( \19928 , \19927 );
or \U$19586 ( \19929 , \19866 , \19928 );
not \U$19587 ( \19930 , \19923 );
nand \U$19588 ( \19931 , \19930 , \19867 );
nand \U$19589 ( \19932 , \19929 , \19931 );
not \U$19590 ( \19933 , \19932 );
and \U$19591 ( \19934 , \19846 , \19933 );
not \U$19592 ( \19935 , \19846 );
and \U$19593 ( \19936 , \19935 , \19932 );
nor \U$19594 ( \19937 , \19934 , \19936 );
xor \U$19595 ( \19938 , \18770 , \18437 );
xor \U$19596 ( \19939 , \19938 , \18765 );
xor \U$19597 ( \19940 , \19937 , \19939 );
not \U$19598 ( \19941 , \19940 );
xor \U$19599 ( \19942 , \17059 , \17179 );
xor \U$19600 ( \19943 , \19942 , \17319 );
not \U$19601 ( \19944 , \19943 );
not \U$19602 ( \19945 , \19457 );
not \U$19603 ( \19946 , \19945 );
not \U$19604 ( \19947 , \19332 );
or \U$19605 ( \19948 , \19946 , \19947 );
not \U$19606 ( \19949 , \19354 );
nand \U$19607 ( \19950 , \19949 , \19453 );
nand \U$19608 ( \19951 , \19948 , \19950 );
not \U$19609 ( \19952 , \19951 );
and \U$19610 ( \19953 , \19863 , \19864 );
and \U$19611 ( \19954 , \19852 , \19862 );
nor \U$19612 ( \19955 , \19953 , \19954 );
not \U$19613 ( \19956 , \19955 );
or \U$19614 ( \19957 , \19952 , \19956 );
or \U$19615 ( \19958 , \19955 , \19951 );
nand \U$19616 ( \19959 , \19957 , \19958 );
not \U$19617 ( \19960 , \19959 );
not \U$19618 ( \19961 , \19960 );
or \U$19619 ( \19962 , \19944 , \19961 );
not \U$19620 ( \19963 , \19943 );
nand \U$19621 ( \19964 , \19963 , \19959 );
nand \U$19622 ( \19965 , \19962 , \19964 );
not \U$19623 ( \19966 , \19087 );
and \U$19624 ( \19967 , \19108 , \19079 );
not \U$19625 ( \19968 , \19108 );
and \U$19626 ( \19969 , \19968 , \19078 );
nor \U$19627 ( \19970 , \19967 , \19969 );
not \U$19628 ( \19971 , \19970 );
and \U$19629 ( \19972 , \19966 , \19971 );
and \U$19630 ( \19973 , \19087 , \19970 );
nor \U$19631 ( \19974 , \19972 , \19973 );
not \U$19632 ( \19975 , \19053 );
not \U$19633 ( \19976 , \19018 );
and \U$19634 ( \19977 , \19975 , \19976 );
and \U$19635 ( \19978 , \19053 , \19018 );
nor \U$19636 ( \19979 , \19977 , \19978 );
not \U$19637 ( \19980 , \19979 );
not \U$19638 ( \19981 , \19980 );
nand \U$19639 ( \19982 , \19349 , \19339 );
not \U$19640 ( \19983 , \19982 );
not \U$19641 ( \19984 , \19353 );
or \U$19642 ( \19985 , \19983 , \19984 );
not \U$19643 ( \19986 , \19339 );
nand \U$19644 ( \19987 , \19986 , \19350 );
nand \U$19645 ( \19988 , \19985 , \19987 );
not \U$19646 ( \19989 , \19988 );
not \U$19647 ( \19990 , \19989 );
or \U$19648 ( \19991 , \19981 , \19990 );
nand \U$19649 ( \19992 , \19979 , \19988 );
nand \U$19650 ( \19993 , \19991 , \19992 );
not \U$19651 ( \19994 , \19993 );
xor \U$19652 ( \19995 , \19974 , \19994 );
xor \U$19653 ( \19996 , \18334 , \18316 );
xnor \U$19654 ( \19997 , \19996 , \18299 );
not \U$19655 ( \19998 , \19997 );
not \U$19656 ( \19999 , \18122 );
not \U$19657 ( \20000 , \18136 );
not \U$19658 ( \20001 , \18103 );
or \U$19659 ( \20002 , \20000 , \20001 );
or \U$19660 ( \20003 , \18103 , \18136 );
nand \U$19661 ( \20004 , \20002 , \20003 );
not \U$19662 ( \20005 , \20004 );
or \U$19663 ( \20006 , \19999 , \20005 );
or \U$19664 ( \20007 , \20004 , \18122 );
nand \U$19665 ( \20008 , \20006 , \20007 );
not \U$19666 ( \20009 , \20008 );
or \U$19667 ( \20010 , \19998 , \20009 );
xor \U$19668 ( \20011 , \19884 , \19889 );
and \U$19669 ( \20012 , \20011 , \19893 );
and \U$19670 ( \20013 , \19884 , \19889 );
or \U$19671 ( \20014 , \20012 , \20013 );
nand \U$19672 ( \20015 , \20010 , \20014 );
not \U$19673 ( \20016 , \20008 );
not \U$19674 ( \20017 , \19997 );
nand \U$19675 ( \20018 , \20016 , \20017 );
and \U$19676 ( \20019 , \20015 , \20018 );
buf \U$19677 ( \20020 , \19678 );
not \U$19678 ( \20021 , \20020 );
not \U$19679 ( \20022 , \19691 );
or \U$19680 ( \20023 , \20021 , \20022 );
nand \U$19681 ( \20024 , \19677 , \19672 );
nand \U$19682 ( \20025 , \20023 , \20024 );
not \U$19683 ( \20026 , \20025 );
not \U$19684 ( \20027 , \796 );
not \U$19685 ( \20028 , \18294 );
or \U$19686 ( \20029 , \20027 , \20028 );
nand \U$19687 ( \20030 , \19705 , \791 );
nand \U$19688 ( \20031 , \20029 , \20030 );
not \U$19689 ( \20032 , \20031 );
not \U$19690 ( \20033 , \2087 );
not \U$19691 ( \20034 , \18113 );
or \U$19692 ( \20035 , \20033 , \20034 );
nand \U$19693 ( \20036 , \19712 , \2072 );
nand \U$19694 ( \20037 , \20035 , \20036 );
not \U$19695 ( \20038 , \20037 );
or \U$19696 ( \20039 , \20032 , \20038 );
or \U$19697 ( \20040 , \20037 , \20031 );
not \U$19698 ( \20041 , \3170 );
not \U$19699 ( \20042 , \18100 );
or \U$19700 ( \20043 , \20041 , \20042 );
nand \U$19701 ( \20044 , \19510 , \13033 );
nand \U$19702 ( \20045 , \20043 , \20044 );
nand \U$19703 ( \20046 , \20040 , \20045 );
nand \U$19704 ( \20047 , \20039 , \20046 );
not \U$19705 ( \20048 , \20047 );
or \U$19706 ( \20049 , \20026 , \20048 );
not \U$19707 ( \20050 , \20025 );
not \U$19708 ( \20051 , \20050 );
not \U$19709 ( \20052 , \20047 );
not \U$19710 ( \20053 , \20052 );
or \U$19711 ( \20054 , \20051 , \20053 );
and \U$19712 ( \20055 , \19566 , \13409 );
and \U$19713 ( \20056 , \18132 , \3467 );
nor \U$19714 ( \20057 , \20055 , \20056 );
not \U$19715 ( \20058 , \20057 );
not \U$19716 ( \20059 , \20058 );
not \U$19717 ( \20060 , \5047 );
not \U$19718 ( \20061 , \18253 );
or \U$19719 ( \20062 , \20060 , \20061 );
nand \U$19720 ( \20063 , \19768 , \4919 );
nand \U$19721 ( \20064 , \20062 , \20063 );
not \U$19722 ( \20065 , \20064 );
not \U$19723 ( \20066 , \18719 );
not \U$19724 ( \20067 , \18707 );
not \U$19725 ( \20068 , \20067 );
not \U$19726 ( \20069 , \18728 );
or \U$19727 ( \20070 , \20068 , \20069 );
or \U$19728 ( \20071 , \18728 , \20067 );
nand \U$19729 ( \20072 , \20070 , \20071 );
not \U$19730 ( \20073 , \20072 );
or \U$19731 ( \20074 , \20066 , \20073 );
nand \U$19732 ( \20075 , \18728 , \18707 );
nand \U$19733 ( \20076 , \20074 , \20075 );
not \U$19734 ( \20077 , \20076 );
not \U$19735 ( \20078 , \20077 );
or \U$19736 ( \20079 , \20065 , \20078 );
or \U$19737 ( \20080 , \20064 , \20077 );
nand \U$19738 ( \20081 , \20079 , \20080 );
not \U$19739 ( \20082 , \20081 );
or \U$19740 ( \20083 , \20059 , \20082 );
not \U$19741 ( \20084 , \20064 );
not \U$19742 ( \20085 , \20084 );
nand \U$19743 ( \20086 , \20085 , \20076 );
nand \U$19744 ( \20087 , \20083 , \20086 );
nand \U$19745 ( \20088 , \20054 , \20087 );
nand \U$19746 ( \20089 , \20049 , \20088 );
not \U$19747 ( \20090 , \20089 );
xor \U$19748 ( \20091 , \20019 , \20090 );
xor \U$19749 ( \20092 , \18592 , \18623 );
and \U$19750 ( \20093 , \20092 , \18597 );
and \U$19751 ( \20094 , \18592 , \18623 );
nor \U$19752 ( \20095 , \20093 , \20094 );
and \U$19753 ( \20096 , \20091 , \20095 );
and \U$19754 ( \20097 , \20019 , \20090 );
or \U$19755 ( \20098 , \20096 , \20097 );
xnor \U$19756 ( \20099 , \19995 , \20098 );
not \U$19757 ( \20100 , \18370 );
not \U$19758 ( \20101 , \18289 );
or \U$19759 ( \20102 , \20100 , \20101 );
nand \U$19760 ( \20103 , \18337 , \18369 );
nand \U$19761 ( \20104 , \20102 , \20103 );
not \U$19762 ( \20105 , \20104 );
not \U$19763 ( \20106 , \20105 );
not \U$19764 ( \20107 , \18139 );
not \U$19765 ( \20108 , \18265 );
or \U$19766 ( \20109 , \20107 , \20108 );
nand \U$19767 ( \20110 , \18264 , \18185 );
nand \U$19768 ( \20111 , \20109 , \20110 );
not \U$19769 ( \20112 , \20111 );
or \U$19770 ( \20113 , \20106 , \20112 );
or \U$19771 ( \20114 , \20111 , \20105 );
nand \U$19772 ( \20115 , \20113 , \20114 );
not \U$19773 ( \20116 , \19263 );
not \U$19774 ( \20117 , \20116 );
xor \U$19775 ( \20118 , \19286 , \19331 );
not \U$19776 ( \20119 , \20118 );
or \U$19777 ( \20120 , \20117 , \20119 );
nand \U$19778 ( \20121 , \19331 , \19286 );
nand \U$19779 ( \20122 , \20120 , \20121 );
xor \U$19780 ( \20123 , \20115 , \20122 );
xor \U$19781 ( \20124 , \20099 , \20123 );
not \U$19782 ( \20125 , \20124 );
not \U$19783 ( \20126 , \20045 );
not \U$19784 ( \20127 , \20126 );
not \U$19785 ( \20128 , \20037 );
not \U$19786 ( \20129 , \20031 );
not \U$19787 ( \20130 , \20129 );
or \U$19788 ( \20131 , \20128 , \20130 );
or \U$19789 ( \20132 , \20129 , \20037 );
nand \U$19790 ( \20133 , \20131 , \20132 );
not \U$19791 ( \20134 , \20133 );
or \U$19792 ( \20135 , \20127 , \20134 );
or \U$19793 ( \20136 , \20133 , \20126 );
nand \U$19794 ( \20137 , \20135 , \20136 );
xor \U$19795 ( \20138 , \20077 , \20057 );
xnor \U$19796 ( \20139 , \20138 , \20084 );
xor \U$19797 ( \20140 , \20137 , \20139 );
not \U$19798 ( \20141 , \18957 );
not \U$19799 ( \20142 , \19808 );
or \U$19800 ( \20143 , \20141 , \20142 );
nand \U$19801 ( \20144 , \18016 , \17234 );
nand \U$19802 ( \20145 , \20143 , \20144 );
not \U$19803 ( \20146 , \20145 );
buf \U$19804 ( \20147 , \19045 );
not \U$19805 ( \20148 , \20147 );
not \U$19806 ( \20149 , \19363 );
or \U$19807 ( \20150 , \20148 , \20149 );
not \U$19808 ( \20151 , RI98734e0_189);
not \U$19809 ( \20152 , \1096 );
or \U$19810 ( \20153 , \20151 , \20152 );
or \U$19811 ( \20154 , \1096 , RI98734e0_189);
nand \U$19812 ( \20155 , \20153 , \20154 );
nand \U$19813 ( \20156 , \20155 , \19036 );
nand \U$19814 ( \20157 , \20150 , \20156 );
not \U$19815 ( \20158 , \20157 );
nand \U$19816 ( \20159 , \19788 , \8819 );
nand \U$19817 ( \20160 , \18028 , \8802 );
and \U$19818 ( \20161 , \20159 , \20160 );
not \U$19819 ( \20162 , \20161 );
or \U$19820 ( \20163 , \20158 , \20162 );
or \U$19821 ( \20164 , \20161 , \20157 );
nand \U$19822 ( \20165 , \20163 , \20164 );
not \U$19823 ( \20166 , \20165 );
or \U$19824 ( \20167 , \20146 , \20166 );
not \U$19825 ( \20168 , \20159 );
not \U$19826 ( \20169 , \20160 );
or \U$19827 ( \20170 , \20168 , \20169 );
nand \U$19828 ( \20171 , \20170 , \20157 );
nand \U$19829 ( \20172 , \20167 , \20171 );
and \U$19830 ( \20173 , \20140 , \20172 );
and \U$19831 ( \20174 , \20137 , \20139 );
or \U$19832 ( \20175 , \20173 , \20174 );
not \U$19833 ( \20176 , \20175 );
not \U$19834 ( \20177 , \19734 );
not \U$19835 ( \20178 , \19692 );
or \U$19836 ( \20179 , \20177 , \20178 );
not \U$19837 ( \20180 , \19680 );
xor \U$19838 ( \20181 , \20020 , \19691 );
nand \U$19839 ( \20182 , \20180 , \20181 );
nand \U$19840 ( \20183 , \20179 , \20182 );
or \U$19841 ( \20184 , \19559 , \19575 );
nand \U$19842 ( \20185 , \20184 , \19512 );
nand \U$19843 ( \20186 , \19559 , \19575 );
nand \U$19844 ( \20187 , \20185 , \20186 );
not \U$19845 ( \20188 , \20187 );
not \U$19846 ( \20189 , \19758 );
and \U$19847 ( \20190 , \19770 , \19748 );
not \U$19848 ( \20191 , \19770 );
not \U$19849 ( \20192 , \19748 );
and \U$19850 ( \20193 , \20191 , \20192 );
nor \U$19851 ( \20194 , \20190 , \20193 );
not \U$19852 ( \20195 , \20194 );
or \U$19853 ( \20196 , \20189 , \20195 );
nand \U$19854 ( \20197 , \19771 , \19748 );
nand \U$19855 ( \20198 , \20196 , \20197 );
xor \U$19856 ( \20199 , \19599 , \19610 );
and \U$19857 ( \20200 , \20199 , \19621 );
and \U$19858 ( \20201 , \19599 , \19610 );
or \U$19859 ( \20202 , \20200 , \20201 );
or \U$19860 ( \20203 , \20198 , \20202 );
not \U$19861 ( \20204 , \20203 );
or \U$19862 ( \20205 , \20188 , \20204 );
nand \U$19863 ( \20206 , \20198 , \20202 );
nand \U$19864 ( \20207 , \20205 , \20206 );
xor \U$19865 ( \20208 , \20183 , \20207 );
not \U$19866 ( \20209 , \20208 );
or \U$19867 ( \20210 , \20176 , \20209 );
nand \U$19868 ( \20211 , \20207 , \20183 );
nand \U$19869 ( \20212 , \20210 , \20211 );
not \U$19870 ( \20213 , \20212 );
xor \U$19871 ( \20214 , \20019 , \20090 );
xor \U$19872 ( \20215 , \20214 , \20095 );
nand \U$19873 ( \20216 , \20213 , \20215 );
not \U$19874 ( \20217 , \19997 );
not \U$19875 ( \20218 , \20016 );
or \U$19876 ( \20219 , \20217 , \20218 );
not \U$19877 ( \20220 , \19997 );
nand \U$19878 ( \20221 , \20220 , \20008 );
nand \U$19879 ( \20222 , \20219 , \20221 );
xor \U$19880 ( \20223 , \20222 , \20014 );
not \U$19881 ( \20224 , \20223 );
xor \U$19882 ( \20225 , \20025 , \20052 );
xor \U$19883 ( \20226 , \20225 , \20087 );
not \U$19884 ( \20227 , \20226 );
or \U$19885 ( \20228 , \20224 , \20227 );
or \U$19886 ( \20229 , \20226 , \20223 );
nand \U$19887 ( \20230 , \20228 , \20229 );
not \U$19888 ( \20231 , \20230 );
xor \U$19889 ( \20232 , \17996 , \18038 );
xor \U$19890 ( \20233 , \20232 , \18084 );
not \U$19891 ( \20234 , \20233 );
or \U$19892 ( \20235 , \20231 , \20234 );
not \U$19893 ( \20236 , \20226 );
nand \U$19894 ( \20237 , \20236 , \20223 );
nand \U$19895 ( \20238 , \20235 , \20237 );
and \U$19896 ( \20239 , \20216 , \20238 );
not \U$19897 ( \20240 , \20212 );
nor \U$19898 ( \20241 , \20240 , \20215 );
nor \U$19899 ( \20242 , \20239 , \20241 );
not \U$19900 ( \20243 , \20242 );
and \U$19901 ( \20244 , \20125 , \20243 );
and \U$19902 ( \20245 , \20124 , \20242 );
nor \U$19903 ( \20246 , \20244 , \20245 );
xor \U$19904 ( \20247 , \19965 , \20246 );
not \U$19905 ( \20248 , \20247 );
xor \U$19906 ( \20249 , \19927 , \19865 );
not \U$19907 ( \20250 , \20249 );
xor \U$19908 ( \20251 , \18505 , \18494 );
xnor \U$19909 ( \20252 , \20251 , \18524 );
xor \U$19910 ( \20253 , \18459 , \18469 );
xor \U$19911 ( \20254 , \20253 , \18479 );
not \U$19912 ( \20255 , \20254 );
nand \U$19913 ( \20256 , \20252 , \20255 );
not \U$19914 ( \20257 , \20256 );
not \U$19915 ( \20258 , \18583 );
not \U$19916 ( \20259 , \18560 );
not \U$19917 ( \20260 , \20259 );
or \U$19918 ( \20261 , \20258 , \20260 );
not \U$19919 ( \20262 , \18583 );
nand \U$19920 ( \20263 , \20262 , \18560 );
nand \U$19921 ( \20264 , \20261 , \20263 );
not \U$19922 ( \20265 , \20264 );
or \U$19923 ( \20266 , \20257 , \20265 );
not \U$19924 ( \20267 , \20255 );
not \U$19925 ( \20268 , \20252 );
nand \U$19926 ( \20269 , \20267 , \20268 );
nand \U$19927 ( \20270 , \20266 , \20269 );
xor \U$19928 ( \20271 , \20145 , \20165 );
not \U$19929 ( \20272 , \20271 );
xor \U$19930 ( \20273 , \18643 , \18674 );
xor \U$19931 ( \20274 , \20273 , \18660 );
not \U$19932 ( \20275 , \1518 );
and \U$19933 ( \20276 , RI9871c80_137, \19595 );
not \U$19934 ( \20277 , RI9871c80_137);
and \U$19935 ( \20278 , \20277 , \13281 );
or \U$19936 ( \20279 , \20276 , \20278 );
not \U$19937 ( \20280 , \20279 );
or \U$19938 ( \20281 , \20275 , \20280 );
not \U$19939 ( \20282 , \1800 );
not \U$19940 ( \20283 , \13625 );
or \U$19941 ( \20284 , \20282 , \20283 );
nand \U$19942 ( \20285 , \18350 , RI9871c80_137);
nand \U$19943 ( \20286 , \20284 , \20285 );
nand \U$19944 ( \20287 , \20286 , \1500 );
nand \U$19945 ( \20288 , \20281 , \20287 );
not \U$19946 ( \20289 , \20288 );
not \U$19947 ( \20290 , \1455 );
not \U$19948 ( \20291 , \1619 );
not \U$19949 ( \20292 , \10064 );
not \U$19950 ( \20293 , \20292 );
or \U$19951 ( \20294 , \20291 , \20293 );
nand \U$19952 ( \20295 , \17767 , RI9871c08_136);
nand \U$19953 ( \20296 , \20294 , \20295 );
not \U$19954 ( \20297 , \20296 );
or \U$19955 ( \20298 , \20290 , \20297 );
not \U$19956 ( \20299 , \1850 );
not \U$19957 ( \20300 , \9138 );
or \U$19958 ( \20301 , \20299 , \20300 );
not \U$19959 ( \20302 , \17756 );
not \U$19960 ( \20303 , \20302 );
nand \U$19961 ( \20304 , \20303 , RI9871c08_136);
nand \U$19962 ( \20305 , \20301 , \20304 );
nand \U$19963 ( \20306 , \20305 , \1429 );
nand \U$19964 ( \20307 , \20298 , \20306 );
not \U$19965 ( \20308 , \20307 );
or \U$19966 ( \20309 , \20289 , \20308 );
or \U$19967 ( \20310 , \20307 , \20288 );
not \U$19968 ( \20311 , \1292 );
not \U$19969 ( \20312 , \1283 );
not \U$19970 ( \20313 , \14193 );
or \U$19971 ( \20314 , \20312 , \20313 );
nand \U$19972 ( \20315 , \12773 , RI9871b18_134);
nand \U$19973 ( \20316 , \20314 , \20315 );
not \U$19974 ( \20317 , \20316 );
or \U$19975 ( \20318 , \20311 , \20317 );
and \U$19976 ( \20319 , RI9871b18_134, \12788 );
not \U$19977 ( \20320 , RI9871b18_134);
and \U$19978 ( \20321 , \20320 , \12783 );
or \U$19979 ( \20322 , \20319 , \20321 );
nand \U$19980 ( \20323 , \20322 , \1323 );
nand \U$19981 ( \20324 , \20318 , \20323 );
nand \U$19982 ( \20325 , \20310 , \20324 );
nand \U$19983 ( \20326 , \20309 , \20325 );
xor \U$19984 ( \20327 , \19524 , \19554 );
xor \U$19985 ( \20328 , \20327 , \19535 );
xor \U$19986 ( \20329 , \20326 , \20328 );
not \U$19987 ( \20330 , \6286 );
not \U$19988 ( \20331 , \18635 );
or \U$19989 ( \20332 , \20330 , \20331 );
not \U$19990 ( \20333 , RI98728b0_163);
not \U$19991 ( \20334 , \4985 );
or \U$19992 ( \20335 , \20333 , \20334 );
or \U$19993 ( \20336 , \5736 , RI98728b0_163);
nand \U$19994 ( \20337 , \20335 , \20336 );
nand \U$19995 ( \20338 , \20337 , \6284 );
nand \U$19996 ( \20339 , \20332 , \20338 );
and \U$19997 ( \20340 , \20329 , \20339 );
and \U$19998 ( \20341 , \20326 , \20328 );
or \U$19999 ( \20342 , \20340 , \20341 );
nor \U$20000 ( \20343 , \20274 , \20342 );
or \U$20001 ( \20344 , \20272 , \20343 );
nand \U$20002 ( \20345 , \20274 , \20342 );
nand \U$20003 ( \20346 , \20344 , \20345 );
xor \U$20004 ( \20347 , \20270 , \20346 );
xor \U$20005 ( \20348 , \20137 , \20139 );
xor \U$20006 ( \20349 , \20348 , \20172 );
and \U$20007 ( \20350 , \20347 , \20349 );
and \U$20008 ( \20351 , \20270 , \20346 );
or \U$20009 ( \20352 , \20350 , \20351 );
not \U$20010 ( \20353 , \20352 );
not \U$20011 ( \20354 , \20207 );
xor \U$20012 ( \20355 , \20183 , \20354 );
xnor \U$20013 ( \20356 , \20355 , \20175 );
not \U$20014 ( \20357 , \20356 );
or \U$20015 ( \20358 , \20353 , \20357 );
or \U$20016 ( \20359 , \20352 , \20356 );
not \U$20017 ( \20360 , \5796 );
not \U$20018 ( \20361 , \19727 );
or \U$20019 ( \20362 , \20360 , \20361 );
not \U$20020 ( \20363 , RI9872478_154);
not \U$20021 ( \20364 , \8053 );
or \U$20022 ( \20365 , \20363 , \20364 );
or \U$20023 ( \20366 , \8053 , RI9872478_154);
nand \U$20024 ( \20367 , \20365 , \20366 );
nand \U$20025 ( \20368 , \20367 , \5034 );
nand \U$20026 ( \20369 , \20362 , \20368 );
not \U$20027 ( \20370 , \1135 );
not \U$20028 ( \20371 , \18503 );
or \U$20029 ( \20372 , \20370 , \20371 );
and \U$20030 ( \20373 , RI98718c0_129, \12460 );
not \U$20031 ( \20374 , RI98718c0_129);
and \U$20032 ( \20375 , \20374 , \8708 );
or \U$20033 ( \20376 , \20373 , \20375 );
nand \U$20034 ( \20377 , \20376 , \1083 );
nand \U$20035 ( \20378 , \20372 , \20377 );
or \U$20036 ( \20379 , \20369 , \20378 );
not \U$20037 ( \20380 , \6144 );
not \U$20038 ( \20381 , \19698 );
or \U$20039 ( \20382 , \20380 , \20381 );
and \U$20040 ( \20383 , RI98719b0_131, \18498 );
not \U$20041 ( \20384 , RI98719b0_131);
not \U$20042 ( \20385 , \8722 );
not \U$20043 ( \20386 , \20385 );
and \U$20044 ( \20387 , \20384 , \20386 );
or \U$20045 ( \20388 , \20383 , \20387 );
nand \U$20046 ( \20389 , \20388 , \11432 );
nand \U$20047 ( \20390 , \20382 , \20389 );
and \U$20048 ( \20391 , \20379 , \20390 );
and \U$20049 ( \20392 , \20369 , \20378 );
nor \U$20050 ( \20393 , \20391 , \20392 );
not \U$20051 ( \20394 , \20393 );
not \U$20052 ( \20395 , \20394 );
not \U$20053 ( \20396 , \2087 );
not \U$20054 ( \20397 , \19719 );
or \U$20055 ( \20398 , \20396 , \20397 );
and \U$20056 ( \20399 , RI9871aa0_133, \8841 );
not \U$20057 ( \20400 , RI9871aa0_133);
and \U$20058 ( \20401 , \20400 , \18312 );
or \U$20059 ( \20402 , \20399 , \20401 );
nand \U$20060 ( \20403 , \20402 , \2071 );
nand \U$20061 ( \20404 , \20398 , \20403 );
not \U$20062 ( \20405 , \20404 );
not \U$20063 ( \20406 , \20405 );
not \U$20064 ( \20407 , \3170 );
not \U$20065 ( \20408 , \19504 );
or \U$20066 ( \20409 , \20407 , \20408 );
not \U$20067 ( \20410 , \8660 );
not \U$20068 ( \20411 , \8662 );
and \U$20069 ( \20412 , \20410 , \20411 );
and \U$20070 ( \20413 , \8660 , \8662 );
nor \U$20071 ( \20414 , \20412 , \20413 );
and \U$20072 ( \20415 , \20414 , \3154 );
not \U$20073 ( \20416 , \20414 );
and \U$20074 ( \20417 , \20416 , RI9872310_151);
nor \U$20075 ( \20418 , \20415 , \20417 );
nand \U$20076 ( \20419 , \20418 , \3163 );
nand \U$20077 ( \20420 , \20409 , \20419 );
not \U$20078 ( \20421 , \20420 );
not \U$20079 ( \20422 , \20421 );
or \U$20080 ( \20423 , \20406 , \20422 );
not \U$20081 ( \20424 , \3467 );
not \U$20082 ( \20425 , \19573 );
or \U$20083 ( \20426 , \20424 , \20425 );
not \U$20084 ( \20427 , RI98726d0_159);
not \U$20085 ( \20428 , \12716 );
or \U$20086 ( \20429 , \20427 , \20428 );
not \U$20087 ( \20430 , \8877 );
or \U$20088 ( \20431 , \20430 , RI98726d0_159);
nand \U$20089 ( \20432 , \20429 , \20431 );
nand \U$20090 ( \20433 , \20432 , \3464 );
nand \U$20091 ( \20434 , \20426 , \20433 );
nand \U$20092 ( \20435 , \20423 , \20434 );
nand \U$20093 ( \20436 , \20420 , \20404 );
nand \U$20094 ( \20437 , \20435 , \20436 );
not \U$20095 ( \20438 , \8790 );
xor \U$20096 ( \20439 , \8916 , RI98725e0_157);
not \U$20097 ( \20440 , \20439 );
or \U$20098 ( \20441 , \20438 , \20440 );
nand \U$20099 ( \20442 , \19754 , \17098 );
nand \U$20100 ( \20443 , \20441 , \20442 );
not \U$20101 ( \20444 , \20443 );
not \U$20102 ( \20445 , \875 );
not \U$20103 ( \20446 , RI9872130_147);
not \U$20104 ( \20447 , \13934 );
or \U$20105 ( \20448 , \20446 , \20447 );
not \U$20106 ( \20449 , \17003 );
buf \U$20107 ( \20450 , \20449 );
or \U$20108 ( \20451 , \20450 , RI9872130_147);
nand \U$20109 ( \20452 , \20448 , \20451 );
not \U$20110 ( \20453 , \20452 );
or \U$20111 ( \20454 , \20445 , \20453 );
not \U$20112 ( \20455 , \919 );
not \U$20113 ( \20456 , \13860 );
not \U$20114 ( \20457 , \20456 );
or \U$20115 ( \20458 , \20455 , \20457 );
or \U$20116 ( \20459 , \17883 , \919 );
nand \U$20117 ( \20460 , \20458 , \20459 );
nand \U$20118 ( \20461 , \20460 , \924 );
nand \U$20119 ( \20462 , \20454 , \20461 );
not \U$20120 ( \20463 , \20462 );
not \U$20121 ( \20464 , \1013 );
not \U$20122 ( \20465 , \19549 );
or \U$20123 ( \20466 , \20464 , \20465 );
not \U$20124 ( \20467 , \18194 );
not \U$20125 ( \20468 , \1157 );
or \U$20126 ( \20469 , \20467 , \20468 );
or \U$20127 ( \20470 , \1042 , \18194 );
nand \U$20128 ( \20471 , \20469 , \20470 );
nand \U$20129 ( \20472 , \20471 , \1016 );
nand \U$20130 ( \20473 , \20466 , \20472 );
not \U$20131 ( \20474 , \858 );
xnor \U$20132 ( \20475 , RI9871d70_139, \19411 );
not \U$20133 ( \20476 , \20475 );
or \U$20134 ( \20477 , \20474 , \20476 );
nand \U$20135 ( \20478 , \19395 , \832 );
nand \U$20136 ( \20479 , \20477 , \20478 );
xor \U$20137 ( \20480 , \20473 , \20479 );
not \U$20138 ( \20481 , \20480 );
or \U$20139 ( \20482 , \20463 , \20481 );
nand \U$20140 ( \20483 , \20479 , \20473 );
nand \U$20141 ( \20484 , \20482 , \20483 );
not \U$20142 ( \20485 , \1351 );
not \U$20143 ( \20486 , \1367 );
not \U$20144 ( \20487 , \17702 );
or \U$20145 ( \20488 , \20486 , \20487 );
not \U$20146 ( \20489 , \17701 );
buf \U$20147 ( \20490 , \20489 );
nand \U$20148 ( \20491 , \20490 , RI9871e60_141);
nand \U$20149 ( \20492 , \20488 , \20491 );
not \U$20150 ( \20493 , \20492 );
or \U$20151 ( \20494 , \20485 , \20493 );
not \U$20152 ( \20495 , \19542 );
not \U$20153 ( \20496 , RI9871e60_141);
and \U$20154 ( \20497 , \20495 , \20496 );
and \U$20155 ( \20498 , \19542 , RI9871e60_141);
nor \U$20156 ( \20499 , \20497 , \20498 );
not \U$20157 ( \20500 , \20499 );
nand \U$20158 ( \20501 , \20500 , \1379 );
nand \U$20159 ( \20502 , \20494 , \20501 );
nand \U$20160 ( \20503 , \5621 , \1009 );
and \U$20161 ( \20504 , \18705 , \20503 );
and \U$20162 ( \20505 , RI9871e60_141, RI9871f50_143);
nor \U$20163 ( \20506 , \20504 , \20505 );
and \U$20164 ( \20507 , \13385 , \20506 );
and \U$20165 ( \20508 , \20502 , \20507 );
not \U$20166 ( \20509 , \20508 );
not \U$20167 ( \20510 , \1351 );
not \U$20168 ( \20511 , \19521 );
or \U$20169 ( \20512 , \20510 , \20511 );
nand \U$20170 ( \20513 , \20492 , \1379 );
nand \U$20171 ( \20514 , \20512 , \20513 );
not \U$20172 ( \20515 , \20514 );
not \U$20173 ( \20516 , \1218 );
nand \U$20174 ( \20517 , \20516 , \19383 );
not \U$20175 ( \20518 , \20517 );
or \U$20176 ( \20519 , \20515 , \20518 );
or \U$20177 ( \20520 , \20517 , \20514 );
nand \U$20178 ( \20521 , \20519 , \20520 );
not \U$20179 ( \20522 , \20521 );
or \U$20180 ( \20523 , \20509 , \20522 );
nand \U$20181 ( \20524 , \1220 , \20514 , \19383 );
nand \U$20182 ( \20525 , \20523 , \20524 );
xor \U$20183 ( \20526 , \20484 , \20525 );
not \U$20184 ( \20527 , \20526 );
or \U$20185 ( \20528 , \20444 , \20527 );
nand \U$20186 ( \20529 , \20525 , \20484 );
nand \U$20187 ( \20530 , \20528 , \20529 );
xor \U$20188 ( \20531 , \20437 , \20530 );
not \U$20189 ( \20532 , \20531 );
or \U$20190 ( \20533 , \20395 , \20532 );
not \U$20191 ( \20534 , \20436 );
not \U$20192 ( \20535 , \20435 );
or \U$20193 ( \20536 , \20534 , \20535 );
nand \U$20194 ( \20537 , \20536 , \20530 );
nand \U$20195 ( \20538 , \20533 , \20537 );
not \U$20196 ( \20539 , \20538 );
xor \U$20197 ( \20540 , \19386 , \19397 );
not \U$20198 ( \20541 , \924 );
not \U$20199 ( \20542 , \19582 );
or \U$20200 ( \20543 , \20541 , \20542 );
nand \U$20201 ( \20544 , \20460 , \875 );
nand \U$20202 ( \20545 , \20543 , \20544 );
or \U$20203 ( \20546 , \20540 , \20545 );
not \U$20204 ( \20547 , \1517 );
not \U$20205 ( \20548 , \19604 );
or \U$20206 ( \20549 , \20547 , \20548 );
nand \U$20207 ( \20550 , \20279 , \1500 );
nand \U$20208 ( \20551 , \20549 , \20550 );
nand \U$20209 ( \20552 , \20546 , \20551 );
nand \U$20210 ( \20553 , \20540 , \20545 );
nand \U$20211 ( \20554 , \20552 , \20553 );
not \U$20212 ( \20555 , \20554 );
not \U$20213 ( \20556 , \19398 );
not \U$20214 ( \20557 , \19422 );
xnor \U$20215 ( \20558 , \20556 , \20557 );
not \U$20216 ( \20559 , \20558 );
or \U$20217 ( \20560 , \20555 , \20559 );
or \U$20218 ( \20561 , \20554 , \20558 );
nand \U$20219 ( \20562 , \20560 , \20561 );
not \U$20220 ( \20563 , \20562 );
not \U$20221 ( \20564 , \1455 );
not \U$20222 ( \20565 , \20305 );
or \U$20223 ( \20566 , \20564 , \20565 );
nand \U$20224 ( \20567 , \19617 , \1428 );
nand \U$20225 ( \20568 , \20566 , \20567 );
not \U$20226 ( \20569 , \1323 );
not \U$20227 ( \20570 , \19744 );
or \U$20228 ( \20571 , \20569 , \20570 );
nand \U$20229 ( \20572 , \20322 , \1292 );
nand \U$20230 ( \20573 , \20571 , \20572 );
xor \U$20231 ( \20574 , \20568 , \20573 );
not \U$20232 ( \20575 , \20574 );
not \U$20233 ( \20576 , \4923 );
not \U$20234 ( \20577 , \19761 );
or \U$20235 ( \20578 , \20576 , \20577 );
not \U$20236 ( \20579 , RI9872388_152);
not \U$20237 ( \20580 , \10581 );
not \U$20238 ( \20581 , \20580 );
or \U$20239 ( \20582 , \20579 , \20581 );
not \U$20240 ( \20583 , \10581 );
or \U$20241 ( \20584 , \20583 , RI9872388_152);
nand \U$20242 ( \20585 , \20582 , \20584 );
nand \U$20243 ( \20586 , \20585 , \4919 );
nand \U$20244 ( \20587 , \20578 , \20586 );
not \U$20245 ( \20588 , \20587 );
or \U$20246 ( \20589 , \20575 , \20588 );
nand \U$20247 ( \20590 , \20573 , \20568 );
nand \U$20248 ( \20591 , \20589 , \20590 );
not \U$20249 ( \20592 , \20591 );
or \U$20250 ( \20593 , \20563 , \20592 );
not \U$20251 ( \20594 , \20558 );
nand \U$20252 ( \20595 , \20594 , \20554 );
nand \U$20253 ( \20596 , \20593 , \20595 );
not \U$20254 ( \20597 , \20596 );
not \U$20255 ( \20598 , \20597 );
not \U$20256 ( \20599 , \8028 );
xor \U$20257 ( \20600 , RI9872a18_166, \4174 );
not \U$20258 ( \20601 , \20600 );
or \U$20259 ( \20602 , \20599 , \20601 );
nand \U$20260 ( \20603 , \18694 , \8039 );
nand \U$20261 ( \20604 , \20602 , \20603 );
not \U$20262 ( \20605 , \9937 );
not \U$20263 ( \20606 , \18671 );
or \U$20264 ( \20607 , \20605 , \20606 );
and \U$20265 ( \20608 , \1333 , \1335 );
not \U$20266 ( \20609 , \1333 );
not \U$20267 ( \20610 , \1335 );
and \U$20268 ( \20611 , \20609 , \20610 );
nor \U$20269 ( \20612 , \20608 , \20611 );
xnor \U$20270 ( \20613 , RI9873030_179, \20612 );
nand \U$20271 ( \20614 , \20613 , \18672 );
nand \U$20272 ( \20615 , \20607 , \20614 );
xor \U$20273 ( \20616 , \20604 , \20615 );
not \U$20274 ( \20617 , \7338 );
not \U$20275 ( \20618 , \18658 );
or \U$20276 ( \20619 , \20617 , \20618 );
xor \U$20277 ( \20620 , RI98729a0_165, \4710 );
nand \U$20278 ( \20621 , \20620 , \7325 );
nand \U$20279 ( \20622 , \20619 , \20621 );
and \U$20280 ( \20623 , \20616 , \20622 );
and \U$20281 ( \20624 , \20604 , \20615 );
or \U$20282 ( \20625 , \20623 , \20624 );
buf \U$20283 ( \20626 , \18615 );
not \U$20284 ( \20627 , \20626 );
xor \U$20285 ( \20628 , RI9873558_190, \1125 );
not \U$20286 ( \20629 , \20628 );
or \U$20287 ( \20630 , \20627 , \20629 );
nand \U$20288 ( \20631 , \18547 , RI9873648_192);
nand \U$20289 ( \20632 , \20630 , \20631 );
not \U$20290 ( \20633 , \20632 );
not \U$20291 ( \20634 , \10331 );
not \U$20292 ( \20635 , \18574 );
or \U$20293 ( \20636 , \20634 , \20635 );
not \U$20294 ( \20637 , \1208 );
not \U$20295 ( \20638 , \20637 );
and \U$20296 ( \20639 , \9694 , \20638 );
not \U$20297 ( \20640 , \9694 );
and \U$20298 ( \20641 , \20640 , \3126 );
nor \U$20299 ( \20642 , \20639 , \20641 );
nand \U$20300 ( \20643 , \20642 , \9686 );
nand \U$20301 ( \20644 , \20636 , \20643 );
not \U$20302 ( \20645 , \20644 );
or \U$20303 ( \20646 , \20633 , \20645 );
or \U$20304 ( \20647 , \20644 , \20632 );
not \U$20305 ( \20648 , \19046 );
not \U$20306 ( \20649 , \20155 );
or \U$20307 ( \20650 , \20648 , \20649 );
xor \U$20308 ( \20651 , RI98734e0_189, \1415 );
nand \U$20309 ( \20652 , \20651 , \19244 );
nand \U$20310 ( \20653 , \20650 , \20652 );
nand \U$20311 ( \20654 , \20647 , \20653 );
nand \U$20312 ( \20655 , \20646 , \20654 );
xor \U$20313 ( \20656 , \20625 , \20655 );
not \U$20314 ( \20657 , \12868 );
not \U$20315 ( \20658 , \18739 );
or \U$20316 ( \20659 , \20657 , \20658 );
not \U$20317 ( \20660 , \13022 );
not \U$20318 ( \20661 , \943 );
or \U$20319 ( \20662 , \20660 , \20661 );
or \U$20320 ( \20663 , \11283 , \13022 );
nand \U$20321 ( \20664 , \20662 , \20663 );
nand \U$20322 ( \20665 , \20664 , \13020 );
nand \U$20323 ( \20666 , \20659 , \20665 );
not \U$20324 ( \20667 , \20666 );
not \U$20325 ( \20668 , \9214 );
not \U$20326 ( \20669 , \18467 );
or \U$20327 ( \20670 , \20668 , \20669 );
not \U$20328 ( \20671 , \3537 );
not \U$20329 ( \20672 , RI9872b80_169);
and \U$20330 ( \20673 , \20671 , \20672 );
and \U$20331 ( \20674 , \6718 , RI9872b80_169);
nor \U$20332 ( \20675 , \20673 , \20674 );
nand \U$20333 ( \20676 , \20675 , \9196 );
nand \U$20334 ( \20677 , \20670 , \20676 );
not \U$20335 ( \20678 , \20677 );
nand \U$20336 ( \20679 , \18477 , \19282 );
not \U$20337 ( \20680 , RI98733f0_187);
not \U$20338 ( \20681 , \1318 );
or \U$20339 ( \20682 , \20680 , \20681 );
nand \U$20340 ( \20683 , \1306 , \17539 );
nand \U$20341 ( \20684 , \20682 , \20683 );
nand \U$20342 ( \20685 , \20684 , \17251 );
and \U$20343 ( \20686 , \20679 , \20685 );
not \U$20344 ( \20687 , \20686 );
or \U$20345 ( \20688 , \20678 , \20687 );
not \U$20346 ( \20689 , \20685 );
not \U$20347 ( \20690 , \20679 );
or \U$20348 ( \20691 , \20689 , \20690 );
not \U$20349 ( \20692 , \20677 );
nand \U$20350 ( \20693 , \20691 , \20692 );
nand \U$20351 ( \20694 , \20688 , \20693 );
not \U$20352 ( \20695 , \20694 );
or \U$20353 ( \20696 , \20667 , \20695 );
not \U$20354 ( \20697 , \20685 );
not \U$20355 ( \20698 , \20679 );
or \U$20356 ( \20699 , \20697 , \20698 );
nand \U$20357 ( \20700 , \20699 , \20677 );
nand \U$20358 ( \20701 , \20696 , \20700 );
and \U$20359 ( \20702 , \20656 , \20701 );
and \U$20360 ( \20703 , \20625 , \20655 );
or \U$20361 ( \20704 , \20702 , \20703 );
not \U$20362 ( \20705 , \20704 );
or \U$20363 ( \20706 , \20598 , \20705 );
or \U$20364 ( \20707 , \20704 , \20597 );
nand \U$20365 ( \20708 , \20706 , \20707 );
not \U$20366 ( \20709 , \20708 );
or \U$20367 ( \20710 , \20539 , \20709 );
not \U$20368 ( \20711 , \20597 );
nand \U$20369 ( \20712 , \20711 , \20704 );
nand \U$20370 ( \20713 , \20710 , \20712 );
nand \U$20371 ( \20714 , \20359 , \20713 );
nand \U$20372 ( \20715 , \20358 , \20714 );
not \U$20373 ( \20716 , \20715 );
xor \U$20374 ( \20717 , \20215 , \20212 );
xor \U$20375 ( \20718 , \20717 , \20238 );
not \U$20376 ( \20719 , \20718 );
or \U$20377 ( \20720 , \20716 , \20719 );
or \U$20378 ( \20721 , \20718 , \20715 );
nand \U$20379 ( \20722 , \20720 , \20721 );
not \U$20380 ( \20723 , \20722 );
or \U$20381 ( \20724 , \20250 , \20723 );
not \U$20382 ( \20725 , \20718 );
nand \U$20383 ( \20726 , \20725 , \20715 );
nand \U$20384 ( \20727 , \20724 , \20726 );
not \U$20385 ( \20728 , \20727 );
or \U$20386 ( \20729 , \20248 , \20728 );
or \U$20387 ( \20730 , \20727 , \20247 );
nand \U$20388 ( \20731 , \20729 , \20730 );
not \U$20389 ( \20732 , \20731 );
or \U$20390 ( \20733 , \19941 , \20732 );
not \U$20391 ( \20734 , \20247 );
nand \U$20392 ( \20735 , \20734 , \20727 );
nand \U$20393 ( \20736 , \20733 , \20735 );
not \U$20394 ( \20737 , \20736 );
xor \U$20395 ( \20738 , \19229 , \20737 );
not \U$20396 ( \20739 , \20124 );
nand \U$20397 ( \20740 , \20739 , \20242 );
not \U$20398 ( \20741 , \20740 );
not \U$20399 ( \20742 , \19965 );
or \U$20400 ( \20743 , \20741 , \20742 );
not \U$20401 ( \20744 , \20242 );
nand \U$20402 ( \20745 , \20744 , \20124 );
nand \U$20403 ( \20746 , \20743 , \20745 );
not \U$20404 ( \20747 , \20122 );
not \U$20405 ( \20748 , \20115 );
or \U$20406 ( \20749 , \20747 , \20748 );
nand \U$20407 ( \20750 , \20111 , \20104 );
nand \U$20408 ( \20751 , \20749 , \20750 );
not \U$20409 ( \20752 , \20751 );
not \U$20410 ( \20753 , \19974 );
not \U$20411 ( \20754 , \20753 );
not \U$20412 ( \20755 , \19993 );
or \U$20413 ( \20756 , \20754 , \20755 );
nand \U$20414 ( \20757 , \19988 , \19980 );
nand \U$20415 ( \20758 , \20756 , \20757 );
not \U$20416 ( \20759 , \20758 );
and \U$20417 ( \20760 , \17682 , \17727 );
not \U$20418 ( \20761 , \18842 );
not \U$20419 ( \20762 , \9429 );
or \U$20420 ( \20763 , \20761 , \20762 );
not \U$20421 ( \20764 , \13933 );
buf \U$20422 ( \20765 , \20764 );
and \U$20423 ( \20766 , \20765 , \9120 );
not \U$20424 ( \20767 , \20765 );
and \U$20425 ( \20768 , \20767 , \17682 );
nor \U$20426 ( \20769 , \20766 , \20768 );
nand \U$20427 ( \20770 , \20769 , \1220 );
nand \U$20428 ( \20771 , \20763 , \20770 );
not \U$20429 ( \20772 , \20771 );
xor \U$20430 ( \20773 , \20760 , \20772 );
xor \U$20431 ( \20774 , \9139 , RI9872130_147);
not \U$20432 ( \20775 , \20774 );
not \U$20433 ( \20776 , \875 );
or \U$20434 ( \20777 , \20775 , \20776 );
not \U$20435 ( \20778 , RI9872130_147);
not \U$20436 ( \20779 , \9114 );
or \U$20437 ( \20780 , \20778 , \20779 );
or \U$20438 ( \20781 , \9722 , RI9872130_147);
nand \U$20439 ( \20782 , \20780 , \20781 );
nand \U$20440 ( \20783 , \20782 , \924 );
nand \U$20441 ( \20784 , \20777 , \20783 );
xor \U$20442 ( \20785 , \20773 , \20784 );
not \U$20443 ( \20786 , \1013 );
not \U$20444 ( \20787 , \13623 );
and \U$20445 ( \20788 , \20787 , \1146 );
not \U$20446 ( \20789 , \20787 );
and \U$20447 ( \20790 , \20789 , \8085 );
nor \U$20448 ( \20791 , \20788 , \20790 );
not \U$20449 ( \20792 , \20791 );
or \U$20450 ( \20793 , \20786 , \20792 );
nand \U$20451 ( \20794 , \17019 , \1018 );
nand \U$20452 ( \20795 , \20793 , \20794 );
not \U$20453 ( \20796 , \1352 );
and \U$20454 ( \20797 , \12774 , RI9871e60_141);
not \U$20455 ( \20798 , \12774 );
and \U$20456 ( \20799 , \20798 , \17844 );
nor \U$20457 ( \20800 , \20797 , \20799 );
not \U$20458 ( \20801 , \20800 );
or \U$20459 ( \20802 , \20796 , \20801 );
nand \U$20460 ( \20803 , \18999 , \1380 );
nand \U$20461 ( \20804 , \20802 , \20803 );
not \U$20462 ( \20805 , \20804 );
xor \U$20463 ( \20806 , \20795 , \20805 );
not \U$20464 ( \20807 , \832 );
and \U$20465 ( \20808 , RI9871d70_139, \10064 );
not \U$20466 ( \20809 , RI9871d70_139);
and \U$20467 ( \20810 , \20809 , \20292 );
or \U$20468 ( \20811 , \20808 , \20810 );
not \U$20469 ( \20812 , \20811 );
or \U$20470 ( \20813 , \20807 , \20812 );
nand \U$20471 ( \20814 , \18991 , \859 );
nand \U$20472 ( \20815 , \20813 , \20814 );
xnor \U$20473 ( \20816 , \20806 , \20815 );
xor \U$20474 ( \20817 , \20785 , \20816 );
xor \U$20475 ( \20818 , \18785 , \17021 );
not \U$20476 ( \20819 , \20818 );
not \U$20477 ( \20820 , \17051 );
or \U$20478 ( \20821 , \20819 , \20820 );
xor \U$20479 ( \20822 , \20818 , \17051 );
nand \U$20480 ( \20823 , \20822 , \17037 );
nand \U$20481 ( \20824 , \20821 , \20823 );
xnor \U$20482 ( \20825 , \20817 , \20824 );
not \U$20483 ( \20826 , \16985 );
not \U$20484 ( \20827 , \20826 );
not \U$20485 ( \20828 , \17053 );
or \U$20486 ( \20829 , \20827 , \20828 );
not \U$20487 ( \20830 , \17052 );
not \U$20488 ( \20831 , \16985 );
or \U$20489 ( \20832 , \20830 , \20831 );
nand \U$20490 ( \20833 , \20832 , \16933 );
nand \U$20491 ( \20834 , \20829 , \20833 );
not \U$20492 ( \20835 , \20834 );
xor \U$20493 ( \20836 , \20825 , \20835 );
not \U$20494 ( \20837 , \18982 );
not \U$20495 ( \20838 , \20837 );
not \U$20496 ( \20839 , \19008 );
or \U$20497 ( \20840 , \20838 , \20839 );
nand \U$20498 ( \20841 , \18993 , \19003 );
nand \U$20499 ( \20842 , \20840 , \20841 );
not \U$20500 ( \20843 , \20842 );
or \U$20501 ( \20844 , \16950 , \16980 );
nand \U$20502 ( \20845 , \20844 , \16961 );
nand \U$20503 ( \20846 , \16950 , \16980 );
nand \U$20504 ( \20847 , \20845 , \20846 );
xor \U$20505 ( \20848 , \20843 , \20847 );
xor \U$20506 ( \20849 , \17455 , \17465 );
and \U$20507 ( \20850 , \20849 , \17475 );
and \U$20508 ( \20851 , \17455 , \17465 );
or \U$20509 ( \20852 , \20850 , \20851 );
xor \U$20510 ( \20853 , \20848 , \20852 );
xnor \U$20511 ( \20854 , \20836 , \20853 );
not \U$20512 ( \20855 , \20854 );
not \U$20513 ( \20856 , \20855 );
or \U$20514 ( \20857 , \20759 , \20856 );
not \U$20515 ( \20858 , \20758 );
nand \U$20516 ( \20859 , \20858 , \20854 );
nand \U$20517 ( \20860 , \20857 , \20859 );
not \U$20518 ( \20861 , \20860 );
xor \U$20519 ( \20862 , \20752 , \20861 );
not \U$20520 ( \20863 , \20123 );
not \U$20521 ( \20864 , \20099 );
or \U$20522 ( \20865 , \20863 , \20864 );
not \U$20523 ( \20866 , \20098 );
and \U$20524 ( \20867 , \19993 , \19974 );
not \U$20525 ( \20868 , \19993 );
and \U$20526 ( \20869 , \20868 , \20753 );
or \U$20527 ( \20870 , \20867 , \20869 );
nand \U$20528 ( \20871 , \20866 , \20870 );
nand \U$20529 ( \20872 , \20865 , \20871 );
not \U$20530 ( \20873 , \20872 );
xnor \U$20531 ( \20874 , \20862 , \20873 );
not \U$20532 ( \20875 , \19943 );
not \U$20533 ( \20876 , \19959 );
or \U$20534 ( \20877 , \20875 , \20876 );
not \U$20535 ( \20878 , \19955 );
nand \U$20536 ( \20879 , \20878 , \19951 );
nand \U$20537 ( \20880 , \20877 , \20879 );
not \U$20538 ( \20881 , \20880 );
and \U$20539 ( \20882 , \20874 , \20881 );
not \U$20540 ( \20883 , \20874 );
and \U$20541 ( \20884 , \20883 , \20880 );
or \U$20542 ( \20885 , \20882 , \20884 );
xor \U$20543 ( \20886 , \20746 , \20885 );
not \U$20544 ( \20887 , \19939 );
not \U$20545 ( \20888 , \19937 );
or \U$20546 ( \20889 , \20887 , \20888 );
not \U$20547 ( \20890 , \19845 );
not \U$20548 ( \20891 , \19843 );
or \U$20549 ( \20892 , \20890 , \20891 );
nand \U$20550 ( \20893 , \20892 , \19932 );
nand \U$20551 ( \20894 , \20889 , \20893 );
xnor \U$20552 ( \20895 , \20886 , \20894 );
and \U$20553 ( \20896 , \20738 , \20895 );
and \U$20554 ( \20897 , \19229 , \20737 );
or \U$20555 ( \20898 , \20896 , \20897 );
not \U$20556 ( \20899 , \20898 );
not \U$20557 ( \20900 , \20899 );
or \U$20558 ( \20901 , \20816 , \20785 );
nand \U$20559 ( \20902 , \20901 , \20824 );
nand \U$20560 ( \20903 , \20816 , \20785 );
nand \U$20561 ( \20904 , \20902 , \20903 );
not \U$20562 ( \20905 , \17356 );
not \U$20563 ( \20906 , \17433 );
not \U$20564 ( \20907 , \20906 );
or \U$20565 ( \20908 , \20905 , \20907 );
nand \U$20566 ( \20909 , \17398 , \17428 );
nand \U$20567 ( \20910 , \20908 , \20909 );
xor \U$20568 ( \20911 , \20904 , \20910 );
xor \U$20569 ( \20912 , \17607 , \17635 );
and \U$20570 ( \20913 , \20912 , \17675 );
and \U$20571 ( \20914 , \17607 , \17635 );
or \U$20572 ( \20915 , \20913 , \20914 );
xor \U$20573 ( \20916 , \20911 , \20915 );
not \U$20574 ( \20917 , \832 );
and \U$20575 ( \20918 , \13070 , RI9871d70_139);
not \U$20576 ( \20919 , \13070 );
and \U$20577 ( \20920 , \20919 , \2243 );
nor \U$20578 ( \20921 , \20918 , \20920 );
not \U$20579 ( \20922 , \20921 );
or \U$20580 ( \20923 , \20917 , \20922 );
nand \U$20581 ( \20924 , \20811 , \859 );
nand \U$20582 ( \20925 , \20923 , \20924 );
xor \U$20583 ( \20926 , \20771 , \20925 );
not \U$20584 ( \20927 , \1013 );
not \U$20585 ( \20928 , \13281 );
and \U$20586 ( \20929 , \12592 , \20928 );
not \U$20587 ( \20930 , \12592 );
and \U$20588 ( \20931 , \20930 , \13281 );
nor \U$20589 ( \20932 , \20929 , \20931 );
not \U$20590 ( \20933 , \20932 );
or \U$20591 ( \20934 , \20927 , \20933 );
not \U$20592 ( \20935 , \20791 );
or \U$20593 ( \20936 , \20935 , \1612 );
nand \U$20594 ( \20937 , \20934 , \20936 );
xor \U$20595 ( \20938 , \20926 , \20937 );
and \U$20596 ( \20939 , \19147 , \19157 );
and \U$20597 ( \20940 , \19136 , \19146 );
nor \U$20598 ( \20941 , \20939 , \20940 );
xor \U$20599 ( \20942 , \20938 , \20941 );
xor \U$20600 ( \20943 , \19167 , \19178 );
and \U$20601 ( \20944 , \20943 , \19191 );
and \U$20602 ( \20945 , \19167 , \19178 );
or \U$20603 ( \20946 , \20944 , \20945 );
xnor \U$20604 ( \20947 , \20942 , \20946 );
xor \U$20605 ( \20948 , \18910 , \18920 );
and \U$20606 ( \20949 , \20948 , \18930 );
and \U$20607 ( \20950 , \18910 , \18920 );
or \U$20608 ( \20951 , \20949 , \20950 );
or \U$20609 ( \20952 , \18953 , \18968 );
nand \U$20610 ( \20953 , \20952 , \18955 );
xor \U$20611 ( \20954 , \20951 , \20953 );
not \U$20612 ( \20955 , \19202 );
and \U$20613 ( \20956 , \19224 , \19212 );
not \U$20614 ( \20957 , \19224 );
not \U$20615 ( \20958 , \19212 );
and \U$20616 ( \20959 , \20957 , \20958 );
nor \U$20617 ( \20960 , \20956 , \20959 );
not \U$20618 ( \20961 , \20960 );
or \U$20619 ( \20962 , \20955 , \20961 );
nand \U$20620 ( \20963 , \19224 , \19212 );
nand \U$20621 ( \20964 , \20962 , \20963 );
xor \U$20622 ( \20965 , \20954 , \20964 );
xor \U$20623 ( \20966 , \20947 , \20965 );
not \U$20624 ( \20967 , \18931 );
xor \U$20625 ( \20968 , \18967 , \18899 );
xor \U$20626 ( \20969 , \20968 , \18956 );
not \U$20627 ( \20970 , \20969 );
or \U$20628 ( \20971 , \20967 , \20970 );
not \U$20629 ( \20972 , \18899 );
nand \U$20630 ( \20973 , \20972 , \18972 );
nand \U$20631 ( \20974 , \20971 , \20973 );
xor \U$20632 ( \20975 , \20966 , \20974 );
xor \U$20633 ( \20976 , \20916 , \20975 );
or \U$20634 ( \20977 , \18826 , \18822 );
and \U$20635 ( \20978 , \20977 , \18869 );
and \U$20636 ( \20979 , \18822 , \18826 );
nor \U$20637 ( \20980 , \20978 , \20979 );
not \U$20638 ( \20981 , \1083 );
not \U$20639 ( \20982 , \17604 );
or \U$20640 ( \20983 , \20981 , \20982 );
and \U$20641 ( \20984 , RI98718c0_129, \10601 );
not \U$20642 ( \20985 , RI98718c0_129);
and \U$20643 ( \20986 , \20985 , \8624 );
nor \U$20644 ( \20987 , \20984 , \20986 );
nand \U$20645 ( \20988 , \20987 , \6672 );
nand \U$20646 ( \20989 , \20983 , \20988 );
not \U$20647 ( \20990 , \1456 );
not \U$20648 ( \20991 , \17630 );
or \U$20649 ( \20992 , \20990 , \20991 );
not \U$20650 ( \20993 , RI9871c08_136);
not \U$20651 ( \20994 , \8857 );
or \U$20652 ( \20995 , \20993 , \20994 );
nand \U$20653 ( \20996 , \9885 , \1850 );
nand \U$20654 ( \20997 , \20995 , \20996 );
nand \U$20655 ( \20998 , \20997 , \1429 );
nand \U$20656 ( \20999 , \20992 , \20998 );
xor \U$20657 ( \21000 , \20989 , \20999 );
not \U$20658 ( \21001 , \12720 );
not \U$20659 ( \21002 , \17612 );
or \U$20660 ( \21003 , \21001 , \21002 );
and \U$20661 ( \21004 , RI9871b18_134, \8575 );
not \U$20662 ( \21005 , RI9871b18_134);
and \U$20663 ( \21006 , \21005 , \8579 );
nor \U$20664 ( \21007 , \21004 , \21006 );
nand \U$20665 ( \21008 , \21007 , \1323 );
nand \U$20666 ( \21009 , \21003 , \21008 );
xor \U$20667 ( \21010 , \21000 , \21009 );
not \U$20668 ( \21011 , \6145 );
and \U$20669 ( \21012 , RI98719b0_131, \8334 );
not \U$20670 ( \21013 , RI98719b0_131);
and \U$20671 ( \21014 , \21013 , \8916 );
or \U$20672 ( \21015 , \21012 , \21014 );
not \U$20673 ( \21016 , \21015 );
or \U$20674 ( \21017 , \21011 , \21016 );
nand \U$20675 ( \21018 , \17577 , \793 );
nand \U$20676 ( \21019 , \21017 , \21018 );
not \U$20677 ( \21020 , \2087 );
not \U$20678 ( \21021 , RI9871aa0_133);
not \U$20679 ( \21022 , \10583 );
or \U$20680 ( \21023 , \21021 , \21022 );
or \U$20681 ( \21024 , \10583 , RI9871aa0_133);
nand \U$20682 ( \21025 , \21023 , \21024 );
not \U$20683 ( \21026 , \21025 );
or \U$20684 ( \21027 , \21020 , \21026 );
nand \U$20685 ( \21028 , \17587 , \2072 );
nand \U$20686 ( \21029 , \21027 , \21028 );
xor \U$20687 ( \21030 , \21019 , \21029 );
not \U$20688 ( \21031 , \3170 );
not \U$20689 ( \21032 , \3154 );
not \U$20690 ( \21033 , \12802 );
or \U$20691 ( \21034 , \21032 , \21033 );
nand \U$20692 ( \21035 , \8054 , RI9872310_151);
nand \U$20693 ( \21036 , \21034 , \21035 );
not \U$20694 ( \21037 , \21036 );
or \U$20695 ( \21038 , \21031 , \21037 );
not \U$20696 ( \21039 , \18796 );
or \U$20697 ( \21040 , \21039 , \10947 );
nand \U$20698 ( \21041 , \21038 , \21040 );
xor \U$20699 ( \21042 , \21030 , \21041 );
xor \U$20700 ( \21043 , \21010 , \21042 );
not \U$20701 ( \21044 , \1162 );
not \U$20702 ( \21045 , \20769 );
or \U$20703 ( \21046 , \21044 , \21045 );
and \U$20704 ( \21047 , \17883 , \17682 );
not \U$20705 ( \21048 , \17883 );
and \U$20706 ( \21049 , \21048 , \12780 );
nor \U$20707 ( \21050 , \21047 , \21049 );
nand \U$20708 ( \21051 , \1220 , \21050 );
nand \U$20709 ( \21052 , \21046 , \21051 );
nand \U$20710 ( \21053 , RI9873468_188, RI98734e0_189);
and \U$20711 ( \21054 , \21053 , RI98733f0_187);
not \U$20712 ( \21055 , \21054 );
and \U$20713 ( \21056 , \17744 , \8678 );
not \U$20714 ( \21057 , \21056 );
or \U$20715 ( \21058 , \21055 , \21057 );
or \U$20716 ( \21059 , \21056 , \21054 );
nand \U$20717 ( \21060 , \21058 , \21059 );
xnor \U$20718 ( \21061 , \21052 , \21060 );
not \U$20719 ( \21062 , \5796 );
not \U$20720 ( \21063 , RI9872478_154);
not \U$20721 ( \21064 , \14562 );
or \U$20722 ( \21065 , \21063 , \21064 );
or \U$20723 ( \21066 , \12616 , RI9872478_154);
nand \U$20724 ( \21067 , \21065 , \21066 );
not \U$20725 ( \21068 , \21067 );
or \U$20726 ( \21069 , \21062 , \21068 );
nand \U$20727 ( \21070 , \18852 , \5034 );
nand \U$20728 ( \21071 , \21069 , \21070 );
xor \U$20729 ( \21072 , \21061 , \21071 );
not \U$20730 ( \21073 , \9273 );
not \U$20731 ( \21074 , RI9872e50_175);
not \U$20732 ( \21075 , \820 );
or \U$20733 ( \21076 , \21074 , \21075 );
nand \U$20734 ( \21077 , \6219 , \9694 );
nand \U$20735 ( \21078 , \21076 , \21077 );
not \U$20736 ( \21079 , \21078 );
or \U$20737 ( \21080 , \21073 , \21079 );
nand \U$20738 ( \21081 , \18864 , \9686 );
nand \U$20739 ( \21082 , \21080 , \21081 );
xnor \U$20740 ( \21083 , \21072 , \21082 );
xor \U$20741 ( \21084 , \21043 , \21083 );
xor \U$20742 ( \21085 , \20980 , \21084 );
not \U$20743 ( \21086 , \19192 );
xor \U$20744 ( \21087 , \19203 , \19158 );
xor \U$20745 ( \21088 , \21087 , \20960 );
not \U$20746 ( \21089 , \21088 );
or \U$20747 ( \21090 , \21086 , \21089 );
not \U$20748 ( \21091 , \19158 );
nand \U$20749 ( \21092 , \21091 , \19225 );
nand \U$20750 ( \21093 , \21090 , \21092 );
xnor \U$20751 ( \21094 , \21085 , \21093 );
xor \U$20752 ( \21095 , \20976 , \21094 );
xor \U$20753 ( \21096 , \18888 , \18894 );
and \U$20754 ( \21097 , \21096 , \19227 );
and \U$20755 ( \21098 , \18888 , \18894 );
or \U$20756 ( \21099 , \21097 , \21098 );
xor \U$20757 ( \21100 , \21095 , \21099 );
xor \U$20758 ( \21101 , \18870 , \18878 );
and \U$20759 ( \21102 , \21101 , \18887 );
and \U$20760 ( \21103 , \18870 , \18878 );
or \U$20761 ( \21104 , \21102 , \21103 );
not \U$20762 ( \21105 , \19118 );
not \U$20763 ( \21106 , \19122 );
or \U$20764 ( \21107 , \21105 , \21106 );
nand \U$20765 ( \21108 , \19113 , \19058 );
nand \U$20766 ( \21109 , \21107 , \21108 );
and \U$20767 ( \21110 , RI9871c80_137, \12470 );
not \U$20768 ( \21111 , RI9871c80_137);
and \U$20769 ( \21112 , \21111 , \18498 );
nor \U$20770 ( \21113 , \21110 , \21112 );
and \U$20771 ( \21114 , \21113 , \1518 );
and \U$20772 ( \21115 , \1501 , \19132 );
nor \U$20773 ( \21116 , \21114 , \21115 );
not \U$20774 ( \21117 , \21116 );
not \U$20775 ( \21118 , \4919 );
not \U$20776 ( \21119 , \19142 );
or \U$20777 ( \21120 , \21118 , \21119 );
not \U$20778 ( \21121 , \4902 );
not \U$20779 ( \21122 , \4472 );
or \U$20780 ( \21123 , \21121 , \21122 );
nand \U$20781 ( \21124 , \4470 , RI9872388_152);
nand \U$20782 ( \21125 , \21123 , \21124 );
nand \U$20783 ( \21126 , \21125 , \4925 );
nand \U$20784 ( \21127 , \21120 , \21126 );
not \U$20785 ( \21128 , \21127 );
or \U$20786 ( \21129 , \21117 , \21128 );
or \U$20787 ( \21130 , \21127 , \21116 );
nand \U$20788 ( \21131 , \21129 , \21130 );
not \U$20789 ( \21132 , \10242 );
not \U$20790 ( \21133 , \8807 );
not \U$20791 ( \21134 , \8165 );
or \U$20792 ( \21135 , \21133 , \21134 );
or \U$20793 ( \21136 , \944 , \8811 );
nand \U$20794 ( \21137 , \21135 , \21136 );
not \U$20795 ( \21138 , \21137 );
or \U$20796 ( \21139 , \21132 , \21138 );
nand \U$20797 ( \21140 , \19155 , \10251 );
nand \U$20798 ( \21141 , \21139 , \21140 );
xor \U$20799 ( \21142 , \21131 , \21141 );
not \U$20800 ( \21143 , \21142 );
xor \U$20801 ( \21144 , \18850 , \18868 );
nand \U$20802 ( \21145 , \21144 , \18856 );
not \U$20803 ( \21146 , \21145 );
and \U$20804 ( \21147 , \18850 , \18868 );
nor \U$20805 ( \21148 , \21146 , \21147 );
not \U$20806 ( \21149 , \21148 );
or \U$20807 ( \21150 , \21143 , \21149 );
not \U$20808 ( \21151 , \21147 );
not \U$20809 ( \21152 , \21151 );
not \U$20810 ( \21153 , \21145 );
or \U$20811 ( \21154 , \21152 , \21153 );
not \U$20812 ( \21155 , \21142 );
nand \U$20813 ( \21156 , \21154 , \21155 );
nand \U$20814 ( \21157 , \21150 , \21156 );
not \U$20815 ( \21158 , \5642 );
not \U$20816 ( \21159 , \19200 );
or \U$20817 ( \21160 , \21158 , \21159 );
not \U$20818 ( \21161 , \5644 );
not \U$20819 ( \21162 , \6718 );
or \U$20820 ( \21163 , \21161 , \21162 );
or \U$20821 ( \21164 , \3543 , \5644 );
nand \U$20822 ( \21165 , \21163 , \21164 );
nand \U$20823 ( \21166 , \21165 , \7188 );
nand \U$20824 ( \21167 , \21160 , \21166 );
not \U$20825 ( \21168 , \6611 );
not \U$20826 ( \21169 , RI98728b0_163);
not \U$20827 ( \21170 , \3691 );
or \U$20828 ( \21171 , \21169 , \21170 );
or \U$20829 ( \21172 , \3691 , RI98728b0_163);
nand \U$20830 ( \21173 , \21171 , \21172 );
not \U$20831 ( \21174 , \21173 );
or \U$20832 ( \21175 , \21168 , \21174 );
nand \U$20833 ( \21176 , \19208 , \6284 );
nand \U$20834 ( \21177 , \21175 , \21176 );
xor \U$20835 ( \21178 , \21167 , \21177 );
not \U$20836 ( \21179 , \9527 );
not \U$20837 ( \21180 , \19220 );
or \U$20838 ( \21181 , \21179 , \21180 );
and \U$20839 ( \21182 , \916 , \14080 );
not \U$20840 ( \21183 , \916 );
and \U$20841 ( \21184 , \21183 , RI9872f40_177);
nor \U$20842 ( \21185 , \21182 , \21184 );
nand \U$20843 ( \21186 , \21185 , \11199 );
nand \U$20844 ( \21187 , \21181 , \21186 );
xor \U$20845 ( \21188 , \21178 , \21187 );
not \U$20846 ( \21189 , \21188 );
and \U$20847 ( \21190 , \21157 , \21189 );
not \U$20848 ( \21191 , \21157 );
and \U$20849 ( \21192 , \21191 , \21188 );
nor \U$20850 ( \21193 , \21190 , \21192 );
not \U$20851 ( \21194 , \21193 );
not \U$20852 ( \21195 , \17098 );
and \U$20853 ( \21196 , RI98725e0_157, \4986 );
not \U$20854 ( \21197 , RI98725e0_157);
and \U$20855 ( \21198 , \21197 , \9374 );
or \U$20856 ( \21199 , \21196 , \21198 );
not \U$20857 ( \21200 , \21199 );
or \U$20858 ( \21201 , \21195 , \21200 );
nand \U$20859 ( \21202 , \19162 , \18171 );
nand \U$20860 ( \21203 , \21201 , \21202 );
not \U$20861 ( \21204 , \9670 );
not \U$20862 ( \21205 , \19176 );
or \U$20863 ( \21206 , \21204 , \21205 );
not \U$20864 ( \21207 , \9185 );
not \U$20865 ( \21208 , \9834 );
or \U$20866 ( \21209 , \21207 , \21208 );
nand \U$20867 ( \21210 , \17363 , RI9872bf8_170);
nand \U$20868 ( \21211 , \21209 , \21210 );
nand \U$20869 ( \21212 , \21211 , \9668 );
nand \U$20870 ( \21213 , \21206 , \21212 );
xor \U$20871 ( \21214 , \21203 , \21213 );
not \U$20872 ( \21215 , \18508 );
not \U$20873 ( \21216 , \19184 );
or \U$20874 ( \21217 , \21215 , \21216 );
and \U$20875 ( \21218 , RI9873288_184, \7330 );
not \U$20876 ( \21219 , RI9873288_184);
and \U$20877 ( \21220 , \21219 , \2360 );
nor \U$20878 ( \21221 , \21218 , \21220 );
nand \U$20879 ( \21222 , \21221 , \18522 );
nand \U$20880 ( \21223 , \21217 , \21222 );
xor \U$20881 ( \21224 , \21214 , \21223 );
not \U$20882 ( \21225 , \7338 );
and \U$20883 ( \21226 , RI98729a0_165, \2116 );
not \U$20884 ( \21227 , RI98729a0_165);
and \U$20885 ( \21228 , \21227 , \3275 );
or \U$20886 ( \21229 , \21226 , \21228 );
not \U$20887 ( \21230 , \21229 );
or \U$20888 ( \21231 , \21225 , \21230 );
nand \U$20889 ( \21232 , \18950 , \7325 );
nand \U$20890 ( \21233 , \21231 , \21232 );
not \U$20891 ( \21234 , \17234 );
and \U$20892 ( \21235 , RI9873210_183, \1724 );
not \U$20893 ( \21236 , RI9873210_183);
and \U$20894 ( \21237 , \21236 , \1126 );
or \U$20895 ( \21238 , \21235 , \21237 );
not \U$20896 ( \21239 , \21238 );
or \U$20897 ( \21240 , \21234 , \21239 );
nand \U$20898 ( \21241 , \18965 , \18957 );
nand \U$20899 ( \21242 , \21240 , \21241 );
xor \U$20900 ( \21243 , \21233 , \21242 );
not \U$20901 ( \21244 , \8029 );
not \U$20902 ( \21245 , \18939 );
or \U$20903 ( \21246 , \21244 , \21245 );
not \U$20904 ( \21247 , RI9872a18_166);
not \U$20905 ( \21248 , \3127 );
or \U$20906 ( \21249 , \21247 , \21248 );
nand \U$20907 ( \21250 , \11114 , \8031 );
nand \U$20908 ( \21251 , \21249 , \21250 );
nand \U$20909 ( \21252 , \21251 , \8041 );
nand \U$20910 ( \21253 , \21246 , \21252 );
xor \U$20911 ( \21254 , \21243 , \21253 );
xor \U$20912 ( \21255 , \21224 , \21254 );
not \U$20913 ( \21256 , \11350 );
not \U$20914 ( \21257 , \18928 );
or \U$20915 ( \21258 , \21256 , \21257 );
not \U$20916 ( \21259 , \6692 );
xor \U$20917 ( \21260 , RI98730a8_180, \21259 );
nand \U$20918 ( \21261 , \21260 , \12868 );
nand \U$20919 ( \21262 , \21258 , \21261 );
not \U$20920 ( \21263 , \13109 );
not \U$20921 ( \21264 , \18916 );
or \U$20922 ( \21265 , \21263 , \21264 );
not \U$20923 ( \21266 , RI9873030_179);
not \U$20924 ( \21267 , \9230 );
or \U$20925 ( \21268 , \21266 , \21267 );
or \U$20926 ( \21269 , \1320 , RI9873030_179);
nand \U$20927 ( \21270 , \21268 , \21269 );
nand \U$20928 ( \21271 , \21270 , \9937 );
nand \U$20929 ( \21272 , \21265 , \21271 );
not \U$20930 ( \21273 , \21272 );
xor \U$20931 ( \21274 , \21262 , \21273 );
not \U$20932 ( \21275 , \9196 );
not \U$20933 ( \21276 , \18906 );
or \U$20934 ( \21277 , \21275 , \21276 );
not \U$20935 ( \21278 , \9198 );
not \U$20936 ( \21279 , \1713 );
or \U$20937 ( \21280 , \21278 , \21279 );
or \U$20938 ( \21281 , \10133 , \9198 );
nand \U$20939 ( \21282 , \21280 , \21281 );
nand \U$20940 ( \21283 , \21282 , \9214 );
nand \U$20941 ( \21284 , \21277 , \21283 );
not \U$20942 ( \21285 , \21284 );
and \U$20943 ( \21286 , \21274 , \21285 );
not \U$20944 ( \21287 , \21274 );
and \U$20945 ( \21288 , \21287 , \21284 );
nor \U$20946 ( \21289 , \21286 , \21288 );
xor \U$20947 ( \21290 , \21255 , \21289 );
not \U$20948 ( \21291 , \21290 );
or \U$20949 ( \21292 , \21194 , \21291 );
or \U$20950 ( \21293 , \21290 , \21193 );
nand \U$20951 ( \21294 , \21292 , \21293 );
xor \U$20952 ( \21295 , \21109 , \21294 );
xor \U$20953 ( \21296 , \21104 , \21295 );
not \U$20954 ( \21297 , \19127 );
xor \U$20955 ( \21298 , \19226 , \18973 );
not \U$20956 ( \21299 , \21298 );
or \U$20957 ( \21300 , \21297 , \21299 );
nand \U$20958 ( \21301 , \19226 , \18973 );
nand \U$20959 ( \21302 , \21300 , \21301 );
xnor \U$20960 ( \21303 , \21296 , \21302 );
xor \U$20961 ( \21304 , \21100 , \21303 );
not \U$20962 ( \21305 , \21304 );
not \U$20963 ( \21306 , \20894 );
not \U$20964 ( \21307 , \20746 );
not \U$20965 ( \21308 , \21307 );
not \U$20966 ( \21309 , \20885 );
or \U$20967 ( \21310 , \21308 , \21309 );
or \U$20968 ( \21311 , \20885 , \21307 );
nand \U$20969 ( \21312 , \21310 , \21311 );
not \U$20970 ( \21313 , \21312 );
or \U$20971 ( \21314 , \21306 , \21313 );
nand \U$20972 ( \21315 , \20885 , \20746 );
nand \U$20973 ( \21316 , \21314 , \21315 );
not \U$20974 ( \21317 , \21316 );
or \U$20975 ( \21318 , \21305 , \21317 );
or \U$20976 ( \21319 , \21316 , \21304 );
nand \U$20977 ( \21320 , \21318 , \21319 );
not \U$20978 ( \21321 , \20880 );
not \U$20979 ( \21322 , \20874 );
or \U$20980 ( \21323 , \21321 , \21322 );
nand \U$20981 ( \21324 , \20860 , \20752 );
not \U$20982 ( \21325 , \21324 );
nand \U$20983 ( \21326 , \20861 , \20751 );
not \U$20984 ( \21327 , \21326 );
or \U$20985 ( \21328 , \21325 , \21327 );
nand \U$20986 ( \21329 , \21328 , \20872 );
nand \U$20987 ( \21330 , \21323 , \21329 );
not \U$20988 ( \21331 , \21330 );
not \U$20989 ( \21332 , \20751 );
not \U$20990 ( \21333 , \20860 );
or \U$20991 ( \21334 , \21332 , \21333 );
nand \U$20992 ( \21335 , \20854 , \20758 );
nand \U$20993 ( \21336 , \21334 , \21335 );
not \U$20994 ( \21337 , \18817 );
not \U$20995 ( \21338 , \18804 );
or \U$20996 ( \21339 , \21337 , \21338 );
not \U$20997 ( \21340 , \18787 );
nand \U$20998 ( \21341 , \21340 , \18800 );
nand \U$20999 ( \21342 , \21339 , \21341 );
not \U$21000 ( \21343 , \20795 );
not \U$21001 ( \21344 , \20815 );
nand \U$21002 ( \21345 , \21344 , \20805 );
not \U$21003 ( \21346 , \21345 );
or \U$21004 ( \21347 , \21343 , \21346 );
nand \U$21005 ( \21348 , \20815 , \20804 );
nand \U$21006 ( \21349 , \21347 , \21348 );
xor \U$21007 ( \21350 , \20760 , \20772 );
and \U$21008 ( \21351 , \21350 , \20784 );
and \U$21009 ( \21352 , \20760 , \20772 );
or \U$21010 ( \21353 , \21351 , \21352 );
nor \U$21011 ( \21354 , \21349 , \21353 );
not \U$21012 ( \21355 , \21354 );
nand \U$21013 ( \21356 , \21353 , \21349 );
nand \U$21014 ( \21357 , \21355 , \21356 );
not \U$21015 ( \21358 , \21357 );
and \U$21016 ( \21359 , \21342 , \21358 );
not \U$21017 ( \21360 , \21342 );
and \U$21018 ( \21361 , \21360 , \21357 );
nor \U$21019 ( \21362 , \21359 , \21361 );
not \U$21020 ( \21363 , \17606 );
not \U$21021 ( \21364 , \17596 );
or \U$21022 ( \21365 , \21363 , \21364 );
not \U$21023 ( \21366 , \17594 );
nand \U$21024 ( \21367 , \21366 , \17581 );
nand \U$21025 ( \21368 , \21365 , \21367 );
not \U$21026 ( \21369 , \3465 );
not \U$21027 ( \21370 , \18813 );
or \U$21028 ( \21371 , \21369 , \21370 );
and \U$21029 ( \21372 , RI98726d0_159, \7541 );
not \U$21030 ( \21373 , RI98726d0_159);
and \U$21031 ( \21374 , \21373 , \6059 );
nor \U$21032 ( \21375 , \21372 , \21374 );
nand \U$21033 ( \21376 , \21375 , \3467 );
nand \U$21034 ( \21377 , \21371 , \21376 );
not \U$21035 ( \21378 , \21377 );
not \U$21036 ( \21379 , \875 );
not \U$21037 ( \21380 , \20782 );
or \U$21038 ( \21381 , \21379 , \21380 );
not \U$21039 ( \21382 , RI9872130_147);
not \U$21040 ( \21383 , \12460 );
or \U$21041 ( \21384 , \21382 , \21383 );
or \U$21042 ( \21385 , \9850 , RI9872130_147);
nand \U$21043 ( \21386 , \21384 , \21385 );
nand \U$21044 ( \21387 , \21386 , \924 );
nand \U$21045 ( \21388 , \21381 , \21387 );
not \U$21046 ( \21389 , \20800 );
not \U$21047 ( \21390 , \1379 );
or \U$21048 ( \21391 , \21389 , \21390 );
not \U$21049 ( \21392 , \11453 );
not \U$21050 ( \21393 , \21392 );
and \U$21051 ( \21394 , RI9871e60_141, \21393 );
not \U$21052 ( \21395 , RI9871e60_141);
and \U$21053 ( \21396 , \21395 , \12783 );
or \U$21054 ( \21397 , \21394 , \21396 );
nand \U$21055 ( \21398 , \21397 , \1352 );
nand \U$21056 ( \21399 , \21391 , \21398 );
xnor \U$21057 ( \21400 , \21388 , \21399 );
not \U$21058 ( \21401 , \21400 );
and \U$21059 ( \21402 , \21378 , \21401 );
and \U$21060 ( \21403 , \21377 , \21400 );
nor \U$21061 ( \21404 , \21402 , \21403 );
not \U$21062 ( \21405 , \21404 );
and \U$21063 ( \21406 , \21368 , \21405 );
not \U$21064 ( \21407 , \21368 );
and \U$21065 ( \21408 , \21407 , \21404 );
nor \U$21066 ( \21409 , \21406 , \21408 );
xor \U$21067 ( \21410 , \17616 , \17623 );
and \U$21068 ( \21411 , \21410 , \17634 );
and \U$21069 ( \21412 , \17616 , \17623 );
or \U$21070 ( \21413 , \21411 , \21412 );
and \U$21071 ( \21414 , \21409 , \21413 );
not \U$21072 ( \21415 , \21409 );
not \U$21073 ( \21416 , \21413 );
and \U$21074 ( \21417 , \21415 , \21416 );
nor \U$21075 ( \21418 , \21414 , \21417 );
xor \U$21076 ( \21419 , \21362 , \21418 );
not \U$21077 ( \21420 , \20847 );
not \U$21078 ( \21421 , \20843 );
not \U$21079 ( \21422 , \20852 );
or \U$21080 ( \21423 , \21421 , \21422 );
or \U$21081 ( \21424 , \20852 , \20843 );
nand \U$21082 ( \21425 , \21423 , \21424 );
not \U$21083 ( \21426 , \21425 );
or \U$21084 ( \21427 , \21420 , \21426 );
not \U$21085 ( \21428 , \20843 );
nand \U$21086 ( \21429 , \21428 , \20852 );
nand \U$21087 ( \21430 , \21427 , \21429 );
xor \U$21088 ( \21431 , \21419 , \21430 );
xor \U$21089 ( \21432 , \20835 , \20825 );
and \U$21090 ( \21433 , \21432 , \20853 );
and \U$21091 ( \21434 , \20835 , \20825 );
nor \U$21092 ( \21435 , \21433 , \21434 );
nor \U$21093 ( \21436 , \21431 , \21435 );
not \U$21094 ( \21437 , \21436 );
nand \U$21095 ( \21438 , \21435 , \21431 );
nand \U$21096 ( \21439 , \21437 , \21438 );
xor \U$21097 ( \21440 , \17437 , \17570 );
and \U$21098 ( \21441 , \21440 , \17676 );
and \U$21099 ( \21442 , \17437 , \17570 );
or \U$21100 ( \21443 , \21441 , \21442 );
not \U$21101 ( \21444 , \21443 );
and \U$21102 ( \21445 , \21439 , \21444 );
not \U$21103 ( \21446 , \21439 );
and \U$21104 ( \21447 , \21446 , \21443 );
nor \U$21105 ( \21448 , \21445 , \21447 );
xor \U$21106 ( \21449 , \21336 , \21448 );
not \U$21107 ( \21450 , \21449 );
xor \U$21108 ( \21451 , \17322 , \17943 );
and \U$21109 ( \21452 , \21451 , \17677 );
and \U$21110 ( \21453 , \17322 , \17943 );
nor \U$21111 ( \21454 , \21452 , \21453 );
not \U$21112 ( \21455 , \21454 );
and \U$21113 ( \21456 , \21450 , \21455 );
and \U$21114 ( \21457 , \21449 , \21454 );
nor \U$21115 ( \21458 , \21456 , \21457 );
not \U$21116 ( \21459 , \21458 );
or \U$21117 ( \21460 , \21331 , \21459 );
or \U$21118 ( \21461 , \21330 , \21458 );
nand \U$21119 ( \21462 , \21460 , \21461 );
buf \U$21120 ( \21463 , \21462 );
or \U$21121 ( \21464 , \19228 , \17945 );
nand \U$21122 ( \21465 , \21464 , \18780 );
nand \U$21123 ( \21466 , \19228 , \17945 );
nand \U$21124 ( \21467 , \21465 , \21466 );
buf \U$21125 ( \21468 , \21467 );
not \U$21126 ( \21469 , \21468 );
and \U$21127 ( \21470 , \21463 , \21469 );
not \U$21128 ( \21471 , \21463 );
and \U$21129 ( \21472 , \21471 , \21468 );
nor \U$21130 ( \21473 , \21470 , \21472 );
nor \U$21131 ( \21474 , \21320 , \21473 );
not \U$21132 ( \21475 , \21474 );
nand \U$21133 ( \21476 , \21320 , \21473 );
nand \U$21134 ( \21477 , \21475 , \21476 );
not \U$21135 ( \21478 , \21477 );
or \U$21136 ( \21479 , \20900 , \21478 );
xor \U$21137 ( \21480 , \19229 , \20737 );
xor \U$21138 ( \21481 , \21480 , \20895 );
buf \U$21139 ( \21482 , \19837 );
not \U$21140 ( \21483 , \19842 );
and \U$21141 ( \21484 , \21482 , \21483 );
not \U$21142 ( \21485 , \21482 );
and \U$21143 ( \21486 , \21485 , \19842 );
nor \U$21144 ( \21487 , \21484 , \21486 );
not \U$21145 ( \21488 , \21487 );
not \U$21146 ( \21489 , \21488 );
xor \U$21147 ( \21490 , \19475 , \19493 );
xnor \U$21148 ( \21491 , \21490 , \19831 );
not \U$21149 ( \21492 , \21491 );
not \U$21150 ( \21493 , \21492 );
not \U$21151 ( \21494 , \20233 );
and \U$21152 ( \21495 , \20230 , \21494 );
not \U$21153 ( \21496 , \20230 );
and \U$21154 ( \21497 , \21496 , \20233 );
nor \U$21155 ( \21498 , \21495 , \21497 );
not \U$21156 ( \21499 , \21498 );
xor \U$21157 ( \21500 , \19903 , \19918 );
xnor \U$21158 ( \21501 , \21500 , \19921 );
not \U$21159 ( \21502 , \21501 );
or \U$21160 ( \21503 , \21499 , \21502 );
or \U$21161 ( \21504 , \21501 , \21498 );
nand \U$21162 ( \21505 , \21503 , \21504 );
not \U$21163 ( \21506 , \21505 );
or \U$21164 ( \21507 , \21493 , \21506 );
not \U$21165 ( \21508 , \21498 );
nand \U$21166 ( \21509 , \21508 , \21501 );
nand \U$21167 ( \21510 , \21507 , \21509 );
not \U$21168 ( \21511 , \21510 );
xnor \U$21169 ( \21512 , \20562 , \20591 );
not \U$21170 ( \21513 , \21512 );
not \U$21171 ( \21514 , \5847 );
not \U$21172 ( \21515 , \20439 );
or \U$21173 ( \21516 , \21514 , \21515 );
not \U$21174 ( \21517 , RI98725e0_157);
not \U$21175 ( \21518 , \9598 );
not \U$21176 ( \21519 , \21518 );
or \U$21177 ( \21520 , \21517 , \21519 );
or \U$21178 ( \21521 , \8074 , RI98725e0_157);
nand \U$21179 ( \21522 , \21520 , \21521 );
nand \U$21180 ( \21523 , \21522 , \18171 );
nand \U$21181 ( \21524 , \21516 , \21523 );
not \U$21182 ( \21525 , \21524 );
not \U$21183 ( \21526 , \924 );
not \U$21184 ( \21527 , \20452 );
or \U$21185 ( \21528 , \21526 , \21527 );
buf \U$21186 ( \21529 , \17741 );
and \U$21187 ( \21530 , RI9872130_147, \21529 );
not \U$21188 ( \21531 , RI9872130_147);
and \U$21189 ( \21532 , \21531 , \17912 );
or \U$21190 ( \21533 , \21530 , \21532 );
nand \U$21191 ( \21534 , \21533 , \875 );
nand \U$21192 ( \21535 , \21528 , \21534 );
not \U$21193 ( \21536 , \21535 );
not \U$21194 ( \21537 , \19383 );
not \U$21195 ( \21538 , \1043 );
or \U$21196 ( \21539 , \21537 , \21538 );
or \U$21197 ( \21540 , \18218 , \19383 );
nand \U$21198 ( \21541 , \21539 , \21540 );
not \U$21199 ( \21542 , \21541 );
not \U$21200 ( \21543 , \1016 );
or \U$21201 ( \21544 , \21542 , \21543 );
nand \U$21202 ( \21545 , \20471 , \1013 );
nand \U$21203 ( \21546 , \21544 , \21545 );
not \U$21204 ( \21547 , \832 );
not \U$21205 ( \21548 , \20475 );
or \U$21206 ( \21549 , \21547 , \21548 );
not \U$21207 ( \21550 , RI9871d70_139);
not \U$21208 ( \21551 , \16996 );
or \U$21209 ( \21552 , \21550 , \21551 );
not \U$21210 ( \21553 , \16995 );
or \U$21211 ( \21554 , \21553 , RI9871d70_139);
nand \U$21212 ( \21555 , \21552 , \21554 );
nand \U$21213 ( \21556 , \21555 , \859 );
nand \U$21214 ( \21557 , \21549 , \21556 );
xor \U$21215 ( \21558 , \21546 , \21557 );
not \U$21216 ( \21559 , \21558 );
or \U$21217 ( \21560 , \21536 , \21559 );
nand \U$21218 ( \21561 , \21546 , \21557 );
nand \U$21219 ( \21562 , \21560 , \21561 );
not \U$21220 ( \21563 , \21562 );
not \U$21221 ( \21564 , \21563 );
not \U$21222 ( \21565 , \3464 );
not \U$21223 ( \21566 , RI98726d0_159);
not \U$21224 ( \21567 , \18110 );
or \U$21225 ( \21568 , \21566 , \21567 );
or \U$21226 ( \21569 , \8607 , RI98726d0_159);
nand \U$21227 ( \21570 , \21568 , \21569 );
not \U$21228 ( \21571 , \21570 );
or \U$21229 ( \21572 , \21565 , \21571 );
nand \U$21230 ( \21573 , \20432 , \3467 );
nand \U$21231 ( \21574 , \21572 , \21573 );
not \U$21232 ( \21575 , \21574 );
or \U$21233 ( \21576 , \21564 , \21575 );
or \U$21234 ( \21577 , \21574 , \21563 );
nand \U$21235 ( \21578 , \21576 , \21577 );
not \U$21236 ( \21579 , \21578 );
or \U$21237 ( \21580 , \21525 , \21579 );
not \U$21238 ( \21581 , \21563 );
nand \U$21239 ( \21582 , \21581 , \21574 );
nand \U$21240 ( \21583 , \21580 , \21582 );
not \U$21241 ( \21584 , \2071 );
not \U$21242 ( \21585 , RI9871aa0_133);
not \U$21243 ( \21586 , \10369 );
or \U$21244 ( \21587 , \21585 , \21586 );
or \U$21245 ( \21588 , \13298 , RI9871aa0_133);
nand \U$21246 ( \21589 , \21587 , \21588 );
not \U$21247 ( \21590 , \21589 );
or \U$21248 ( \21591 , \21584 , \21590 );
nand \U$21249 ( \21592 , \20402 , \2087 );
nand \U$21250 ( \21593 , \21591 , \21592 );
not \U$21251 ( \21594 , \21593 );
not \U$21252 ( \21595 , \6144 );
not \U$21253 ( \21596 , \20388 );
or \U$21254 ( \21597 , \21595 , \21596 );
not \U$21255 ( \21598 , \1078 );
not \U$21256 ( \21599 , \8695 );
or \U$21257 ( \21600 , \21598 , \21599 );
or \U$21258 ( \21601 , \9750 , \1078 );
nand \U$21259 ( \21602 , \21600 , \21601 );
nand \U$21260 ( \21603 , \21602 , \11432 );
nand \U$21261 ( \21604 , \21597 , \21603 );
not \U$21262 ( \21605 , \21604 );
not \U$21263 ( \21606 , \21605 );
not \U$21264 ( \21607 , \3163 );
not \U$21265 ( \21608 , RI9872310_151);
not \U$21266 ( \21609 , \11406 );
or \U$21267 ( \21610 , \21608 , \21609 );
or \U$21268 ( \21611 , \11406 , RI9872310_151);
nand \U$21269 ( \21612 , \21610 , \21611 );
not \U$21270 ( \21613 , \21612 );
or \U$21271 ( \21614 , \21607 , \21613 );
nand \U$21272 ( \21615 , \20418 , \12514 );
nand \U$21273 ( \21616 , \21614 , \21615 );
not \U$21274 ( \21617 , \21616 );
or \U$21275 ( \21618 , \21606 , \21617 );
or \U$21276 ( \21619 , \21616 , \21605 );
nand \U$21277 ( \21620 , \21618 , \21619 );
not \U$21278 ( \21621 , \21620 );
or \U$21279 ( \21622 , \21594 , \21621 );
nand \U$21280 ( \21623 , \21616 , \21604 );
nand \U$21281 ( \21624 , \21622 , \21623 );
or \U$21282 ( \21625 , \21583 , \21624 );
not \U$21283 ( \21626 , \1083 );
and \U$21284 ( \21627 , RI98718c0_129, \9114 );
not \U$21285 ( \21628 , RI98718c0_129);
and \U$21286 ( \21629 , \21628 , \18344 );
or \U$21287 ( \21630 , \21627 , \21629 );
not \U$21288 ( \21631 , \21630 );
or \U$21289 ( \21632 , \21626 , \21631 );
nand \U$21290 ( \21633 , \20376 , \1135 );
nand \U$21291 ( \21634 , \21632 , \21633 );
not \U$21292 ( \21635 , \21634 );
not \U$21293 ( \21636 , \21635 );
not \U$21294 ( \21637 , \4919 );
not \U$21295 ( \21638 , RI9872388_152);
not \U$21296 ( \21639 , \7466 );
or \U$21297 ( \21640 , \21638 , \21639 );
not \U$21298 ( \21641 , \7465 );
not \U$21299 ( \21642 , \21641 );
or \U$21300 ( \21643 , \21642 , RI9872388_152);
nand \U$21301 ( \21644 , \21640 , \21643 );
not \U$21302 ( \21645 , \21644 );
or \U$21303 ( \21646 , \21637 , \21645 );
nand \U$21304 ( \21647 , \20585 , \4923 );
nand \U$21305 ( \21648 , \21646 , \21647 );
not \U$21306 ( \21649 , \21648 );
not \U$21307 ( \21650 , \21649 );
or \U$21308 ( \21651 , \21636 , \21650 );
not \U$21309 ( \21652 , \5034 );
not \U$21310 ( \21653 , \5025 );
not \U$21311 ( \21654 , \18793 );
or \U$21312 ( \21655 , \21653 , \21654 );
or \U$21313 ( \21656 , \5025 , \6528 );
nand \U$21314 ( \21657 , \21655 , \21656 );
not \U$21315 ( \21658 , \21657 );
or \U$21316 ( \21659 , \21652 , \21658 );
nand \U$21317 ( \21660 , \20367 , \5796 );
nand \U$21318 ( \21661 , \21659 , \21660 );
nand \U$21319 ( \21662 , \21651 , \21661 );
nand \U$21320 ( \21663 , \21648 , \21634 );
nand \U$21321 ( \21664 , \21662 , \21663 );
nand \U$21322 ( \21665 , \21625 , \21664 );
nand \U$21323 ( \21666 , \21583 , \21624 );
nand \U$21324 ( \21667 , \21665 , \21666 );
not \U$21325 ( \21668 , \21667 );
not \U$21326 ( \21669 , \21668 );
or \U$21327 ( \21670 , \21513 , \21669 );
xor \U$21328 ( \21671 , \18696 , \18729 );
xnor \U$21329 ( \21672 , \21671 , \18741 );
not \U$21330 ( \21673 , \21672 );
nand \U$21331 ( \21674 , \21670 , \21673 );
not \U$21332 ( \21675 , \21512 );
nand \U$21333 ( \21676 , \21675 , \21667 );
nand \U$21334 ( \21677 , \21674 , \21676 );
xor \U$21335 ( \21678 , \19906 , \19912 );
xor \U$21336 ( \21679 , \21678 , \19915 );
xor \U$21337 ( \21680 , \21677 , \21679 );
xor \U$21338 ( \21681 , \19894 , \19897 );
xor \U$21339 ( \21682 , \21681 , \19896 );
and \U$21340 ( \21683 , \21680 , \21682 );
and \U$21341 ( \21684 , \21677 , \21679 );
or \U$21342 ( \21685 , \21683 , \21684 );
not \U$21343 ( \21686 , \21685 );
not \U$21344 ( \21687 , \18754 );
not \U$21345 ( \21688 , \18628 );
and \U$21346 ( \21689 , \21687 , \21688 );
and \U$21347 ( \21690 , \18754 , \18628 );
nor \U$21348 ( \21691 , \21689 , \21690 );
not \U$21349 ( \21692 , \21691 );
xor \U$21350 ( \21693 , \18632 , \18680 );
xnor \U$21351 ( \21694 , \21693 , \18749 );
not \U$21352 ( \21695 , \21694 );
not \U$21353 ( \21696 , \18528 );
not \U$21354 ( \21697 , \18483 );
or \U$21355 ( \21698 , \21696 , \21697 );
nand \U$21356 ( \21699 , \18529 , \18482 );
nand \U$21357 ( \21700 , \21698 , \21699 );
xor \U$21358 ( \21701 , \21700 , \18587 );
not \U$21359 ( \21702 , \21701 );
xor \U$21360 ( \21703 , \20202 , \20187 );
xnor \U$21361 ( \21704 , \21703 , \20198 );
nand \U$21362 ( \21705 , \21702 , \21704 );
not \U$21363 ( \21706 , \21705 );
or \U$21364 ( \21707 , \21695 , \21706 );
not \U$21365 ( \21708 , \21704 );
nand \U$21366 ( \21709 , \21708 , \21701 );
nand \U$21367 ( \21710 , \21707 , \21709 );
not \U$21368 ( \21711 , \21710 );
and \U$21369 ( \21712 , \21692 , \21711 );
and \U$21370 ( \21713 , \21710 , \21691 );
nor \U$21371 ( \21714 , \21712 , \21713 );
not \U$21372 ( \21715 , \21714 );
not \U$21373 ( \21716 , \21715 );
or \U$21374 ( \21717 , \21686 , \21716 );
not \U$21375 ( \21718 , \21691 );
nand \U$21376 ( \21719 , \21718 , \21710 );
nand \U$21377 ( \21720 , \21717 , \21719 );
not \U$21378 ( \21721 , \21720 );
not \U$21379 ( \21722 , \21721 );
or \U$21380 ( \21723 , \21511 , \21722 );
or \U$21381 ( \21724 , \21721 , \21510 );
nand \U$21382 ( \21725 , \21723 , \21724 );
not \U$21383 ( \21726 , \21725 );
or \U$21384 ( \21727 , \21489 , \21726 );
nand \U$21385 ( \21728 , \21720 , \21510 );
nand \U$21386 ( \21729 , \21727 , \21728 );
not \U$21387 ( \21730 , \19940 );
not \U$21388 ( \21731 , \20731 );
not \U$21389 ( \21732 , \21731 );
or \U$21390 ( \21733 , \21730 , \21732 );
not \U$21391 ( \21734 , \19940 );
nand \U$21392 ( \21735 , \21734 , \20731 );
nand \U$21393 ( \21736 , \21733 , \21735 );
xor \U$21394 ( \21737 , \21729 , \21736 );
xor \U$21395 ( \21738 , \21704 , \21701 );
xor \U$21396 ( \21739 , \21694 , \21738 );
not \U$21397 ( \21740 , \21739 );
not \U$21398 ( \21741 , \21740 );
xor \U$21399 ( \21742 , \20254 , \20264 );
xor \U$21400 ( \21743 , \21742 , \20268 );
xor \U$21401 ( \21744 , \20342 , \20274 );
xnor \U$21402 ( \21745 , \21744 , \20272 );
xor \U$21403 ( \21746 , \21743 , \21745 );
xor \U$21404 ( \21747 , \19783 , \19797 );
xnor \U$21405 ( \21748 , \21747 , \19817 );
not \U$21406 ( \21749 , \21748 );
not \U$21407 ( \21750 , \21749 );
xor \U$21408 ( \21751 , \20288 , \20324 );
xnor \U$21409 ( \21752 , \21751 , \20307 );
not \U$21410 ( \21753 , \21752 );
xor \U$21411 ( \21754 , \20502 , \20507 );
not \U$21412 ( \21755 , \832 );
not \U$21413 ( \21756 , \21555 );
or \U$21414 ( \21757 , \21755 , \21756 );
not \U$21415 ( \21758 , \8859 );
not \U$21416 ( \21759 , \17702 );
or \U$21417 ( \21760 , \21758 , \21759 );
nand \U$21418 ( \21761 , \20490 , RI9871d70_139);
nand \U$21419 ( \21762 , \21760 , \21761 );
nand \U$21420 ( \21763 , \21762 , \858 );
nand \U$21421 ( \21764 , \21757 , \21763 );
not \U$21422 ( \21765 , \21764 );
not \U$21423 ( \21766 , \20499 );
not \U$21424 ( \21767 , \1374 );
and \U$21425 ( \21768 , \21766 , \21767 );
not \U$21426 ( \21769 , RI9871e60_141);
not \U$21427 ( \21770 , \18193 );
or \U$21428 ( \21771 , \21769 , \21770 );
buf \U$21429 ( \21772 , \18192 );
buf \U$21430 ( \21773 , \21772 );
or \U$21431 ( \21774 , \21773 , RI9871e60_141);
nand \U$21432 ( \21775 , \21771 , \21774 );
and \U$21433 ( \21776 , \21775 , \1379 );
nor \U$21434 ( \21777 , \21768 , \21776 );
not \U$21435 ( \21778 , \18704 );
not \U$21436 ( \21779 , \21778 );
and \U$21437 ( \21780 , \21779 , \1013 );
not \U$21438 ( \21781 , \21780 );
and \U$21439 ( \21782 , \21777 , \21781 );
not \U$21440 ( \21783 , \21777 );
and \U$21441 ( \21784 , \21783 , \21780 );
nor \U$21442 ( \21785 , \21782 , \21784 );
not \U$21443 ( \21786 , \21785 );
or \U$21444 ( \21787 , \21765 , \21786 );
not \U$21445 ( \21788 , \21777 );
nand \U$21446 ( \21789 , \21788 , \21780 );
nand \U$21447 ( \21790 , \21787 , \21789 );
xor \U$21448 ( \21791 , \21754 , \21790 );
not \U$21449 ( \21792 , \21791 );
not \U$21450 ( \21793 , \1323 );
not \U$21451 ( \21794 , \20316 );
or \U$21452 ( \21795 , \21793 , \21794 );
not \U$21453 ( \21796 , RI9871b18_134);
not \U$21454 ( \21797 , \17090 );
or \U$21455 ( \21798 , \21796 , \21797 );
nand \U$21456 ( \21799 , \13281 , \2479 );
nand \U$21457 ( \21800 , \21798 , \21799 );
nand \U$21458 ( \21801 , \21800 , \1292 );
nand \U$21459 ( \21802 , \21795 , \21801 );
not \U$21460 ( \21803 , \21802 );
or \U$21461 ( \21804 , \21792 , \21803 );
nand \U$21462 ( \21805 , \21790 , \21754 );
nand \U$21463 ( \21806 , \21804 , \21805 );
not \U$21464 ( \21807 , \21806 );
not \U$21465 ( \21808 , \21807 );
or \U$21466 ( \21809 , \21753 , \21808 );
not \U$21467 ( \21810 , \1136 );
not \U$21468 ( \21811 , \21630 );
or \U$21469 ( \21812 , \21810 , \21811 );
and \U$21470 ( \21813 , RI98718c0_129, \12597 );
not \U$21471 ( \21814 , RI98718c0_129);
and \U$21472 ( \21815 , \21814 , \12594 );
or \U$21473 ( \21816 , \21813 , \21815 );
nand \U$21474 ( \21817 , \21816 , \1083 );
nand \U$21475 ( \21818 , \21812 , \21817 );
not \U$21476 ( \21819 , \21818 );
not \U$21477 ( \21820 , \1518 );
not \U$21478 ( \21821 , \20286 );
or \U$21479 ( \21822 , \21820 , \21821 );
not \U$21480 ( \21823 , RI9871c80_137);
not \U$21481 ( \21824 , \17013 );
or \U$21482 ( \21825 , \21823 , \21824 );
or \U$21483 ( \21826 , \13860 , RI9871c80_137);
nand \U$21484 ( \21827 , \21825 , \21826 );
nand \U$21485 ( \21828 , \21827 , \1500 );
nand \U$21486 ( \21829 , \21822 , \21828 );
not \U$21487 ( \21830 , \21829 );
nand \U$21488 ( \21831 , \20296 , \1429 );
xor \U$21489 ( \21832 , RI9871c08_136, \12787 );
nand \U$21490 ( \21833 , \21832 , \1455 );
nand \U$21491 ( \21834 , \21831 , \21833 );
not \U$21492 ( \21835 , \21834 );
not \U$21493 ( \21836 , \21835 );
or \U$21494 ( \21837 , \21830 , \21836 );
not \U$21495 ( \21838 , \21833 );
not \U$21496 ( \21839 , \21831 );
or \U$21497 ( \21840 , \21838 , \21839 );
not \U$21498 ( \21841 , \21829 );
nand \U$21499 ( \21842 , \21840 , \21841 );
nand \U$21500 ( \21843 , \21837 , \21842 );
not \U$21501 ( \21844 , \21843 );
or \U$21502 ( \21845 , \21819 , \21844 );
nand \U$21503 ( \21846 , \21834 , \21829 );
nand \U$21504 ( \21847 , \21845 , \21846 );
nand \U$21505 ( \21848 , \21809 , \21847 );
not \U$21506 ( \21849 , \21752 );
nand \U$21507 ( \21850 , \21849 , \21806 );
and \U$21508 ( \21851 , \21848 , \21850 );
xor \U$21509 ( \21852 , \20666 , \21851 );
xnor \U$21510 ( \21853 , \21852 , \20694 );
not \U$21511 ( \21854 , \21853 );
or \U$21512 ( \21855 , \21750 , \21854 );
not \U$21513 ( \21856 , \20694 );
not \U$21514 ( \21857 , \20666 );
not \U$21515 ( \21858 , \21857 );
and \U$21516 ( \21859 , \21856 , \21858 );
and \U$21517 ( \21860 , \20694 , \21857 );
nor \U$21518 ( \21861 , \21859 , \21860 );
or \U$21519 ( \21862 , \21851 , \21861 );
nand \U$21520 ( \21863 , \21855 , \21862 );
and \U$21521 ( \21864 , \21746 , \21863 );
and \U$21522 ( \21865 , \21743 , \21745 );
or \U$21523 ( \21866 , \21864 , \21865 );
not \U$21524 ( \21867 , \21866 );
or \U$21525 ( \21868 , \21741 , \21867 );
xor \U$21526 ( \21869 , \21677 , \21679 );
xor \U$21527 ( \21870 , \21869 , \21682 );
not \U$21528 ( \21871 , \21866 );
nand \U$21529 ( \21872 , \21871 , \21739 );
nand \U$21530 ( \21873 , \21870 , \21872 );
nand \U$21531 ( \21874 , \21868 , \21873 );
not \U$21532 ( \21875 , \21874 );
xor \U$21533 ( \21876 , \19738 , \19772 );
xor \U$21534 ( \21877 , \21876 , \19819 );
and \U$21535 ( \21878 , \19512 , \19623 );
not \U$21536 ( \21879 , \19512 );
and \U$21537 ( \21880 , \21879 , \19622 );
nor \U$21538 ( \21881 , \21878 , \21880 );
xnor \U$21539 ( \21882 , \19575 , \19559 );
xor \U$21540 ( \21883 , \21881 , \21882 );
not \U$21541 ( \21884 , \21883 );
and \U$21542 ( \21885 , \19661 , \21884 );
not \U$21543 ( \21886 , \19661 );
and \U$21544 ( \21887 , \21886 , \21883 );
nor \U$21545 ( \21888 , \21885 , \21887 );
not \U$21546 ( \21889 , \21888 );
or \U$21547 ( \21890 , \21877 , \21889 );
not \U$21548 ( \21891 , \20434 );
not \U$21549 ( \21892 , \20421 );
or \U$21550 ( \21893 , \21891 , \21892 );
or \U$21551 ( \21894 , \20421 , \20434 );
nand \U$21552 ( \21895 , \21893 , \21894 );
buf \U$21553 ( \21896 , \20404 );
and \U$21554 ( \21897 , \21895 , \21896 );
not \U$21555 ( \21898 , \21895 );
not \U$21556 ( \21899 , \21896 );
and \U$21557 ( \21900 , \21898 , \21899 );
nor \U$21558 ( \21901 , \21897 , \21900 );
not \U$21559 ( \21902 , \21901 );
xor \U$21560 ( \21903 , \20443 , \20526 );
not \U$21561 ( \21904 , \21903 );
or \U$21562 ( \21905 , \21902 , \21904 );
or \U$21563 ( \21906 , \21901 , \21903 );
xor \U$21564 ( \21907 , \20326 , \20328 );
xor \U$21565 ( \21908 , \21907 , \20339 );
nand \U$21566 ( \21909 , \21906 , \21908 );
nand \U$21567 ( \21910 , \21905 , \21909 );
nand \U$21568 ( \21911 , \21890 , \21910 );
nand \U$21569 ( \21912 , \21877 , \21889 );
nand \U$21570 ( \21913 , \21911 , \21912 );
not \U$21571 ( \21914 , \19643 );
not \U$21572 ( \21915 , \19659 );
not \U$21573 ( \21916 , \19655 );
and \U$21574 ( \21917 , \21915 , \21916 );
and \U$21575 ( \21918 , \19655 , \19659 );
nor \U$21576 ( \21919 , \21917 , \21918 );
not \U$21577 ( \21920 , \21919 );
and \U$21578 ( \21921 , \21914 , \21920 );
and \U$21579 ( \21922 , \19643 , \21919 );
nor \U$21580 ( \21923 , \21921 , \21922 );
not \U$21581 ( \21924 , \21923 );
xor \U$21582 ( \21925 , \20604 , \20615 );
xor \U$21583 ( \21926 , \21925 , \20622 );
or \U$21584 ( \21927 , \21924 , \21926 );
xor \U$21585 ( \21928 , \20644 , \20653 );
xor \U$21586 ( \21929 , \21928 , \20632 );
nand \U$21587 ( \21930 , \21927 , \21929 );
nand \U$21588 ( \21931 , \21926 , \21924 );
nand \U$21589 ( \21932 , \21930 , \21931 );
not \U$21590 ( \21933 , \21932 );
xor \U$21591 ( \21934 , \20625 , \20655 );
xor \U$21592 ( \21935 , \21934 , \20701 );
xor \U$21593 ( \21936 , \20574 , \20587 );
xor \U$21594 ( \21937 , \20545 , \20551 );
xnor \U$21595 ( \21938 , \21937 , \20540 );
xnor \U$21596 ( \21939 , \21936 , \21938 );
not \U$21597 ( \21940 , \21939 );
not \U$21598 ( \21941 , \9527 );
and \U$21599 ( \21942 , \6333 , \8732 );
not \U$21600 ( \21943 , \6333 );
and \U$21601 ( \21944 , \21943 , RI9872f40_177);
nor \U$21602 ( \21945 , \21942 , \21944 );
not \U$21603 ( \21946 , \21945 );
or \U$21604 ( \21947 , \21941 , \21946 );
nand \U$21605 ( \21948 , \19653 , \8752 );
nand \U$21606 ( \21949 , \21947 , \21948 );
not \U$21607 ( \21950 , \21949 );
not \U$21608 ( \21951 , \9320 );
not \U$21609 ( \21952 , RI9872568_156);
not \U$21610 ( \21953 , \11435 );
or \U$21611 ( \21954 , \21952 , \21953 );
not \U$21612 ( \21955 , \5703 );
not \U$21613 ( \21956 , \21955 );
nand \U$21614 ( \21957 , \21956 , \5644 );
nand \U$21615 ( \21958 , \21954 , \21957 );
not \U$21616 ( \21959 , \21958 );
or \U$21617 ( \21960 , \21951 , \21959 );
nand \U$21618 ( \21961 , \19632 , \5653 );
nand \U$21619 ( \21962 , \21960 , \21961 );
xor \U$21620 ( \21963 , \20521 , \20508 );
and \U$21621 ( \21964 , \21962 , \21963 );
not \U$21622 ( \21965 , \21962 );
not \U$21623 ( \21966 , \21963 );
and \U$21624 ( \21967 , \21965 , \21966 );
nor \U$21625 ( \21968 , \21964 , \21967 );
not \U$21626 ( \21969 , \21968 );
or \U$21627 ( \21970 , \21950 , \21969 );
nand \U$21628 ( \21971 , \21962 , \21963 );
nand \U$21629 ( \21972 , \21970 , \21971 );
not \U$21630 ( \21973 , \21972 );
or \U$21631 ( \21974 , \21940 , \21973 );
not \U$21632 ( \21975 , \20587 );
nor \U$21633 ( \21976 , \21975 , \20574 );
not \U$21634 ( \21977 , \20574 );
nor \U$21635 ( \21978 , \21977 , \20587 );
or \U$21636 ( \21979 , \21976 , \21978 );
not \U$21637 ( \21980 , \21938 );
nand \U$21638 ( \21981 , \21979 , \21980 );
nand \U$21639 ( \21982 , \21974 , \21981 );
and \U$21640 ( \21983 , \21935 , \21982 );
not \U$21641 ( \21984 , \21935 );
not \U$21642 ( \21985 , \21982 );
and \U$21643 ( \21986 , \21984 , \21985 );
nor \U$21644 ( \21987 , \21983 , \21986 );
not \U$21645 ( \21988 , \21987 );
or \U$21646 ( \21989 , \21933 , \21988 );
nand \U$21647 ( \21990 , \21935 , \21982 );
nand \U$21648 ( \21991 , \21989 , \21990 );
xor \U$21649 ( \21992 , \21913 , \21991 );
xor \U$21650 ( \21993 , \20270 , \20346 );
xor \U$21651 ( \21994 , \21993 , \20349 );
and \U$21652 ( \21995 , \21992 , \21994 );
and \U$21653 ( \21996 , \21913 , \21991 );
or \U$21654 ( \21997 , \21995 , \21996 );
not \U$21655 ( \21998 , \21997 );
nand \U$21656 ( \21999 , \21875 , \21998 );
not \U$21657 ( \22000 , \21999 );
not \U$21658 ( \22001 , \21491 );
not \U$21659 ( \22002 , \21505 );
or \U$21660 ( \22003 , \22001 , \22002 );
or \U$21661 ( \22004 , \21505 , \21491 );
nand \U$21662 ( \22005 , \22003 , \22004 );
not \U$21663 ( \22006 , \22005 );
or \U$21664 ( \22007 , \22000 , \22006 );
nand \U$21665 ( \22008 , \21874 , \21997 );
nand \U$21666 ( \22009 , \22007 , \22008 );
not \U$21667 ( \22010 , \22009 );
xor \U$21668 ( \22011 , \20713 , \20356 );
xnor \U$21669 ( \22012 , \22011 , \20352 );
not \U$21670 ( \22013 , \22012 );
not \U$21671 ( \22014 , \21714 );
not \U$21672 ( \22015 , \21685 );
and \U$21673 ( \22016 , \22014 , \22015 );
and \U$21674 ( \22017 , \21714 , \21685 );
nor \U$21675 ( \22018 , \22016 , \22017 );
not \U$21676 ( \22019 , \22018 );
or \U$21677 ( \22020 , \22013 , \22019 );
and \U$21678 ( \22021 , \19826 , \19666 );
not \U$21679 ( \22022 , \19826 );
not \U$21680 ( \22023 , \19666 );
and \U$21681 ( \22024 , \22022 , \22023 );
nor \U$21682 ( \22025 , \22021 , \22024 );
not \U$21683 ( \22026 , \22025 );
not \U$21684 ( \22027 , \6282 );
not \U$21685 ( \22028 , RI98728b0_163);
not \U$21686 ( \22029 , \5775 );
or \U$21687 ( \22030 , \22028 , \22029 );
or \U$21688 ( \22031 , \5775 , RI98728b0_163);
nand \U$21689 ( \22032 , \22030 , \22031 );
not \U$21690 ( \22033 , \22032 );
or \U$21691 ( \22034 , \22027 , \22033 );
nand \U$21692 ( \22035 , \20337 , \6285 );
nand \U$21693 ( \22036 , \22034 , \22035 );
not \U$21694 ( \22037 , \9072 );
not \U$21695 ( \22038 , \20600 );
or \U$21696 ( \22039 , \22037 , \22038 );
not \U$21697 ( \22040 , \8031 );
not \U$21698 ( \22041 , \4407 );
or \U$21699 ( \22042 , \22040 , \22041 );
not \U$21700 ( \22043 , \5205 );
or \U$21701 ( \22044 , \22043 , \8031 );
nand \U$21702 ( \22045 , \22042 , \22044 );
nand \U$21703 ( \22046 , \22045 , \8028 );
nand \U$21704 ( \22047 , \22039 , \22046 );
xor \U$21705 ( \22048 , \22036 , \22047 );
not \U$21706 ( \22049 , \12868 );
not \U$21707 ( \22050 , \20664 );
or \U$21708 ( \22051 , \22049 , \22050 );
xnor \U$21709 ( \22052 , RI98730a8_180, \18668 );
nand \U$21710 ( \22053 , \22052 , \13020 );
nand \U$21711 ( \22054 , \22051 , \22053 );
and \U$21712 ( \22055 , \22048 , \22054 );
and \U$21713 ( \22056 , \22036 , \22047 );
or \U$21714 ( \22057 , \22055 , \22056 );
not \U$21715 ( \22058 , \9312 );
not \U$21716 ( \22059 , RI9872d60_173);
not \U$21717 ( \22060 , \9162 );
or \U$21718 ( \22061 , \22059 , \22060 );
or \U$21719 ( \22062 , \6378 , RI9872d60_173);
nand \U$21720 ( \22063 , \22061 , \22062 );
not \U$21721 ( \22064 , \22063 );
or \U$21722 ( \22065 , \22058 , \22064 );
nand \U$21723 ( \22066 , \19795 , \10624 );
nand \U$21724 ( \22067 , \22065 , \22066 );
not \U$21725 ( \22068 , RI9873648_192);
not \U$21726 ( \22069 , \20628 );
or \U$21727 ( \22070 , \22068 , \22069 );
xor \U$21728 ( \22071 , RI9873558_190, \1105 );
nand \U$21729 ( \22072 , \22071 , \20626 );
nand \U$21730 ( \22073 , \22070 , \22072 );
xor \U$21731 ( \22074 , \22067 , \22073 );
not \U$21732 ( \22075 , \13484 );
not \U$21733 ( \22076 , \19815 );
or \U$21734 ( \22077 , \22075 , \22076 );
and \U$21735 ( \22078 , RI9873210_183, \846 );
not \U$21736 ( \22079 , RI9873210_183);
and \U$21737 ( \22080 , \22079 , \2215 );
nor \U$21738 ( \22081 , \22078 , \22080 );
nand \U$21739 ( \22082 , \22081 , \13476 );
nand \U$21740 ( \22083 , \22077 , \22082 );
and \U$21741 ( \22084 , \22074 , \22083 );
and \U$21742 ( \22085 , \22067 , \22073 );
or \U$21743 ( \22086 , \22084 , \22085 );
or \U$21744 ( \22087 , \22057 , \22086 );
not \U$21745 ( \22088 , \19036 );
not \U$21746 ( \22089 , RI98734e0_189);
not \U$21747 ( \22090 , \1446 );
or \U$21748 ( \22091 , \22089 , \22090 );
or \U$21749 ( \22092 , \1446 , RI98734e0_189);
nand \U$21750 ( \22093 , \22091 , \22092 );
not \U$21751 ( \22094 , \22093 );
or \U$21752 ( \22095 , \22088 , \22094 );
nand \U$21753 ( \22096 , \20651 , \20147 );
nand \U$21754 ( \22097 , \22095 , \22096 );
not \U$21755 ( \22098 , \22097 );
not \U$21756 ( \22099 , \18562 );
xnor \U$21757 ( \22100 , RI9872e50_175, \1190 );
not \U$21758 ( \22101 , \22100 );
or \U$21759 ( \22102 , \22099 , \22101 );
nand \U$21760 ( \22103 , \20642 , \10331 );
nand \U$21761 ( \22104 , \22102 , \22103 );
not \U$21762 ( \22105 , \22104 );
or \U$21763 ( \22106 , \22098 , \22105 );
or \U$21764 ( \22107 , \22097 , \22104 );
not \U$21765 ( \22108 , \18508 );
and \U$21766 ( \22109 , RI9873288_184, \9205 );
not \U$21767 ( \22110 , RI9873288_184);
and \U$21768 ( \22111 , \22110 , \6442 );
nor \U$21769 ( \22112 , \22109 , \22111 );
not \U$21770 ( \22113 , \22112 );
or \U$21771 ( \22114 , \22108 , \22113 );
nand \U$21772 ( \22115 , \19640 , \18522 );
nand \U$21773 ( \22116 , \22114 , \22115 );
nand \U$21774 ( \22117 , \22107 , \22116 );
nand \U$21775 ( \22118 , \22106 , \22117 );
nand \U$21776 ( \22119 , \22087 , \22118 );
nand \U$21777 ( \22120 , \22086 , \22057 );
nand \U$21778 ( \22121 , \22119 , \22120 );
not \U$21779 ( \22122 , \22121 );
xor \U$21780 ( \22123 , \20462 , \20480 );
not \U$21781 ( \22124 , \7325 );
xor \U$21782 ( \22125 , RI98729a0_165, \4959 );
not \U$21783 ( \22126 , \22125 );
or \U$21784 ( \22127 , \22124 , \22126 );
nand \U$21785 ( \22128 , \20620 , \7338 );
nand \U$21786 ( \22129 , \22127 , \22128 );
xor \U$21787 ( \22130 , \22123 , \22129 );
not \U$21788 ( \22131 , \19321 );
xor \U$21789 ( \22132 , RI9873030_179, \1365 );
not \U$21790 ( \22133 , \22132 );
or \U$21791 ( \22134 , \22131 , \22133 );
nand \U$21792 ( \22135 , \20613 , \9937 );
nand \U$21793 ( \22136 , \22134 , \22135 );
and \U$21794 ( \22137 , \22130 , \22136 );
and \U$21795 ( \22138 , \22123 , \22129 );
or \U$21796 ( \22139 , \22137 , \22138 );
not \U$21797 ( \22140 , \20369 );
xor \U$21798 ( \22141 , \20390 , \20378 );
not \U$21799 ( \22142 , \22141 );
and \U$21800 ( \22143 , \22140 , \22142 );
and \U$21801 ( \22144 , \20369 , \22141 );
nor \U$21802 ( \22145 , \22143 , \22144 );
xor \U$21803 ( \22146 , \22139 , \22145 );
not \U$21804 ( \22147 , \9196 );
not \U$21805 ( \22148 , \9198 );
not \U$21806 ( \22149 , \10698 );
or \U$21807 ( \22150 , \22148 , \22149 );
nand \U$21808 ( \22151 , \14930 , RI9872b80_169);
nand \U$21809 ( \22152 , \22150 , \22151 );
not \U$21810 ( \22153 , \22152 );
or \U$21811 ( \22154 , \22147 , \22153 );
nand \U$21812 ( \22155 , \20675 , \9214 );
nand \U$21813 ( \22156 , \22154 , \22155 );
not \U$21814 ( \22157 , \22156 );
not \U$21815 ( \22158 , \22157 );
not \U$21816 ( \22159 , \9249 );
not \U$21817 ( \22160 , RI9872bf8_170);
not \U$21818 ( \22161 , \3859 );
or \U$21819 ( \22162 , \22160 , \22161 );
or \U$21820 ( \22163 , \3859 , RI9872bf8_170);
nand \U$21821 ( \22164 , \22162 , \22163 );
not \U$21822 ( \22165 , \22164 );
or \U$21823 ( \22166 , \22159 , \22165 );
buf \U$21824 ( \22167 , \9226 );
nand \U$21825 ( \22168 , \19779 , \22167 );
nand \U$21826 ( \22169 , \22166 , \22168 );
not \U$21827 ( \22170 , \22169 );
not \U$21828 ( \22171 , \22170 );
or \U$21829 ( \22172 , \22158 , \22171 );
not \U$21830 ( \22173 , \17371 );
not \U$21831 ( \22174 , RI98733f0_187);
not \U$21832 ( \22175 , \1581 );
or \U$21833 ( \22176 , \22174 , \22175 );
or \U$21834 ( \22177 , \1581 , RI98733f0_187);
nand \U$21835 ( \22178 , \22176 , \22177 );
not \U$21836 ( \22179 , \22178 );
or \U$21837 ( \22180 , \22173 , \22179 );
nand \U$21838 ( \22181 , \20684 , \17263 );
nand \U$21839 ( \22182 , \22180 , \22181 );
nand \U$21840 ( \22183 , \22172 , \22182 );
nand \U$21841 ( \22184 , \22169 , \22156 );
nand \U$21842 ( \22185 , \22183 , \22184 );
and \U$21843 ( \22186 , \22146 , \22185 );
and \U$21844 ( \22187 , \22139 , \22145 );
or \U$21845 ( \22188 , \22186 , \22187 );
not \U$21846 ( \22189 , \22188 );
not \U$21847 ( \22190 , \20393 );
not \U$21848 ( \22191 , \20531 );
or \U$21849 ( \22192 , \22190 , \22191 );
or \U$21850 ( \22193 , \20531 , \20393 );
nand \U$21851 ( \22194 , \22192 , \22193 );
not \U$21852 ( \22195 , \22194 );
not \U$21853 ( \22196 , \22195 );
or \U$21854 ( \22197 , \22189 , \22196 );
not \U$21855 ( \22198 , \22188 );
nand \U$21856 ( \22199 , \22194 , \22198 );
nand \U$21857 ( \22200 , \22197 , \22199 );
not \U$21858 ( \22201 , \22200 );
or \U$21859 ( \22202 , \22122 , \22201 );
nand \U$21860 ( \22203 , \22194 , \22188 );
nand \U$21861 ( \22204 , \22202 , \22203 );
not \U$21862 ( \22205 , \22204 );
not \U$21863 ( \22206 , \22205 );
xor \U$21864 ( \22207 , \20597 , \20538 );
xnor \U$21865 ( \22208 , \22207 , \20704 );
not \U$21866 ( \22209 , \22208 );
or \U$21867 ( \22210 , \22206 , \22209 );
or \U$21868 ( \22211 , \22208 , \22205 );
nand \U$21869 ( \22212 , \22210 , \22211 );
not \U$21870 ( \22213 , \22212 );
or \U$21871 ( \22214 , \22026 , \22213 );
nand \U$21872 ( \22215 , \22208 , \22204 );
nand \U$21873 ( \22216 , \22214 , \22215 );
buf \U$21874 ( \22217 , \22216 );
nand \U$21875 ( \22218 , \22020 , \22217 );
not \U$21876 ( \22219 , \22012 );
not \U$21877 ( \22220 , \22018 );
nand \U$21878 ( \22221 , \22219 , \22220 );
nand \U$21879 ( \22222 , \22218 , \22221 );
not \U$21880 ( \22223 , \22222 );
or \U$21881 ( \22224 , \22010 , \22223 );
and \U$21882 ( \22225 , \22009 , \22222 );
not \U$21883 ( \22226 , \22009 );
and \U$21884 ( \22227 , \22221 , \22218 );
and \U$21885 ( \22228 , \22226 , \22227 );
nor \U$21886 ( \22229 , \22225 , \22228 );
xor \U$21887 ( \22230 , \20722 , \20249 );
nand \U$21888 ( \22231 , \22229 , \22230 );
nand \U$21889 ( \22232 , \22224 , \22231 );
and \U$21890 ( \22233 , \21737 , \22232 );
and \U$21891 ( \22234 , \21729 , \21736 );
or \U$21892 ( \22235 , \22233 , \22234 );
not \U$21893 ( \22236 , \22235 );
or \U$21894 ( \22237 , \21481 , \22236 );
xor \U$21895 ( \22238 , \21729 , \21736 );
xor \U$21896 ( \22239 , \22238 , \22232 );
not \U$21897 ( \22240 , \21725 );
not \U$21898 ( \22241 , \21487 );
and \U$21899 ( \22242 , \22240 , \22241 );
and \U$21900 ( \22243 , \21725 , \21487 );
nor \U$21901 ( \22244 , \22242 , \22243 );
not \U$21902 ( \22245 , \22244 );
not \U$21903 ( \22246 , \22230 );
and \U$21904 ( \22247 , \22229 , \22246 );
not \U$21905 ( \22248 , \22229 );
and \U$21906 ( \22249 , \22248 , \22230 );
nor \U$21907 ( \22250 , \22247 , \22249 );
not \U$21908 ( \22251 , \22250 );
or \U$21909 ( \22252 , \22245 , \22251 );
and \U$21910 ( \22253 , \21739 , \21866 );
not \U$21911 ( \22254 , \21739 );
and \U$21912 ( \22255 , \22254 , \21871 );
nor \U$21913 ( \22256 , \22253 , \22255 );
xnor \U$21914 ( \22257 , \22256 , \21870 );
not \U$21915 ( \22258 , \22257 );
not \U$21916 ( \22259 , \21932 );
not \U$21917 ( \22260 , \22259 );
not \U$21918 ( \22261 , \21987 );
or \U$21919 ( \22262 , \22260 , \22261 );
or \U$21920 ( \22263 , \21987 , \22259 );
nand \U$21921 ( \22264 , \22262 , \22263 );
not \U$21922 ( \22265 , \22264 );
xor \U$21923 ( \22266 , \21877 , \21910 );
xor \U$21924 ( \22267 , \22266 , \21888 );
nand \U$21925 ( \22268 , \22265 , \22267 );
not \U$21926 ( \22269 , \22268 );
nand \U$21927 ( \22270 , \18704 , \1349 );
nand \U$21928 ( \22271 , \22270 , \1350 , RI9871e60_141);
not \U$21929 ( \22272 , \22271 );
not \U$21930 ( \22273 , \1351 );
not \U$21931 ( \22274 , \21775 );
or \U$21932 ( \22275 , \22273 , \22274 );
and \U$21933 ( \22276 , RI9871e60_141, \18704 );
not \U$21934 ( \22277 , RI9871e60_141);
not \U$21935 ( \22278 , \18704 );
and \U$21936 ( \22279 , \22277 , \22278 );
nor \U$21937 ( \22280 , \22276 , \22279 );
nand \U$21938 ( \22281 , \22280 , \1379 );
nand \U$21939 ( \22282 , \22275 , \22281 );
nand \U$21940 ( \22283 , \22272 , \22282 );
not \U$21941 ( \22284 , \875 );
not \U$21942 ( \22285 , \17868 );
and \U$21943 ( \22286 , \22285 , \919 );
not \U$21944 ( \22287 , \22285 );
and \U$21945 ( \22288 , \22287 , RI9872130_147);
or \U$21946 ( \22289 , \22286 , \22288 );
not \U$21947 ( \22290 , \22289 );
or \U$21948 ( \22291 , \22284 , \22290 );
nand \U$21949 ( \22292 , \21533 , \924 );
nand \U$21950 ( \22293 , \22291 , \22292 );
xor \U$21951 ( \22294 , \22283 , \22293 );
not \U$21952 ( \22295 , \1500 );
not \U$21953 ( \22296 , RI9871c80_137);
not \U$21954 ( \22297 , \13934 );
or \U$21955 ( \22298 , \22296 , \22297 );
or \U$21956 ( \22299 , \20765 , RI9871c80_137);
nand \U$21957 ( \22300 , \22298 , \22299 );
not \U$21958 ( \22301 , \22300 );
or \U$21959 ( \22302 , \22295 , \22301 );
nand \U$21960 ( \22303 , \21827 , \1518 );
nand \U$21961 ( \22304 , \22302 , \22303 );
xnor \U$21962 ( \22305 , \22294 , \22304 );
not \U$21963 ( \22306 , \7326 );
and \U$21964 ( \22307 , \6185 , RI98729a0_165);
not \U$21965 ( \22308 , \6185 );
and \U$21966 ( \22309 , \22308 , \7333 );
nor \U$21967 ( \22310 , \22307 , \22309 );
not \U$21968 ( \22311 , \22310 );
or \U$21969 ( \22312 , \22306 , \22311 );
not \U$21970 ( \22313 , RI98729a0_165);
xor \U$21971 ( \22314 , \4978 , \4980 );
not \U$21972 ( \22315 , \22314 );
or \U$21973 ( \22316 , \22313 , \22315 );
or \U$21974 ( \22317 , \22314 , RI98729a0_165);
nand \U$21975 ( \22318 , \22316 , \22317 );
nand \U$21976 ( \22319 , \22318 , \7338 );
nand \U$21977 ( \22320 , \22312 , \22319 );
xor \U$21978 ( \22321 , \22305 , \22320 );
not \U$21979 ( \22322 , \8029 );
not \U$21980 ( \22323 , RI9872a18_166);
not \U$21981 ( \22324 , \7007 );
or \U$21982 ( \22325 , \22323 , \22324 );
nand \U$21983 ( \22326 , \4960 , \8031 );
nand \U$21984 ( \22327 , \22325 , \22326 );
not \U$21985 ( \22328 , \22327 );
or \U$21986 ( \22329 , \22322 , \22328 );
and \U$21987 ( \22330 , RI9872a18_166, \4469 );
not \U$21988 ( \22331 , RI9872a18_166);
and \U$21989 ( \22332 , \22331 , \4710 );
or \U$21990 ( \22333 , \22330 , \22332 );
nand \U$21991 ( \22334 , \22333 , \13017 );
nand \U$21992 ( \22335 , \22329 , \22334 );
and \U$21993 ( \22336 , \22321 , \22335 );
and \U$21994 ( \22337 , \22305 , \22320 );
nor \U$21995 ( \22338 , \22336 , \22337 );
not \U$21996 ( \22339 , \22338 );
not \U$21997 ( \22340 , \22339 );
xor \U$21998 ( \22341 , \21843 , \21818 );
not \U$21999 ( \22342 , \4084 );
not \U$22000 ( \22343 , \21522 );
or \U$22001 ( \22344 , \22342 , \22343 );
and \U$22002 ( \22345 , RI98725e0_157, \8873 );
not \U$22003 ( \22346 , RI98725e0_157);
not \U$22004 ( \22347 , \8619 );
and \U$22005 ( \22348 , \22346 , \22347 );
nor \U$22006 ( \22349 , \22345 , \22348 );
nand \U$22007 ( \22350 , \22349 , \4101 );
nand \U$22008 ( \22351 , \22344 , \22350 );
not \U$22009 ( \22352 , \22351 );
not \U$22010 ( \22353 , \3467 );
not \U$22011 ( \22354 , \21570 );
or \U$22012 ( \22355 , \22353 , \22354 );
not \U$22013 ( \22356 , RI98726d0_159);
not \U$22014 ( \22357 , \8667 );
or \U$22015 ( \22358 , \22356 , \22357 );
or \U$22016 ( \22359 , \9880 , RI98726d0_159);
nand \U$22017 ( \22360 , \22358 , \22359 );
nand \U$22018 ( \22361 , \22360 , \3464 );
nand \U$22019 ( \22362 , \22355 , \22361 );
not \U$22020 ( \22363 , \22362 );
not \U$22021 ( \22364 , \22363 );
or \U$22022 ( \22365 , \22352 , \22364 );
not \U$22023 ( \22366 , \22351 );
nand \U$22024 ( \22367 , \22366 , \22362 );
nand \U$22025 ( \22368 , \22365 , \22367 );
not \U$22026 ( \22369 , \3170 );
not \U$22027 ( \22370 , \21612 );
or \U$22028 ( \22371 , \22369 , \22370 );
not \U$22029 ( \22372 , RI9872310_151);
not \U$22030 ( \22373 , \12847 );
or \U$22031 ( \22374 , \22372 , \22373 );
or \U$22032 ( \22375 , \8579 , RI9872310_151);
nand \U$22033 ( \22376 , \22374 , \22375 );
nand \U$22034 ( \22377 , \22376 , \6653 );
nand \U$22035 ( \22378 , \22371 , \22377 );
and \U$22036 ( \22379 , \22368 , \22378 );
not \U$22037 ( \22380 , \22368 );
not \U$22038 ( \22381 , \22378 );
and \U$22039 ( \22382 , \22380 , \22381 );
nor \U$22040 ( \22383 , \22379 , \22382 );
xor \U$22041 ( \22384 , \22341 , \22383 );
not \U$22042 ( \22385 , \22384 );
or \U$22043 ( \22386 , \22340 , \22385 );
nand \U$22044 ( \22387 , \22383 , \22341 );
nand \U$22045 ( \22388 , \22386 , \22387 );
not \U$22046 ( \22389 , \22388 );
not \U$22047 ( \22390 , \1292 );
not \U$22048 ( \22391 , \18350 );
not \U$22049 ( \22392 , \22391 );
and \U$22050 ( \22393 , RI9871b18_134, \22392 );
not \U$22051 ( \22394 , RI9871b18_134);
not \U$22052 ( \22395 , \18350 );
and \U$22053 ( \22396 , \22394 , \22395 );
or \U$22054 ( \22397 , \22393 , \22396 );
not \U$22055 ( \22398 , \22397 );
or \U$22056 ( \22399 , \22390 , \22398 );
nand \U$22057 ( \22400 , \21800 , \1323 );
nand \U$22058 ( \22401 , \22399 , \22400 );
not \U$22059 ( \22402 , \791 );
xor \U$22060 ( \22403 , RI98719b0_131, \18344 );
not \U$22061 ( \22404 , \22403 );
or \U$22062 ( \22405 , \22402 , \22404 );
and \U$22063 ( \22406 , RI98719b0_131, \9849 );
not \U$22064 ( \22407 , RI98719b0_131);
and \U$22065 ( \22408 , \22407 , \8708 );
or \U$22066 ( \22409 , \22406 , \22408 );
nand \U$22067 ( \22410 , \22409 , \796 );
nand \U$22068 ( \22411 , \22405 , \22410 );
xor \U$22069 ( \22412 , \22401 , \22411 );
not \U$22070 ( \22413 , \22412 );
not \U$22071 ( \22414 , \6284 );
not \U$22072 ( \22415 , RI98728b0_163);
not \U$22073 ( \22416 , \7111 );
or \U$22074 ( \22417 , \22415 , \22416 );
or \U$22075 ( \22418 , \9556 , RI98728b0_163);
nand \U$22076 ( \22419 , \22417 , \22418 );
not \U$22077 ( \22420 , \22419 );
or \U$22078 ( \22421 , \22414 , \22420 );
and \U$22079 ( \22422 , RI98728b0_163, \5763 );
not \U$22080 ( \22423 , RI98728b0_163);
and \U$22081 ( \22424 , \22423 , \5766 );
or \U$22082 ( \22425 , \22422 , \22424 );
nand \U$22083 ( \22426 , \22425 , \6610 );
nand \U$22084 ( \22427 , \22421 , \22426 );
not \U$22085 ( \22428 , \22427 );
or \U$22086 ( \22429 , \22413 , \22428 );
nand \U$22087 ( \22430 , \22411 , \22401 );
nand \U$22088 ( \22431 , \22429 , \22430 );
not \U$22089 ( \22432 , \22431 );
not \U$22090 ( \22433 , \4923 );
and \U$22091 ( \22434 , \8334 , RI9872388_152);
not \U$22092 ( \22435 , \8334 );
and \U$22093 ( \22436 , \22435 , \4902 );
or \U$22094 ( \22437 , \22434 , \22436 );
not \U$22095 ( \22438 , \22437 );
or \U$22096 ( \22439 , \22433 , \22438 );
and \U$22097 ( \22440 , RI9872388_152, \10391 );
not \U$22098 ( \22441 , RI9872388_152);
and \U$22099 ( \22442 , \22441 , \21518 );
nor \U$22100 ( \22443 , \22440 , \22442 );
nand \U$22101 ( \22444 , \22443 , \4919 );
nand \U$22102 ( \22445 , \22439 , \22444 );
not \U$22103 ( \22446 , \22445 );
not \U$22104 ( \22447 , \5034 );
not \U$22105 ( \22448 , RI9872478_154);
not \U$22106 ( \22449 , \7465 );
or \U$22107 ( \22450 , \22448 , \22449 );
or \U$22108 ( \22451 , \7465 , RI9872478_154);
nand \U$22109 ( \22452 , \22450 , \22451 );
not \U$22110 ( \22453 , \22452 );
or \U$22111 ( \22454 , \22447 , \22453 );
and \U$22112 ( \22455 , RI9872478_154, \10581 );
not \U$22113 ( \22456 , RI9872478_154);
and \U$22114 ( \22457 , \22456 , \7002 );
nor \U$22115 ( \22458 , \22455 , \22457 );
buf \U$22116 ( \22459 , \5035 );
nand \U$22117 ( \22460 , \22458 , \22459 );
nand \U$22118 ( \22461 , \22454 , \22460 );
not \U$22119 ( \22462 , \832 );
not \U$22120 ( \22463 , \21762 );
or \U$22121 ( \22464 , \22462 , \22463 );
not \U$22122 ( \22465 , RI9871d70_139);
buf \U$22123 ( \22466 , \19542 );
not \U$22124 ( \22467 , \22466 );
or \U$22125 ( \22468 , \22465 , \22467 );
or \U$22126 ( \22469 , \22466 , RI9871d70_139);
nand \U$22127 ( \22470 , \22468 , \22469 );
nand \U$22128 ( \22471 , \22470 , \858 );
nand \U$22129 ( \22472 , \22464 , \22471 );
not \U$22130 ( \22473 , \22472 );
not \U$22131 ( \22474 , \22282 );
not \U$22132 ( \22475 , \22271 );
and \U$22133 ( \22476 , \22474 , \22475 );
and \U$22134 ( \22477 , \22282 , \22271 );
nor \U$22135 ( \22478 , \22476 , \22477 );
not \U$22136 ( \22479 , \22478 );
or \U$22137 ( \22480 , \22473 , \22479 );
or \U$22138 ( \22481 , \22478 , \22472 );
nand \U$22139 ( \22482 , \22480 , \22481 );
not \U$22140 ( \22483 , \22482 );
not \U$22141 ( \22484 , \1517 );
not \U$22142 ( \22485 , \22300 );
or \U$22143 ( \22486 , \22484 , \22485 );
not \U$22144 ( \22487 , RI9871c80_137);
not \U$22145 ( \22488 , \17741 );
or \U$22146 ( \22489 , \22487 , \22488 );
or \U$22147 ( \22490 , \17911 , RI9871c80_137);
nand \U$22148 ( \22491 , \22489 , \22490 );
nand \U$22149 ( \22492 , \22491 , \1500 );
nand \U$22150 ( \22493 , \22486 , \22492 );
not \U$22151 ( \22494 , \22493 );
or \U$22152 ( \22495 , \22483 , \22494 );
not \U$22153 ( \22496 , \22478 );
nand \U$22154 ( \22497 , \22496 , \22472 );
nand \U$22155 ( \22498 , \22495 , \22497 );
xor \U$22156 ( \22499 , \22461 , \22498 );
not \U$22157 ( \22500 , \22499 );
or \U$22158 ( \22501 , \22446 , \22500 );
nand \U$22159 ( \22502 , \22461 , \22498 );
nand \U$22160 ( \22503 , \22501 , \22502 );
not \U$22161 ( \22504 , \22503 );
nand \U$22162 ( \22505 , \22432 , \22504 );
not \U$22163 ( \22506 , \22505 );
not \U$22164 ( \22507 , \5642 );
not \U$22165 ( \22508 , \5644 );
not \U$22166 ( \22509 , \18793 );
or \U$22167 ( \22510 , \22508 , \22509 );
or \U$22168 ( \22511 , \6528 , \5644 );
nand \U$22169 ( \22512 , \22510 , \22511 );
not \U$22170 ( \22513 , \22512 );
or \U$22171 ( \22514 , \22507 , \22513 );
not \U$22172 ( \22515 , \5648 );
buf \U$22173 ( \22516 , \6296 );
not \U$22174 ( \22517 , \22516 );
or \U$22175 ( \22518 , \22515 , \22517 );
nand \U$22176 ( \22519 , \8053 , RI9872568_156);
nand \U$22177 ( \22520 , \22518 , \22519 );
nand \U$22178 ( \22521 , \22520 , \5653 );
nand \U$22179 ( \22522 , \22514 , \22521 );
not \U$22180 ( \22523 , \8790 );
not \U$22181 ( \22524 , \8606 );
and \U$22182 ( \22525 , RI98725e0_157, \22524 );
not \U$22183 ( \22526 , RI98725e0_157);
and \U$22184 ( \22527 , \22526 , \8597 );
or \U$22185 ( \22528 , \22525 , \22527 );
not \U$22186 ( \22529 , \22528 );
or \U$22187 ( \22530 , \22523 , \22529 );
nand \U$22188 ( \22531 , \22349 , \5847 );
nand \U$22189 ( \22532 , \22530 , \22531 );
xor \U$22190 ( \22533 , \22522 , \22532 );
not \U$22191 ( \22534 , \3163 );
not \U$22192 ( \22535 , RI9872310_151);
not \U$22193 ( \22536 , \8554 );
or \U$22194 ( \22537 , \22535 , \22536 );
or \U$22195 ( \22538 , \8554 , RI9872310_151);
nand \U$22196 ( \22539 , \22537 , \22538 );
not \U$22197 ( \22540 , \22539 );
or \U$22198 ( \22541 , \22534 , \22540 );
nand \U$22199 ( \22542 , \22376 , \3170 );
nand \U$22200 ( \22543 , \22541 , \22542 );
not \U$22201 ( \22544 , \22543 );
not \U$22202 ( \22545 , \22544 );
and \U$22203 ( \22546 , \22533 , \22545 );
and \U$22204 ( \22547 , \22522 , \22532 );
or \U$22205 ( \22548 , \22546 , \22547 );
not \U$22206 ( \22549 , \22548 );
or \U$22207 ( \22550 , \22506 , \22549 );
nand \U$22208 ( \22551 , \22431 , \22503 );
nand \U$22209 ( \22552 , \22550 , \22551 );
not \U$22210 ( \22553 , \22552 );
xor \U$22211 ( \22554 , \21807 , \21849 );
not \U$22212 ( \22555 , \21847 );
xnor \U$22213 ( \22556 , \22554 , \22555 );
and \U$22214 ( \22557 , \22553 , \22556 );
not \U$22215 ( \22558 , \22553 );
not \U$22216 ( \22559 , \22556 );
and \U$22217 ( \22560 , \22558 , \22559 );
nor \U$22218 ( \22561 , \22557 , \22560 );
not \U$22219 ( \22562 , \22561 );
or \U$22220 ( \22563 , \22389 , \22562 );
not \U$22221 ( \22564 , \22553 );
nand \U$22222 ( \22565 , \22564 , \22559 );
nand \U$22223 ( \22566 , \22563 , \22565 );
not \U$22224 ( \22567 , \22566 );
not \U$22225 ( \22568 , \21923 );
not \U$22226 ( \22569 , \21926 );
or \U$22227 ( \22570 , \22568 , \22569 );
or \U$22228 ( \22571 , \21926 , \21923 );
nand \U$22229 ( \22572 , \22570 , \22571 );
not \U$22230 ( \22573 , \21929 );
and \U$22231 ( \22574 , \22572 , \22573 );
not \U$22232 ( \22575 , \22572 );
and \U$22233 ( \22576 , \22575 , \21929 );
nor \U$22234 ( \22577 , \22574 , \22576 );
not \U$22235 ( \22578 , \22577 );
and \U$22236 ( \22579 , \22567 , \22578 );
and \U$22237 ( \22580 , \22566 , \22577 );
nor \U$22238 ( \22581 , \22579 , \22580 );
not \U$22239 ( \22582 , \22581 );
not \U$22240 ( \22583 , \22582 );
not \U$22241 ( \22584 , \9214 );
not \U$22242 ( \22585 , RI9872b80_169);
not \U$22243 ( \22586 , \12616 );
or \U$22244 ( \22587 , \22585 , \22586 );
or \U$22245 ( \22588 , \18647 , RI9872b80_169);
nand \U$22246 ( \22589 , \22587 , \22588 );
not \U$22247 ( \22590 , \22589 );
or \U$22248 ( \22591 , \22584 , \22590 );
and \U$22249 ( \22592 , RI9872b80_169, \4408 );
not \U$22250 ( \22593 , RI9872b80_169);
and \U$22251 ( \22594 , \22593 , \22043 );
or \U$22252 ( \22595 , \22592 , \22594 );
nand \U$22253 ( \22596 , \22595 , \10679 );
nand \U$22254 ( \22597 , \22591 , \22596 );
not \U$22255 ( \22598 , \22597 );
not \U$22256 ( \22599 , \18239 );
not \U$22257 ( \22600 , \6164 );
or \U$22258 ( \22601 , \22599 , \22600 );
not \U$22259 ( \22602 , \18239 );
nand \U$22260 ( \22603 , \22602 , \1446 );
nand \U$22261 ( \22604 , \22601 , \22603 );
nand \U$22262 ( \22605 , \22604 , \20626 );
xor \U$22263 ( \22606 , RI9873558_190, \1415 );
nand \U$22264 ( \22607 , \22606 , RI9873648_192);
nand \U$22265 ( \22608 , \22605 , \22607 );
not \U$22266 ( \22609 , \13020 );
xor \U$22267 ( \22610 , RI98730a8_180, \1365 );
not \U$22268 ( \22611 , \22610 );
or \U$22269 ( \22612 , \22609 , \22611 );
and \U$22270 ( \22613 , RI98730a8_180, \1339 );
not \U$22271 ( \22614 , RI98730a8_180);
not \U$22272 ( \22615 , \20612 );
and \U$22273 ( \22616 , \22614 , \22615 );
or \U$22274 ( \22617 , \22613 , \22616 );
buf \U$22275 ( \22618 , \11342 );
nand \U$22276 ( \22619 , \22617 , \22618 );
nand \U$22277 ( \22620 , \22612 , \22619 );
not \U$22278 ( \22621 , \22620 );
and \U$22279 ( \22622 , \22608 , \22621 );
not \U$22280 ( \22623 , \22608 );
and \U$22281 ( \22624 , \22623 , \22620 );
or \U$22282 ( \22625 , \22622 , \22624 );
not \U$22283 ( \22626 , \22625 );
or \U$22284 ( \22627 , \22598 , \22626 );
not \U$22285 ( \22628 , \22607 );
not \U$22286 ( \22629 , \22605 );
or \U$22287 ( \22630 , \22628 , \22629 );
nand \U$22288 ( \22631 , \22630 , \22620 );
nand \U$22289 ( \22632 , \22627 , \22631 );
not \U$22290 ( \22633 , \22632 );
not \U$22291 ( \22634 , \22633 );
not \U$22292 ( \22635 , \22634 );
not \U$22293 ( \22636 , \9670 );
not \U$22294 ( \22637 , \3568 );
not \U$22295 ( \22638 , RI9872bf8_170);
or \U$22296 ( \22639 , \22637 , \22638 );
or \U$22297 ( \22640 , \14930 , RI9872bf8_170);
nand \U$22298 ( \22641 , \22639 , \22640 );
not \U$22299 ( \22642 , \22641 );
or \U$22300 ( \22643 , \22636 , \22642 );
not \U$22301 ( \22644 , \9244 );
not \U$22302 ( \22645 , \3537 );
or \U$22303 ( \22646 , \22644 , \22645 );
or \U$22304 ( \22647 , \6718 , \9244 );
nand \U$22305 ( \22648 , \22646 , \22647 );
nand \U$22306 ( \22649 , \22648 , \9668 );
nand \U$22307 ( \22650 , \22643 , \22649 );
not \U$22308 ( \22651 , \22650 );
not \U$22309 ( \22652 , \22651 );
not \U$22310 ( \22653 , \8802 );
and \U$22311 ( \22654 , RI9872d60_173, \2947 );
not \U$22312 ( \22655 , RI9872d60_173);
and \U$22313 ( \22656 , \22655 , \5884 );
or \U$22314 ( \22657 , \22654 , \22656 );
not \U$22315 ( \22658 , \22657 );
or \U$22316 ( \22659 , \22653 , \22658 );
and \U$22317 ( \22660 , \3859 , \8807 );
not \U$22318 ( \22661 , \3859 );
and \U$22319 ( \22662 , \22661 , RI9872d60_173);
nor \U$22320 ( \22663 , \22660 , \22662 );
buf \U$22321 ( \22664 , \8817 );
nand \U$22322 ( \22665 , \22663 , \22664 );
nand \U$22323 ( \22666 , \22659 , \22665 );
not \U$22324 ( \22667 , \22666 );
not \U$22325 ( \22668 , \22667 );
or \U$22326 ( \22669 , \22652 , \22668 );
buf \U$22327 ( \22670 , \13483 );
not \U$22328 ( \22671 , \22670 );
not \U$22329 ( \22672 , \18012 );
not \U$22330 ( \22673 , \943 );
or \U$22331 ( \22674 , \22672 , \22673 );
not \U$22332 ( \22675 , RI9873210_183);
or \U$22333 ( \22676 , \6651 , \22675 );
nand \U$22334 ( \22677 , \22674 , \22676 );
not \U$22335 ( \22678 , \22677 );
or \U$22336 ( \22679 , \22671 , \22678 );
and \U$22337 ( \22680 , RI9873210_183, \5719 );
not \U$22338 ( \22681 , RI9873210_183);
and \U$22339 ( \22682 , \22681 , \7019 );
nor \U$22340 ( \22683 , \22680 , \22682 );
nand \U$22341 ( \22684 , \22683 , \13476 );
nand \U$22342 ( \22685 , \22679 , \22684 );
nand \U$22343 ( \22686 , \22669 , \22685 );
nand \U$22344 ( \22687 , \22666 , \22650 );
and \U$22345 ( \22688 , \22686 , \22687 );
not \U$22346 ( \22689 , \22688 );
not \U$22347 ( \22690 , \18563 );
xnor \U$22348 ( \22691 , \6378 , RI9872e50_175);
not \U$22349 ( \22692 , \22691 );
or \U$22350 ( \22693 , \22690 , \22692 );
not \U$22351 ( \22694 , RI9872e50_175);
not \U$22352 ( \22695 , \1485 );
or \U$22353 ( \22696 , \22694 , \22695 );
nand \U$22354 ( \22697 , \1486 , \9694 );
nand \U$22355 ( \22698 , \22696 , \22697 );
nand \U$22356 ( \22699 , \22698 , \10333 );
nand \U$22357 ( \22700 , \22693 , \22699 );
not \U$22358 ( \22701 , \22700 );
not \U$22359 ( \22702 , \19046 );
xor \U$22360 ( \22703 , RI98734e0_189, \1306 );
not \U$22361 ( \22704 , \22703 );
or \U$22362 ( \22705 , \22702 , \22704 );
not \U$22363 ( \22706 , \16999 );
not \U$22364 ( \22707 , \1273 );
or \U$22365 ( \22708 , \22706 , \22707 );
not \U$22366 ( \22709 , RI98734e0_189);
or \U$22367 ( \22710 , \22709 , \1273 );
nand \U$22368 ( \22711 , \22708 , \22710 );
nand \U$22369 ( \22712 , \22711 , \19036 );
nand \U$22370 ( \22713 , \22705 , \22712 );
not \U$22371 ( \22714 , \18522 );
not \U$22372 ( \22715 , RI9873288_184);
not \U$22373 ( \22716 , \22715 );
not \U$22374 ( \22717 , \8004 );
or \U$22375 ( \22718 , \22716 , \22717 );
not \U$22376 ( \22719 , RI9873288_184);
or \U$22377 ( \22720 , \8004 , \22719 );
nand \U$22378 ( \22721 , \22718 , \22720 );
not \U$22379 ( \22722 , \22721 );
or \U$22380 ( \22723 , \22714 , \22722 );
not \U$22381 ( \22724 , RI9873288_184);
not \U$22382 ( \22725 , \16923 );
or \U$22383 ( \22726 , \22724 , \22725 );
not \U$22384 ( \22727 , RI9873288_184);
nand \U$22385 ( \22728 , \22727 , \845 );
nand \U$22386 ( \22729 , \22726 , \22728 );
nand \U$22387 ( \22730 , \22729 , \17545 );
nand \U$22388 ( \22731 , \22723 , \22730 );
xor \U$22389 ( \22732 , \22713 , \22731 );
not \U$22390 ( \22733 , \22732 );
or \U$22391 ( \22734 , \22701 , \22733 );
not \U$22392 ( \22735 , \22713 );
not \U$22393 ( \22736 , \22735 );
nand \U$22394 ( \22737 , \22736 , \22731 );
nand \U$22395 ( \22738 , \22734 , \22737 );
not \U$22396 ( \22739 , \22738 );
or \U$22397 ( \22740 , \22689 , \22739 );
or \U$22398 ( \22741 , \22738 , \22688 );
nand \U$22399 ( \22742 , \22740 , \22741 );
not \U$22400 ( \22743 , \22742 );
or \U$22401 ( \22744 , \22635 , \22743 );
not \U$22402 ( \22745 , \22688 );
nand \U$22403 ( \22746 , \22745 , \22738 );
nand \U$22404 ( \22747 , \22744 , \22746 );
not \U$22405 ( \22748 , \22747 );
not \U$22406 ( \22749 , \2087 );
not \U$22407 ( \22750 , \21589 );
or \U$22408 ( \22751 , \22749 , \22750 );
not \U$22409 ( \22752 , \8722 );
and \U$22410 ( \22753 , RI9871aa0_133, \22752 );
not \U$22411 ( \22754 , RI9871aa0_133);
and \U$22412 ( \22755 , \22754 , \12470 );
or \U$22413 ( \22756 , \22753 , \22755 );
nand \U$22414 ( \22757 , \22756 , \2071 );
nand \U$22415 ( \22758 , \22751 , \22757 );
not \U$22416 ( \22759 , \22758 );
and \U$22417 ( \22760 , \21602 , \796 );
and \U$22418 ( \22761 , \22409 , \11432 );
nor \U$22419 ( \22762 , \22760 , \22761 );
nand \U$22420 ( \22763 , \22759 , \22762 );
not \U$22421 ( \22764 , \22763 );
not \U$22422 ( \22765 , \5653 );
not \U$22423 ( \22766 , \21958 );
or \U$22424 ( \22767 , \22765 , \22766 );
nand \U$22425 ( \22768 , \22520 , \5642 );
nand \U$22426 ( \22769 , \22767 , \22768 );
not \U$22427 ( \22770 , \22769 );
or \U$22428 ( \22771 , \22764 , \22770 );
not \U$22429 ( \22772 , \22762 );
nand \U$22430 ( \22773 , \22772 , \22758 );
nand \U$22431 ( \22774 , \22771 , \22773 );
not \U$22432 ( \22775 , \22774 );
not \U$22433 ( \22776 , \22378 );
not \U$22434 ( \22777 , \22368 );
or \U$22435 ( \22778 , \22776 , \22777 );
nand \U$22436 ( \22779 , \22362 , \22351 );
nand \U$22437 ( \22780 , \22778 , \22779 );
xor \U$22438 ( \22781 , \22775 , \22780 );
not \U$22439 ( \22782 , \4923 );
not \U$22440 ( \22783 , \21644 );
or \U$22441 ( \22784 , \22782 , \22783 );
nand \U$22442 ( \22785 , \22437 , \4918 );
nand \U$22443 ( \22786 , \22784 , \22785 );
not \U$22444 ( \22787 , \22786 );
not \U$22445 ( \22788 , \22283 );
nand \U$22446 ( \22789 , \22788 , \22293 );
not \U$22447 ( \22790 , \22789 );
not \U$22448 ( \22791 , \22304 );
not \U$22449 ( \22792 , \22791 );
or \U$22450 ( \22793 , \22790 , \22792 );
not \U$22451 ( \22794 , \22293 );
nand \U$22452 ( \22795 , \22794 , \22283 );
nand \U$22453 ( \22796 , \22793 , \22795 );
not \U$22454 ( \22797 , \5035 );
not \U$22455 ( \22798 , \21657 );
or \U$22456 ( \22799 , \22797 , \22798 );
nand \U$22457 ( \22800 , \22458 , \5034 );
nand \U$22458 ( \22801 , \22799 , \22800 );
not \U$22459 ( \22802 , \22801 );
xor \U$22460 ( \22803 , \22796 , \22802 );
nand \U$22461 ( \22804 , \22787 , \22803 );
buf \U$22462 ( \22805 , \22801 );
not \U$22463 ( \22806 , \22805 );
nand \U$22464 ( \22807 , \22806 , \22796 );
nand \U$22465 ( \22808 , \22804 , \22807 );
xnor \U$22466 ( \22809 , \22781 , \22808 );
not \U$22467 ( \22810 , \22809 );
xor \U$22468 ( \22811 , \22762 , \22758 );
not \U$22469 ( \22812 , \22769 );
xor \U$22470 ( \22813 , \22811 , \22812 );
xor \U$22471 ( \22814 , \22796 , \22786 );
xnor \U$22472 ( \22815 , \22814 , \22805 );
xor \U$22473 ( \22816 , \22813 , \22815 );
not \U$22474 ( \22817 , \3465 );
not \U$22475 ( \22818 , RI98726d0_159);
not \U$22476 ( \22819 , \8650 );
or \U$22477 ( \22820 , \22818 , \22819 );
or \U$22478 ( \22821 , \8650 , RI98726d0_159);
nand \U$22479 ( \22822 , \22820 , \22821 );
not \U$22480 ( \22823 , \22822 );
or \U$22481 ( \22824 , \22817 , \22823 );
nand \U$22482 ( \22825 , \22360 , \3467 );
nand \U$22483 ( \22826 , \22824 , \22825 );
not \U$22484 ( \22827 , \2072 );
and \U$22485 ( \22828 , \8695 , RI9871aa0_133);
not \U$22486 ( \22829 , \8695 );
and \U$22487 ( \22830 , \22829 , \2076 );
nor \U$22488 ( \22831 , \22828 , \22830 );
not \U$22489 ( \22832 , \22831 );
or \U$22490 ( \22833 , \22827 , \22832 );
nand \U$22491 ( \22834 , \22756 , \2087 );
nand \U$22492 ( \22835 , \22833 , \22834 );
or \U$22493 ( \22836 , \22826 , \22835 );
not \U$22494 ( \22837 , \22836 );
not \U$22495 ( \22838 , \8732 );
not \U$22496 ( \22839 , \11755 );
or \U$22497 ( \22840 , \22838 , \22839 );
nand \U$22498 ( \22841 , \5946 , RI9872f40_177);
nand \U$22499 ( \22842 , \22840 , \22841 );
not \U$22500 ( \22843 , \22842 );
not \U$22501 ( \22844 , \9527 );
or \U$22502 ( \22845 , \22843 , \22844 );
not \U$22503 ( \22846 , RI9872f40_177);
not \U$22504 ( \22847 , \3127 );
or \U$22505 ( \22848 , \22846 , \22847 );
or \U$22506 ( \22849 , \6021 , RI9872f40_177);
nand \U$22507 ( \22850 , \22848 , \22849 );
nand \U$22508 ( \22851 , \22850 , \8752 );
nand \U$22509 ( \22852 , \22845 , \22851 );
not \U$22510 ( \22853 , \22852 );
or \U$22511 ( \22854 , \22837 , \22853 );
nand \U$22512 ( \22855 , \22826 , \22835 );
nand \U$22513 ( \22856 , \22854 , \22855 );
and \U$22514 ( \22857 , \22816 , \22856 );
and \U$22515 ( \22858 , \22813 , \22815 );
or \U$22516 ( \22859 , \22857 , \22858 );
not \U$22517 ( \22860 , \22859 );
or \U$22518 ( \22861 , \22810 , \22860 );
or \U$22519 ( \22862 , \22859 , \22809 );
nand \U$22520 ( \22863 , \22861 , \22862 );
not \U$22521 ( \22864 , \22863 );
or \U$22522 ( \22865 , \22748 , \22864 );
not \U$22523 ( \22866 , \22809 );
nand \U$22524 ( \22867 , \22866 , \22859 );
nand \U$22525 ( \22868 , \22865 , \22867 );
not \U$22526 ( \22869 , \22868 );
or \U$22527 ( \22870 , \22583 , \22869 );
not \U$22528 ( \22871 , \22577 );
nand \U$22529 ( \22872 , \22871 , \22566 );
nand \U$22530 ( \22873 , \22870 , \22872 );
not \U$22531 ( \22874 , \22873 );
or \U$22532 ( \22875 , \22269 , \22874 );
not \U$22533 ( \22876 , \22267 );
nand \U$22534 ( \22877 , \22876 , \22264 );
nand \U$22535 ( \22878 , \22875 , \22877 );
xor \U$22536 ( \22879 , \21913 , \21991 );
xor \U$22537 ( \22880 , \22879 , \21994 );
or \U$22538 ( \22881 , \22878 , \22880 );
not \U$22539 ( \22882 , \22881 );
or \U$22540 ( \22883 , \22258 , \22882 );
nand \U$22541 ( \22884 , \22878 , \22880 );
nand \U$22542 ( \22885 , \22883 , \22884 );
not \U$22543 ( \22886 , \22885 );
not \U$22544 ( \22887 , \22216 );
not \U$22545 ( \22888 , \22012 );
or \U$22546 ( \22889 , \22887 , \22888 );
or \U$22547 ( \22890 , \22216 , \22012 );
nand \U$22548 ( \22891 , \22889 , \22890 );
and \U$22549 ( \22892 , \22891 , \22220 );
not \U$22550 ( \22893 , \22891 );
and \U$22551 ( \22894 , \22893 , \22018 );
nor \U$22552 ( \22895 , \22892 , \22894 );
xor \U$22553 ( \22896 , \22205 , \22025 );
xor \U$22554 ( \22897 , \22896 , \22208 );
not \U$22555 ( \22898 , \22897 );
not \U$22556 ( \22899 , \22898 );
xor \U$22557 ( \22900 , \21583 , \21624 );
not \U$22558 ( \22901 , \21664 );
xor \U$22559 ( \22902 , \22900 , \22901 );
not \U$22560 ( \22903 , \22902 );
xor \U$22561 ( \22904 , \21635 , \21649 );
xnor \U$22562 ( \22905 , \22904 , \21661 );
not \U$22563 ( \22906 , \21524 );
and \U$22564 ( \22907 , \21578 , \22906 );
not \U$22565 ( \22908 , \21578 );
and \U$22566 ( \22909 , \22908 , \21524 );
nor \U$22567 ( \22910 , \22907 , \22909 );
nand \U$22568 ( \22911 , \22905 , \22910 );
not \U$22569 ( \22912 , \22911 );
not \U$22570 ( \22913 , \13020 );
not \U$22571 ( \22914 , \22617 );
or \U$22572 ( \22915 , \22913 , \22914 );
nand \U$22573 ( \22916 , \22052 , \22618 );
nand \U$22574 ( \22917 , \22915 , \22916 );
not \U$22575 ( \22918 , \9196 );
not \U$22576 ( \22919 , \22589 );
or \U$22577 ( \22920 , \22918 , \22919 );
nand \U$22578 ( \22921 , \22152 , \9214 );
nand \U$22579 ( \22922 , \22920 , \22921 );
xor \U$22580 ( \22923 , \22917 , \22922 );
not \U$22581 ( \22924 , \17263 );
not \U$22582 ( \22925 , \22178 );
or \U$22583 ( \22926 , \22924 , \22925 );
not \U$22584 ( \22927 , RI98733f0_187);
not \U$22585 ( \22928 , \6585 );
or \U$22586 ( \22929 , \22927 , \22928 );
or \U$22587 ( \22930 , \915 , RI98733f0_187);
nand \U$22588 ( \22931 , \22929 , \22930 );
nand \U$22589 ( \22932 , \22931 , \17252 );
nand \U$22590 ( \22933 , \22926 , \22932 );
and \U$22591 ( \22934 , \22923 , \22933 );
and \U$22592 ( \22935 , \22917 , \22922 );
or \U$22593 ( \22936 , \22934 , \22935 );
not \U$22594 ( \22937 , \22936 );
or \U$22595 ( \22938 , \22912 , \22937 );
not \U$22596 ( \22939 , \22905 );
not \U$22597 ( \22940 , \22910 );
nand \U$22598 ( \22941 , \22939 , \22940 );
nand \U$22599 ( \22942 , \22938 , \22941 );
not \U$22600 ( \22943 , \22942 );
or \U$22601 ( \22944 , \22903 , \22943 );
or \U$22602 ( \22945 , \22942 , \22902 );
nand \U$22603 ( \22946 , \22944 , \22945 );
not \U$22604 ( \22947 , \22946 );
not \U$22605 ( \22948 , \9668 );
not \U$22606 ( \22949 , \22164 );
or \U$22607 ( \22950 , \22948 , \22949 );
nand \U$22608 ( \22951 , \22648 , \9249 );
nand \U$22609 ( \22952 , \22950 , \22951 );
not \U$22610 ( \22953 , \10251 );
not \U$22611 ( \22954 , \22657 );
or \U$22612 ( \22955 , \22953 , \22954 );
nand \U$22613 ( \22956 , \22063 , \8801 );
nand \U$22614 ( \22957 , \22955 , \22956 );
xor \U$22615 ( \22958 , \22952 , \22957 );
not \U$22616 ( \22959 , \13484 );
not \U$22617 ( \22960 , \22081 );
or \U$22618 ( \22961 , \22959 , \22960 );
nand \U$22619 ( \22962 , \22677 , \13477 );
nand \U$22620 ( \22963 , \22961 , \22962 );
and \U$22621 ( \22964 , \22958 , \22963 );
and \U$22622 ( \22965 , \22952 , \22957 );
or \U$22623 ( \22966 , \22964 , \22965 );
not \U$22624 ( \22967 , \22966 );
not \U$22625 ( \22968 , \8752 );
not \U$22626 ( \22969 , \21945 );
or \U$22627 ( \22970 , \22968 , \22969 );
nand \U$22628 ( \22971 , \22850 , \8743 );
nand \U$22629 ( \22972 , \22970 , \22971 );
not \U$22630 ( \22973 , \22972 );
xor \U$22631 ( \22974 , \21558 , \21535 );
not \U$22632 ( \22975 , \22974 );
not \U$22633 ( \22976 , \19243 );
not \U$22634 ( \22977 , \22703 );
or \U$22635 ( \22978 , \22976 , \22977 );
nand \U$22636 ( \22979 , \22093 , \19046 );
nand \U$22637 ( \22980 , \22978 , \22979 );
not \U$22638 ( \22981 , \22980 );
not \U$22639 ( \22982 , \22981 );
or \U$22640 ( \22983 , \22975 , \22982 );
or \U$22641 ( \22984 , \22981 , \22974 );
nand \U$22642 ( \22985 , \22983 , \22984 );
not \U$22643 ( \22986 , \22985 );
or \U$22644 ( \22987 , \22973 , \22986 );
nand \U$22645 ( \22988 , \22980 , \22974 );
nand \U$22646 ( \22989 , \22987 , \22988 );
not \U$22647 ( \22990 , \9273 );
not \U$22648 ( \22991 , \22100 );
or \U$22649 ( \22992 , \22990 , \22991 );
nand \U$22650 ( \22993 , \22698 , \18563 );
nand \U$22651 ( \22994 , \22992 , \22993 );
not \U$22652 ( \22995 , \22994 );
not \U$22653 ( \22996 , \17528 );
not \U$22654 ( \22997 , \22112 );
or \U$22655 ( \22998 , \22996 , \22997 );
nand \U$22656 ( \22999 , \22721 , \18508 );
nand \U$22657 ( \23000 , \22998 , \22999 );
not \U$22658 ( \23001 , RI9873648_192);
not \U$22659 ( \23002 , \22071 );
or \U$22660 ( \23003 , \23001 , \23002 );
nand \U$22661 ( \23004 , \22606 , \18545 );
nand \U$22662 ( \23005 , \23003 , \23004 );
xor \U$22663 ( \23006 , \23000 , \23005 );
not \U$22664 ( \23007 , \23006 );
or \U$22665 ( \23008 , \22995 , \23007 );
nand \U$22666 ( \23009 , \23000 , \23005 );
nand \U$22667 ( \23010 , \23008 , \23009 );
xor \U$22668 ( \23011 , \22989 , \23010 );
not \U$22669 ( \23012 , \23011 );
or \U$22670 ( \23013 , \22967 , \23012 );
nand \U$22671 ( \23014 , \23010 , \22989 );
nand \U$22672 ( \23015 , \23013 , \23014 );
not \U$22673 ( \23016 , \23015 );
or \U$22674 ( \23017 , \22947 , \23016 );
not \U$22675 ( \23018 , \22902 );
nand \U$22676 ( \23019 , \23018 , \22942 );
nand \U$22677 ( \23020 , \23017 , \23019 );
buf \U$22678 ( \23021 , \21968 );
not \U$22679 ( \23022 , \21949 );
and \U$22680 ( \23023 , \23021 , \23022 );
not \U$22681 ( \23024 , \23021 );
and \U$22682 ( \23025 , \23024 , \21949 );
nor \U$22683 ( \23026 , \23023 , \23025 );
not \U$22684 ( \23027 , \23026 );
not \U$22685 ( \23028 , \23027 );
xor \U$22686 ( \23029 , \21604 , \21593 );
xnor \U$22687 ( \23030 , \23029 , \21616 );
not \U$22688 ( \23031 , \23030 );
not \U$22689 ( \23032 , \23031 );
not \U$22690 ( \23033 , \7338 );
not \U$22691 ( \23034 , \22125 );
or \U$22692 ( \23035 , \23033 , \23034 );
nand \U$22693 ( \23036 , \22318 , \7325 );
nand \U$22694 ( \23037 , \23035 , \23036 );
not \U$22695 ( \23038 , \9937 );
not \U$22696 ( \23039 , \22132 );
or \U$22697 ( \23040 , \23038 , \23039 );
and \U$22698 ( \23041 , RI9873030_179, \1061 );
not \U$22699 ( \23042 , RI9873030_179);
not \U$22700 ( \23043 , \1061 );
and \U$22701 ( \23044 , \23042 , \23043 );
nor \U$22702 ( \23045 , \23041 , \23044 );
nand \U$22703 ( \23046 , \23045 , \9952 );
nand \U$22704 ( \23047 , \23040 , \23046 );
xor \U$22705 ( \23048 , \23037 , \23047 );
not \U$22706 ( \23049 , \13017 );
not \U$22707 ( \23050 , \22045 );
or \U$22708 ( \23051 , \23049 , \23050 );
nand \U$22709 ( \23052 , \22333 , \8027 );
nand \U$22710 ( \23053 , \23051 , \23052 );
nand \U$22711 ( \23054 , \23048 , \23053 );
not \U$22712 ( \23055 , \23054 );
and \U$22713 ( \23056 , \23037 , \23047 );
nor \U$22714 ( \23057 , \23055 , \23056 );
not \U$22715 ( \23058 , \23057 );
or \U$22716 ( \23059 , \23032 , \23058 );
not \U$22717 ( \23060 , \23056 );
not \U$22718 ( \23061 , \23060 );
not \U$22719 ( \23062 , \23054 );
or \U$22720 ( \23063 , \23061 , \23062 );
nand \U$22721 ( \23064 , \23063 , \23030 );
nand \U$22722 ( \23065 , \23059 , \23064 );
not \U$22723 ( \23066 , \23065 );
or \U$22724 ( \23067 , \23028 , \23066 );
not \U$22725 ( \23068 , \23060 );
not \U$22726 ( \23069 , \23054 );
or \U$22727 ( \23070 , \23068 , \23069 );
nand \U$22728 ( \23071 , \23070 , \23031 );
nand \U$22729 ( \23072 , \23067 , \23071 );
not \U$22730 ( \23073 , \23072 );
not \U$22731 ( \23074 , \22808 );
not \U$22732 ( \23075 , \23074 );
not \U$22733 ( \23076 , \22774 );
or \U$22734 ( \23077 , \23075 , \23076 );
not \U$22735 ( \23078 , \22775 );
not \U$22736 ( \23079 , \22808 );
or \U$22737 ( \23080 , \23078 , \23079 );
nand \U$22738 ( \23081 , \23080 , \22780 );
nand \U$22739 ( \23082 , \23077 , \23081 );
xor \U$22740 ( \23083 , \21939 , \21972 );
and \U$22741 ( \23084 , \23082 , \23083 );
not \U$22742 ( \23085 , \23082 );
not \U$22743 ( \23086 , \23083 );
and \U$22744 ( \23087 , \23085 , \23086 );
nor \U$22745 ( \23088 , \23084 , \23087 );
not \U$22746 ( \23089 , \23088 );
or \U$22747 ( \23090 , \23073 , \23089 );
nand \U$22748 ( \23091 , \23083 , \23082 );
nand \U$22749 ( \23092 , \23090 , \23091 );
not \U$22750 ( \23093 , \23092 );
and \U$22751 ( \23094 , \21512 , \21673 );
not \U$22752 ( \23095 , \21512 );
and \U$22753 ( \23096 , \23095 , \21672 );
nor \U$22754 ( \23097 , \23094 , \23096 );
xnor \U$22755 ( \23098 , \23097 , \21668 );
nand \U$22756 ( \23099 , \23093 , \23098 );
nand \U$22757 ( \23100 , \23020 , \23099 );
not \U$22758 ( \23101 , \23098 );
nand \U$22759 ( \23102 , \23101 , \23092 );
nand \U$22760 ( \23103 , \23100 , \23102 );
not \U$22761 ( \23104 , \22121 );
not \U$22762 ( \23105 , \22200 );
not \U$22763 ( \23106 , \23105 );
or \U$22764 ( \23107 , \23104 , \23106 );
not \U$22765 ( \23108 , \22121 );
nand \U$22766 ( \23109 , \23108 , \22200 );
nand \U$22767 ( \23110 , \23107 , \23109 );
not \U$22768 ( \23111 , \23110 );
not \U$22769 ( \23112 , \23111 );
not \U$22770 ( \23113 , \23112 );
xor \U$22771 ( \23114 , \22057 , \22118 );
xnor \U$22772 ( \23115 , \23114 , \22086 );
xor \U$22773 ( \23116 , \21903 , \21901 );
xnor \U$22774 ( \23117 , \23116 , \21908 );
nand \U$22775 ( \23118 , \23115 , \23117 );
xor \U$22776 ( \23119 , \22036 , \22047 );
xor \U$22777 ( \23120 , \23119 , \22054 );
not \U$22778 ( \23121 , \23120 );
not \U$22779 ( \23122 , \21791 );
not \U$22780 ( \23123 , \21802 );
not \U$22781 ( \23124 , \23123 );
or \U$22782 ( \23125 , \23122 , \23124 );
or \U$22783 ( \23126 , \23123 , \21791 );
nand \U$22784 ( \23127 , \23125 , \23126 );
not \U$22785 ( \23128 , \1083 );
and \U$22786 ( \23129 , \13391 , \1111 );
not \U$22787 ( \23130 , \13391 );
and \U$22788 ( \23131 , \23130 , RI98718c0_129);
nor \U$22789 ( \23132 , \23129 , \23131 );
not \U$22790 ( \23133 , \23132 );
or \U$22791 ( \23134 , \23128 , \23133 );
nand \U$22792 ( \23135 , \21816 , \1135 );
nand \U$22793 ( \23136 , \23134 , \23135 );
not \U$22794 ( \23137 , \23136 );
not \U$22795 ( \23138 , RI9871c08_136);
not \U$22796 ( \23139 , \12772 );
or \U$22797 ( \23140 , \23138 , \23139 );
nand \U$22798 ( \23141 , \17081 , \1850 );
nand \U$22799 ( \23142 , \23140 , \23141 );
nand \U$22800 ( \23143 , \23142 , \1455 );
nand \U$22801 ( \23144 , \21832 , \1428 );
nand \U$22802 ( \23145 , \23143 , \23144 );
xor \U$22803 ( \23146 , \21764 , \21785 );
xor \U$22804 ( \23147 , \23145 , \23146 );
not \U$22805 ( \23148 , \23147 );
or \U$22806 ( \23149 , \23137 , \23148 );
not \U$22807 ( \23150 , \23144 );
not \U$22808 ( \23151 , \23143 );
or \U$22809 ( \23152 , \23150 , \23151 );
nand \U$22810 ( \23153 , \23152 , \23146 );
nand \U$22811 ( \23154 , \23149 , \23153 );
xor \U$22812 ( \23155 , \23127 , \23154 );
not \U$22813 ( \23156 , \22032 );
not \U$22814 ( \23157 , \6286 );
or \U$22815 ( \23158 , \23156 , \23157 );
not \U$22816 ( \23159 , \22425 );
or \U$22817 ( \23160 , \23159 , \6283 );
nand \U$22818 ( \23161 , \23158 , \23160 );
and \U$22819 ( \23162 , \23155 , \23161 );
and \U$22820 ( \23163 , \23127 , \23154 );
nor \U$22821 ( \23164 , \23162 , \23163 );
not \U$22822 ( \23165 , \23164 );
xor \U$22823 ( \23166 , \22123 , \22129 );
xor \U$22824 ( \23167 , \23166 , \22136 );
not \U$22825 ( \23168 , \23167 );
or \U$22826 ( \23169 , \23165 , \23168 );
or \U$22827 ( \23170 , \23167 , \23164 );
nand \U$22828 ( \23171 , \23169 , \23170 );
not \U$22829 ( \23172 , \23171 );
or \U$22830 ( \23173 , \23121 , \23172 );
not \U$22831 ( \23174 , \23164 );
nand \U$22832 ( \23175 , \23174 , \23167 );
nand \U$22833 ( \23176 , \23173 , \23175 );
and \U$22834 ( \23177 , \23118 , \23176 );
nor \U$22835 ( \23178 , \23115 , \23117 );
nor \U$22836 ( \23179 , \23177 , \23178 );
not \U$22837 ( \23180 , \23179 );
not \U$22838 ( \23181 , \23180 );
or \U$22839 ( \23182 , \23113 , \23181 );
not \U$22840 ( \23183 , \23111 );
not \U$22841 ( \23184 , \23179 );
or \U$22842 ( \23185 , \23183 , \23184 );
xor \U$22843 ( \23186 , \21851 , \21861 );
xnor \U$22844 ( \23187 , \23186 , \21748 );
not \U$22845 ( \23188 , \23187 );
xor \U$22846 ( \23189 , \22139 , \22145 );
xor \U$22847 ( \23190 , \23189 , \22185 );
not \U$22848 ( \23191 , \23190 );
xor \U$22849 ( \23192 , \22156 , \22169 );
xnor \U$22850 ( \23193 , \23192 , \22182 );
not \U$22851 ( \23194 , \23193 );
xor \U$22852 ( \23195 , \22097 , \22104 );
xnor \U$22853 ( \23196 , \23195 , \22116 );
not \U$22854 ( \23197 , \23196 );
or \U$22855 ( \23198 , \23194 , \23197 );
xor \U$22856 ( \23199 , \22067 , \22073 );
xor \U$22857 ( \23200 , \23199 , \22083 );
nand \U$22858 ( \23201 , \23198 , \23200 );
not \U$22859 ( \23202 , \23193 );
not \U$22860 ( \23203 , \23196 );
nand \U$22861 ( \23204 , \23202 , \23203 );
nand \U$22862 ( \23205 , \23191 , \23201 , \23204 );
not \U$22863 ( \23206 , \23205 );
or \U$22864 ( \23207 , \23188 , \23206 );
nand \U$22865 ( \23208 , \23201 , \23204 );
nand \U$22866 ( \23209 , \23208 , \23190 );
nand \U$22867 ( \23210 , \23207 , \23209 );
nand \U$22868 ( \23211 , \23185 , \23210 );
nand \U$22869 ( \23212 , \23182 , \23211 );
xor \U$22870 ( \23213 , \23103 , \23212 );
not \U$22871 ( \23214 , \23213 );
or \U$22872 ( \23215 , \22899 , \23214 );
not \U$22873 ( \23216 , \23102 );
not \U$22874 ( \23217 , \23100 );
or \U$22875 ( \23218 , \23216 , \23217 );
nand \U$22876 ( \23219 , \23218 , \23212 );
nand \U$22877 ( \23220 , \23215 , \23219 );
and \U$22878 ( \23221 , \22895 , \23220 );
not \U$22879 ( \23222 , \22895 );
not \U$22880 ( \23223 , \23220 );
and \U$22881 ( \23224 , \23222 , \23223 );
nor \U$22882 ( \23225 , \23221 , \23224 );
not \U$22883 ( \23226 , \23225 );
or \U$22884 ( \23227 , \22886 , \23226 );
nand \U$22885 ( \23228 , \23220 , \22895 );
nand \U$22886 ( \23229 , \23227 , \23228 );
nand \U$22887 ( \23230 , \22252 , \23229 );
or \U$22888 ( \23231 , \22250 , \22244 );
nand \U$22889 ( \23232 , \23230 , \23231 );
nand \U$22890 ( \23233 , \22239 , \23232 );
nand \U$22891 ( \23234 , \22237 , \23233 );
not \U$22892 ( \23235 , \21474 );
nand \U$22893 ( \23236 , \23235 , \21476 , \20898 );
nand \U$22894 ( \23237 , \21481 , \22236 );
nand \U$22895 ( \23238 , \23234 , \23236 , \23237 );
nand \U$22896 ( \23239 , \21479 , \23238 );
xor \U$22897 ( \23240 , \20916 , \20975 );
and \U$22898 ( \23241 , \23240 , \21094 );
and \U$22899 ( \23242 , \20916 , \20975 );
or \U$22900 ( \23243 , \23241 , \23242 );
not \U$22901 ( \23244 , \21203 );
xor \U$22902 ( \23245 , \21223 , \21213 );
not \U$22903 ( \23246 , \23245 );
or \U$22904 ( \23247 , \23244 , \23246 );
nand \U$22905 ( \23248 , \21223 , \21213 );
nand \U$22906 ( \23249 , \23247 , \23248 );
xor \U$22907 ( \23250 , \21233 , \21242 );
and \U$22908 ( \23251 , \23250 , \21253 );
and \U$22909 ( \23252 , \21233 , \21242 );
or \U$22910 ( \23253 , \23251 , \23252 );
xor \U$22911 ( \23254 , \23249 , \23253 );
xor \U$22912 ( \23255 , \21167 , \21177 );
and \U$22913 ( \23256 , \23255 , \21187 );
and \U$22914 ( \23257 , \21167 , \21177 );
or \U$22915 ( \23258 , \23256 , \23257 );
xor \U$22916 ( \23259 , \23254 , \23258 );
not \U$22917 ( \23260 , \23259 );
xor \U$22918 ( \23261 , \21224 , \21254 );
and \U$22919 ( \23262 , \23261 , \21289 );
and \U$22920 ( \23263 , \21224 , \21254 );
or \U$22921 ( \23264 , \23262 , \23263 );
not \U$22922 ( \23265 , \23264 );
not \U$22923 ( \23266 , \23265 );
or \U$22924 ( \23267 , \23260 , \23266 );
or \U$22925 ( \23268 , \23259 , \23265 );
nand \U$22926 ( \23269 , \23267 , \23268 );
not \U$22927 ( \23270 , \21188 );
not \U$22928 ( \23271 , \21157 );
or \U$22929 ( \23272 , \23270 , \23271 );
not \U$22930 ( \23273 , \21151 );
not \U$22931 ( \23274 , \21145 );
or \U$22932 ( \23275 , \23273 , \23274 );
nand \U$22933 ( \23276 , \23275 , \21142 );
nand \U$22934 ( \23277 , \23272 , \23276 );
not \U$22935 ( \23278 , \23277 );
and \U$22936 ( \23279 , \23269 , \23278 );
not \U$22937 ( \23280 , \23269 );
and \U$22938 ( \23281 , \23280 , \23277 );
nor \U$22939 ( \23282 , \23279 , \23281 );
not \U$22940 ( \23283 , \21109 );
not \U$22941 ( \23284 , \21294 );
or \U$22942 ( \23285 , \23283 , \23284 );
not \U$22943 ( \23286 , \21193 );
nand \U$22944 ( \23287 , \23286 , \21290 );
nand \U$22945 ( \23288 , \23285 , \23287 );
xnor \U$22946 ( \23289 , \23282 , \23288 );
not \U$22947 ( \23290 , \23289 );
not \U$22948 ( \23291 , \2087 );
not \U$22949 ( \23292 , \13895 );
or \U$22950 ( \23293 , \23291 , \23292 );
nand \U$22951 ( \23294 , \21025 , \2071 );
nand \U$22952 ( \23295 , \23293 , \23294 );
not \U$22953 ( \23296 , \21060 );
not \U$22954 ( \23297 , \21052 );
or \U$22955 ( \23298 , \23296 , \23297 );
not \U$22956 ( \23299 , \21054 );
nand \U$22957 ( \23300 , \23299 , \21056 );
nand \U$22958 ( \23301 , \23298 , \23300 );
not \U$22959 ( \23302 , \23301 );
not \U$22960 ( \23303 , \23302 );
not \U$22961 ( \23304 , \11433 );
not \U$22962 ( \23305 , \21015 );
or \U$22963 ( \23306 , \23304 , \23305 );
nand \U$22964 ( \23307 , \13826 , \6145 );
nand \U$22965 ( \23308 , \23306 , \23307 );
not \U$22966 ( \23309 , \23308 );
or \U$22967 ( \23310 , \23303 , \23309 );
or \U$22968 ( \23311 , \23308 , \23302 );
nand \U$22969 ( \23312 , \23310 , \23311 );
xor \U$22970 ( \23313 , \23295 , \23312 );
not \U$22971 ( \23314 , \5653 );
not \U$22972 ( \23315 , RI9872568_156);
not \U$22973 ( \23316 , \4370 );
or \U$22974 ( \23317 , \23315 , \23316 );
or \U$22975 ( \23318 , \3861 , RI9872568_156);
nand \U$22976 ( \23319 , \23317 , \23318 );
not \U$22977 ( \23320 , \23319 );
or \U$22978 ( \23321 , \23314 , \23320 );
nand \U$22979 ( \23322 , \21165 , \5642 );
nand \U$22980 ( \23323 , \23321 , \23322 );
not \U$22981 ( \23324 , \5034 );
not \U$22982 ( \23325 , \21067 );
or \U$22983 ( \23326 , \23324 , \23325 );
and \U$22984 ( \23327 , \4154 , \5025 );
not \U$22985 ( \23328 , \4154 );
and \U$22986 ( \23329 , \23328 , RI9872478_154);
nor \U$22987 ( \23330 , \23327 , \23329 );
nand \U$22988 ( \23331 , \5036 , \23330 );
nand \U$22989 ( \23332 , \23326 , \23331 );
xor \U$22990 ( \23333 , \23323 , \23332 );
not \U$22991 ( \23334 , \10242 );
not \U$22992 ( \23335 , RI9872d60_173);
not \U$22993 ( \23336 , \6225 );
or \U$22994 ( \23337 , \23335 , \23336 );
or \U$22995 ( \23338 , \2216 , RI9872d60_173);
nand \U$22996 ( \23339 , \23337 , \23338 );
not \U$22997 ( \23340 , \23339 );
or \U$22998 ( \23341 , \23334 , \23340 );
nand \U$22999 ( \23342 , \10251 , \21137 );
nand \U$23000 ( \23343 , \23341 , \23342 );
xor \U$23001 ( \23344 , \23333 , \23343 );
xor \U$23002 ( \23345 , \23313 , \23344 );
not \U$23003 ( \23346 , \9214 );
and \U$23004 ( \23347 , RI9872b80_169, \1603 );
not \U$23005 ( \23348 , RI9872b80_169);
and \U$23006 ( \23349 , \23348 , \1370 );
or \U$23007 ( \23350 , \23347 , \23349 );
not \U$23008 ( \23351 , \23350 );
or \U$23009 ( \23352 , \23346 , \23351 );
nand \U$23010 ( \23353 , \21282 , \10679 );
nand \U$23011 ( \23354 , \23352 , \23353 );
not \U$23012 ( \23355 , \18957 );
not \U$23013 ( \23356 , \21238 );
or \U$23014 ( \23357 , \23355 , \23356 );
not \U$23015 ( \23358 , \22675 );
not \U$23016 ( \23359 , \2982 );
or \U$23017 ( \23360 , \23358 , \23359 );
or \U$23018 ( \23361 , \2982 , \18012 );
nand \U$23019 ( \23362 , \23360 , \23361 );
nand \U$23020 ( \23363 , \23362 , \13484 );
nand \U$23021 ( \23364 , \23357 , \23363 );
xor \U$23022 ( \23365 , \23354 , \23364 );
not \U$23023 ( \23366 , \9952 );
not \U$23024 ( \23367 , \21270 );
or \U$23025 ( \23368 , \23366 , \23367 );
not \U$23026 ( \23369 , \14132 );
not \U$23027 ( \23370 , \10674 );
or \U$23028 ( \23371 , \23369 , \23370 );
nand \U$23029 ( \23372 , \7092 , RI9873030_179);
nand \U$23030 ( \23373 , \23371 , \23372 );
nand \U$23031 ( \23374 , \23373 , \9937 );
nand \U$23032 ( \23375 , \23368 , \23374 );
xor \U$23033 ( \23376 , \23365 , \23375 );
xnor \U$23034 ( \23377 , \23345 , \23376 );
not \U$23035 ( \23378 , \23377 );
not \U$23036 ( \23379 , \23378 );
not \U$23037 ( \23380 , \3467 );
not \U$23038 ( \23381 , RI98726d0_159);
not \U$23039 ( \23382 , \5776 );
or \U$23040 ( \23383 , \23381 , \23382 );
nand \U$23041 ( \23384 , \7028 , \3593 );
nand \U$23042 ( \23385 , \23383 , \23384 );
not \U$23043 ( \23386 , \23385 );
or \U$23044 ( \23387 , \23380 , \23386 );
nand \U$23045 ( \23388 , \21375 , \3465 );
nand \U$23046 ( \23389 , \23387 , \23388 );
not \U$23047 ( \23390 , \5847 );
not \U$23048 ( \23391 , \4960 );
and \U$23049 ( \23392 , \23391 , \4088 );
not \U$23050 ( \23393 , \23391 );
and \U$23051 ( \23394 , \23393 , RI98725e0_157);
nor \U$23052 ( \23395 , \23392 , \23394 );
not \U$23053 ( \23396 , \23395 );
or \U$23054 ( \23397 , \23390 , \23396 );
nand \U$23055 ( \23398 , \21199 , \4101 );
nand \U$23056 ( \23399 , \23397 , \23398 );
xor \U$23057 ( \23400 , \23389 , \23399 );
not \U$23058 ( \23401 , \9227 );
and \U$23059 ( \23402 , RI9872bf8_170, \11559 );
not \U$23060 ( \23403 , RI9872bf8_170);
and \U$23061 ( \23404 , \23403 , \1658 );
nor \U$23062 ( \23405 , \23402 , \23404 );
not \U$23063 ( \23406 , \23405 );
or \U$23064 ( \23407 , \23401 , \23406 );
nand \U$23065 ( \23408 , \21211 , \9670 );
nand \U$23066 ( \23409 , \23407 , \23408 );
xor \U$23067 ( \23410 , \23400 , \23409 );
not \U$23068 ( \23411 , \9072 );
and \U$23069 ( \23412 , \18904 , \7901 );
not \U$23070 ( \23413 , \18904 );
and \U$23071 ( \23414 , \23413 , RI9872a18_166);
nor \U$23072 ( \23415 , \23412 , \23414 );
not \U$23073 ( \23416 , \23415 );
or \U$23074 ( \23417 , \23411 , \23416 );
nand \U$23075 ( \23418 , \21251 , \9079 );
nand \U$23076 ( \23419 , \23417 , \23418 );
not \U$23077 ( \23420 , \8752 );
and \U$23078 ( \23421 , \1274 , RI9872f40_177);
not \U$23079 ( \23422 , \1274 );
and \U$23080 ( \23423 , \23422 , \8732 );
nor \U$23081 ( \23424 , \23421 , \23423 );
not \U$23082 ( \23425 , \23424 );
or \U$23083 ( \23426 , \23420 , \23425 );
nand \U$23084 ( \23427 , \21185 , \8743 );
nand \U$23085 ( \23428 , \23426 , \23427 );
xor \U$23086 ( \23429 , \23419 , \23428 );
not \U$23087 ( \23430 , \7338 );
and \U$23088 ( \23431 , \1191 , \7333 );
not \U$23089 ( \23432 , \1191 );
and \U$23090 ( \23433 , \23432 , RI98729a0_165);
nor \U$23091 ( \23434 , \23431 , \23433 );
not \U$23092 ( \23435 , \23434 );
or \U$23093 ( \23436 , \23430 , \23435 );
nand \U$23094 ( \23437 , \21229 , \7326 );
nand \U$23095 ( \23438 , \23436 , \23437 );
xnor \U$23096 ( \23439 , \23429 , \23438 );
xor \U$23097 ( \23440 , \23410 , \23439 );
not \U$23098 ( \23441 , \6284 );
not \U$23099 ( \23442 , \21173 );
or \U$23100 ( \23443 , \23441 , \23442 );
and \U$23101 ( \23444 , \2111 , RI98728b0_163);
not \U$23102 ( \23445 , \2111 );
and \U$23103 ( \23446 , \23445 , \5632 );
nor \U$23104 ( \23447 , \23444 , \23446 );
nand \U$23105 ( \23448 , \23447 , \6611 );
nand \U$23106 ( \23449 , \23443 , \23448 );
not \U$23107 ( \23450 , \11350 );
not \U$23108 ( \23451 , \21260 );
or \U$23109 ( \23452 , \23450 , \23451 );
and \U$23110 ( \23453 , RI98730a8_180, \1106 );
not \U$23111 ( \23454 , RI98730a8_180);
and \U$23112 ( \23455 , \23454 , \1097 );
nor \U$23113 ( \23456 , \23453 , \23455 );
nand \U$23114 ( \23457 , \23456 , \12868 );
nand \U$23115 ( \23458 , \23452 , \23457 );
xor \U$23116 ( \23459 , \23449 , \23458 );
not \U$23117 ( \23460 , \9273 );
not \U$23118 ( \23461 , RI9872e50_175);
not \U$23119 ( \23462 , \6443 );
or \U$23120 ( \23463 , \23461 , \23462 );
or \U$23121 ( \23464 , \19218 , RI9872e50_175);
nand \U$23122 ( \23465 , \23463 , \23464 );
not \U$23123 ( \23466 , \23465 );
or \U$23124 ( \23467 , \23460 , \23466 );
nand \U$23125 ( \23468 , \21078 , \9686 );
nand \U$23126 ( \23469 , \23467 , \23468 );
xor \U$23127 ( \23470 , \23459 , \23469 );
xnor \U$23128 ( \23471 , \23440 , \23470 );
not \U$23129 ( \23472 , \23471 );
not \U$23130 ( \23473 , \23472 );
or \U$23131 ( \23474 , \23379 , \23473 );
nand \U$23132 ( \23475 , \23471 , \23377 );
nand \U$23133 ( \23476 , \23474 , \23475 );
xor \U$23134 ( \23477 , \20904 , \20910 );
and \U$23135 ( \23478 , \23477 , \20915 );
and \U$23136 ( \23479 , \20904 , \20910 );
or \U$23137 ( \23480 , \23478 , \23479 );
not \U$23138 ( \23481 , \23480 );
and \U$23139 ( \23482 , \23476 , \23481 );
not \U$23140 ( \23483 , \23476 );
and \U$23141 ( \23484 , \23483 , \23480 );
nor \U$23142 ( \23485 , \23482 , \23484 );
not \U$23143 ( \23486 , \23485 );
and \U$23144 ( \23487 , \23290 , \23486 );
and \U$23145 ( \23488 , \23289 , \23485 );
nor \U$23146 ( \23489 , \23487 , \23488 );
xor \U$23147 ( \23490 , \23243 , \23489 );
not \U$23148 ( \23491 , \21295 );
not \U$23149 ( \23492 , \21104 );
not \U$23150 ( \23493 , \23492 );
not \U$23151 ( \23494 , \21302 );
or \U$23152 ( \23495 , \23493 , \23494 );
or \U$23153 ( \23496 , \21302 , \23492 );
nand \U$23154 ( \23497 , \23495 , \23496 );
not \U$23155 ( \23498 , \23497 );
or \U$23156 ( \23499 , \23491 , \23498 );
nand \U$23157 ( \23500 , \21302 , \21104 );
nand \U$23158 ( \23501 , \23499 , \23500 );
xor \U$23159 ( \23502 , \23490 , \23501 );
not \U$23160 ( \23503 , \21454 );
not \U$23161 ( \23504 , \23503 );
not \U$23162 ( \23505 , \21449 );
or \U$23163 ( \23506 , \23504 , \23505 );
nand \U$23164 ( \23507 , \21336 , \21448 );
nand \U$23165 ( \23508 , \23506 , \23507 );
not \U$23166 ( \23509 , \23508 );
not \U$23167 ( \23510 , \23509 );
xor \U$23168 ( \23511 , \21362 , \21418 );
and \U$23169 ( \23512 , \23511 , \21430 );
and \U$23170 ( \23513 , \21362 , \21418 );
or \U$23171 ( \23514 , \23512 , \23513 );
not \U$23172 ( \23515 , \23514 );
not \U$23173 ( \23516 , \20937 );
not \U$23174 ( \23517 , \20926 );
or \U$23175 ( \23518 , \23516 , \23517 );
nand \U$23176 ( \23519 , \20925 , \20771 );
nand \U$23177 ( \23520 , \23518 , \23519 );
not \U$23178 ( \23521 , \23520 );
not \U$23179 ( \23522 , \4925 );
not \U$23180 ( \23523 , \4902 );
not \U$23181 ( \23524 , \13058 );
or \U$23182 ( \23525 , \23523 , \23524 );
nand \U$23183 ( \23526 , \5206 , RI9872388_152);
nand \U$23184 ( \23527 , \23525 , \23526 );
not \U$23185 ( \23528 , \23527 );
or \U$23186 ( \23529 , \23522 , \23528 );
nand \U$23187 ( \23530 , \21125 , \4919 );
nand \U$23188 ( \23531 , \23529 , \23530 );
not \U$23189 ( \23532 , \23531 );
not \U$23190 ( \23533 , \23532 );
or \U$23191 ( \23534 , \23521 , \23533 );
or \U$23192 ( \23535 , \23532 , \23520 );
nand \U$23193 ( \23536 , \23534 , \23535 );
not \U$23194 ( \23537 , \21400 );
not \U$23195 ( \23538 , \23537 );
not \U$23196 ( \23539 , \21377 );
or \U$23197 ( \23540 , \23538 , \23539 );
nand \U$23198 ( \23541 , \21388 , \21399 );
nand \U$23199 ( \23542 , \23540 , \23541 );
xor \U$23200 ( \23543 , \23536 , \23542 );
not \U$23201 ( \23544 , \21354 );
not \U$23202 ( \23545 , \23544 );
not \U$23203 ( \23546 , \21342 );
or \U$23204 ( \23547 , \23545 , \23546 );
nand \U$23205 ( \23548 , \23547 , \21356 );
and \U$23206 ( \23549 , \23543 , \23548 );
not \U$23207 ( \23550 , \23543 );
not \U$23208 ( \23551 , \23548 );
and \U$23209 ( \23552 , \23550 , \23551 );
nor \U$23210 ( \23553 , \23549 , \23552 );
not \U$23211 ( \23554 , \21413 );
not \U$23212 ( \23555 , \21409 );
or \U$23213 ( \23556 , \23554 , \23555 );
nand \U$23214 ( \23557 , \21368 , \21405 );
nand \U$23215 ( \23558 , \23556 , \23557 );
not \U$23216 ( \23559 , \23558 );
and \U$23217 ( \23560 , \23553 , \23559 );
not \U$23218 ( \23561 , \23553 );
and \U$23219 ( \23562 , \23561 , \23558 );
nor \U$23220 ( \23563 , \23560 , \23562 );
not \U$23221 ( \23564 , \23563 );
or \U$23222 ( \23565 , \23515 , \23564 );
or \U$23223 ( \23566 , \23514 , \23563 );
nand \U$23224 ( \23567 , \23565 , \23566 );
xor \U$23225 ( \23568 , \20951 , \20953 );
and \U$23226 ( \23569 , \23568 , \20964 );
and \U$23227 ( \23570 , \20951 , \20953 );
or \U$23228 ( \23571 , \23569 , \23570 );
buf \U$23229 ( \23572 , \23571 );
not \U$23230 ( \23573 , \20938 );
nand \U$23231 ( \23574 , \20941 , \23573 );
and \U$23232 ( \23575 , \23574 , \20946 );
nor \U$23233 ( \23576 , \23573 , \20941 );
nor \U$23234 ( \23577 , \23575 , \23576 );
not \U$23235 ( \23578 , \23577 );
xor \U$23236 ( \23579 , \21019 , \21029 );
and \U$23237 ( \23580 , \23579 , \21041 );
and \U$23238 ( \23581 , \21019 , \21029 );
or \U$23239 ( \23582 , \23580 , \23581 );
not \U$23240 ( \23583 , \23582 );
not \U$23241 ( \23584 , \20989 );
not \U$23242 ( \23585 , \20999 );
or \U$23243 ( \23586 , \23584 , \23585 );
or \U$23244 ( \23587 , \20999 , \20989 );
nand \U$23245 ( \23588 , \23587 , \21009 );
nand \U$23246 ( \23589 , \23586 , \23588 );
not \U$23247 ( \23590 , \1013 );
not \U$23248 ( \23591 , \14195 );
or \U$23249 ( \23592 , \23590 , \23591 );
nand \U$23250 ( \23593 , \20932 , \1018 );
nand \U$23251 ( \23594 , \23592 , \23593 );
nor \U$23252 ( \23595 , \23594 , \13935 );
not \U$23253 ( \23596 , \23595 );
nand \U$23254 ( \23597 , \23594 , \13935 );
nand \U$23255 ( \23598 , \23596 , \23597 );
not \U$23256 ( \23599 , \3170 );
not \U$23257 ( \23600 , \13905 );
or \U$23258 ( \23601 , \23599 , \23600 );
nand \U$23259 ( \23602 , \21036 , \3163 );
nand \U$23260 ( \23603 , \23601 , \23602 );
xnor \U$23261 ( \23604 , \23598 , \23603 );
xor \U$23262 ( \23605 , \23589 , \23604 );
not \U$23263 ( \23606 , \23605 );
not \U$23264 ( \23607 , \23606 );
or \U$23265 ( \23608 , \23583 , \23607 );
not \U$23266 ( \23609 , \23582 );
nand \U$23267 ( \23610 , \23609 , \23605 );
nand \U$23268 ( \23611 , \23608 , \23610 );
not \U$23269 ( \23612 , \23611 );
or \U$23270 ( \23613 , \23578 , \23612 );
or \U$23271 ( \23614 , \23611 , \23577 );
nand \U$23272 ( \23615 , \23613 , \23614 );
not \U$23273 ( \23616 , \23615 );
and \U$23274 ( \23617 , \23572 , \23616 );
not \U$23275 ( \23618 , \23572 );
and \U$23276 ( \23619 , \23618 , \23615 );
nor \U$23277 ( \23620 , \23617 , \23619 );
and \U$23278 ( \23621 , \23567 , \23620 );
not \U$23279 ( \23622 , \23567 );
not \U$23280 ( \23623 , \23620 );
and \U$23281 ( \23624 , \23622 , \23623 );
nor \U$23282 ( \23625 , \23621 , \23624 );
not \U$23283 ( \23626 , \21438 );
not \U$23284 ( \23627 , \21444 );
or \U$23285 ( \23628 , \23626 , \23627 );
not \U$23286 ( \23629 , \21436 );
nand \U$23287 ( \23630 , \23628 , \23629 );
xor \U$23288 ( \23631 , \23625 , \23630 );
buf \U$23289 ( \23632 , \23631 );
not \U$23290 ( \23633 , \23632 );
xor \U$23291 ( \23634 , \20947 , \20965 );
and \U$23292 ( \23635 , \23634 , \20974 );
and \U$23293 ( \23636 , \20947 , \20965 );
or \U$23294 ( \23637 , \23635 , \23636 );
not \U$23295 ( \23638 , \23637 );
not \U$23296 ( \23639 , \23638 );
not \U$23297 ( \23640 , \21272 );
not \U$23298 ( \23641 , \21284 );
or \U$23299 ( \23642 , \23640 , \23641 );
not \U$23300 ( \23643 , \21285 );
not \U$23301 ( \23644 , \21273 );
or \U$23302 ( \23645 , \23643 , \23644 );
nand \U$23303 ( \23646 , \23645 , \21262 );
nand \U$23304 ( \23647 , \23642 , \23646 );
not \U$23305 ( \23648 , \23647 );
not \U$23306 ( \23649 , \23648 );
not \U$23307 ( \23650 , \21050 );
not \U$23308 ( \23651 , \9429 );
or \U$23309 ( \23652 , \23650 , \23651 );
nand \U$23310 ( \23653 , \6316 , \14183 );
nand \U$23311 ( \23654 , \23652 , \23653 );
not \U$23312 ( \23655 , \1352 );
not \U$23313 ( \23656 , \13880 );
or \U$23314 ( \23657 , \23655 , \23656 );
nand \U$23315 ( \23658 , \21397 , \1380 );
nand \U$23316 ( \23659 , \23657 , \23658 );
xor \U$23317 ( \23660 , \23654 , \23659 );
not \U$23318 ( \23661 , \859 );
not \U$23319 ( \23662 , \20921 );
or \U$23320 ( \23663 , \23661 , \23662 );
nand \U$23321 ( \23664 , \832 , \14205 );
nand \U$23322 ( \23665 , \23663 , \23664 );
xor \U$23323 ( \23666 , \23660 , \23665 );
not \U$23324 ( \23667 , \23666 );
not \U$23325 ( \23668 , \21141 );
not \U$23326 ( \23669 , \21131 );
or \U$23327 ( \23670 , \23668 , \23669 );
not \U$23328 ( \23671 , \21116 );
nand \U$23329 ( \23672 , \23671 , \21127 );
nand \U$23330 ( \23673 , \23670 , \23672 );
not \U$23331 ( \23674 , \23673 );
not \U$23332 ( \23675 , \23674 );
or \U$23333 ( \23676 , \23667 , \23675 );
not \U$23334 ( \23677 , \23666 );
nand \U$23335 ( \23678 , \23677 , \23673 );
nand \U$23336 ( \23679 , \23676 , \23678 );
not \U$23337 ( \23680 , \23679 );
or \U$23338 ( \23681 , \23649 , \23680 );
or \U$23339 ( \23682 , \23679 , \23648 );
nand \U$23340 ( \23683 , \23681 , \23682 );
not \U$23341 ( \23684 , \1323 );
not \U$23342 ( \23685 , RI9871b18_134);
not \U$23343 ( \23686 , \11406 );
or \U$23344 ( \23687 , \23685 , \23686 );
or \U$23345 ( \23688 , \11406 , RI9871b18_134);
nand \U$23346 ( \23689 , \23687 , \23688 );
not \U$23347 ( \23690 , \23689 );
or \U$23348 ( \23691 , \23684 , \23690 );
not \U$23349 ( \23692 , \1293 );
nand \U$23350 ( \23693 , \23692 , \21007 );
nand \U$23351 ( \23694 , \23691 , \23693 );
not \U$23352 ( \23695 , \6673 );
not \U$23353 ( \23696 , \13846 );
or \U$23354 ( \23697 , \23695 , \23696 );
nand \U$23355 ( \23698 , \20987 , \1083 );
nand \U$23356 ( \23699 , \23697 , \23698 );
xor \U$23357 ( \23700 , \23694 , \23699 );
not \U$23358 ( \23701 , \1430 );
not \U$23359 ( \23702 , \13834 );
or \U$23360 ( \23703 , \23701 , \23702 );
not \U$23361 ( \23704 , \20997 );
or \U$23362 ( \23705 , \23704 , \1457 );
nand \U$23363 ( \23706 , \23703 , \23705 );
xor \U$23364 ( \23707 , \23700 , \23706 );
not \U$23365 ( \23708 , \919 );
not \U$23366 ( \23709 , \9750 );
or \U$23367 ( \23710 , \23708 , \23709 );
not \U$23368 ( \23711 , \18328 );
buf \U$23369 ( \23712 , \23711 );
not \U$23370 ( \23713 , \23712 );
nand \U$23371 ( \23714 , \23713 , RI9872130_147);
nand \U$23372 ( \23715 , \23710 , \23714 );
and \U$23373 ( \23716 , \23715 , \924 );
not \U$23374 ( \23717 , \21386 );
nor \U$23375 ( \23718 , \23717 , \7927 );
nor \U$23376 ( \23719 , \23716 , \23718 );
and \U$23377 ( \23720 , RI9871c80_137, \8554 );
not \U$23378 ( \23721 , RI9871c80_137);
and \U$23379 ( \23722 , \23721 , \9764 );
or \U$23380 ( \23723 , \23720 , \23722 );
not \U$23381 ( \23724 , \23723 );
nor \U$23382 ( \23725 , \23724 , \1746 );
not \U$23383 ( \23726 , \21113 );
nor \U$23384 ( \23727 , \23726 , \1591 );
or \U$23385 ( \23728 , \23725 , \23727 );
xor \U$23386 ( \23729 , \23719 , \23728 );
not \U$23387 ( \23730 , \18508 );
not \U$23388 ( \23731 , \21221 );
or \U$23389 ( \23732 , \23730 , \23731 );
nand \U$23390 ( \23733 , \17528 , RI9873288_184);
nand \U$23391 ( \23734 , \23732 , \23733 );
buf \U$23392 ( \23735 , \23734 );
xnor \U$23393 ( \23736 , \23729 , \23735 );
xor \U$23394 ( \23737 , \23707 , \23736 );
not \U$23395 ( \23738 , \21071 );
not \U$23396 ( \23739 , \21061 );
not \U$23397 ( \23740 , \21082 );
or \U$23398 ( \23741 , \23739 , \23740 );
or \U$23399 ( \23742 , \21082 , \21061 );
nand \U$23400 ( \23743 , \23741 , \23742 );
not \U$23401 ( \23744 , \23743 );
or \U$23402 ( \23745 , \23738 , \23744 );
not \U$23403 ( \23746 , \21061 );
nand \U$23404 ( \23747 , \23746 , \21082 );
nand \U$23405 ( \23748 , \23745 , \23747 );
xor \U$23406 ( \23749 , \23737 , \23748 );
xor \U$23407 ( \23750 , \23683 , \23749 );
xor \U$23408 ( \23751 , \21010 , \21042 );
and \U$23409 ( \23752 , \23751 , \21083 );
and \U$23410 ( \23753 , \21010 , \21042 );
or \U$23411 ( \23754 , \23752 , \23753 );
xor \U$23412 ( \23755 , \23750 , \23754 );
not \U$23413 ( \23756 , \23755 );
and \U$23414 ( \23757 , \23639 , \23756 );
and \U$23415 ( \23758 , \23638 , \23755 );
nor \U$23416 ( \23759 , \23757 , \23758 );
not \U$23417 ( \23760 , \23759 );
xor \U$23418 ( \23761 , \21093 , \21084 );
not \U$23419 ( \23762 , \20980 );
and \U$23420 ( \23763 , \23761 , \23762 );
and \U$23421 ( \23764 , \21093 , \21084 );
or \U$23422 ( \23765 , \23763 , \23764 );
not \U$23423 ( \23766 , \23765 );
not \U$23424 ( \23767 , \23766 );
or \U$23425 ( \23768 , \23760 , \23767 );
or \U$23426 ( \23769 , \23766 , \23759 );
nand \U$23427 ( \23770 , \23768 , \23769 );
not \U$23428 ( \23771 , \23770 );
not \U$23429 ( \23772 , \23771 );
or \U$23430 ( \23773 , \23633 , \23772 );
not \U$23431 ( \23774 , \23631 );
nand \U$23432 ( \23775 , \23774 , \23770 );
nand \U$23433 ( \23776 , \23773 , \23775 );
not \U$23434 ( \23777 , \23776 );
not \U$23435 ( \23778 , \23777 );
or \U$23436 ( \23779 , \23510 , \23778 );
nand \U$23437 ( \23780 , \23776 , \23508 );
nand \U$23438 ( \23781 , \23779 , \23780 );
xor \U$23439 ( \23782 , \23502 , \23781 );
not \U$23440 ( \23783 , \23782 );
not \U$23441 ( \23784 , \21099 );
not \U$23442 ( \23785 , \21095 );
nand \U$23443 ( \23786 , \23785 , \21303 );
not \U$23444 ( \23787 , \23786 );
or \U$23445 ( \23788 , \23784 , \23787 );
not \U$23446 ( \23789 , \21303 );
nand \U$23447 ( \23790 , \23789 , \21095 );
nand \U$23448 ( \23791 , \23788 , \23790 );
not \U$23449 ( \23792 , \21467 );
not \U$23450 ( \23793 , \21462 );
or \U$23451 ( \23794 , \23792 , \23793 );
not \U$23452 ( \23795 , \21458 );
nand \U$23453 ( \23796 , \23795 , \21330 );
nand \U$23454 ( \23797 , \23794 , \23796 );
xor \U$23455 ( \23798 , \23791 , \23797 );
not \U$23456 ( \23799 , \23798 );
or \U$23457 ( \23800 , \23783 , \23799 );
not \U$23458 ( \23801 , \23782 );
not \U$23459 ( \23802 , \23801 );
or \U$23460 ( \23803 , \23798 , \23802 );
nand \U$23461 ( \23804 , \23800 , \23803 );
not \U$23462 ( \23805 , \21473 );
not \U$23463 ( \23806 , \23805 );
not \U$23464 ( \23807 , \21320 );
or \U$23465 ( \23808 , \23806 , \23807 );
not \U$23466 ( \23809 , \21304 );
nand \U$23467 ( \23810 , \23809 , \21316 );
nand \U$23468 ( \23811 , \23808 , \23810 );
nor \U$23469 ( \23812 , \23804 , \23811 );
not \U$23470 ( \23813 , \23812 );
nand \U$23471 ( \23814 , \23239 , \23813 );
xor \U$23472 ( \23815 , \22244 , \23229 );
xnor \U$23473 ( \23816 , \23815 , \22250 );
buf \U$23474 ( \23817 , \22005 );
and \U$23475 ( \23818 , \21874 , \21997 );
not \U$23476 ( \23819 , \21874 );
and \U$23477 ( \23820 , \23819 , \21998 );
nor \U$23478 ( \23821 , \23818 , \23820 );
xnor \U$23479 ( \23822 , \23817 , \23821 );
not \U$23480 ( \23823 , \23822 );
not \U$23481 ( \23824 , \23823 );
not \U$23482 ( \23825 , \22885 );
not \U$23483 ( \23826 , \23225 );
not \U$23484 ( \23827 , \23826 );
or \U$23485 ( \23828 , \23825 , \23827 );
not \U$23486 ( \23829 , \22885 );
nand \U$23487 ( \23830 , \23829 , \23225 );
nand \U$23488 ( \23831 , \23828 , \23830 );
not \U$23489 ( \23832 , \23831 );
or \U$23490 ( \23833 , \23824 , \23832 );
not \U$23491 ( \23834 , \23213 );
not \U$23492 ( \23835 , \22897 );
and \U$23493 ( \23836 , \23834 , \23835 );
and \U$23494 ( \23837 , \23213 , \22897 );
nor \U$23495 ( \23838 , \23836 , \23837 );
not \U$23496 ( \23839 , \23838 );
not \U$23497 ( \23840 , \23839 );
not \U$23498 ( \23841 , \23115 );
not \U$23499 ( \23842 , \23841 );
xor \U$23500 ( \23843 , \23176 , \23117 );
not \U$23501 ( \23844 , \23843 );
or \U$23502 ( \23845 , \23842 , \23844 );
or \U$23503 ( \23846 , \23843 , \23841 );
nand \U$23504 ( \23847 , \23845 , \23846 );
not \U$23505 ( \23848 , \23847 );
xor \U$23506 ( \23849 , \23190 , \23208 );
xnor \U$23507 ( \23850 , \23849 , \23187 );
nand \U$23508 ( \23851 , \23848 , \23850 );
not \U$23509 ( \23852 , \23851 );
xor \U$23510 ( \23853 , \22952 , \22957 );
xor \U$23511 ( \23854 , \23853 , \22963 );
not \U$23512 ( \23855 , \23854 );
xor \U$23513 ( \23856 , \23005 , \22994 );
xnor \U$23514 ( \23857 , \23856 , \23000 );
nand \U$23515 ( \23858 , \23855 , \23857 );
xor \U$23516 ( \23859 , \22972 , \22985 );
and \U$23517 ( \23860 , \23858 , \23859 );
not \U$23518 ( \23861 , \23854 );
nor \U$23519 ( \23862 , \23861 , \23857 );
nor \U$23520 ( \23863 , \23860 , \23862 );
not \U$23521 ( \23864 , \23863 );
xor \U$23522 ( \23865 , \23193 , \23203 );
xnor \U$23523 ( \23866 , \23865 , \23200 );
not \U$23524 ( \23867 , \23866 );
xor \U$23525 ( \23868 , \23065 , \23026 );
nand \U$23526 ( \23869 , \23867 , \23868 );
nand \U$23527 ( \23870 , \23864 , \23869 );
not \U$23528 ( \23871 , \23868 );
nand \U$23529 ( \23872 , \23871 , \23866 );
nand \U$23530 ( \23873 , \23870 , \23872 );
not \U$23531 ( \23874 , \23873 );
or \U$23532 ( \23875 , \23852 , \23874 );
not \U$23533 ( \23876 , \23850 );
nand \U$23534 ( \23877 , \23876 , \23847 );
nand \U$23535 ( \23878 , \23875 , \23877 );
not \U$23536 ( \23879 , \23878 );
xor \U$23537 ( \23880 , \23110 , \23180 );
xnor \U$23538 ( \23881 , \23880 , \23210 );
nand \U$23539 ( \23882 , \23879 , \23881 );
not \U$23540 ( \23883 , \23882 );
xor \U$23541 ( \23884 , \22264 , \22267 );
xnor \U$23542 ( \23885 , \23884 , \22873 );
not \U$23543 ( \23886 , \23885 );
or \U$23544 ( \23887 , \23883 , \23886 );
not \U$23545 ( \23888 , \23881 );
buf \U$23546 ( \23889 , \23878 );
nand \U$23547 ( \23890 , \23888 , \23889 );
nand \U$23548 ( \23891 , \23887 , \23890 );
not \U$23549 ( \23892 , \23891 );
or \U$23550 ( \23893 , \23840 , \23892 );
not \U$23551 ( \23894 , \23891 );
not \U$23552 ( \23895 , \23894 );
not \U$23553 ( \23896 , \23838 );
or \U$23554 ( \23897 , \23895 , \23896 );
xor \U$23555 ( \23898 , \21743 , \21745 );
xor \U$23556 ( \23899 , \23898 , \21863 );
not \U$23557 ( \23900 , \23098 );
not \U$23558 ( \23901 , \23092 );
not \U$23559 ( \23902 , \23901 );
or \U$23560 ( \23903 , \23900 , \23902 );
nand \U$23561 ( \23904 , \23903 , \23102 );
not \U$23562 ( \23905 , \23020 );
and \U$23563 ( \23906 , \23904 , \23905 );
not \U$23564 ( \23907 , \23904 );
and \U$23565 ( \23908 , \23907 , \23020 );
nor \U$23566 ( \23909 , \23906 , \23908 );
xor \U$23567 ( \23910 , \23899 , \23909 );
xnor \U$23568 ( \23911 , \23088 , \23072 );
not \U$23569 ( \23912 , \23911 );
xnor \U$23570 ( \23913 , \23015 , \22946 );
not \U$23571 ( \23914 , \23913 );
or \U$23572 ( \23915 , \23912 , \23914 );
xor \U$23573 ( \23916 , \22917 , \22922 );
xor \U$23574 ( \23917 , \23916 , \22933 );
not \U$23575 ( \23918 , \924 );
not \U$23576 ( \23919 , \22289 );
or \U$23577 ( \23920 , \23918 , \23919 );
not \U$23578 ( \23921 , RI9872130_147);
not \U$23579 ( \23922 , \18216 );
or \U$23580 ( \23923 , \23921 , \23922 );
not \U$23581 ( \23924 , \19519 );
or \U$23582 ( \23925 , \23924 , RI9872130_147);
nand \U$23583 ( \23926 , \23923 , \23925 );
nand \U$23584 ( \23927 , \23926 , \875 );
nand \U$23585 ( \23928 , \23920 , \23927 );
not \U$23586 ( \23929 , \23928 );
not \U$23587 ( \23930 , \924 );
not \U$23588 ( \23931 , \23926 );
or \U$23589 ( \23932 , \23930 , \23931 );
buf \U$23590 ( \23933 , \17701 );
not \U$23591 ( \23934 , \23933 );
and \U$23592 ( \23935 , RI9872130_147, \23934 );
not \U$23593 ( \23936 , RI9872130_147);
and \U$23594 ( \23937 , \23936 , \17703 );
or \U$23595 ( \23938 , \23935 , \23937 );
nand \U$23596 ( \23939 , \23938 , \875 );
nand \U$23597 ( \23940 , \23932 , \23939 );
not \U$23598 ( \23941 , \23940 );
and \U$23599 ( \23942 , \19383 , \1351 );
not \U$23600 ( \23943 , \832 );
not \U$23601 ( \23944 , \22470 );
or \U$23602 ( \23945 , \23943 , \23944 );
not \U$23603 ( \23946 , RI9871d70_139);
buf \U$23604 ( \23947 , \18192 );
not \U$23605 ( \23948 , \23947 );
not \U$23606 ( \23949 , \23948 );
not \U$23607 ( \23950 , \23949 );
or \U$23608 ( \23951 , \23946 , \23950 );
not \U$23609 ( \23952 , \23947 );
not \U$23610 ( \23953 , \23952 );
or \U$23611 ( \23954 , \23953 , RI9871d70_139);
nand \U$23612 ( \23955 , \23951 , \23954 );
nand \U$23613 ( \23956 , \23955 , \858 );
nand \U$23614 ( \23957 , \23945 , \23956 );
xor \U$23615 ( \23958 , \23942 , \23957 );
not \U$23616 ( \23959 , \23958 );
or \U$23617 ( \23960 , \23941 , \23959 );
nand \U$23618 ( \23961 , \23957 , \23942 );
nand \U$23619 ( \23962 , \23960 , \23961 );
not \U$23620 ( \23963 , \23962 );
not \U$23621 ( \23964 , \23963 );
or \U$23622 ( \23965 , \23929 , \23964 );
not \U$23623 ( \23966 , \23928 );
nand \U$23624 ( \23967 , \23966 , \23962 );
nand \U$23625 ( \23968 , \23965 , \23967 );
not \U$23626 ( \23969 , \23968 );
not \U$23627 ( \23970 , \1135 );
not \U$23628 ( \23971 , \23132 );
or \U$23629 ( \23972 , \23970 , \23971 );
not \U$23630 ( \23973 , \1111 );
not \U$23631 ( \23974 , \18152 );
or \U$23632 ( \23975 , \23973 , \23974 );
nand \U$23633 ( \23976 , \21393 , RI98718c0_129);
nand \U$23634 ( \23977 , \23975 , \23976 );
nand \U$23635 ( \23978 , \23977 , \1083 );
nand \U$23636 ( \23979 , \23972 , \23978 );
not \U$23637 ( \23980 , \23979 );
or \U$23638 ( \23981 , \23969 , \23980 );
nand \U$23639 ( \23982 , \23962 , \23928 );
nand \U$23640 ( \23983 , \23981 , \23982 );
not \U$23641 ( \23984 , \23983 );
and \U$23642 ( \23985 , RI9873030_179, \6333 );
not \U$23643 ( \23986 , RI9873030_179);
and \U$23644 ( \23987 , \23986 , \1038 );
or \U$23645 ( \23988 , \23985 , \23987 );
and \U$23646 ( \23989 , \23988 , \13109 );
not \U$23647 ( \23990 , \23045 );
nor \U$23648 ( \23991 , \23990 , \11581 );
nor \U$23649 ( \23992 , \23989 , \23991 );
not \U$23650 ( \23993 , \23992 );
not \U$23651 ( \23994 , \23993 );
or \U$23652 ( \23995 , \23984 , \23994 );
not \U$23653 ( \23996 , \23983 );
not \U$23654 ( \23997 , \23996 );
not \U$23655 ( \23998 , \23992 );
or \U$23656 ( \23999 , \23997 , \23998 );
not \U$23657 ( \24000 , \17371 );
xor \U$23658 ( \24001 , RI98733f0_187, \9205 );
not \U$23659 ( \24002 , \24001 );
or \U$23660 ( \24003 , \24000 , \24002 );
nand \U$23661 ( \24004 , \22931 , \17263 );
nand \U$23662 ( \24005 , \24003 , \24004 );
nand \U$23663 ( \24006 , \23999 , \24005 );
nand \U$23664 ( \24007 , \23995 , \24006 );
or \U$23665 ( \24008 , \23917 , \24007 );
xor \U$23666 ( \24009 , \23037 , \23053 );
xor \U$23667 ( \24010 , \24009 , \23047 );
nand \U$23668 ( \24011 , \24008 , \24010 );
nand \U$23669 ( \24012 , \23917 , \24007 );
nand \U$23670 ( \24013 , \24011 , \24012 );
not \U$23671 ( \24014 , \24013 );
nand \U$23672 ( \24015 , \22941 , \22911 );
and \U$23673 ( \24016 , \24015 , \22936 );
not \U$23674 ( \24017 , \24015 );
not \U$23675 ( \24018 , \22936 );
and \U$23676 ( \24019 , \24017 , \24018 );
nor \U$23677 ( \24020 , \24016 , \24019 );
nand \U$23678 ( \24021 , \24014 , \24020 );
not \U$23679 ( \24022 , \24021 );
xor \U$23680 ( \24023 , \22966 , \22989 );
xor \U$23681 ( \24024 , \24023 , \23010 );
not \U$23682 ( \24025 , \24024 );
or \U$23683 ( \24026 , \24022 , \24025 );
not \U$23684 ( \24027 , \24020 );
nand \U$23685 ( \24028 , \24027 , \24013 );
nand \U$23686 ( \24029 , \24026 , \24028 );
nand \U$23687 ( \24030 , \23915 , \24029 );
or \U$23688 ( \24031 , \23913 , \23911 );
nand \U$23689 ( \24032 , \24030 , \24031 );
and \U$23690 ( \24033 , \23910 , \24032 );
and \U$23691 ( \24034 , \23899 , \23909 );
or \U$23692 ( \24035 , \24033 , \24034 );
buf \U$23693 ( \24036 , \24035 );
nand \U$23694 ( \24037 , \23897 , \24036 );
nand \U$23695 ( \24038 , \23893 , \24037 );
not \U$23696 ( \24039 , \24038 );
nand \U$23697 ( \24040 , \23833 , \24039 );
not \U$23698 ( \24041 , \23831 );
nand \U$23699 ( \24042 , \24041 , \23822 );
nand \U$23700 ( \24043 , \24040 , \24042 );
nand \U$23701 ( \24044 , \23816 , \24043 );
not \U$23702 ( \24045 , \24044 );
xor \U$23703 ( \24046 , \22880 , \22257 );
xor \U$23704 ( \24047 , \24046 , \22878 );
xor \U$23705 ( \24048 , \24035 , \23894 );
xnor \U$23706 ( \24049 , \24048 , \23839 );
xor \U$23707 ( \24050 , \24047 , \24049 );
xor \U$23708 ( \24051 , \23847 , \23850 );
xnor \U$23709 ( \24052 , \24051 , \23873 );
not \U$23710 ( \24053 , \24052 );
xor \U$23711 ( \24054 , \23854 , \23859 );
xnor \U$23712 ( \24055 , \24054 , \23857 );
not \U$23713 ( \24056 , \24055 );
xor \U$23714 ( \24057 , \23983 , \23993 );
xnor \U$23715 ( \24058 , \24057 , \24005 );
xor \U$23716 ( \24059 , \22445 , \22499 );
not \U$23717 ( \24060 , \24059 );
nand \U$23718 ( \24061 , \24058 , \24060 );
not \U$23719 ( \24062 , \22842 );
not \U$23720 ( \24063 , \8752 );
or \U$23721 ( \24064 , \24062 , \24063 );
and \U$23722 ( \24065 , RI9872f40_177, \1485 );
not \U$23723 ( \24066 , RI9872f40_177);
and \U$23724 ( \24067 , \24066 , \6382 );
or \U$23725 ( \24068 , \24065 , \24067 );
nand \U$23726 ( \24069 , \24068 , \8743 );
nand \U$23727 ( \24070 , \24064 , \24069 );
not \U$23728 ( \24071 , \24070 );
not \U$23729 ( \24072 , \20147 );
not \U$23730 ( \24073 , \22711 );
or \U$23731 ( \24074 , \24072 , \24073 );
xnor \U$23732 ( \24075 , RI98734e0_189, \914 );
buf \U$23733 ( \24076 , \19034 );
nand \U$23734 ( \24077 , \24075 , \24076 );
nand \U$23735 ( \24078 , \24074 , \24077 );
not \U$23736 ( \24079 , \24078 );
not \U$23737 ( \24080 , \24079 );
buf \U$23738 ( \24081 , \22482 );
xor \U$23739 ( \24082 , \22493 , \24081 );
not \U$23740 ( \24083 , \24082 );
and \U$23741 ( \24084 , \24080 , \24083 );
and \U$23742 ( \24085 , \24079 , \24082 );
nor \U$23743 ( \24086 , \24084 , \24085 );
not \U$23744 ( \24087 , \24086 );
not \U$23745 ( \24088 , \24087 );
or \U$23746 ( \24089 , \24071 , \24088 );
nand \U$23747 ( \24090 , \24078 , \24082 );
nand \U$23748 ( \24091 , \24089 , \24090 );
and \U$23749 ( \24092 , \24061 , \24091 );
nor \U$23750 ( \24093 , \24058 , \24060 );
nor \U$23751 ( \24094 , \24092 , \24093 );
not \U$23752 ( \24095 , \24094 );
xor \U$23753 ( \24096 , \22688 , \22633 );
not \U$23754 ( \24097 , \22738 );
xnor \U$23755 ( \24098 , \24096 , \24097 );
not \U$23756 ( \24099 , \24098 );
or \U$23757 ( \24100 , \24095 , \24099 );
or \U$23758 ( \24101 , \24098 , \24094 );
nand \U$23759 ( \24102 , \24100 , \24101 );
not \U$23760 ( \24103 , \24102 );
or \U$23761 ( \24104 , \24056 , \24103 );
not \U$23762 ( \24105 , \24094 );
nand \U$23763 ( \24106 , \24105 , \24098 );
nand \U$23764 ( \24107 , \24104 , \24106 );
not \U$23765 ( \24108 , \24107 );
xor \U$23766 ( \24109 , \23868 , \23863 );
xnor \U$23767 ( \24110 , \24109 , \23866 );
not \U$23768 ( \24111 , \24013 );
not \U$23769 ( \24112 , \24020 );
and \U$23770 ( \24113 , \24111 , \24112 );
and \U$23771 ( \24114 , \24013 , \24020 );
nor \U$23772 ( \24115 , \24113 , \24114 );
xor \U$23773 ( \24116 , \24024 , \24115 );
nand \U$23774 ( \24117 , \24110 , \24116 );
not \U$23775 ( \24118 , \24117 );
or \U$23776 ( \24119 , \24108 , \24118 );
not \U$23777 ( \24120 , \24110 );
not \U$23778 ( \24121 , \24116 );
nand \U$23779 ( \24122 , \24120 , \24121 );
nand \U$23780 ( \24123 , \24119 , \24122 );
not \U$23781 ( \24124 , \24123 );
xor \U$23782 ( \24125 , \23911 , \24029 );
xnor \U$23783 ( \24126 , \24125 , \23913 );
not \U$23784 ( \24127 , \24126 );
or \U$23785 ( \24128 , \24124 , \24127 );
or \U$23786 ( \24129 , \24123 , \24126 );
nand \U$23787 ( \24130 , \24128 , \24129 );
not \U$23788 ( \24131 , \24130 );
or \U$23789 ( \24132 , \24053 , \24131 );
not \U$23790 ( \24133 , \24126 );
nand \U$23791 ( \24134 , \24133 , \24123 );
nand \U$23792 ( \24135 , \24132 , \24134 );
not \U$23793 ( \24136 , \24135 );
xor \U$23794 ( \24137 , \23899 , \23909 );
xor \U$23795 ( \24138 , \24137 , \24032 );
xnor \U$23796 ( \24139 , \22747 , \22863 );
not \U$23797 ( \24140 , \24139 );
xor \U$23798 ( \24141 , \22341 , \22383 );
xnor \U$23799 ( \24142 , \24141 , \22338 );
xor \U$23800 ( \24143 , \22813 , \22815 );
xor \U$23801 ( \24144 , \24143 , \22856 );
xor \U$23802 ( \24145 , \24142 , \24144 );
xor \U$23803 ( \24146 , \22700 , \22735 );
xnor \U$23804 ( \24147 , \24146 , \22731 );
not \U$23805 ( \24148 , \24147 );
not \U$23806 ( \24149 , \22321 );
not \U$23807 ( \24150 , \22335 );
not \U$23808 ( \24151 , \24150 );
and \U$23809 ( \24152 , \24149 , \24151 );
and \U$23810 ( \24153 , \22321 , \24150 );
nor \U$23811 ( \24154 , \24152 , \24153 );
xor \U$23812 ( \24155 , \22597 , \24154 );
xnor \U$23813 ( \24156 , \24155 , \22625 );
not \U$23814 ( \24157 , \24156 );
or \U$23815 ( \24158 , \24148 , \24157 );
not \U$23816 ( \24159 , \24154 );
not \U$23817 ( \24160 , \22597 );
not \U$23818 ( \24161 , \22625 );
not \U$23819 ( \24162 , \24161 );
or \U$23820 ( \24163 , \24160 , \24162 );
not \U$23821 ( \24164 , \22597 );
nand \U$23822 ( \24165 , \24164 , \22625 );
nand \U$23823 ( \24166 , \24163 , \24165 );
nand \U$23824 ( \24167 , \24159 , \24166 );
nand \U$23825 ( \24168 , \24158 , \24167 );
and \U$23826 ( \24169 , \24145 , \24168 );
and \U$23827 ( \24170 , \24142 , \24144 );
or \U$23828 ( \24171 , \24169 , \24170 );
nand \U$23829 ( \24172 , \24140 , \24171 );
not \U$23830 ( \24173 , \24172 );
not \U$23831 ( \24174 , \24171 );
not \U$23832 ( \24175 , \24174 );
not \U$23833 ( \24176 , \24139 );
or \U$23834 ( \24177 , \24175 , \24176 );
xor \U$23835 ( \24178 , \22543 , \22532 );
xor \U$23836 ( \24179 , \24178 , \22522 );
not \U$23837 ( \24180 , \9072 );
not \U$23838 ( \24181 , \22327 );
or \U$23839 ( \24182 , \24180 , \24181 );
and \U$23840 ( \24183 , RI9872a18_166, \5736 );
not \U$23841 ( \24184 , RI9872a18_166);
not \U$23842 ( \24185 , \4984 );
and \U$23843 ( \24186 , \24184 , \24185 );
or \U$23844 ( \24187 , \24183 , \24186 );
nand \U$23845 ( \24188 , \24187 , \8028 );
nand \U$23846 ( \24189 , \24182 , \24188 );
not \U$23847 ( \24190 , \24189 );
not \U$23848 ( \24191 , \9214 );
not \U$23849 ( \24192 , \22595 );
or \U$23850 ( \24193 , \24191 , \24192 );
not \U$23851 ( \24194 , RI9872b80_169);
not \U$23852 ( \24195 , \4470 );
or \U$23853 ( \24196 , \24194 , \24195 );
or \U$23854 ( \24197 , \4470 , RI9872b80_169);
nand \U$23855 ( \24198 , \24196 , \24197 );
nand \U$23856 ( \24199 , \24198 , \9196 );
nand \U$23857 ( \24200 , \24193 , \24199 );
not \U$23858 ( \24201 , \22618 );
not \U$23859 ( \24202 , \22610 );
or \U$23860 ( \24203 , \24201 , \24202 );
not \U$23861 ( \24204 , \13022 );
not \U$23862 ( \24205 , \1061 );
or \U$23863 ( \24206 , \24204 , \24205 );
or \U$23864 ( \24207 , \6573 , \13022 );
nand \U$23865 ( \24208 , \24206 , \24207 );
buf \U$23866 ( \24209 , \11350 );
nand \U$23867 ( \24210 , \24208 , \24209 );
nand \U$23868 ( \24211 , \24203 , \24210 );
xor \U$23869 ( \24212 , \24200 , \24211 );
not \U$23870 ( \24213 , \24212 );
or \U$23871 ( \24214 , \24190 , \24213 );
nand \U$23872 ( \24215 , \24200 , \24211 );
nand \U$23873 ( \24216 , \24214 , \24215 );
xor \U$23874 ( \24217 , \24179 , \24216 );
xor \U$23875 ( \24218 , \22826 , \22835 );
xor \U$23876 ( \24219 , \22852 , \24218 );
and \U$23877 ( \24220 , \24217 , \24219 );
and \U$23878 ( \24221 , \24179 , \24216 );
or \U$23879 ( \24222 , \24220 , \24221 );
not \U$23880 ( \24223 , \24222 );
xor \U$23881 ( \24224 , \22431 , \22503 );
xnor \U$23882 ( \24225 , \24224 , \22548 );
nand \U$23883 ( \24226 , \24223 , \24225 );
not \U$23884 ( \24227 , \24226 );
not \U$23885 ( \24228 , \17371 );
not \U$23886 ( \24229 , RI98733f0_187);
not \U$23887 ( \24230 , \8006 );
or \U$23888 ( \24231 , \24229 , \24230 );
nand \U$23889 ( \24232 , \8005 , \17539 );
nand \U$23890 ( \24233 , \24231 , \24232 );
not \U$23891 ( \24234 , \24233 );
or \U$23892 ( \24235 , \24228 , \24234 );
nand \U$23893 ( \24236 , \24001 , \17263 );
nand \U$23894 ( \24237 , \24235 , \24236 );
not \U$23895 ( \24238 , \24237 );
and \U$23896 ( \24239 , \22310 , \7338 );
not \U$23897 ( \24240 , RI98729a0_165);
not \U$23898 ( \24241 , \5761 );
or \U$23899 ( \24242 , \24240 , \24241 );
or \U$23900 ( \24243 , \6481 , RI98729a0_165);
nand \U$23901 ( \24244 , \24242 , \24243 );
and \U$23902 ( \24245 , \24244 , \7325 );
nor \U$23903 ( \24246 , \24239 , \24245 );
not \U$23904 ( \24247 , \24246 );
not \U$23905 ( \24248 , \9937 );
not \U$23906 ( \24249 , \23988 );
or \U$23907 ( \24250 , \24248 , \24249 );
not \U$23908 ( \24251 , \14132 );
not \U$23909 ( \24252 , \1211 );
or \U$23910 ( \24253 , \24251 , \24252 );
nand \U$23911 ( \24254 , \1210 , RI9873030_179);
nand \U$23912 ( \24255 , \24253 , \24254 );
nand \U$23913 ( \24256 , \24255 , \13109 );
nand \U$23914 ( \24257 , \24250 , \24256 );
not \U$23915 ( \24258 , \24257 );
or \U$23916 ( \24259 , \24247 , \24258 );
or \U$23917 ( \24260 , \24257 , \24246 );
nand \U$23918 ( \24261 , \24259 , \24260 );
not \U$23919 ( \24262 , \24261 );
or \U$23920 ( \24263 , \24238 , \24262 );
not \U$23921 ( \24264 , \24246 );
nand \U$23922 ( \24265 , \24264 , \24257 );
nand \U$23923 ( \24266 , \24263 , \24265 );
not \U$23924 ( \24267 , \24266 );
not \U$23925 ( \24268 , \17234 );
not \U$23926 ( \24269 , \22683 );
or \U$23927 ( \24270 , \24268 , \24269 );
not \U$23928 ( \24271 , RI9873210_183);
not \U$23929 ( \24272 , \17363 );
or \U$23930 ( \24273 , \24271 , \24272 );
or \U$23931 ( \24274 , \1340 , RI9873210_183);
nand \U$23932 ( \24275 , \24273 , \24274 );
nand \U$23933 ( \24276 , \24275 , \13477 );
nand \U$23934 ( \24277 , \24270 , \24276 );
not \U$23935 ( \24278 , \22604 );
not \U$23936 ( \24279 , RI9873648_192);
or \U$23937 ( \24280 , \24278 , \24279 );
not \U$23938 ( \24281 , \18239 );
not \U$23939 ( \24282 , \1306 );
or \U$23940 ( \24283 , \24281 , \24282 );
or \U$23941 ( \24284 , \1306 , \18239 );
nand \U$23942 ( \24285 , \24283 , \24284 );
nand \U$23943 ( \24286 , \24285 , \18545 );
nand \U$23944 ( \24287 , \24280 , \24286 );
xor \U$23945 ( \24288 , \24277 , \24287 );
not \U$23946 ( \24289 , \9670 );
and \U$23947 ( \24290 , \18647 , \9185 );
not \U$23948 ( \24291 , \18647 );
and \U$23949 ( \24292 , \24291 , RI9872bf8_170);
nor \U$23950 ( \24293 , \24290 , \24292 );
not \U$23951 ( \24294 , \24293 );
or \U$23952 ( \24295 , \24289 , \24294 );
nand \U$23953 ( \24296 , \22641 , \9227 );
nand \U$23954 ( \24297 , \24295 , \24296 );
and \U$23955 ( \24298 , \24288 , \24297 );
and \U$23956 ( \24299 , \24277 , \24287 );
or \U$23957 ( \24300 , \24298 , \24299 );
nand \U$23958 ( \24301 , \22729 , \17528 );
not \U$23959 ( \24302 , \22727 );
not \U$23960 ( \24303 , \942 );
or \U$23961 ( \24304 , \24302 , \24303 );
not \U$23962 ( \24305 , RI9873288_184);
or \U$23963 ( \24306 , \5908 , \24305 );
nand \U$23964 ( \24307 , \24304 , \24306 );
nand \U$23965 ( \24308 , \24307 , \19641 );
nand \U$23966 ( \24309 , \24301 , \24308 );
not \U$23967 ( \24310 , \8801 );
not \U$23968 ( \24311 , \22663 );
or \U$23969 ( \24312 , \24310 , \24311 );
not \U$23970 ( \24313 , \8811 );
not \U$23971 ( \24314 , \18685 );
or \U$23972 ( \24315 , \24313 , \24314 );
or \U$23973 ( \24316 , \18685 , \8811 );
nand \U$23974 ( \24317 , \24315 , \24316 );
nand \U$23975 ( \24318 , \24317 , \8819 );
nand \U$23976 ( \24319 , \24312 , \24318 );
xor \U$23977 ( \24320 , \24309 , \24319 );
not \U$23978 ( \24321 , \10333 );
not \U$23979 ( \24322 , \22691 );
or \U$23980 ( \24323 , \24321 , \24322 );
not \U$23981 ( \24324 , RI9872e50_175);
not \U$23982 ( \24325 , \2947 );
or \U$23983 ( \24326 , \24324 , \24325 );
or \U$23984 ( \24327 , \2947 , RI9872e50_175);
nand \U$23985 ( \24328 , \24326 , \24327 );
nand \U$23986 ( \24329 , \24328 , \18563 );
nand \U$23987 ( \24330 , \24323 , \24329 );
nand \U$23988 ( \24331 , \24320 , \24330 );
not \U$23989 ( \24332 , \24308 );
not \U$23990 ( \24333 , \24301 );
or \U$23991 ( \24334 , \24332 , \24333 );
nand \U$23992 ( \24335 , \24334 , \24319 );
nand \U$23993 ( \24336 , \24331 , \24335 );
xor \U$23994 ( \24337 , \24300 , \24336 );
not \U$23995 ( \24338 , \24337 );
or \U$23996 ( \24339 , \24267 , \24338 );
not \U$23997 ( \24340 , \24335 );
not \U$23998 ( \24341 , \24331 );
or \U$23999 ( \24342 , \24340 , \24341 );
nand \U$24000 ( \24343 , \24342 , \24300 );
nand \U$24001 ( \24344 , \24339 , \24343 );
not \U$24002 ( \24345 , \24344 );
or \U$24003 ( \24346 , \24227 , \24345 );
not \U$24004 ( \24347 , \24225 );
nand \U$24005 ( \24348 , \24347 , \24222 );
nand \U$24006 ( \24349 , \24346 , \24348 );
nand \U$24007 ( \24350 , \24177 , \24349 );
not \U$24008 ( \24351 , \24350 );
or \U$24009 ( \24352 , \24173 , \24351 );
not \U$24010 ( \24353 , \22388 );
and \U$24011 ( \24354 , \22561 , \24353 );
not \U$24012 ( \24355 , \22561 );
and \U$24013 ( \24356 , \24355 , \22388 );
nor \U$24014 ( \24357 , \24354 , \24356 );
not \U$24015 ( \24358 , \24357 );
not \U$24016 ( \24359 , \24358 );
xnor \U$24017 ( \24360 , \23171 , \23120 );
not \U$24018 ( \24361 , \24360 );
not \U$24019 ( \24362 , \3467 );
not \U$24020 ( \24363 , \22822 );
or \U$24021 ( \24364 , \24362 , \24363 );
not \U$24022 ( \24365 , RI98726d0_159);
not \U$24023 ( \24366 , \8842 );
or \U$24024 ( \24367 , \24365 , \24366 );
not \U$24025 ( \24368 , \9911 );
nand \U$24026 ( \24369 , \24368 , \3593 );
nand \U$24027 ( \24370 , \24367 , \24369 );
nand \U$24028 ( \24371 , \24370 , \13409 );
nand \U$24029 ( \24372 , \24364 , \24371 );
not \U$24030 ( \24373 , \24372 );
not \U$24031 ( \24374 , \3169 );
not \U$24032 ( \24375 , \22539 );
or \U$24033 ( \24376 , \24374 , \24375 );
and \U$24034 ( \24377 , RI9872310_151, \8722 );
not \U$24035 ( \24378 , RI9872310_151);
and \U$24036 ( \24379 , \24378 , \22752 );
nor \U$24037 ( \24380 , \24377 , \24379 );
nand \U$24038 ( \24381 , \24380 , \3163 );
nand \U$24039 ( \24382 , \24376 , \24381 );
not \U$24040 ( \24383 , \24382 );
not \U$24041 ( \24384 , \2087 );
not \U$24042 ( \24385 , \22831 );
or \U$24043 ( \24386 , \24384 , \24385 );
not \U$24044 ( \24387 , RI9871aa0_133);
not \U$24045 ( \24388 , \12460 );
or \U$24046 ( \24389 , \24387 , \24388 );
or \U$24047 ( \24390 , \12460 , RI9871aa0_133);
nand \U$24048 ( \24391 , \24389 , \24390 );
nand \U$24049 ( \24392 , \24391 , \2072 );
nand \U$24050 ( \24393 , \24386 , \24392 );
not \U$24051 ( \24394 , \24393 );
and \U$24052 ( \24395 , \24383 , \24394 );
not \U$24053 ( \24396 , \24383 );
and \U$24054 ( \24397 , \24396 , \24393 );
nor \U$24055 ( \24398 , \24395 , \24397 );
not \U$24056 ( \24399 , \24398 );
or \U$24057 ( \24400 , \24373 , \24399 );
nand \U$24058 ( \24401 , \24382 , \24393 );
nand \U$24059 ( \24402 , \24400 , \24401 );
not \U$24060 ( \24403 , \24402 );
not \U$24061 ( \24404 , \23136 );
not \U$24062 ( \24405 , \24404 );
not \U$24063 ( \24406 , \23147 );
and \U$24064 ( \24407 , \24405 , \24406 );
and \U$24065 ( \24408 , \23147 , \24404 );
nor \U$24066 ( \24409 , \24407 , \24408 );
xor \U$24067 ( \24410 , \22412 , \24409 );
xnor \U$24068 ( \24411 , \24410 , \22427 );
not \U$24069 ( \24412 , \24411 );
or \U$24070 ( \24413 , \24403 , \24412 );
not \U$24071 ( \24414 , \24409 );
xor \U$24072 ( \24415 , \22412 , \22427 );
nand \U$24073 ( \24416 , \24414 , \24415 );
nand \U$24074 ( \24417 , \24413 , \24416 );
not \U$24075 ( \24418 , \24417 );
xnor \U$24076 ( \24419 , \23155 , \23161 );
not \U$24077 ( \24420 , \24419 );
not \U$24078 ( \24421 , \6286 );
not \U$24079 ( \24422 , \22419 );
or \U$24080 ( \24423 , \24421 , \24422 );
not \U$24081 ( \24424 , \12805 );
xor \U$24082 ( \24425 , RI98728b0_163, \24424 );
nand \U$24083 ( \24426 , \24425 , \6284 );
nand \U$24084 ( \24427 , \24423 , \24426 );
not \U$24085 ( \24428 , \24427 );
not \U$24086 ( \24429 , \1292 );
not \U$24087 ( \24430 , RI9871b18_134);
not \U$24088 ( \24431 , \18710 );
or \U$24089 ( \24432 , \24430 , \24431 );
or \U$24090 ( \24433 , \20765 , RI9871b18_134);
nand \U$24091 ( \24434 , \24432 , \24433 );
not \U$24092 ( \24435 , \24434 );
or \U$24093 ( \24436 , \24429 , \24435 );
and \U$24094 ( \24437 , RI9871b18_134, \17013 );
not \U$24095 ( \24438 , RI9871b18_134);
not \U$24096 ( \24439 , \13860 );
and \U$24097 ( \24440 , \24438 , \24439 );
or \U$24098 ( \24441 , \24437 , \24440 );
nand \U$24099 ( \24442 , \24441 , \1323 );
nand \U$24100 ( \24443 , \24436 , \24442 );
not \U$24101 ( \24444 , \24443 );
or \U$24102 ( \24445 , \919 , \829 );
not \U$24103 ( \24446 , \829 );
not \U$24104 ( \24447 , \919 );
or \U$24105 ( \24448 , \24446 , \24447 );
not \U$24106 ( \24449 , \18704 );
not \U$24107 ( \24450 , \24449 );
nand \U$24108 ( \24451 , \24448 , \24450 );
nand \U$24109 ( \24452 , \24445 , \24451 , RI9871d70_139);
not \U$24110 ( \24453 , \24452 );
not \U$24111 ( \24454 , \832 );
not \U$24112 ( \24455 , \23955 );
or \U$24113 ( \24456 , \24454 , \24455 );
not \U$24114 ( \24457 , \8859 );
not \U$24115 ( \24458 , \21779 );
or \U$24116 ( \24459 , \24457 , \24458 );
or \U$24117 ( \24460 , \18704 , \1347 );
nand \U$24118 ( \24461 , \24459 , \24460 );
nand \U$24119 ( \24462 , \24461 , \858 );
nand \U$24120 ( \24463 , \24456 , \24462 );
nand \U$24121 ( \24464 , \24453 , \24463 );
not \U$24122 ( \24465 , \24464 );
not \U$24123 ( \24466 , \1500 );
not \U$24124 ( \24467 , RI9871c80_137);
not \U$24125 ( \24468 , \17868 );
or \U$24126 ( \24469 , \24467 , \24468 );
not \U$24127 ( \24470 , \19412 );
or \U$24128 ( \24471 , \24470 , RI9871c80_137);
nand \U$24129 ( \24472 , \24469 , \24471 );
not \U$24130 ( \24473 , \24472 );
or \U$24131 ( \24474 , \24466 , \24473 );
nand \U$24132 ( \24475 , \22491 , \1493 );
nand \U$24133 ( \24476 , \24474 , \24475 );
not \U$24134 ( \24477 , \24476 );
or \U$24135 ( \24478 , \24465 , \24477 );
or \U$24136 ( \24479 , \24476 , \24464 );
nand \U$24137 ( \24480 , \24478 , \24479 );
not \U$24138 ( \24481 , \24480 );
or \U$24139 ( \24482 , \24444 , \24481 );
not \U$24140 ( \24483 , \24464 );
nand \U$24141 ( \24484 , \24483 , \24476 );
nand \U$24142 ( \24485 , \24482 , \24484 );
not \U$24143 ( \24486 , \5034 );
not \U$24144 ( \24487 , \8915 );
xor \U$24145 ( \24488 , RI9872478_154, \24487 );
not \U$24146 ( \24489 , \24488 );
or \U$24147 ( \24490 , \24486 , \24489 );
nand \U$24148 ( \24491 , \22452 , \22459 );
nand \U$24149 ( \24492 , \24490 , \24491 );
xor \U$24150 ( \24493 , \24485 , \24492 );
not \U$24151 ( \24494 , \24493 );
or \U$24152 ( \24495 , \24428 , \24494 );
nand \U$24153 ( \24496 , \24492 , \24485 );
nand \U$24154 ( \24497 , \24495 , \24496 );
not \U$24155 ( \24498 , \24497 );
not \U$24156 ( \24499 , \791 );
not \U$24157 ( \24500 , \1078 );
not \U$24158 ( \24501 , \13065 );
not \U$24159 ( \24502 , \24501 );
not \U$24160 ( \24503 , \24502 );
or \U$24161 ( \24504 , \24500 , \24503 );
or \U$24162 ( \24505 , \13067 , \1078 );
nand \U$24163 ( \24506 , \24504 , \24505 );
not \U$24164 ( \24507 , \24506 );
or \U$24165 ( \24508 , \24499 , \24507 );
nand \U$24166 ( \24509 , \22403 , \6144 );
nand \U$24167 ( \24510 , \24508 , \24509 );
not \U$24168 ( \24511 , \24510 );
not \U$24169 ( \24512 , \1323 );
not \U$24170 ( \24513 , \22397 );
or \U$24171 ( \24514 , \24512 , \24513 );
nand \U$24172 ( \24515 , \24441 , \1292 );
nand \U$24173 ( \24516 , \24514 , \24515 );
not \U$24174 ( \24517 , \1429 );
not \U$24175 ( \24518 , \23142 );
or \U$24176 ( \24519 , \24517 , \24518 );
not \U$24177 ( \24520 , RI9871c08_136);
not \U$24178 ( \24521 , \17090 );
or \U$24179 ( \24522 , \24520 , \24521 );
not \U$24180 ( \24523 , \13281 );
or \U$24181 ( \24524 , \24523 , RI9871c08_136);
nand \U$24182 ( \24525 , \24522 , \24524 );
nand \U$24183 ( \24526 , \24525 , \1455 );
nand \U$24184 ( \24527 , \24519 , \24526 );
xor \U$24185 ( \24528 , \24516 , \24527 );
not \U$24186 ( \24529 , \24528 );
or \U$24187 ( \24530 , \24511 , \24529 );
nand \U$24188 ( \24531 , \24527 , \24516 );
nand \U$24189 ( \24532 , \24530 , \24531 );
not \U$24190 ( \24533 , \24532 );
nand \U$24191 ( \24534 , \24498 , \24533 );
not \U$24192 ( \24535 , \24534 );
not \U$24193 ( \24536 , \17098 );
not \U$24194 ( \24537 , \22528 );
or \U$24195 ( \24538 , \24536 , \24537 );
and \U$24196 ( \24539 , RI98725e0_157, \9881 );
not \U$24197 ( \24540 , RI98725e0_157);
and \U$24198 ( \24541 , \24540 , \9880 );
nor \U$24199 ( \24542 , \24539 , \24541 );
nand \U$24200 ( \24543 , \24542 , \8790 );
nand \U$24201 ( \24544 , \24538 , \24543 );
not \U$24202 ( \24545 , \24544 );
not \U$24203 ( \24546 , \4923 );
not \U$24204 ( \24547 , \22443 );
or \U$24205 ( \24548 , \24546 , \24547 );
not \U$24206 ( \24549 , \22347 );
xor \U$24207 ( \24550 , RI9872388_152, \24549 );
nand \U$24208 ( \24551 , \24550 , \4918 );
nand \U$24209 ( \24552 , \24548 , \24551 );
not \U$24210 ( \24553 , \5653 );
not \U$24211 ( \24554 , \22512 );
or \U$24212 ( \24555 , \24553 , \24554 );
not \U$24213 ( \24556 , RI9872568_156);
not \U$24214 ( \24557 , \20580 );
or \U$24215 ( \24558 , \24556 , \24557 );
or \U$24216 ( \24559 , \10582 , RI9872568_156);
nand \U$24217 ( \24560 , \24558 , \24559 );
nand \U$24218 ( \24561 , \24560 , \5642 );
nand \U$24219 ( \24562 , \24555 , \24561 );
xor \U$24220 ( \24563 , \24552 , \24562 );
not \U$24221 ( \24564 , \24563 );
or \U$24222 ( \24565 , \24545 , \24564 );
nand \U$24223 ( \24566 , \24562 , \24552 );
nand \U$24224 ( \24567 , \24565 , \24566 );
not \U$24225 ( \24568 , \24567 );
or \U$24226 ( \24569 , \24535 , \24568 );
buf \U$24227 ( \24570 , \24497 );
nand \U$24228 ( \24571 , \24570 , \24532 );
nand \U$24229 ( \24572 , \24569 , \24571 );
not \U$24230 ( \24573 , \24572 );
or \U$24231 ( \24574 , \24420 , \24573 );
or \U$24232 ( \24575 , \24572 , \24419 );
nand \U$24233 ( \24576 , \24574 , \24575 );
not \U$24234 ( \24577 , \24576 );
or \U$24235 ( \24578 , \24418 , \24577 );
not \U$24236 ( \24579 , \24419 );
nand \U$24237 ( \24580 , \24579 , \24572 );
nand \U$24238 ( \24581 , \24578 , \24580 );
not \U$24239 ( \24582 , \24581 );
or \U$24240 ( \24583 , \24361 , \24582 );
or \U$24241 ( \24584 , \24581 , \24360 );
nand \U$24242 ( \24585 , \24583 , \24584 );
not \U$24243 ( \24586 , \24585 );
or \U$24244 ( \24587 , \24359 , \24586 );
not \U$24245 ( \24588 , \24360 );
nand \U$24246 ( \24589 , \24588 , \24581 );
nand \U$24247 ( \24590 , \24587 , \24589 );
not \U$24248 ( \24591 , \24590 );
nand \U$24249 ( \24592 , \24352 , \24591 );
not \U$24250 ( \24593 , \24592 );
nand \U$24251 ( \24594 , \24350 , \24172 , \24590 );
not \U$24252 ( \24595 , \24594 );
or \U$24253 ( \24596 , \24593 , \24595 );
not \U$24254 ( \24597 , \22868 );
not \U$24255 ( \24598 , \22581 );
and \U$24256 ( \24599 , \24597 , \24598 );
and \U$24257 ( \24600 , \22868 , \22581 );
nor \U$24258 ( \24601 , \24599 , \24600 );
not \U$24259 ( \24602 , \24601 );
nand \U$24260 ( \24603 , \24596 , \24602 );
not \U$24261 ( \24604 , \24172 );
not \U$24262 ( \24605 , \24350 );
or \U$24263 ( \24606 , \24604 , \24605 );
not \U$24264 ( \24607 , \24591 );
nand \U$24265 ( \24608 , \24606 , \24607 );
nand \U$24266 ( \24609 , \24603 , \24608 );
xor \U$24267 ( \24610 , \24138 , \24609 );
not \U$24268 ( \24611 , \24610 );
or \U$24269 ( \24612 , \24136 , \24611 );
not \U$24270 ( \24613 , \24608 );
not \U$24271 ( \24614 , \24603 );
or \U$24272 ( \24615 , \24613 , \24614 );
nand \U$24273 ( \24616 , \24615 , \24138 );
nand \U$24274 ( \24617 , \24612 , \24616 );
xor \U$24275 ( \24618 , \24050 , \24617 );
xor \U$24276 ( \24619 , \23881 , \23889 );
xnor \U$24277 ( \24620 , \24619 , \23885 );
and \U$24278 ( \24621 , \24320 , \24330 );
not \U$24279 ( \24622 , \24320 );
not \U$24280 ( \24623 , \24330 );
and \U$24281 ( \24624 , \24622 , \24623 );
nor \U$24282 ( \24625 , \24621 , \24624 );
not \U$24283 ( \24626 , \24625 );
buf \U$24284 ( \24627 , \8742 );
not \U$24285 ( \24628 , \24627 );
xor \U$24286 ( \24629 , \2110 , RI9872f40_177);
not \U$24287 ( \24630 , \24629 );
or \U$24288 ( \24631 , \24628 , \24630 );
nand \U$24289 ( \24632 , \24068 , \13214 );
nand \U$24290 ( \24633 , \24631 , \24632 );
not \U$24291 ( \24634 , \24633 );
not \U$24292 ( \24635 , \9273 );
not \U$24293 ( \24636 , \24328 );
or \U$24294 ( \24637 , \24635 , \24636 );
not \U$24295 ( \24638 , RI9872e50_175);
not \U$24296 ( \24639 , \3859 );
or \U$24297 ( \24640 , \24638 , \24639 );
or \U$24298 ( \24641 , \3859 , RI9872e50_175);
nand \U$24299 ( \24642 , \24640 , \24641 );
nand \U$24300 ( \24643 , \24642 , \18563 );
nand \U$24301 ( \24644 , \24637 , \24643 );
not \U$24302 ( \24645 , \24644 );
or \U$24303 ( \24646 , \24634 , \24645 );
or \U$24304 ( \24647 , \24644 , \24633 );
not \U$24305 ( \24648 , \17528 );
not \U$24306 ( \24649 , \24307 );
or \U$24307 ( \24650 , \24648 , \24649 );
and \U$24308 ( \24651 , RI9873288_184, \5720 );
not \U$24309 ( \24652 , RI9873288_184);
and \U$24310 ( \24653 , \24652 , \11559 );
or \U$24311 ( \24654 , \24651 , \24653 );
nand \U$24312 ( \24655 , \24654 , \17545 );
nand \U$24313 ( \24656 , \24650 , \24655 );
nand \U$24314 ( \24657 , \24647 , \24656 );
nand \U$24315 ( \24658 , \24646 , \24657 );
not \U$24316 ( \24659 , \24658 );
xor \U$24317 ( \24660 , \24544 , \24552 );
xnor \U$24318 ( \24661 , \24660 , \24562 );
not \U$24319 ( \24662 , \24661 );
or \U$24320 ( \24663 , \24659 , \24662 );
or \U$24321 ( \24664 , \24658 , \24661 );
nand \U$24322 ( \24665 , \24663 , \24664 );
not \U$24323 ( \24666 , \24665 );
or \U$24324 ( \24667 , \24626 , \24666 );
not \U$24325 ( \24668 , \24661 );
nand \U$24326 ( \24669 , \24668 , \24658 );
nand \U$24327 ( \24670 , \24667 , \24669 );
not \U$24328 ( \24671 , \24670 );
not \U$24329 ( \24672 , \24091 );
xor \U$24330 ( \24673 , \24532 , \24570 );
xnor \U$24331 ( \24674 , \24673 , \24567 );
xor \U$24332 ( \24675 , \24672 , \24674 );
xor \U$24333 ( \24676 , \23993 , \24059 );
and \U$24334 ( \24677 , \24005 , \23996 );
not \U$24335 ( \24678 , \24005 );
and \U$24336 ( \24679 , \24678 , \23983 );
or \U$24337 ( \24680 , \24677 , \24679 );
xnor \U$24338 ( \24681 , \24676 , \24680 );
xnor \U$24339 ( \24682 , \24675 , \24681 );
not \U$24340 ( \24683 , \24682 );
or \U$24341 ( \24684 , \24671 , \24683 );
xor \U$24342 ( \24685 , \23993 , \24672 );
not \U$24343 ( \24686 , \24059 );
not \U$24344 ( \24687 , \24680 );
or \U$24345 ( \24688 , \24686 , \24687 );
or \U$24346 ( \24689 , \24680 , \24059 );
nand \U$24347 ( \24690 , \24688 , \24689 );
xnor \U$24348 ( \24691 , \24685 , \24690 );
or \U$24349 ( \24692 , \24691 , \24674 );
nand \U$24350 ( \24693 , \24684 , \24692 );
not \U$24351 ( \24694 , \24693 );
not \U$24352 ( \24695 , \24417 );
not \U$24353 ( \24696 , \24695 );
buf \U$24354 ( \24697 , \24576 );
not \U$24355 ( \24698 , \24697 );
or \U$24356 ( \24699 , \24696 , \24698 );
or \U$24357 ( \24700 , \24697 , \24695 );
nand \U$24358 ( \24701 , \24699 , \24700 );
not \U$24359 ( \24702 , \24701 );
not \U$24360 ( \24703 , \24222 );
not \U$24361 ( \24704 , \24225 );
and \U$24362 ( \24705 , \24703 , \24704 );
and \U$24363 ( \24706 , \24222 , \24225 );
nor \U$24364 ( \24707 , \24705 , \24706 );
and \U$24365 ( \24708 , \24707 , \24344 );
not \U$24366 ( \24709 , \24707 );
not \U$24367 ( \24710 , \24344 );
and \U$24368 ( \24711 , \24709 , \24710 );
nor \U$24369 ( \24712 , \24708 , \24711 );
not \U$24370 ( \24713 , \24712 );
or \U$24371 ( \24714 , \24702 , \24713 );
or \U$24372 ( \24715 , \24712 , \24701 );
nand \U$24373 ( \24716 , \24714 , \24715 );
not \U$24374 ( \24717 , \24716 );
or \U$24375 ( \24718 , \24694 , \24717 );
not \U$24376 ( \24719 , \24712 );
nand \U$24377 ( \24720 , \24719 , \24701 );
nand \U$24378 ( \24721 , \24718 , \24720 );
not \U$24379 ( \24722 , \24721 );
not \U$24380 ( \24723 , \23968 );
xor \U$24381 ( \24724 , \23979 , \24723 );
xor \U$24382 ( \24725 , \23940 , \23958 );
not \U$24383 ( \24726 , \2072 );
and \U$24384 ( \24727 , RI9871aa0_133, \11370 );
not \U$24385 ( \24728 , RI9871aa0_133);
not \U$24386 ( \24729 , \18344 );
and \U$24387 ( \24730 , \24728 , \24729 );
nor \U$24388 ( \24731 , \24727 , \24730 );
not \U$24389 ( \24732 , \24731 );
or \U$24390 ( \24733 , \24726 , \24732 );
nand \U$24391 ( \24734 , \24391 , \2087 );
nand \U$24392 ( \24735 , \24733 , \24734 );
xor \U$24393 ( \24736 , \24725 , \24735 );
not \U$24394 ( \24737 , \791 );
not \U$24395 ( \24738 , RI98719b0_131);
not \U$24396 ( \24739 , \10064 );
or \U$24397 ( \24740 , \24738 , \24739 );
or \U$24398 ( \24741 , \17767 , RI98719b0_131);
nand \U$24399 ( \24742 , \24740 , \24741 );
not \U$24400 ( \24743 , \24742 );
or \U$24401 ( \24744 , \24737 , \24743 );
nand \U$24402 ( \24745 , \24506 , \6144 );
nand \U$24403 ( \24746 , \24744 , \24745 );
and \U$24404 ( \24747 , \24736 , \24746 );
and \U$24405 ( \24748 , \24725 , \24735 );
or \U$24406 ( \24749 , \24747 , \24748 );
not \U$24407 ( \24750 , \24749 );
xor \U$24408 ( \24751 , \24724 , \24750 );
not \U$24409 ( \24752 , \1455 );
not \U$24410 ( \24753 , RI9871c08_136);
not \U$24411 ( \24754 , \13623 );
not \U$24412 ( \24755 , \24754 );
or \U$24413 ( \24756 , \24753 , \24755 );
not \U$24414 ( \24757 , \18350 );
not \U$24415 ( \24758 , \24757 );
or \U$24416 ( \24759 , \24758 , RI9871c08_136);
nand \U$24417 ( \24760 , \24756 , \24759 );
not \U$24418 ( \24761 , \24760 );
or \U$24419 ( \24762 , \24752 , \24761 );
nand \U$24420 ( \24763 , \24525 , \1429 );
nand \U$24421 ( \24764 , \24762 , \24763 );
not \U$24422 ( \24765 , \1083 );
not \U$24423 ( \24766 , \1111 );
not \U$24424 ( \24767 , \12774 );
or \U$24425 ( \24768 , \24766 , \24767 );
nand \U$24426 ( \24769 , \12773 , RI98718c0_129);
nand \U$24427 ( \24770 , \24768 , \24769 );
not \U$24428 ( \24771 , \24770 );
or \U$24429 ( \24772 , \24765 , \24771 );
nand \U$24430 ( \24773 , \23977 , \1134 );
nand \U$24431 ( \24774 , \24772 , \24773 );
xor \U$24432 ( \24775 , \24764 , \24774 );
not \U$24433 ( \24776 , \5034 );
and \U$24434 ( \24777 , RI9872478_154, \8074 );
not \U$24435 ( \24778 , RI9872478_154);
not \U$24436 ( \24779 , \21518 );
and \U$24437 ( \24780 , \24778 , \24779 );
or \U$24438 ( \24781 , \24777 , \24780 );
not \U$24439 ( \24782 , \24781 );
or \U$24440 ( \24783 , \24776 , \24782 );
nand \U$24441 ( \24784 , \24488 , \5035 );
nand \U$24442 ( \24785 , \24783 , \24784 );
and \U$24443 ( \24786 , \24775 , \24785 );
and \U$24444 ( \24787 , \24764 , \24774 );
nor \U$24445 ( \24788 , \24786 , \24787 );
and \U$24446 ( \24789 , \24751 , \24788 );
and \U$24447 ( \24790 , \24724 , \24750 );
or \U$24448 ( \24791 , \24789 , \24790 );
not \U$24449 ( \24792 , \24791 );
and \U$24450 ( \24793 , \22650 , \22666 );
not \U$24451 ( \24794 , \22650 );
and \U$24452 ( \24795 , \24794 , \22667 );
nor \U$24453 ( \24796 , \24793 , \24795 );
xnor \U$24454 ( \24797 , \24796 , \22685 );
not \U$24455 ( \24798 , \24797 );
or \U$24456 ( \24799 , \24792 , \24798 );
xor \U$24457 ( \24800 , \24528 , \24510 );
not \U$24458 ( \24801 , \3169 );
not \U$24459 ( \24802 , \24380 );
or \U$24460 ( \24803 , \24801 , \24802 );
not \U$24461 ( \24804 , \3154 );
not \U$24462 ( \24805 , \9750 );
or \U$24463 ( \24806 , \24804 , \24805 );
not \U$24464 ( \24807 , \8694 );
not \U$24465 ( \24808 , \24807 );
or \U$24466 ( \24809 , \24808 , \3154 );
nand \U$24467 ( \24810 , \24806 , \24809 );
nand \U$24468 ( \24811 , \24810 , \3163 );
nand \U$24469 ( \24812 , \24803 , \24811 );
not \U$24470 ( \24813 , \5642 );
not \U$24471 ( \24814 , RI9872568_156);
not \U$24472 ( \24815 , \18128 );
or \U$24473 ( \24816 , \24814 , \24815 );
or \U$24474 ( \24817 , \8924 , RI9872568_156);
nand \U$24475 ( \24818 , \24816 , \24817 );
not \U$24476 ( \24819 , \24818 );
or \U$24477 ( \24820 , \24813 , \24819 );
nand \U$24478 ( \24821 , \24560 , \7188 );
nand \U$24479 ( \24822 , \24820 , \24821 );
xor \U$24480 ( \24823 , \24812 , \24822 );
not \U$24481 ( \24824 , \7333 );
not \U$24482 ( \24825 , \5703 );
or \U$24483 ( \24826 , \24824 , \24825 );
or \U$24484 ( \24827 , \18808 , \16892 );
nand \U$24485 ( \24828 , \24826 , \24827 );
not \U$24486 ( \24829 , \24828 );
not \U$24487 ( \24830 , \7325 );
or \U$24488 ( \24831 , \24829 , \24830 );
nand \U$24489 ( \24832 , \24244 , \7338 );
nand \U$24490 ( \24833 , \24831 , \24832 );
and \U$24491 ( \24834 , \24823 , \24833 );
and \U$24492 ( \24835 , \24812 , \24822 );
or \U$24493 ( \24836 , \24834 , \24835 );
xor \U$24494 ( \24837 , \24800 , \24836 );
not \U$24495 ( \24838 , \4919 );
not \U$24496 ( \24839 , RI9872388_152);
not \U$24497 ( \24840 , \18111 );
or \U$24498 ( \24841 , \24839 , \24840 );
buf \U$24499 ( \24842 , \18107 );
or \U$24500 ( \24843 , \24842 , RI9872388_152);
nand \U$24501 ( \24844 , \24841 , \24843 );
not \U$24502 ( \24845 , \24844 );
or \U$24503 ( \24846 , \24838 , \24845 );
nand \U$24504 ( \24847 , \24550 , \4925 );
nand \U$24505 ( \24848 , \24846 , \24847 );
not \U$24506 ( \24849 , \24848 );
xor \U$24507 ( \24850 , \24452 , \24463 );
not \U$24508 ( \24851 , \924 );
not \U$24509 ( \24852 , \23938 );
or \U$24510 ( \24853 , \24851 , \24852 );
buf \U$24511 ( \24854 , \17862 );
and \U$24512 ( \24855 , \24854 , RI9872130_147);
not \U$24513 ( \24856 , \24854 );
and \U$24514 ( \24857 , \24856 , \919 );
nor \U$24515 ( \24858 , \24855 , \24857 );
nand \U$24516 ( \24859 , \24858 , \875 );
nand \U$24517 ( \24860 , \24853 , \24859 );
xnor \U$24518 ( \24861 , \24850 , \24860 );
not \U$24519 ( \24862 , \1517 );
not \U$24520 ( \24863 , \24472 );
or \U$24521 ( \24864 , \24862 , \24863 );
and \U$24522 ( \24865 , RI9871c80_137, \18216 );
not \U$24523 ( \24866 , RI9871c80_137);
not \U$24524 ( \24867 , \16995 );
not \U$24525 ( \24868 , \24867 );
and \U$24526 ( \24869 , \24866 , \24868 );
or \U$24527 ( \24870 , \24865 , \24869 );
not \U$24528 ( \24871 , \24870 );
or \U$24529 ( \24872 , \24871 , \1499 );
nand \U$24530 ( \24873 , \24864 , \24872 );
nand \U$24531 ( \24874 , \24861 , \24873 );
xnor \U$24532 ( \24875 , \24452 , \24463 );
nand \U$24533 ( \24876 , \24860 , \24875 );
and \U$24534 ( \24877 , \24874 , \24876 );
not \U$24535 ( \24878 , \8790 );
and \U$24536 ( \24879 , \8650 , \6042 );
not \U$24537 ( \24880 , \8650 );
and \U$24538 ( \24881 , \24880 , RI98725e0_157);
nor \U$24539 ( \24882 , \24879 , \24881 );
not \U$24540 ( \24883 , \24882 );
or \U$24541 ( \24884 , \24878 , \24883 );
nand \U$24542 ( \24885 , \24542 , \5847 );
nand \U$24543 ( \24886 , \24884 , \24885 );
xnor \U$24544 ( \24887 , \24877 , \24886 );
not \U$24545 ( \24888 , \24887 );
or \U$24546 ( \24889 , \24849 , \24888 );
not \U$24547 ( \24890 , \24877 );
nand \U$24548 ( \24891 , \24890 , \24886 );
nand \U$24549 ( \24892 , \24889 , \24891 );
and \U$24550 ( \24893 , \24837 , \24892 );
and \U$24551 ( \24894 , \24800 , \24836 );
or \U$24552 ( \24895 , \24893 , \24894 );
nand \U$24553 ( \24896 , \24799 , \24895 );
or \U$24554 ( \24897 , \24797 , \24791 );
nand \U$24555 ( \24898 , \24896 , \24897 );
not \U$24556 ( \24899 , \24898 );
xor \U$24557 ( \24900 , \24010 , \24007 );
xnor \U$24558 ( \24901 , \24900 , \23917 );
nand \U$24559 ( \24902 , \24899 , \24901 );
not \U$24560 ( \24903 , \24902 );
xor \U$24561 ( \24904 , \24372 , \24398 );
not \U$24562 ( \24905 , \13020 );
not \U$24563 ( \24906 , RI98730a8_180);
not \U$24564 ( \24907 , \6330 );
or \U$24565 ( \24908 , \24906 , \24907 );
or \U$24566 ( \24909 , \9326 , RI98730a8_180);
nand \U$24567 ( \24910 , \24908 , \24909 );
not \U$24568 ( \24911 , \24910 );
or \U$24569 ( \24912 , \24905 , \24911 );
nand \U$24570 ( \24913 , \24208 , \17347 );
nand \U$24571 ( \24914 , \24912 , \24913 );
not \U$24572 ( \24915 , \24914 );
not \U$24573 ( \24916 , \13017 );
not \U$24574 ( \24917 , \24187 );
or \U$24575 ( \24918 , \24916 , \24917 );
not \U$24576 ( \24919 , \15389 );
not \U$24577 ( \24920 , \5393 );
or \U$24578 ( \24921 , \24919 , \24920 );
nand \U$24579 ( \24922 , \5775 , RI9872a18_166);
nand \U$24580 ( \24923 , \24921 , \24922 );
nand \U$24581 ( \24924 , \24923 , \8027 );
nand \U$24582 ( \24925 , \24918 , \24924 );
not \U$24583 ( \24926 , \24925 );
not \U$24584 ( \24927 , \24926 );
not \U$24585 ( \24928 , \9196 );
not \U$24586 ( \24929 , RI9872b80_169);
not \U$24587 ( \24930 , \23391 );
or \U$24588 ( \24931 , \24929 , \24930 );
or \U$24589 ( \24932 , \11548 , RI9872b80_169);
nand \U$24590 ( \24933 , \24931 , \24932 );
not \U$24591 ( \24934 , \24933 );
or \U$24592 ( \24935 , \24928 , \24934 );
nand \U$24593 ( \24936 , \24198 , \9214 );
nand \U$24594 ( \24937 , \24935 , \24936 );
not \U$24595 ( \24938 , \24937 );
or \U$24596 ( \24939 , \24927 , \24938 );
or \U$24597 ( \24940 , \24937 , \24926 );
nand \U$24598 ( \24941 , \24939 , \24940 );
not \U$24599 ( \24942 , \24941 );
or \U$24600 ( \24943 , \24915 , \24942 );
nand \U$24601 ( \24944 , \24937 , \24925 );
nand \U$24602 ( \24945 , \24943 , \24944 );
xor \U$24603 ( \24946 , \24904 , \24945 );
not \U$24604 ( \24947 , \13109 );
and \U$24605 ( \24948 , RI9873030_179, \5946 );
not \U$24606 ( \24949 , RI9873030_179);
and \U$24607 ( \24950 , \24949 , \11755 );
or \U$24608 ( \24951 , \24948 , \24950 );
not \U$24609 ( \24952 , \24951 );
or \U$24610 ( \24953 , \24947 , \24952 );
nand \U$24611 ( \24954 , \24255 , \9937 );
nand \U$24612 ( \24955 , \24953 , \24954 );
not \U$24613 ( \24956 , \24955 );
xor \U$24614 ( \24957 , \24480 , \24443 );
not \U$24615 ( \24958 , \24957 );
not \U$24616 ( \24959 , RI9873648_192);
not \U$24617 ( \24960 , \24285 );
or \U$24618 ( \24961 , \24959 , \24960 );
not \U$24619 ( \24962 , \18239 );
not \U$24620 ( \24963 , \1273 );
or \U$24621 ( \24964 , \24962 , \24963 );
or \U$24622 ( \24965 , \18239 , \1273 );
nand \U$24623 ( \24966 , \24964 , \24965 );
nand \U$24624 ( \24967 , \24966 , \18545 );
nand \U$24625 ( \24968 , \24961 , \24967 );
not \U$24626 ( \24969 , \24968 );
not \U$24627 ( \24970 , \24969 );
or \U$24628 ( \24971 , \24958 , \24970 );
or \U$24629 ( \24972 , \24969 , \24957 );
nand \U$24630 ( \24973 , \24971 , \24972 );
not \U$24631 ( \24974 , \24973 );
or \U$24632 ( \24975 , \24956 , \24974 );
nand \U$24633 ( \24976 , \24968 , \24957 );
nand \U$24634 ( \24977 , \24975 , \24976 );
and \U$24635 ( \24978 , \24946 , \24977 );
and \U$24636 ( \24979 , \24904 , \24945 );
or \U$24637 ( \24980 , \24978 , \24979 );
not \U$24638 ( \24981 , \24980 );
xor \U$24639 ( \24982 , \24409 , \24402 );
xnor \U$24640 ( \24983 , \24982 , \24415 );
not \U$24641 ( \24984 , \24983 );
nand \U$24642 ( \24985 , \24981 , \24984 );
not \U$24643 ( \24986 , \24985 );
not \U$24644 ( \24987 , \9312 );
not \U$24645 ( \24988 , \8807 );
not \U$24646 ( \24989 , \3569 );
or \U$24647 ( \24990 , \24988 , \24989 );
nand \U$24648 ( \24991 , \14930 , RI9872d60_173);
nand \U$24649 ( \24992 , \24990 , \24991 );
not \U$24650 ( \24993 , \24992 );
or \U$24651 ( \24994 , \24987 , \24993 );
nand \U$24652 ( \24995 , \24317 , \8802 );
nand \U$24653 ( \24996 , \24994 , \24995 );
not \U$24654 ( \24997 , \24996 );
not \U$24655 ( \24998 , \18957 );
xnor \U$24656 ( \24999 , RI9873210_183, \1366 );
not \U$24657 ( \25000 , \24999 );
or \U$24658 ( \25001 , \24998 , \25000 );
nand \U$24659 ( \25002 , \24275 , \17123 );
nand \U$24660 ( \25003 , \25001 , \25002 );
not \U$24661 ( \25004 , \9668 );
not \U$24662 ( \25005 , \24293 );
or \U$24663 ( \25006 , \25004 , \25005 );
not \U$24664 ( \25007 , \9185 );
not \U$24665 ( \25008 , \15685 );
or \U$24666 ( \25009 , \25007 , \25008 );
nand \U$24667 ( \25010 , \5205 , RI9872bf8_170);
nand \U$24668 ( \25011 , \25009 , \25010 );
nand \U$24669 ( \25012 , \25011 , \9670 );
nand \U$24670 ( \25013 , \25006 , \25012 );
xor \U$24671 ( \25014 , \25003 , \25013 );
not \U$24672 ( \25015 , \25014 );
or \U$24673 ( \25016 , \24997 , \25015 );
nand \U$24674 ( \25017 , \25013 , \25003 );
nand \U$24675 ( \25018 , \25016 , \25017 );
not \U$24676 ( \25019 , \25018 );
not \U$24677 ( \25020 , \5632 );
not \U$24678 ( \25021 , \7905 );
or \U$24679 ( \25022 , \25020 , \25021 );
nand \U$24680 ( \25023 , \18794 , RI98728b0_163);
nand \U$24681 ( \25024 , \25022 , \25023 );
nand \U$24682 ( \25025 , \25024 , \6284 );
buf \U$24683 ( \25026 , \24425 );
nand \U$24684 ( \25027 , \25026 , \6286 );
not \U$24685 ( \25028 , \3465 );
not \U$24686 ( \25029 , \3593 );
not \U$24687 ( \25030 , \10372 );
or \U$24688 ( \25031 , \25029 , \25030 );
nand \U$24689 ( \25032 , \8554 , RI98726d0_159);
nand \U$24690 ( \25033 , \25031 , \25032 );
not \U$24691 ( \25034 , \25033 );
or \U$24692 ( \25035 , \25028 , \25034 );
nand \U$24693 ( \25036 , \24370 , \3467 );
nand \U$24694 ( \25037 , \25035 , \25036 );
not \U$24695 ( \25038 , \25037 );
nand \U$24696 ( \25039 , \25025 , \25027 , \25038 );
not \U$24697 ( \25040 , \25039 );
not \U$24698 ( \25041 , \19036 );
and \U$24699 ( \25042 , RI98734e0_189, \891 );
not \U$24700 ( \25043 , RI98734e0_189);
and \U$24701 ( \25044 , \25043 , \6442 );
nor \U$24702 ( \25045 , \25042 , \25044 );
not \U$24703 ( \25046 , \25045 );
or \U$24704 ( \25047 , \25041 , \25046 );
nand \U$24705 ( \25048 , \24075 , \20147 );
nand \U$24706 ( \25049 , \25047 , \25048 );
not \U$24707 ( \25050 , \25049 );
or \U$24708 ( \25051 , \25040 , \25050 );
nand \U$24709 ( \25052 , \25027 , \25025 );
nand \U$24710 ( \25053 , \25052 , \25037 );
nand \U$24711 ( \25054 , \25051 , \25053 );
xor \U$24712 ( \25055 , \24493 , \24427 );
buf \U$24713 ( \25056 , \25055 );
and \U$24714 ( \25057 , \25054 , \25056 );
not \U$24715 ( \25058 , \25054 );
not \U$24716 ( \25059 , \25056 );
and \U$24717 ( \25060 , \25058 , \25059 );
nor \U$24718 ( \25061 , \25057 , \25060 );
not \U$24719 ( \25062 , \25061 );
or \U$24720 ( \25063 , \25019 , \25062 );
nand \U$24721 ( \25064 , \25054 , \25056 );
nand \U$24722 ( \25065 , \25063 , \25064 );
not \U$24723 ( \25066 , \25065 );
or \U$24724 ( \25067 , \24986 , \25066 );
nand \U$24725 ( \25068 , \24980 , \24983 );
nand \U$24726 ( \25069 , \25067 , \25068 );
not \U$24727 ( \25070 , \25069 );
or \U$24728 ( \25071 , \24903 , \25070 );
not \U$24729 ( \25072 , \24901 );
nand \U$24730 ( \25073 , \25072 , \24898 );
nand \U$24731 ( \25074 , \25071 , \25073 );
not \U$24732 ( \25075 , \25074 );
not \U$24733 ( \25076 , \25075 );
not \U$24734 ( \25077 , \24585 );
not \U$24735 ( \25078 , \24357 );
and \U$24736 ( \25079 , \25077 , \25078 );
and \U$24737 ( \25080 , \24585 , \24357 );
nor \U$24738 ( \25081 , \25079 , \25080 );
not \U$24739 ( \25082 , \25081 );
not \U$24740 ( \25083 , \25082 );
or \U$24741 ( \25084 , \25076 , \25083 );
nand \U$24742 ( \25085 , \25081 , \25074 );
nand \U$24743 ( \25086 , \25084 , \25085 );
not \U$24744 ( \25087 , \25086 );
or \U$24745 ( \25088 , \24722 , \25087 );
not \U$24746 ( \25089 , \25081 );
nand \U$24747 ( \25090 , \25089 , \25074 );
nand \U$24748 ( \25091 , \25088 , \25090 );
not \U$24749 ( \25092 , \25091 );
not \U$24750 ( \25093 , \25092 );
not \U$24751 ( \25094 , \25093 );
xor \U$24752 ( \25095 , \24590 , \24601 );
nand \U$24753 ( \25096 , \24350 , \24172 );
xnor \U$24754 ( \25097 , \25095 , \25096 );
not \U$24755 ( \25098 , \25097 );
or \U$24756 ( \25099 , \25094 , \25098 );
not \U$24757 ( \25100 , \25092 );
not \U$24758 ( \25101 , \25097 );
not \U$24759 ( \25102 , \25101 );
or \U$24760 ( \25103 , \25100 , \25102 );
not \U$24761 ( \25104 , \24052 );
not \U$24762 ( \25105 , \24130 );
not \U$24763 ( \25106 , \25105 );
or \U$24764 ( \25107 , \25104 , \25106 );
not \U$24765 ( \25108 , \24052 );
nand \U$24766 ( \25109 , \25108 , \24130 );
nand \U$24767 ( \25110 , \25107 , \25109 );
nand \U$24768 ( \25111 , \25103 , \25110 );
nand \U$24769 ( \25112 , \25099 , \25111 );
xor \U$24770 ( \25113 , \24620 , \25112 );
xor \U$24771 ( \25114 , \24135 , \24610 );
and \U$24772 ( \25115 , \25113 , \25114 );
and \U$24773 ( \25116 , \24620 , \25112 );
or \U$24774 ( \25117 , \25115 , \25116 );
nor \U$24775 ( \25118 , \24618 , \25117 );
not \U$24776 ( \25119 , \23822 );
not \U$24777 ( \25120 , \24038 );
and \U$24778 ( \25121 , \25119 , \25120 );
and \U$24779 ( \25122 , \24038 , \23822 );
nor \U$24780 ( \25123 , \25121 , \25122 );
not \U$24781 ( \25124 , \25123 );
not \U$24782 ( \25125 , \23831 );
or \U$24783 ( \25126 , \25124 , \25125 );
or \U$24784 ( \25127 , \25123 , \23831 );
nand \U$24785 ( \25128 , \25126 , \25127 );
xor \U$24786 ( \25129 , \24047 , \24049 );
and \U$24787 ( \25130 , \25129 , \24617 );
and \U$24788 ( \25131 , \24047 , \24049 );
or \U$24789 ( \25132 , \25130 , \25131 );
nor \U$24790 ( \25133 , \25128 , \25132 );
nor \U$24791 ( \25134 , \25118 , \25133 );
not \U$24792 ( \25135 , \25134 );
xor \U$24793 ( \25136 , \24620 , \25112 );
xor \U$24794 ( \25137 , \25136 , \25114 );
xor \U$24795 ( \25138 , \24140 , \24349 );
xnor \U$24796 ( \25139 , \25138 , \24174 );
not \U$24797 ( \25140 , \25139 );
nand \U$24798 ( \25141 , \24117 , \24122 );
and \U$24799 ( \25142 , \25141 , \24107 );
not \U$24800 ( \25143 , \25141 );
not \U$24801 ( \25144 , \24107 );
and \U$24802 ( \25145 , \25143 , \25144 );
nor \U$24803 ( \25146 , \25142 , \25145 );
nand \U$24804 ( \25147 , \25140 , \25146 );
not \U$24805 ( \25148 , \25147 );
xor \U$24806 ( \25149 , \24337 , \24266 );
not \U$24807 ( \25150 , \25149 );
xor \U$24808 ( \25151 , \24179 , \24216 );
xor \U$24809 ( \25152 , \25151 , \24219 );
not \U$24810 ( \25153 , \25152 );
not \U$24811 ( \25154 , \24237 );
not \U$24812 ( \25155 , \25154 );
not \U$24813 ( \25156 , \24261 );
or \U$24814 ( \25157 , \25155 , \25156 );
or \U$24815 ( \25158 , \25154 , \24261 );
nand \U$24816 ( \25159 , \25157 , \25158 );
not \U$24817 ( \25160 , \25159 );
and \U$24818 ( \25161 , \21779 , \832 );
not \U$24819 ( \25162 , \924 );
not \U$24820 ( \25163 , \24858 );
or \U$24821 ( \25164 , \25162 , \25163 );
not \U$24822 ( \25165 , RI9872130_147);
not \U$24823 ( \25166 , \18193 );
not \U$24824 ( \25167 , \25166 );
not \U$24825 ( \25168 , \25167 );
or \U$24826 ( \25169 , \25165 , \25168 );
or \U$24827 ( \25170 , \18194 , RI9872130_147);
nand \U$24828 ( \25171 , \25169 , \25170 );
nand \U$24829 ( \25172 , \25171 , \875 );
nand \U$24830 ( \25173 , \25164 , \25172 );
xor \U$24831 ( \25174 , \25161 , \25173 );
not \U$24832 ( \25175 , \1493 );
not \U$24833 ( \25176 , \24870 );
or \U$24834 ( \25177 , \25175 , \25176 );
not \U$24835 ( \25178 , \1584 );
not \U$24836 ( \25179 , \20490 );
not \U$24837 ( \25180 , \25179 );
or \U$24838 ( \25181 , \25178 , \25180 );
nand \U$24839 ( \25182 , \23934 , RI9871c80_137);
nand \U$24840 ( \25183 , \25181 , \25182 );
nand \U$24841 ( \25184 , \25183 , \1500 );
nand \U$24842 ( \25185 , \25177 , \25184 );
and \U$24843 ( \25186 , \25174 , \25185 );
and \U$24844 ( \25187 , \25161 , \25173 );
nor \U$24845 ( \25188 , \25186 , \25187 );
not \U$24846 ( \25189 , \25188 );
not \U$24847 ( \25190 , \1323 );
not \U$24848 ( \25191 , \24434 );
or \U$24849 ( \25192 , \25190 , \25191 );
and \U$24850 ( \25193 , RI9871b18_134, \17908 );
not \U$24851 ( \25194 , RI9871b18_134);
and \U$24852 ( \25195 , \25194 , \17912 );
or \U$24853 ( \25196 , \25193 , \25195 );
nand \U$24854 ( \25197 , \25196 , \1292 );
nand \U$24855 ( \25198 , \25192 , \25197 );
not \U$24856 ( \25199 , \25198 );
or \U$24857 ( \25200 , \25189 , \25199 );
or \U$24858 ( \25201 , \25198 , \25188 );
nand \U$24859 ( \25202 , \25200 , \25201 );
not \U$24860 ( \25203 , \25202 );
not \U$24861 ( \25204 , \6144 );
not \U$24862 ( \25205 , \24742 );
or \U$24863 ( \25206 , \25204 , \25205 );
and \U$24864 ( \25207 , \11455 , \1078 );
not \U$24865 ( \25208 , \11455 );
and \U$24866 ( \25209 , \25208 , RI98719b0_131);
nor \U$24867 ( \25210 , \25207 , \25209 );
nand \U$24868 ( \25211 , \25210 , \793 );
nand \U$24869 ( \25212 , \25206 , \25211 );
not \U$24870 ( \25213 , \25212 );
or \U$24871 ( \25214 , \25203 , \25213 );
not \U$24872 ( \25215 , \25188 );
nand \U$24873 ( \25216 , \25215 , \25198 );
nand \U$24874 ( \25217 , \25214 , \25216 );
not \U$24875 ( \25218 , \25217 );
not \U$24876 ( \25219 , \25218 );
not \U$24877 ( \25220 , \1429 );
not \U$24878 ( \25221 , \24760 );
or \U$24879 ( \25222 , \25220 , \25221 );
not \U$24880 ( \25223 , RI9871c08_136);
not \U$24881 ( \25224 , \13861 );
not \U$24882 ( \25225 , \25224 );
or \U$24883 ( \25226 , \25223 , \25225 );
or \U$24884 ( \25227 , \25224 , RI9871c08_136);
nand \U$24885 ( \25228 , \25226 , \25227 );
nand \U$24886 ( \25229 , \25228 , \1455 );
nand \U$24887 ( \25230 , \25222 , \25229 );
not \U$24888 ( \25231 , \2087 );
not \U$24889 ( \25232 , \24731 );
or \U$24890 ( \25233 , \25231 , \25232 );
xor \U$24891 ( \25234 , RI9871aa0_133, \20302 );
nand \U$24892 ( \25235 , \25234 , \2072 );
nand \U$24893 ( \25236 , \25233 , \25235 );
xor \U$24894 ( \25237 , \25230 , \25236 );
not \U$24895 ( \25238 , \1135 );
not \U$24896 ( \25239 , \24770 );
or \U$24897 ( \25240 , \25238 , \25239 );
and \U$24898 ( \25241 , \13281 , RI98718c0_129);
not \U$24899 ( \25242 , \13281 );
and \U$24900 ( \25243 , \25242 , \1111 );
nor \U$24901 ( \25244 , \25241 , \25243 );
nand \U$24902 ( \25245 , \25244 , \1083 );
nand \U$24903 ( \25246 , \25240 , \25245 );
and \U$24904 ( \25247 , \25237 , \25246 );
and \U$24905 ( \25248 , \25230 , \25236 );
or \U$24906 ( \25249 , \25247 , \25248 );
not \U$24907 ( \25250 , \25249 );
or \U$24908 ( \25251 , \25219 , \25250 );
or \U$24909 ( \25252 , \25249 , \25218 );
nand \U$24910 ( \25253 , \25251 , \25252 );
not \U$24911 ( \25254 , \25253 );
not \U$24912 ( \25255 , \17263 );
not \U$24913 ( \25256 , \24233 );
or \U$24914 ( \25257 , \25255 , \25256 );
not \U$24915 ( \25258 , RI98733f0_187);
not \U$24916 ( \25259 , \18737 );
or \U$24917 ( \25260 , \25258 , \25259 );
or \U$24918 ( \25261 , \18737 , RI98733f0_187);
nand \U$24919 ( \25262 , \25260 , \25261 );
nand \U$24920 ( \25263 , \25262 , \17371 );
nand \U$24921 ( \25264 , \25257 , \25263 );
not \U$24922 ( \25265 , \25264 );
or \U$24923 ( \25266 , \25254 , \25265 );
nand \U$24924 ( \25267 , \25249 , \25217 );
nand \U$24925 ( \25268 , \25266 , \25267 );
not \U$24926 ( \25269 , \25268 );
not \U$24927 ( \25270 , \24087 );
not \U$24928 ( \25271 , \24070 );
not \U$24929 ( \25272 , \25271 );
or \U$24930 ( \25273 , \25270 , \25272 );
nand \U$24931 ( \25274 , \24086 , \24070 );
nand \U$24932 ( \25275 , \25273 , \25274 );
not \U$24933 ( \25276 , \25275 );
not \U$24934 ( \25277 , \25276 );
or \U$24935 ( \25278 , \25269 , \25277 );
not \U$24936 ( \25279 , \25268 );
nand \U$24937 ( \25280 , \25279 , \25275 );
nand \U$24938 ( \25281 , \25278 , \25280 );
not \U$24939 ( \25282 , \25281 );
or \U$24940 ( \25283 , \25160 , \25282 );
nand \U$24941 ( \25284 , \25275 , \25268 );
nand \U$24942 ( \25285 , \25283 , \25284 );
not \U$24943 ( \25286 , \25285 );
not \U$24944 ( \25287 , \25286 );
or \U$24945 ( \25288 , \25153 , \25287 );
or \U$24946 ( \25289 , \25286 , \25152 );
nand \U$24947 ( \25290 , \25288 , \25289 );
not \U$24948 ( \25291 , \25290 );
or \U$24949 ( \25292 , \25150 , \25291 );
nand \U$24950 ( \25293 , \25285 , \25152 );
nand \U$24951 ( \25294 , \25292 , \25293 );
not \U$24952 ( \25295 , \25294 );
xor \U$24953 ( \25296 , \24142 , \24144 );
xor \U$24954 ( \25297 , \25296 , \24168 );
xor \U$24955 ( \25298 , \24055 , \25297 );
buf \U$24956 ( \25299 , \24102 );
xor \U$24957 ( \25300 , \25298 , \25299 );
not \U$24958 ( \25301 , \25300 );
or \U$24959 ( \25302 , \25295 , \25301 );
not \U$24960 ( \25303 , \25299 );
not \U$24961 ( \25304 , \24055 );
not \U$24962 ( \25305 , \25304 );
and \U$24963 ( \25306 , \25303 , \25305 );
and \U$24964 ( \25307 , \25299 , \25304 );
nor \U$24965 ( \25308 , \25306 , \25307 );
not \U$24966 ( \25309 , \25308 );
nand \U$24967 ( \25310 , \25309 , \25297 );
nand \U$24968 ( \25311 , \25302 , \25310 );
not \U$24969 ( \25312 , \25311 );
or \U$24970 ( \25313 , \25148 , \25312 );
not \U$24971 ( \25314 , \25146 );
nand \U$24972 ( \25315 , \25314 , \25139 );
nand \U$24973 ( \25316 , \25313 , \25315 );
xor \U$24974 ( \25317 , \25092 , \25097 );
xnor \U$24975 ( \25318 , \25317 , \25110 );
xor \U$24976 ( \25319 , \25316 , \25318 );
xnor \U$24977 ( \25320 , \24721 , \25086 );
nand \U$24978 ( \25321 , \25073 , \24902 );
xor \U$24979 ( \25322 , \25321 , \25069 );
xor \U$24980 ( \25323 , \24724 , \24750 );
xor \U$24981 ( \25324 , \25323 , \24788 );
not \U$24982 ( \25325 , \25324 );
and \U$24983 ( \25326 , \24212 , \24189 );
not \U$24984 ( \25327 , \24212 );
not \U$24985 ( \25328 , \24189 );
and \U$24986 ( \25329 , \25327 , \25328 );
nor \U$24987 ( \25330 , \25326 , \25329 );
not \U$24988 ( \25331 , \25330 );
not \U$24989 ( \25332 , \25331 );
or \U$24990 ( \25333 , \25325 , \25332 );
xor \U$24991 ( \25334 , \24277 , \24287 );
xor \U$24992 ( \25335 , \25334 , \24297 );
nand \U$24993 ( \25336 , \25333 , \25335 );
not \U$24994 ( \25337 , \25324 );
nand \U$24995 ( \25338 , \25337 , \25330 );
nand \U$24996 ( \25339 , \25336 , \25338 );
not \U$24997 ( \25340 , \25339 );
not \U$24998 ( \25341 , \4084 );
not \U$24999 ( \25342 , \24882 );
or \U$25000 ( \25343 , \25341 , \25342 );
not \U$25001 ( \25344 , RI98725e0_157);
not \U$25002 ( \25345 , \8579 );
or \U$25003 ( \25346 , \25344 , \25345 );
not \U$25004 ( \25347 , \8842 );
nand \U$25005 ( \25348 , \25347 , \4092 );
nand \U$25006 ( \25349 , \25346 , \25348 );
nand \U$25007 ( \25350 , \25349 , \18171 );
nand \U$25008 ( \25351 , \25343 , \25350 );
not \U$25009 ( \25352 , \25351 );
not \U$25010 ( \25353 , \12514 );
not \U$25011 ( \25354 , \24810 );
or \U$25012 ( \25355 , \25353 , \25354 );
and \U$25013 ( \25356 , \3154 , \9849 );
not \U$25014 ( \25357 , \3154 );
and \U$25015 ( \25358 , \25357 , \8707 );
nor \U$25016 ( \25359 , \25356 , \25358 );
nand \U$25017 ( \25360 , \25359 , \3163 );
nand \U$25018 ( \25361 , \25355 , \25360 );
not \U$25019 ( \25362 , \25361 );
and \U$25020 ( \25363 , \7338 , \24828 );
and \U$25021 ( \25364 , RI98729a0_165, \22516 );
not \U$25022 ( \25365 , RI98729a0_165);
and \U$25023 ( \25366 , \25365 , \8903 );
nor \U$25024 ( \25367 , \25364 , \25366 );
and \U$25025 ( \25368 , \25367 , \7326 );
nor \U$25026 ( \25369 , \25363 , \25368 );
not \U$25027 ( \25370 , \25369 );
or \U$25028 ( \25371 , \25362 , \25370 );
or \U$25029 ( \25372 , \25369 , \25361 );
nand \U$25030 ( \25373 , \25371 , \25372 );
not \U$25031 ( \25374 , \25373 );
or \U$25032 ( \25375 , \25352 , \25374 );
not \U$25033 ( \25376 , \25369 );
nand \U$25034 ( \25377 , \25376 , \25361 );
nand \U$25035 ( \25378 , \25375 , \25377 );
not \U$25036 ( \25379 , \1455 );
buf \U$25037 ( \25380 , \13932 );
and \U$25038 ( \25381 , \25380 , \3487 );
not \U$25039 ( \25382 , \25380 );
and \U$25040 ( \25383 , \25382 , RI9871c08_136);
nor \U$25041 ( \25384 , \25381 , \25383 );
not \U$25042 ( \25385 , \25384 );
or \U$25043 ( \25386 , \25379 , \25385 );
nand \U$25044 ( \25387 , \25228 , \1428 );
nand \U$25045 ( \25388 , \25386 , \25387 );
not \U$25046 ( \25389 , \25388 );
not \U$25047 ( \25390 , \25171 );
or \U$25048 ( \25391 , \25390 , \1470 );
and \U$25049 ( \25392 , RI9872130_147, \21778 );
not \U$25050 ( \25393 , RI9872130_147);
not \U$25051 ( \25394 , \22278 );
and \U$25052 ( \25395 , \25393 , \25394 );
nor \U$25053 ( \25396 , \25392 , \25395 );
or \U$25054 ( \25397 , \25396 , \874 );
nand \U$25055 ( \25398 , \25391 , \25397 );
not \U$25056 ( \25399 , \25398 );
or \U$25057 ( \25400 , \1800 , \866 );
or \U$25058 ( \25401 , RI9871c80_137, RI98721a8_148);
nand \U$25059 ( \25402 , \25401 , \24450 );
nand \U$25060 ( \25403 , \25400 , \25402 , RI9872130_147);
nor \U$25061 ( \25404 , \25399 , \25403 );
not \U$25062 ( \25405 , \1290 );
not \U$25063 ( \25406 , \25196 );
or \U$25064 ( \25407 , \25405 , \25406 );
not \U$25065 ( \25408 , \1283 );
not \U$25066 ( \25409 , \17868 );
not \U$25067 ( \25410 , \25409 );
or \U$25068 ( \25411 , \25408 , \25410 );
not \U$25069 ( \25412 , \17725 );
nand \U$25070 ( \25413 , \25412 , RI9871b18_134);
nand \U$25071 ( \25414 , \25411 , \25413 );
nand \U$25072 ( \25415 , \25414 , \1291 );
nand \U$25073 ( \25416 , \25407 , \25415 );
xor \U$25074 ( \25417 , \25404 , \25416 );
not \U$25075 ( \25418 , \25417 );
or \U$25076 ( \25419 , \25389 , \25418 );
nand \U$25077 ( \25420 , \25416 , \25404 );
nand \U$25078 ( \25421 , \25419 , \25420 );
not \U$25079 ( \25422 , \5035 );
not \U$25080 ( \25423 , \24781 );
or \U$25081 ( \25424 , \25422 , \25423 );
not \U$25082 ( \25425 , RI9872478_154);
not \U$25083 ( \25426 , \12716 );
or \U$25084 ( \25427 , \25425 , \25426 );
nand \U$25085 ( \25428 , \16945 , \5025 );
nand \U$25086 ( \25429 , \25427 , \25428 );
nand \U$25087 ( \25430 , \25429 , \5034 );
nand \U$25088 ( \25431 , \25424 , \25430 );
xor \U$25089 ( \25432 , \25421 , \25431 );
not \U$25090 ( \25433 , \4923 );
not \U$25091 ( \25434 , \24844 );
or \U$25092 ( \25435 , \25433 , \25434 );
not \U$25093 ( \25436 , RI9872388_152);
not \U$25094 ( \25437 , \8857 );
or \U$25095 ( \25438 , \25436 , \25437 );
nand \U$25096 ( \25439 , \9881 , \4902 );
nand \U$25097 ( \25440 , \25438 , \25439 );
nand \U$25098 ( \25441 , \25440 , \4919 );
nand \U$25099 ( \25442 , \25435 , \25441 );
and \U$25100 ( \25443 , \25432 , \25442 );
and \U$25101 ( \25444 , \25421 , \25431 );
or \U$25102 ( \25445 , \25443 , \25444 );
or \U$25103 ( \25446 , \25378 , \25445 );
not \U$25104 ( \25447 , \3467 );
not \U$25105 ( \25448 , \25033 );
or \U$25106 ( \25449 , \25447 , \25448 );
and \U$25107 ( \25450 , RI98726d0_159, \20385 );
not \U$25108 ( \25451 , RI98726d0_159);
and \U$25109 ( \25452 , \25451 , \12470 );
or \U$25110 ( \25453 , \25450 , \25452 );
nand \U$25111 ( \25454 , \25453 , \13409 );
nand \U$25112 ( \25455 , \25449 , \25454 );
not \U$25113 ( \25456 , \25455 );
not \U$25114 ( \25457 , \6286 );
not \U$25115 ( \25458 , \25024 );
or \U$25116 ( \25459 , \25457 , \25458 );
not \U$25117 ( \25460 , \5632 );
not \U$25118 ( \25461 , \7003 );
or \U$25119 ( \25462 , \25460 , \25461 );
nand \U$25120 ( \25463 , \10583 , RI98728b0_163);
nand \U$25121 ( \25464 , \25462 , \25463 );
nand \U$25122 ( \25465 , \25464 , \6284 );
nand \U$25123 ( \25466 , \25459 , \25465 );
not \U$25124 ( \25467 , \7188 );
not \U$25125 ( \25468 , \24818 );
or \U$25126 ( \25469 , \25467 , \25468 );
not \U$25127 ( \25470 , \5648 );
not \U$25128 ( \25471 , \12727 );
or \U$25129 ( \25472 , \25470 , \25471 );
nand \U$25130 ( \25473 , RI9872568_156, \8334 );
nand \U$25131 ( \25474 , \25472 , \25473 );
nand \U$25132 ( \25475 , \25474 , \9320 );
nand \U$25133 ( \25476 , \25469 , \25475 );
and \U$25134 ( \25477 , \25466 , \25476 );
not \U$25135 ( \25478 , \25466 );
not \U$25136 ( \25479 , \25476 );
and \U$25137 ( \25480 , \25478 , \25479 );
nor \U$25138 ( \25481 , \25477 , \25480 );
not \U$25139 ( \25482 , \25481 );
or \U$25140 ( \25483 , \25456 , \25482 );
nand \U$25141 ( \25484 , \25466 , \25476 );
nand \U$25142 ( \25485 , \25483 , \25484 );
nand \U$25143 ( \25486 , \25446 , \25485 );
nand \U$25144 ( \25487 , \25378 , \25445 );
nand \U$25145 ( \25488 , \25486 , \25487 );
xor \U$25146 ( \25489 , \24800 , \24836 );
xor \U$25147 ( \25490 , \25489 , \24892 );
nor \U$25148 ( \25491 , \25488 , \25490 );
xor \U$25149 ( \25492 , \24812 , \24822 );
xor \U$25150 ( \25493 , \25492 , \24833 );
xor \U$25151 ( \25494 , \24877 , \24886 );
xnor \U$25152 ( \25495 , \25494 , \24848 );
xor \U$25153 ( \25496 , \25493 , \25495 );
not \U$25154 ( \25497 , \10333 );
not \U$25155 ( \25498 , \24642 );
or \U$25156 ( \25499 , \25497 , \25498 );
not \U$25157 ( \25500 , \9690 );
not \U$25158 ( \25501 , \3537 );
or \U$25159 ( \25502 , \25500 , \25501 );
or \U$25160 ( \25503 , \18685 , \9694 );
nand \U$25161 ( \25504 , \25502 , \25503 );
nand \U$25162 ( \25505 , \25504 , \9686 );
nand \U$25163 ( \25506 , \25499 , \25505 );
not \U$25164 ( \25507 , \25506 );
not \U$25165 ( \25508 , \10251 );
not \U$25166 ( \25509 , RI9872d60_173);
not \U$25167 ( \25510 , \4176 );
or \U$25168 ( \25511 , \25509 , \25510 );
or \U$25169 ( \25512 , \4176 , RI9872d60_173);
nand \U$25170 ( \25513 , \25511 , \25512 );
not \U$25171 ( \25514 , \25513 );
or \U$25172 ( \25515 , \25508 , \25514 );
nand \U$25173 ( \25516 , \24992 , \10624 );
nand \U$25174 ( \25517 , \25515 , \25516 );
not \U$25175 ( \25518 , \25517 );
or \U$25176 ( \25519 , \25507 , \25518 );
or \U$25177 ( \25520 , \25506 , \25517 );
not \U$25178 ( \25521 , \17528 );
not \U$25179 ( \25522 , \24654 );
or \U$25180 ( \25523 , \25521 , \25522 );
not \U$25181 ( \25524 , RI9873288_184);
not \U$25182 ( \25525 , \1344 );
or \U$25183 ( \25526 , \25524 , \25525 );
nand \U$25184 ( \25527 , \5712 , \22727 );
nand \U$25185 ( \25528 , \25526 , \25527 );
nand \U$25186 ( \25529 , \25528 , \17545 );
nand \U$25187 ( \25530 , \25523 , \25529 );
nand \U$25188 ( \25531 , \25520 , \25530 );
nand \U$25189 ( \25532 , \25519 , \25531 );
and \U$25190 ( \25533 , \25496 , \25532 );
and \U$25191 ( \25534 , \25493 , \25495 );
nor \U$25192 ( \25535 , \25533 , \25534 );
or \U$25193 ( \25536 , \25491 , \25535 );
nand \U$25194 ( \25537 , \25488 , \25490 );
nand \U$25195 ( \25538 , \25536 , \25537 );
not \U$25196 ( \25539 , \25538 );
or \U$25197 ( \25540 , \25340 , \25539 );
not \U$25198 ( \25541 , \25339 );
not \U$25199 ( \25542 , \25541 );
not \U$25200 ( \25543 , \25538 );
not \U$25201 ( \25544 , \25543 );
or \U$25202 ( \25545 , \25542 , \25544 );
xor \U$25203 ( \25546 , \24154 , \24166 );
xnor \U$25204 ( \25547 , \25546 , \24147 );
nand \U$25205 ( \25548 , \25545 , \25547 );
nand \U$25206 ( \25549 , \25540 , \25548 );
not \U$25207 ( \25550 , \25549 );
nand \U$25208 ( \25551 , \25322 , \25550 );
not \U$25209 ( \25552 , \25551 );
xor \U$25210 ( \25553 , \24983 , \24981 );
buf \U$25211 ( \25554 , \25065 );
xnor \U$25212 ( \25555 , \25553 , \25554 );
not \U$25213 ( \25556 , \24791 );
not \U$25214 ( \25557 , \24797 );
or \U$25215 ( \25558 , \25556 , \25557 );
nand \U$25216 ( \25559 , \25558 , \24897 );
xnor \U$25217 ( \25560 , \25559 , \24895 );
buf \U$25218 ( \25561 , \25560 );
or \U$25219 ( \25562 , \25555 , \25561 );
xor \U$25220 ( \25563 , \24764 , \24774 );
xor \U$25221 ( \25564 , \25563 , \24785 );
not \U$25222 ( \25565 , \25564 );
xor \U$25223 ( \25566 , \24725 , \24735 );
xor \U$25224 ( \25567 , \25566 , \24746 );
not \U$25225 ( \25568 , \25567 );
nand \U$25226 ( \25569 , \25565 , \25568 );
not \U$25227 ( \25570 , \25569 );
not \U$25228 ( \25571 , \8752 );
not \U$25229 ( \25572 , \24629 );
or \U$25230 ( \25573 , \25571 , \25572 );
and \U$25231 ( \25574 , RI9872f40_177, \5884 );
not \U$25232 ( \25575 , RI9872f40_177);
and \U$25233 ( \25576 , \25575 , \2947 );
nor \U$25234 ( \25577 , \25574 , \25576 );
nand \U$25235 ( \25578 , \25577 , \9527 );
nand \U$25236 ( \25579 , \25573 , \25578 );
not \U$25237 ( \25580 , \25579 );
xor \U$25238 ( \25581 , \24875 , \24860 );
xnor \U$25239 ( \25582 , \25581 , \24873 );
not \U$25240 ( \25583 , \20147 );
not \U$25241 ( \25584 , \25045 );
or \U$25242 ( \25585 , \25583 , \25584 );
and \U$25243 ( \25586 , RI98734e0_189, \6219 );
not \U$25244 ( \25587 , RI98734e0_189);
and \U$25245 ( \25588 , \25587 , \820 );
nor \U$25246 ( \25589 , \25586 , \25588 );
nand \U$25247 ( \25590 , \25589 , \19243 );
nand \U$25248 ( \25591 , \25585 , \25590 );
xnor \U$25249 ( \25592 , \25582 , \25591 );
not \U$25250 ( \25593 , \25592 );
or \U$25251 ( \25594 , \25580 , \25593 );
not \U$25252 ( \25595 , \25582 );
nand \U$25253 ( \25596 , \25595 , \25591 );
nand \U$25254 ( \25597 , \25594 , \25596 );
not \U$25255 ( \25598 , \25597 );
or \U$25256 ( \25599 , \25570 , \25598 );
nand \U$25257 ( \25600 , \25567 , \25564 );
nand \U$25258 ( \25601 , \25599 , \25600 );
not \U$25259 ( \25602 , \25601 );
not \U$25260 ( \25603 , \9214 );
not \U$25261 ( \25604 , \24933 );
or \U$25262 ( \25605 , \25603 , \25604 );
not \U$25263 ( \25606 , RI9872b80_169);
not \U$25264 ( \25607 , \10873 );
or \U$25265 ( \25608 , \25606 , \25607 );
or \U$25266 ( \25609 , \5736 , RI9872b80_169);
nand \U$25267 ( \25610 , \25608 , \25609 );
nand \U$25268 ( \25611 , \25610 , \9196 );
nand \U$25269 ( \25612 , \25605 , \25611 );
not \U$25270 ( \25613 , \9668 );
not \U$25271 ( \25614 , \25011 );
or \U$25272 ( \25615 , \25613 , \25614 );
not \U$25273 ( \25616 , RI9872bf8_170);
not \U$25274 ( \25617 , \4471 );
or \U$25275 ( \25618 , \25616 , \25617 );
or \U$25276 ( \25619 , \12971 , RI9872bf8_170);
nand \U$25277 ( \25620 , \25618 , \25619 );
nand \U$25278 ( \25621 , \25620 , \9670 );
nand \U$25279 ( \25622 , \25615 , \25621 );
or \U$25280 ( \25623 , \25612 , \25622 );
not \U$25281 ( \25624 , \17234 );
not \U$25282 ( \25625 , \24999 );
or \U$25283 ( \25626 , \25624 , \25625 );
xor \U$25284 ( \25627 , RI9873210_183, \1713 );
nand \U$25285 ( \25628 , \25627 , \17243 );
nand \U$25286 ( \25629 , \25626 , \25628 );
nand \U$25287 ( \25630 , \25623 , \25629 );
nand \U$25288 ( \25631 , \25622 , \25612 );
nand \U$25289 ( \25632 , \25630 , \25631 );
not \U$25290 ( \25633 , \24923 );
or \U$25291 ( \25634 , \25633 , \8040 );
and \U$25292 ( \25635 , RI9872a18_166, \5763 );
not \U$25293 ( \25636 , RI9872a18_166);
and \U$25294 ( \25637 , \25636 , \6060 );
nor \U$25295 ( \25638 , \25635 , \25637 );
not \U$25296 ( \25639 , \8028 );
or \U$25297 ( \25640 , \25638 , \25639 );
nand \U$25298 ( \25641 , \25634 , \25640 );
not \U$25299 ( \25642 , \25641 );
not \U$25300 ( \25643 , \12868 );
not \U$25301 ( \25644 , \24910 );
or \U$25302 ( \25645 , \25643 , \25644 );
and \U$25303 ( \25646 , RI98730a8_180, \12393 );
not \U$25304 ( \25647 , RI98730a8_180);
and \U$25305 ( \25648 , \25647 , \6020 );
or \U$25306 ( \25649 , \25646 , \25648 );
nand \U$25307 ( \25650 , \25649 , \13020 );
nand \U$25308 ( \25651 , \25645 , \25650 );
buf \U$25309 ( \25652 , \25651 );
not \U$25310 ( \25653 , \25652 );
or \U$25311 ( \25654 , \25642 , \25653 );
or \U$25312 ( \25655 , \25651 , \25641 );
not \U$25313 ( \25656 , \9937 );
not \U$25314 ( \25657 , \24951 );
or \U$25315 ( \25658 , \25656 , \25657 );
and \U$25316 ( \25659 , \1486 , RI9873030_179);
not \U$25317 ( \25660 , \1486 );
and \U$25318 ( \25661 , \25660 , \14132 );
nor \U$25319 ( \25662 , \25659 , \25661 );
nand \U$25320 ( \25663 , \25662 , \13109 );
nand \U$25321 ( \25664 , \25658 , \25663 );
nand \U$25322 ( \25665 , \25655 , \25664 );
nand \U$25323 ( \25666 , \25654 , \25665 );
xor \U$25324 ( \25667 , \25632 , \25666 );
not \U$25325 ( \25668 , \25038 );
not \U$25326 ( \25669 , \25052 );
or \U$25327 ( \25670 , \25668 , \25669 );
or \U$25328 ( \25671 , \25052 , \25038 );
nand \U$25329 ( \25672 , \25670 , \25671 );
xor \U$25330 ( \25673 , \25049 , \25672 );
and \U$25331 ( \25674 , \25667 , \25673 );
and \U$25332 ( \25675 , \25632 , \25666 );
or \U$25333 ( \25676 , \25674 , \25675 );
not \U$25334 ( \25677 , \25676 );
nand \U$25335 ( \25678 , \25602 , \25677 );
not \U$25336 ( \25679 , \25678 );
and \U$25337 ( \25680 , \24665 , \24625 );
not \U$25338 ( \25681 , \24665 );
not \U$25339 ( \25682 , \24625 );
and \U$25340 ( \25683 , \25681 , \25682 );
nor \U$25341 ( \25684 , \25680 , \25683 );
not \U$25342 ( \25685 , \25684 );
or \U$25343 ( \25686 , \25679 , \25685 );
buf \U$25344 ( \25687 , \25601 );
nand \U$25345 ( \25688 , \25687 , \25676 );
nand \U$25346 ( \25689 , \25686 , \25688 );
nand \U$25347 ( \25690 , \25562 , \25689 );
nand \U$25348 ( \25691 , \25555 , \25561 );
nand \U$25349 ( \25692 , \25690 , \25691 );
not \U$25350 ( \25693 , \25692 );
or \U$25351 ( \25694 , \25552 , \25693 );
or \U$25352 ( \25695 , \25322 , \25550 );
nand \U$25353 ( \25696 , \25694 , \25695 );
not \U$25354 ( \25697 , \25696 );
and \U$25355 ( \25698 , \25320 , \25697 );
not \U$25356 ( \25699 , \25320 );
and \U$25357 ( \25700 , \25699 , \25696 );
nor \U$25358 ( \25701 , \25698 , \25700 );
not \U$25359 ( \25702 , \25701 );
not \U$25360 ( \25703 , \24716 );
not \U$25361 ( \25704 , \25703 );
not \U$25362 ( \25705 , \24693 );
and \U$25363 ( \25706 , \25704 , \25705 );
and \U$25364 ( \25707 , \25703 , \24693 );
nor \U$25365 ( \25708 , \25706 , \25707 );
not \U$25366 ( \25709 , \25708 );
and \U$25367 ( \25710 , \25324 , \25330 );
not \U$25368 ( \25711 , \25324 );
and \U$25369 ( \25712 , \25711 , \25331 );
or \U$25370 ( \25713 , \25710 , \25712 );
and \U$25371 ( \25714 , \25713 , \25335 );
not \U$25372 ( \25715 , \25713 );
not \U$25373 ( \25716 , \25335 );
and \U$25374 ( \25717 , \25715 , \25716 );
nor \U$25375 ( \25718 , \25714 , \25717 );
not \U$25376 ( \25719 , \25718 );
not \U$25377 ( \25720 , \3163 );
not \U$25378 ( \25721 , \9113 );
xor \U$25379 ( \25722 , RI9872310_151, \25721 );
not \U$25380 ( \25723 , \25722 );
or \U$25381 ( \25724 , \25720 , \25723 );
nand \U$25382 ( \25725 , \25359 , \3169 );
nand \U$25383 ( \25726 , \25724 , \25725 );
not \U$25384 ( \25727 , \25726 );
not \U$25385 ( \25728 , \1083 );
and \U$25386 ( \25729 , \20787 , \1111 );
not \U$25387 ( \25730 , \20787 );
and \U$25388 ( \25731 , \25730 , RI98718c0_129);
nor \U$25389 ( \25732 , \25729 , \25731 );
not \U$25390 ( \25733 , \25732 );
or \U$25391 ( \25734 , \25728 , \25733 );
nand \U$25392 ( \25735 , \25244 , \1134 );
nand \U$25393 ( \25736 , \25734 , \25735 );
not \U$25394 ( \25737 , \25736 );
nand \U$25395 ( \25738 , \25727 , \25737 );
not \U$25396 ( \25739 , \25738 );
not \U$25397 ( \25740 , \5035 );
not \U$25398 ( \25741 , \25429 );
or \U$25399 ( \25742 , \25740 , \25741 );
not \U$25400 ( \25743 , \5025 );
not \U$25401 ( \25744 , \8597 );
or \U$25402 ( \25745 , \25743 , \25744 );
or \U$25403 ( \25746 , \8597 , \5025 );
nand \U$25404 ( \25747 , \25745 , \25746 );
nand \U$25405 ( \25748 , \25747 , \5034 );
nand \U$25406 ( \25749 , \25742 , \25748 );
not \U$25407 ( \25750 , \25749 );
or \U$25408 ( \25751 , \25739 , \25750 );
nand \U$25409 ( \25752 , \25726 , \25736 );
nand \U$25410 ( \25753 , \25751 , \25752 );
xor \U$25411 ( \25754 , \25212 , \25202 );
xor \U$25412 ( \25755 , \25753 , \25754 );
not \U$25413 ( \25756 , \25755 );
not \U$25414 ( \25757 , \18171 );
and \U$25415 ( \25758 , RI98725e0_157, \8555 );
not \U$25416 ( \25759 , RI98725e0_157);
and \U$25417 ( \25760 , \25759 , \10372 );
or \U$25418 ( \25761 , \25758 , \25760 );
not \U$25419 ( \25762 , \25761 );
or \U$25420 ( \25763 , \25757 , \25762 );
nand \U$25421 ( \25764 , \25349 , \17098 );
nand \U$25422 ( \25765 , \25763 , \25764 );
not \U$25423 ( \25766 , \25765 );
not \U$25424 ( \25767 , \3464 );
and \U$25425 ( \25768 , \9750 , RI98726d0_159);
not \U$25426 ( \25769 , \9750 );
and \U$25427 ( \25770 , \25769 , \3593 );
nor \U$25428 ( \25771 , \25768 , \25770 );
not \U$25429 ( \25772 , \25771 );
or \U$25430 ( \25773 , \25767 , \25772 );
nand \U$25431 ( \25774 , \25453 , \3467 );
nand \U$25432 ( \25775 , \25773 , \25774 );
not \U$25433 ( \25776 , \4923 );
not \U$25434 ( \25777 , \25440 );
or \U$25435 ( \25778 , \25776 , \25777 );
and \U$25436 ( \25779 , RI9872388_152, \8640 );
not \U$25437 ( \25780 , RI9872388_152);
and \U$25438 ( \25781 , \25780 , \8650 );
nor \U$25439 ( \25782 , \25779 , \25781 );
nand \U$25440 ( \25783 , \25782 , \4919 );
nand \U$25441 ( \25784 , \25778 , \25783 );
xor \U$25442 ( \25785 , \25775 , \25784 );
not \U$25443 ( \25786 , \25785 );
or \U$25444 ( \25787 , \25766 , \25786 );
nand \U$25445 ( \25788 , \25784 , \25775 );
nand \U$25446 ( \25789 , \25787 , \25788 );
not \U$25447 ( \25790 , \25789 );
or \U$25448 ( \25791 , \25756 , \25790 );
nand \U$25449 ( \25792 , \25753 , \25754 );
nand \U$25450 ( \25793 , \25791 , \25792 );
not \U$25451 ( \25794 , \25793 );
xnor \U$25452 ( \25795 , \24941 , \24914 );
xor \U$25453 ( \25796 , \24996 , \25003 );
xor \U$25454 ( \25797 , \25796 , \25013 );
xnor \U$25455 ( \25798 , \25795 , \25797 );
not \U$25456 ( \25799 , \25798 );
or \U$25457 ( \25800 , \25794 , \25799 );
not \U$25458 ( \25801 , \25795 );
nand \U$25459 ( \25802 , \25801 , \25797 );
nand \U$25460 ( \25803 , \25800 , \25802 );
not \U$25461 ( \25804 , \25803 );
not \U$25462 ( \25805 , \25159 );
and \U$25463 ( \25806 , \25281 , \25805 );
not \U$25464 ( \25807 , \25281 );
and \U$25465 ( \25808 , \25807 , \25159 );
nor \U$25466 ( \25809 , \25806 , \25808 );
and \U$25467 ( \25810 , \25804 , \25809 );
not \U$25468 ( \25811 , \25804 );
not \U$25469 ( \25812 , \25809 );
and \U$25470 ( \25813 , \25811 , \25812 );
nor \U$25471 ( \25814 , \25810 , \25813 );
not \U$25472 ( \25815 , \25814 );
or \U$25473 ( \25816 , \25719 , \25815 );
nand \U$25474 ( \25817 , \25803 , \25812 );
nand \U$25475 ( \25818 , \25816 , \25817 );
not \U$25476 ( \25819 , \25818 );
xor \U$25477 ( \25820 , \25055 , \25054 );
xor \U$25478 ( \25821 , \25820 , \25018 );
xor \U$25479 ( \25822 , \24904 , \24945 );
xor \U$25480 ( \25823 , \25822 , \24977 );
nor \U$25481 ( \25824 , \25821 , \25823 );
xor \U$25482 ( \25825 , \24644 , \24633 );
xor \U$25483 ( \25826 , \25825 , \24656 );
not \U$25484 ( \25827 , \25826 );
not \U$25485 ( \25828 , \19282 );
not \U$25486 ( \25829 , \25262 );
or \U$25487 ( \25830 , \25828 , \25829 );
not \U$25488 ( \25831 , \17539 );
not \U$25489 ( \25832 , \5908 );
or \U$25490 ( \25833 , \25831 , \25832 );
or \U$25491 ( \25834 , \6651 , \17539 );
nand \U$25492 ( \25835 , \25833 , \25834 );
nand \U$25493 ( \25836 , \25835 , \17251 );
nand \U$25494 ( \25837 , \25830 , \25836 );
not \U$25495 ( \25838 , \25837 );
nand \U$25496 ( \25839 , \24966 , RI9873648_192);
xnor \U$25497 ( \25840 , RI9873558_190, \914 );
nand \U$25498 ( \25841 , \25840 , \18615 );
and \U$25499 ( \25842 , \25839 , \25841 );
not \U$25500 ( \25843 , \11433 );
not \U$25501 ( \25844 , RI98719b0_131);
not \U$25502 ( \25845 , \12773 );
or \U$25503 ( \25846 , \25844 , \25845 );
not \U$25504 ( \25847 , \17081 );
or \U$25505 ( \25848 , \25847 , RI98719b0_131);
nand \U$25506 ( \25849 , \25846 , \25848 );
not \U$25507 ( \25850 , \25849 );
or \U$25508 ( \25851 , \25843 , \25850 );
nand \U$25509 ( \25852 , \25210 , \796 );
nand \U$25510 ( \25853 , \25851 , \25852 );
not \U$25511 ( \25854 , \25853 );
xnor \U$25512 ( \25855 , \25174 , \25185 );
not \U$25513 ( \25856 , \25855 );
not \U$25514 ( \25857 , \2087 );
not \U$25515 ( \25858 , \25234 );
or \U$25516 ( \25859 , \25857 , \25858 );
and \U$25517 ( \25860 , RI9871aa0_133, \10064 );
not \U$25518 ( \25861 , RI9871aa0_133);
and \U$25519 ( \25862 , \25861 , \11358 );
or \U$25520 ( \25863 , \25860 , \25862 );
nand \U$25521 ( \25864 , \25863 , \2071 );
nand \U$25522 ( \25865 , \25859 , \25864 );
not \U$25523 ( \25866 , \25865 );
or \U$25524 ( \25867 , \25856 , \25866 );
or \U$25525 ( \25868 , \25865 , \25855 );
nand \U$25526 ( \25869 , \25867 , \25868 );
not \U$25527 ( \25870 , \25869 );
or \U$25528 ( \25871 , \25854 , \25870 );
not \U$25529 ( \25872 , \25855 );
nand \U$25530 ( \25873 , \25872 , \25865 );
nand \U$25531 ( \25874 , \25871 , \25873 );
not \U$25532 ( \25875 , \25874 );
and \U$25533 ( \25876 , \25842 , \25875 );
not \U$25534 ( \25877 , \25842 );
and \U$25535 ( \25878 , \25877 , \25874 );
nor \U$25536 ( \25879 , \25876 , \25878 );
not \U$25537 ( \25880 , \25879 );
or \U$25538 ( \25881 , \25838 , \25880 );
not \U$25539 ( \25882 , \25841 );
not \U$25540 ( \25883 , \25839 );
or \U$25541 ( \25884 , \25882 , \25883 );
nand \U$25542 ( \25885 , \25884 , \25874 );
nand \U$25543 ( \25886 , \25881 , \25885 );
not \U$25544 ( \25887 , \25886 );
not \U$25545 ( \25888 , \25887 );
xor \U$25546 ( \25889 , \24973 , \24955 );
not \U$25547 ( \25890 , \25889 );
or \U$25548 ( \25891 , \25888 , \25890 );
or \U$25549 ( \25892 , \25889 , \25887 );
nand \U$25550 ( \25893 , \25891 , \25892 );
not \U$25551 ( \25894 , \25893 );
or \U$25552 ( \25895 , \25827 , \25894 );
not \U$25553 ( \25896 , \25887 );
nand \U$25554 ( \25897 , \25896 , \25889 );
nand \U$25555 ( \25898 , \25895 , \25897 );
not \U$25556 ( \25899 , \25898 );
or \U$25557 ( \25900 , \25824 , \25899 );
not \U$25558 ( \25901 , \25821 );
not \U$25559 ( \25902 , \25823 );
or \U$25560 ( \25903 , \25901 , \25902 );
nand \U$25561 ( \25904 , \25900 , \25903 );
not \U$25562 ( \25905 , \25904 );
xor \U$25563 ( \25906 , \24674 , \24670 );
xor \U$25564 ( \25907 , \25906 , \24691 );
not \U$25565 ( \25908 , \25907 );
not \U$25566 ( \25909 , \25908 );
or \U$25567 ( \25910 , \25905 , \25909 );
not \U$25568 ( \25911 , \25904 );
nand \U$25569 ( \25912 , \25911 , \25907 );
nand \U$25570 ( \25913 , \25910 , \25912 );
not \U$25571 ( \25914 , \25913 );
or \U$25572 ( \25915 , \25819 , \25914 );
nand \U$25573 ( \25916 , \25907 , \25904 );
nand \U$25574 ( \25917 , \25915 , \25916 );
nor \U$25575 ( \25918 , \25709 , \25917 );
not \U$25576 ( \25919 , \25294 );
xor \U$25577 ( \25920 , \25297 , \25919 );
xnor \U$25578 ( \25921 , \25920 , \25308 );
or \U$25579 ( \25922 , \25918 , \25921 );
not \U$25580 ( \25923 , \25708 );
nand \U$25581 ( \25924 , \25923 , \25917 );
nand \U$25582 ( \25925 , \25922 , \25924 );
not \U$25583 ( \25926 , \25925 );
or \U$25584 ( \25927 , \25702 , \25926 );
not \U$25585 ( \25928 , \25320 );
nand \U$25586 ( \25929 , \25928 , \25696 );
nand \U$25587 ( \25930 , \25927 , \25929 );
and \U$25588 ( \25931 , \25319 , \25930 );
and \U$25589 ( \25932 , \25316 , \25318 );
or \U$25590 ( \25933 , \25931 , \25932 );
nand \U$25591 ( \25934 , \25137 , \25933 );
nand \U$25592 ( \25935 , \24618 , \25117 );
nand \U$25593 ( \25936 , \25934 , \25935 );
not \U$25594 ( \25937 , \25936 );
or \U$25595 ( \25938 , \25135 , \25937 );
buf \U$25596 ( \25939 , \25128 );
nand \U$25597 ( \25940 , \25939 , \25132 );
nand \U$25598 ( \25941 , \25938 , \25940 );
not \U$25599 ( \25942 , \25941 );
or \U$25600 ( \25943 , \24045 , \25942 );
not \U$25601 ( \25944 , \23816 );
not \U$25602 ( \25945 , \24043 );
nand \U$25603 ( \25946 , \25944 , \25945 );
nand \U$25604 ( \25947 , \25943 , \25946 );
not \U$25605 ( \25948 , \23236 );
nor \U$25606 ( \25949 , \23812 , \25948 );
and \U$25607 ( \25950 , \21481 , \22236 );
nor \U$25608 ( \25951 , \23232 , \22239 );
nor \U$25609 ( \25952 , \25950 , \25951 );
nand \U$25610 ( \25953 , \25947 , \25949 , \25952 );
buf \U$25611 ( \25954 , \23804 );
nand \U$25612 ( \25955 , \23811 , \25954 );
nand \U$25613 ( \25956 , \23814 , \25953 , \25955 );
not \U$25614 ( \25957 , \23798 );
not \U$25615 ( \25958 , \23801 );
or \U$25616 ( \25959 , \25957 , \25958 );
nand \U$25617 ( \25960 , \23797 , \23791 );
nand \U$25618 ( \25961 , \25959 , \25960 );
not \U$25619 ( \25962 , \25961 );
not \U$25620 ( \25963 , \23558 );
not \U$25621 ( \25964 , \23553 );
or \U$25622 ( \25965 , \25963 , \25964 );
nand \U$25623 ( \25966 , \23548 , \23543 );
nand \U$25624 ( \25967 , \25965 , \25966 );
not \U$25625 ( \25968 , \25967 );
not \U$25626 ( \25969 , \25968 );
not \U$25627 ( \25970 , \3465 );
not \U$25628 ( \25971 , \23385 );
or \U$25629 ( \25972 , \25970 , \25971 );
nand \U$25630 ( \25973 , \14011 , \3467 );
nand \U$25631 ( \25974 , \25972 , \25973 );
not \U$25632 ( \25975 , \4101 );
not \U$25633 ( \25976 , \23395 );
or \U$25634 ( \25977 , \25975 , \25976 );
nand \U$25635 ( \25978 , \14217 , \4084 );
nand \U$25636 ( \25979 , \25977 , \25978 );
not \U$25637 ( \25980 , \25979 );
xor \U$25638 ( \25981 , \25974 , \25980 );
not \U$25639 ( \25982 , \10487 );
not \U$25640 ( \25983 , \14230 );
or \U$25641 ( \25984 , \25982 , \25983 );
nand \U$25642 ( \25985 , \23405 , \9670 );
nand \U$25643 ( \25986 , \25984 , \25985 );
xor \U$25644 ( \25987 , \25981 , \25986 );
not \U$25645 ( \25988 , \9214 );
not \U$25646 ( \25989 , \14021 );
or \U$25647 ( \25990 , \25988 , \25989 );
nand \U$25648 ( \25991 , \23350 , \9196 );
nand \U$25649 ( \25992 , \25990 , \25991 );
not \U$25650 ( \25993 , \17243 );
not \U$25651 ( \25994 , \23362 );
or \U$25652 ( \25995 , \25993 , \25994 );
nand \U$25653 ( \25996 , \13479 , \13484 );
nand \U$25654 ( \25997 , \25995 , \25996 );
xor \U$25655 ( \25998 , \25992 , \25997 );
not \U$25656 ( \25999 , \9937 );
not \U$25657 ( \26000 , \14134 );
or \U$25658 ( \26001 , \25999 , \26000 );
nand \U$25659 ( \26002 , \23373 , \9952 );
nand \U$25660 ( \26003 , \26001 , \26002 );
xnor \U$25661 ( \26004 , \25998 , \26003 );
xor \U$25662 ( \26005 , \25987 , \26004 );
not \U$25663 ( \26006 , \8029 );
not \U$25664 ( \26007 , \23415 );
or \U$25665 ( \26008 , \26006 , \26007 );
nand \U$25666 ( \26009 , \14066 , \8041 );
nand \U$25667 ( \26010 , \26008 , \26009 );
and \U$25668 ( \26011 , \8743 , \23424 );
and \U$25669 ( \26012 , \14084 , \11199 );
nor \U$25670 ( \26013 , \26011 , \26012 );
xor \U$25671 ( \26014 , \26010 , \26013 );
not \U$25672 ( \26015 , \7325 );
not \U$25673 ( \26016 , \23434 );
or \U$25674 ( \26017 , \26015 , \26016 );
nand \U$25675 ( \26018 , \14036 , \7338 );
nand \U$25676 ( \26019 , \26017 , \26018 );
xor \U$25677 ( \26020 , \26014 , \26019 );
xor \U$25678 ( \26021 , \26005 , \26020 );
not \U$25679 ( \26022 , \26021 );
not \U$25680 ( \26023 , \26022 );
or \U$25681 ( \26024 , \25969 , \26023 );
nand \U$25682 ( \26025 , \26021 , \25967 );
nand \U$25683 ( \26026 , \26024 , \26025 );
not \U$25684 ( \26027 , \23419 );
not \U$25685 ( \26028 , \23438 );
or \U$25686 ( \26029 , \26027 , \26028 );
or \U$25687 ( \26030 , \23419 , \23438 );
nand \U$25688 ( \26031 , \26030 , \23428 );
nand \U$25689 ( \26032 , \26029 , \26031 );
not \U$25690 ( \26033 , \5642 );
not \U$25691 ( \26034 , \23319 );
or \U$25692 ( \26035 , \26033 , \26034 );
nand \U$25693 ( \26036 , \14110 , \5653 );
nand \U$25694 ( \26037 , \26035 , \26036 );
not \U$25695 ( \26038 , \5034 );
not \U$25696 ( \26039 , \23330 );
or \U$25697 ( \26040 , \26038 , \26039 );
nand \U$25698 ( \26041 , \14167 , \5036 );
nand \U$25699 ( \26042 , \26040 , \26041 );
not \U$25700 ( \26043 , \26042 );
xor \U$25701 ( \26044 , \26037 , \26043 );
not \U$25702 ( \26045 , \10242 );
not \U$25703 ( \26046 , \14122 );
or \U$25704 ( \26047 , \26045 , \26046 );
nand \U$25705 ( \26048 , \23339 , \10251 );
nand \U$25706 ( \26049 , \26047 , \26048 );
xnor \U$25707 ( \26050 , \26044 , \26049 );
xor \U$25708 ( \26051 , \26032 , \26050 );
not \U$25709 ( \26052 , \6284 );
not \U$25710 ( \26053 , \23447 );
or \U$25711 ( \26054 , \26052 , \26053 );
nand \U$25712 ( \26055 , \14056 , \6611 );
nand \U$25713 ( \26056 , \26054 , \26055 );
not \U$25714 ( \26057 , \12868 );
not \U$25715 ( \26058 , \14073 );
or \U$25716 ( \26059 , \26057 , \26058 );
nand \U$25717 ( \26060 , \23456 , \13020 );
nand \U$25718 ( \26061 , \26059 , \26060 );
xor \U$25719 ( \26062 , \26056 , \26061 );
not \U$25720 ( \26063 , \9686 );
not \U$25721 ( \26064 , \23465 );
or \U$25722 ( \26065 , \26063 , \26064 );
nand \U$25723 ( \26066 , \14046 , \9273 );
nand \U$25724 ( \26067 , \26065 , \26066 );
xnor \U$25725 ( \26068 , \26062 , \26067 );
not \U$25726 ( \26069 , \26068 );
xor \U$25727 ( \26070 , \26051 , \26069 );
not \U$25728 ( \26071 , \26070 );
and \U$25729 ( \26072 , \26026 , \26071 );
not \U$25730 ( \26073 , \26026 );
and \U$25731 ( \26074 , \26073 , \26070 );
nor \U$25732 ( \26075 , \26072 , \26074 );
not \U$25733 ( \26076 , \26075 );
not \U$25734 ( \26077 , \876 );
not \U$25735 ( \26078 , \23715 );
or \U$25736 ( \26079 , \26077 , \26078 );
nand \U$25737 ( \26080 , \13455 , \9876 );
nand \U$25738 ( \26081 , \26079 , \26080 );
not \U$25739 ( \26082 , \1501 );
not \U$25740 ( \26083 , \23723 );
or \U$25741 ( \26084 , \26082 , \26083 );
nand \U$25742 ( \26085 , \13586 , \1518 );
nand \U$25743 ( \26086 , \26084 , \26085 );
xor \U$25744 ( \26087 , \26081 , \26086 );
not \U$25745 ( \26088 , \12720 );
not \U$25746 ( \26089 , \23689 );
or \U$25747 ( \26090 , \26088 , \26089 );
nand \U$25748 ( \26091 , \13566 , \1323 );
nand \U$25749 ( \26092 , \26090 , \26091 );
xor \U$25750 ( \26093 , \26087 , \26092 );
not \U$25751 ( \26094 , \13830 );
not \U$25752 ( \26095 , \13839 );
or \U$25753 ( \26096 , \26094 , \26095 );
nand \U$25754 ( \26097 , \13831 , \13838 );
nand \U$25755 ( \26098 , \26096 , \26097 );
and \U$25756 ( \26099 , \26098 , \13850 );
not \U$25757 ( \26100 , \26098 );
not \U$25758 ( \26101 , \13850 );
and \U$25759 ( \26102 , \26100 , \26101 );
nor \U$25760 ( \26103 , \26099 , \26102 );
xor \U$25761 ( \26104 , \26093 , \26103 );
xor \U$25762 ( \26105 , \13935 , \13914 );
not \U$25763 ( \26106 , \13899 );
xnor \U$25764 ( \26107 , \26105 , \26106 );
xnor \U$25765 ( \26108 , \26104 , \26107 );
not \U$25766 ( \26109 , \26108 );
not \U$25767 ( \26110 , \23313 );
not \U$25768 ( \26111 , \23376 );
or \U$25769 ( \26112 , \26110 , \26111 );
or \U$25770 ( \26113 , \23376 , \23313 );
nand \U$25771 ( \26114 , \26113 , \23344 );
nand \U$25772 ( \26115 , \26112 , \26114 );
not \U$25773 ( \26116 , \26115 );
or \U$25774 ( \26117 , \26109 , \26116 );
or \U$25775 ( \26118 , \26115 , \26108 );
nand \U$25776 ( \26119 , \26117 , \26118 );
xor \U$25777 ( \26120 , \23354 , \23364 );
and \U$25778 ( \26121 , \26120 , \23375 );
and \U$25779 ( \26122 , \23354 , \23364 );
or \U$25780 ( \26123 , \26121 , \26122 );
xor \U$25781 ( \26124 , \23323 , \23332 );
and \U$25782 ( \26125 , \26124 , \23343 );
and \U$25783 ( \26126 , \23323 , \23332 );
or \U$25784 ( \26127 , \26125 , \26126 );
xor \U$25785 ( \26128 , \26123 , \26127 );
xor \U$25786 ( \26129 , \23449 , \23458 );
and \U$25787 ( \26130 , \26129 , \23469 );
and \U$25788 ( \26131 , \23449 , \23458 );
or \U$25789 ( \26132 , \26130 , \26131 );
xor \U$25790 ( \26133 , \26128 , \26132 );
not \U$25791 ( \26134 , \26133 );
and \U$25792 ( \26135 , \26119 , \26134 );
not \U$25793 ( \26136 , \26119 );
and \U$25794 ( \26137 , \26136 , \26133 );
nor \U$25795 ( \26138 , \26135 , \26137 );
not \U$25796 ( \26139 , \26138 );
nand \U$25797 ( \26140 , \26076 , \26139 );
nand \U$25798 ( \26141 , \26075 , \26138 );
nand \U$25799 ( \26142 , \26140 , \26141 );
not \U$25800 ( \26143 , \26142 );
not \U$25801 ( \26144 , \23480 );
not \U$25802 ( \26145 , \23476 );
or \U$25803 ( \26146 , \26144 , \26145 );
or \U$25804 ( \26147 , \23472 , \23377 );
nand \U$25805 ( \26148 , \26146 , \26147 );
not \U$25806 ( \26149 , \26148 );
and \U$25807 ( \26150 , \26143 , \26149 );
and \U$25808 ( \26151 , \26142 , \26148 );
nor \U$25809 ( \26152 , \26150 , \26151 );
not \U$25810 ( \26153 , \23485 );
nand \U$25811 ( \26154 , \23289 , \26153 );
not \U$25812 ( \26155 , \23282 );
nand \U$25813 ( \26156 , \26155 , \23288 );
and \U$25814 ( \26157 , \26154 , \26156 );
xor \U$25815 ( \26158 , \26152 , \26157 );
not \U$25816 ( \26159 , \23755 );
not \U$25817 ( \26160 , \26159 );
not \U$25818 ( \26161 , \23766 );
or \U$25819 ( \26162 , \26160 , \26161 );
nand \U$25820 ( \26163 , \26162 , \23637 );
not \U$25821 ( \26164 , \23766 );
nand \U$25822 ( \26165 , \26164 , \23755 );
and \U$25823 ( \26166 , \26163 , \26165 );
xnor \U$25824 ( \26167 , \26158 , \26166 );
not \U$25825 ( \26168 , \23508 );
not \U$25826 ( \26169 , \23777 );
or \U$25827 ( \26170 , \26168 , \26169 );
nand \U$25828 ( \26171 , \26170 , \23502 );
not \U$25829 ( \26172 , \23508 );
nand \U$25830 ( \26173 , \26172 , \23776 );
nand \U$25831 ( \26174 , \26171 , \26173 );
xor \U$25832 ( \26175 , \26167 , \26174 );
not \U$25833 ( \26176 , \23410 );
not \U$25834 ( \26177 , \23470 );
nand \U$25835 ( \26178 , \26177 , \23439 );
not \U$25836 ( \26179 , \26178 );
or \U$25837 ( \26180 , \26176 , \26179 );
not \U$25838 ( \26181 , \23439 );
nand \U$25839 ( \26182 , \26181 , \23470 );
nand \U$25840 ( \26183 , \26180 , \26182 );
xor \U$25841 ( \26184 , \23249 , \23253 );
and \U$25842 ( \26185 , \26184 , \23258 );
and \U$25843 ( \26186 , \23249 , \23253 );
or \U$25844 ( \26187 , \26185 , \26186 );
not \U$25845 ( \26188 , \23647 );
not \U$25846 ( \26189 , \23679 );
or \U$25847 ( \26190 , \26188 , \26189 );
nand \U$25848 ( \26191 , \23673 , \23666 );
nand \U$25849 ( \26192 , \26190 , \26191 );
xor \U$25850 ( \26193 , \26187 , \26192 );
xnor \U$25851 ( \26194 , \26183 , \26193 );
xor \U$25852 ( \26195 , \23694 , \23699 );
and \U$25853 ( \26196 , \26195 , \23706 );
and \U$25854 ( \26197 , \23694 , \23699 );
or \U$25855 ( \26198 , \26196 , \26197 );
not \U$25856 ( \26199 , \26198 );
nand \U$25857 ( \26200 , \23312 , \23295 );
not \U$25858 ( \26201 , \23302 );
nand \U$25859 ( \26202 , \26201 , \23308 );
nand \U$25860 ( \26203 , \26200 , \26202 );
not \U$25861 ( \26204 , \23595 );
not \U$25862 ( \26205 , \26204 );
not \U$25863 ( \26206 , \23603 );
or \U$25864 ( \26207 , \26205 , \26206 );
nand \U$25865 ( \26208 , \26207 , \23597 );
xor \U$25866 ( \26209 , \26203 , \26208 );
not \U$25867 ( \26210 , \26209 );
not \U$25868 ( \26211 , \26210 );
or \U$25869 ( \26212 , \26199 , \26211 );
not \U$25870 ( \26213 , \26198 );
nand \U$25871 ( \26214 , \26213 , \26209 );
nand \U$25872 ( \26215 , \26212 , \26214 );
xor \U$25873 ( \26216 , \14188 , \14199 );
xor \U$25874 ( \26217 , \26216 , \14209 );
xor \U$25875 ( \26218 , \23389 , \23399 );
and \U$25876 ( \26219 , \26218 , \23409 );
and \U$25877 ( \26220 , \23389 , \23399 );
or \U$25878 ( \26221 , \26219 , \26220 );
xor \U$25879 ( \26222 , \26217 , \26221 );
not \U$25880 ( \26223 , \23728 );
not \U$25881 ( \26224 , \23719 );
and \U$25882 ( \26225 , \23734 , \26224 );
not \U$25883 ( \26226 , \23734 );
and \U$25884 ( \26227 , \26226 , \23719 );
nor \U$25885 ( \26228 , \26225 , \26227 );
not \U$25886 ( \26229 , \26228 );
or \U$25887 ( \26230 , \26223 , \26229 );
nand \U$25888 ( \26231 , \23735 , \26224 );
nand \U$25889 ( \26232 , \26230 , \26231 );
xor \U$25890 ( \26233 , \26222 , \26232 );
xor \U$25891 ( \26234 , \26215 , \26233 );
xor \U$25892 ( \26235 , \23707 , \23736 );
and \U$25893 ( \26236 , \26235 , \23748 );
and \U$25894 ( \26237 , \23707 , \23736 );
or \U$25895 ( \26238 , \26236 , \26237 );
xnor \U$25896 ( \26239 , \26234 , \26238 );
not \U$25897 ( \26240 , \26239 );
not \U$25898 ( \26241 , \23277 );
not \U$25899 ( \26242 , \23259 );
or \U$25900 ( \26243 , \26241 , \26242 );
or \U$25901 ( \26244 , \23259 , \23277 );
nand \U$25902 ( \26245 , \26244 , \23264 );
nand \U$25903 ( \26246 , \26243 , \26245 );
not \U$25904 ( \26247 , \26246 );
or \U$25905 ( \26248 , \26240 , \26247 );
or \U$25906 ( \26249 , \26246 , \26239 );
nand \U$25907 ( \26250 , \26248 , \26249 );
xnor \U$25908 ( \26251 , \26194 , \26250 );
not \U$25909 ( \26252 , \23623 );
not \U$25910 ( \26253 , \23514 );
nand \U$25911 ( \26254 , \26253 , \23563 );
not \U$25912 ( \26255 , \26254 );
or \U$25913 ( \26256 , \26252 , \26255 );
not \U$25914 ( \26257 , \23563 );
nand \U$25915 ( \26258 , \26257 , \23514 );
nand \U$25916 ( \26259 , \26256 , \26258 );
and \U$25917 ( \26260 , \23582 , \23605 );
and \U$25918 ( \26261 , \23589 , \23604 );
nor \U$25919 ( \26262 , \26260 , \26261 );
not \U$25920 ( \26263 , \26262 );
xnor \U$25921 ( \26264 , \13869 , \13882 );
not \U$25922 ( \26265 , \23665 );
not \U$25923 ( \26266 , \23660 );
or \U$25924 ( \26267 , \26265 , \26266 );
nand \U$25925 ( \26268 , \23659 , \23654 );
nand \U$25926 ( \26269 , \26267 , \26268 );
xor \U$25927 ( \26270 , \26264 , \26269 );
not \U$25928 ( \26271 , \4925 );
not \U$25929 ( \26272 , \14175 );
or \U$25930 ( \26273 , \26271 , \26272 );
nand \U$25931 ( \26274 , \23527 , \6553 );
nand \U$25932 ( \26275 , \26273 , \26274 );
xnor \U$25933 ( \26276 , \26270 , \26275 );
not \U$25934 ( \26277 , \26276 );
not \U$25935 ( \26278 , \23542 );
not \U$25936 ( \26279 , \23536 );
or \U$25937 ( \26280 , \26278 , \26279 );
nand \U$25938 ( \26281 , \23531 , \23520 );
nand \U$25939 ( \26282 , \26280 , \26281 );
not \U$25940 ( \26283 , \26282 );
or \U$25941 ( \26284 , \26277 , \26283 );
or \U$25942 ( \26285 , \26282 , \26276 );
nand \U$25943 ( \26286 , \26284 , \26285 );
not \U$25944 ( \26287 , \26286 );
or \U$25945 ( \26288 , \26263 , \26287 );
or \U$25946 ( \26289 , \26286 , \26262 );
nand \U$25947 ( \26290 , \26288 , \26289 );
not \U$25948 ( \26291 , \26290 );
not \U$25949 ( \26292 , \23615 );
not \U$25950 ( \26293 , \23571 );
or \U$25951 ( \26294 , \26292 , \26293 );
not \U$25952 ( \26295 , \23577 );
nand \U$25953 ( \26296 , \26295 , \23611 );
nand \U$25954 ( \26297 , \26294 , \26296 );
not \U$25955 ( \26298 , \26297 );
not \U$25956 ( \26299 , \26298 );
or \U$25957 ( \26300 , \26291 , \26299 );
not \U$25958 ( \26301 , \26290 );
nand \U$25959 ( \26302 , \26301 , \26297 );
nand \U$25960 ( \26303 , \26300 , \26302 );
xor \U$25961 ( \26304 , \23683 , \23749 );
and \U$25962 ( \26305 , \26304 , \23754 );
and \U$25963 ( \26306 , \23683 , \23749 );
or \U$25964 ( \26307 , \26305 , \26306 );
xor \U$25965 ( \26308 , \26303 , \26307 );
xor \U$25966 ( \26309 , \26259 , \26308 );
xor \U$25967 ( \26310 , \26251 , \26309 );
and \U$25968 ( \26311 , \23770 , \23632 );
and \U$25969 ( \26312 , \23625 , \23630 );
nor \U$25970 ( \26313 , \26311 , \26312 );
xor \U$25971 ( \26314 , \26310 , \26313 );
nor \U$25972 ( \26315 , \23501 , \23243 );
or \U$25973 ( \26316 , \26315 , \23489 );
nand \U$25974 ( \26317 , \23501 , \23243 );
nand \U$25975 ( \26318 , \26316 , \26317 );
xor \U$25976 ( \26319 , \26314 , \26318 );
xor \U$25977 ( \26320 , \26175 , \26319 );
nand \U$25978 ( \26321 , \25962 , \26320 );
not \U$25979 ( \26322 , \26319 );
not \U$25980 ( \26323 , \26174 );
nand \U$25981 ( \26324 , \26323 , \26167 );
nand \U$25982 ( \26325 , \26322 , \26324 );
not \U$25983 ( \26326 , \26325 );
not \U$25984 ( \26327 , \26173 );
not \U$25985 ( \26328 , \26171 );
or \U$25986 ( \26329 , \26327 , \26328 );
not \U$25987 ( \26330 , \26167 );
nand \U$25988 ( \26331 , \26329 , \26330 );
not \U$25989 ( \26332 , \26331 );
or \U$25990 ( \26333 , \26326 , \26332 );
nand \U$25991 ( \26334 , \26166 , \26152 );
not \U$25992 ( \26335 , \26157 );
and \U$25993 ( \26336 , \26334 , \26335 );
nor \U$25994 ( \26337 , \26166 , \26152 );
nor \U$25995 ( \26338 , \26336 , \26337 );
not \U$25996 ( \26339 , \26251 );
not \U$25997 ( \26340 , \26309 );
or \U$25998 ( \26341 , \26339 , \26340 );
nand \U$25999 ( \26342 , \26308 , \26259 );
nand \U$26000 ( \26343 , \26341 , \26342 );
not \U$26001 ( \26344 , \26343 );
not \U$26002 ( \26345 , \26307 );
not \U$26003 ( \26346 , \26303 );
or \U$26004 ( \26347 , \26345 , \26346 );
nand \U$26005 ( \26348 , \26290 , \26297 );
nand \U$26006 ( \26349 , \26347 , \26348 );
not \U$26007 ( \26350 , \26133 );
not \U$26008 ( \26351 , \26119 );
or \U$26009 ( \26352 , \26350 , \26351 );
not \U$26010 ( \26353 , \26108 );
nand \U$26011 ( \26354 , \26353 , \26115 );
nand \U$26012 ( \26355 , \26352 , \26354 );
xor \U$26013 ( \26356 , \14068 , \14077 );
xor \U$26014 ( \26357 , \26356 , \14088 );
xor \U$26015 ( \26358 , \13084 , \14169 );
xor \U$26016 ( \26359 , \26358 , \14179 );
or \U$26017 ( \26360 , \26357 , \26359 );
nand \U$26018 ( \26361 , \26357 , \26359 );
nand \U$26019 ( \26362 , \26360 , \26361 );
xor \U$26020 ( \26363 , \14114 , \14138 );
xnor \U$26021 ( \26364 , \26363 , \14124 );
xnor \U$26022 ( \26365 , \26362 , \26364 );
not \U$26023 ( \26366 , \26365 );
or \U$26024 ( \26367 , \26233 , \26215 );
nand \U$26025 ( \26368 , \26367 , \26238 );
nand \U$26026 ( \26369 , \26233 , \26215 );
nand \U$26027 ( \26370 , \26368 , \26369 );
not \U$26028 ( \26371 , \26370 );
or \U$26029 ( \26372 , \26366 , \26371 );
or \U$26030 ( \26373 , \26370 , \26365 );
nand \U$26031 ( \26374 , \26372 , \26373 );
xnor \U$26032 ( \26375 , \26355 , \26374 );
xnor \U$26033 ( \26376 , \26349 , \26375 );
not \U$26034 ( \26377 , \26194 );
not \U$26035 ( \26378 , \26377 );
not \U$26036 ( \26379 , \26250 );
or \U$26037 ( \26380 , \26378 , \26379 );
not \U$26038 ( \26381 , \26239 );
nand \U$26039 ( \26382 , \26381 , \26246 );
nand \U$26040 ( \26383 , \26380 , \26382 );
xnor \U$26041 ( \26384 , \26376 , \26383 );
not \U$26042 ( \26385 , \26384 );
or \U$26043 ( \26386 , \26344 , \26385 );
or \U$26044 ( \26387 , \26343 , \26384 );
nand \U$26045 ( \26388 , \26386 , \26387 );
not \U$26046 ( \26389 , \26388 );
xnor \U$26047 ( \26390 , \13636 , \13606 );
xor \U$26048 ( \26391 , \26081 , \26086 );
and \U$26049 ( \26392 , \26391 , \26092 );
and \U$26050 ( \26393 , \26081 , \26086 );
or \U$26051 ( \26394 , \26392 , \26393 );
xnor \U$26052 ( \26395 , \26390 , \26394 );
not \U$26053 ( \26396 , \26056 );
not \U$26054 ( \26397 , \26067 );
or \U$26055 ( \26398 , \26396 , \26397 );
or \U$26056 ( \26399 , \26067 , \26056 );
nand \U$26057 ( \26400 , \26399 , \26061 );
nand \U$26058 ( \26401 , \26398 , \26400 );
xor \U$26059 ( \26402 , \26395 , \26401 );
not \U$26060 ( \26403 , \13945 );
not \U$26061 ( \26404 , \13888 );
not \U$26062 ( \26405 , \26404 );
and \U$26063 ( \26406 , \26403 , \26405 );
and \U$26064 ( \26407 , \13945 , \26404 );
nor \U$26065 ( \26408 , \26406 , \26407 );
xnor \U$26066 ( \26409 , \26402 , \26408 );
xor \U$26067 ( \26410 , \26123 , \26127 );
and \U$26068 ( \26411 , \26410 , \26132 );
and \U$26069 ( \26412 , \26123 , \26127 );
or \U$26070 ( \26413 , \26411 , \26412 );
not \U$26071 ( \26414 , \26413 );
and \U$26072 ( \26415 , \26409 , \26414 );
not \U$26073 ( \26416 , \26409 );
and \U$26074 ( \26417 , \26416 , \26413 );
nor \U$26075 ( \26418 , \26415 , \26417 );
not \U$26076 ( \26419 , \26418 );
not \U$26077 ( \26420 , \26419 );
and \U$26078 ( \26421 , \25974 , \25979 );
not \U$26079 ( \26422 , \25974 );
nand \U$26080 ( \26423 , \26422 , \25980 );
and \U$26081 ( \26424 , \25986 , \26423 );
nor \U$26082 ( \26425 , \26421 , \26424 );
or \U$26083 ( \26426 , \25992 , \25997 );
nand \U$26084 ( \26427 , \26426 , \26003 );
nand \U$26085 ( \26428 , \25997 , \25992 );
and \U$26086 ( \26429 , \26427 , \26428 );
xor \U$26087 ( \26430 , \26425 , \26429 );
or \U$26088 ( \26431 , \26019 , \26010 );
not \U$26089 ( \26432 , \26013 );
nand \U$26090 ( \26433 , \26431 , \26432 );
nand \U$26091 ( \26434 , \26019 , \26010 );
and \U$26092 ( \26435 , \26433 , \26434 );
xor \U$26093 ( \26436 , \26430 , \26435 );
not \U$26094 ( \26437 , \26436 );
xor \U$26095 ( \26438 , \26217 , \26221 );
and \U$26096 ( \26439 , \26438 , \26232 );
and \U$26097 ( \26440 , \26217 , \26221 );
or \U$26098 ( \26441 , \26439 , \26440 );
not \U$26099 ( \26442 , \26441 );
xor \U$26100 ( \26443 , \26103 , \26107 );
nand \U$26101 ( \26444 , \26443 , \26093 );
not \U$26102 ( \26445 , \26444 );
and \U$26103 ( \26446 , \26103 , \26107 );
nor \U$26104 ( \26447 , \26445 , \26446 );
not \U$26105 ( \26448 , \26447 );
or \U$26106 ( \26449 , \26442 , \26448 );
not \U$26107 ( \26450 , \26446 );
not \U$26108 ( \26451 , \26450 );
not \U$26109 ( \26452 , \26444 );
or \U$26110 ( \26453 , \26451 , \26452 );
not \U$26111 ( \26454 , \26441 );
nand \U$26112 ( \26455 , \26453 , \26454 );
nand \U$26113 ( \26456 , \26449 , \26455 );
not \U$26114 ( \26457 , \26456 );
or \U$26115 ( \26458 , \26437 , \26457 );
or \U$26116 ( \26459 , \26436 , \26456 );
nand \U$26117 ( \26460 , \26458 , \26459 );
not \U$26118 ( \26461 , \26460 );
not \U$26119 ( \26462 , \26461 );
or \U$26120 ( \26463 , \26420 , \26462 );
nand \U$26121 ( \26464 , \26418 , \26460 );
nand \U$26122 ( \26465 , \26463 , \26464 );
not \U$26123 ( \26466 , \26193 );
not \U$26124 ( \26467 , \26183 );
or \U$26125 ( \26468 , \26466 , \26467 );
nand \U$26126 ( \26469 , \26187 , \26192 );
nand \U$26127 ( \26470 , \26468 , \26469 );
not \U$26128 ( \26471 , \26470 );
and \U$26129 ( \26472 , \26465 , \26471 );
not \U$26130 ( \26473 , \26465 );
and \U$26131 ( \26474 , \26473 , \26470 );
nor \U$26132 ( \26475 , \26472 , \26474 );
not \U$26133 ( \26476 , \26475 );
not \U$26134 ( \26477 , \26141 );
not \U$26135 ( \26478 , \26148 );
or \U$26136 ( \26479 , \26477 , \26478 );
nand \U$26137 ( \26480 , \26479 , \26140 );
not \U$26138 ( \26481 , \26480 );
or \U$26139 ( \26482 , \26476 , \26481 );
or \U$26140 ( \26483 , \26475 , \26480 );
nand \U$26141 ( \26484 , \26482 , \26483 );
not \U$26142 ( \26485 , \26022 );
not \U$26143 ( \26486 , \25967 );
or \U$26144 ( \26487 , \26485 , \26486 );
not \U$26145 ( \26488 , \25968 );
not \U$26146 ( \26489 , \26021 );
or \U$26147 ( \26490 , \26488 , \26489 );
nand \U$26148 ( \26491 , \26490 , \26070 );
nand \U$26149 ( \26492 , \26487 , \26491 );
not \U$26150 ( \26493 , \26492 );
not \U$26151 ( \26494 , \26493 );
not \U$26152 ( \26495 , \26050 );
not \U$26153 ( \26496 , \26032 );
nand \U$26154 ( \26497 , \26496 , \26068 );
not \U$26155 ( \26498 , \26497 );
or \U$26156 ( \26499 , \26495 , \26498 );
nand \U$26157 ( \26500 , \26069 , \26032 );
nand \U$26158 ( \26501 , \26499 , \26500 );
and \U$26159 ( \26502 , \13589 , \13568 );
not \U$26160 ( \26503 , \13589 );
not \U$26161 ( \26504 , \13568 );
and \U$26162 ( \26505 , \26503 , \26504 );
nor \U$26163 ( \26506 , \26502 , \26505 );
xor \U$26164 ( \26507 , \13457 , \13468 );
xnor \U$26165 ( \26508 , \26507 , \13494 );
not \U$26166 ( \26509 , \26508 );
and \U$26167 ( \26510 , \26506 , \26509 );
not \U$26168 ( \26511 , \26506 );
and \U$26169 ( \26512 , \26511 , \26508 );
nor \U$26170 ( \26513 , \26510 , \26512 );
not \U$26171 ( \26514 , \26037 );
not \U$26172 ( \26515 , \26043 );
not \U$26173 ( \26516 , \26049 );
or \U$26174 ( \26517 , \26515 , \26516 );
or \U$26175 ( \26518 , \26049 , \26043 );
nand \U$26176 ( \26519 , \26517 , \26518 );
not \U$26177 ( \26520 , \26519 );
or \U$26178 ( \26521 , \26514 , \26520 );
nand \U$26179 ( \26522 , \26049 , \26042 );
nand \U$26180 ( \26523 , \26521 , \26522 );
xnor \U$26181 ( \26524 , \26513 , \26523 );
nor \U$26182 ( \26525 , \26501 , \26524 );
not \U$26183 ( \26526 , \26525 );
nand \U$26184 ( \26527 , \26501 , \26524 );
nand \U$26185 ( \26528 , \26526 , \26527 );
xor \U$26186 ( \26529 , \25987 , \26004 );
and \U$26187 ( \26530 , \26529 , \26020 );
and \U$26188 ( \26531 , \25987 , \26004 );
or \U$26189 ( \26532 , \26530 , \26531 );
and \U$26190 ( \26533 , \26528 , \26532 );
not \U$26191 ( \26534 , \26528 );
not \U$26192 ( \26535 , \26532 );
and \U$26193 ( \26536 , \26534 , \26535 );
nor \U$26194 ( \26537 , \26533 , \26536 );
not \U$26195 ( \26538 , \26537 );
or \U$26196 ( \26539 , \26494 , \26538 );
or \U$26197 ( \26540 , \26537 , \26493 );
nand \U$26198 ( \26541 , \26539 , \26540 );
not \U$26199 ( \26542 , \26262 );
not \U$26200 ( \26543 , \26542 );
not \U$26201 ( \26544 , \26286 );
or \U$26202 ( \26545 , \26543 , \26544 );
not \U$26203 ( \26546 , \26276 );
nand \U$26204 ( \26547 , \26546 , \26282 );
nand \U$26205 ( \26548 , \26545 , \26547 );
xor \U$26206 ( \26549 , \14212 , \14219 );
xor \U$26207 ( \26550 , \26549 , \14232 );
not \U$26208 ( \26551 , \26550 );
buf \U$26209 ( \26552 , \13652 );
not \U$26210 ( \26553 , \26552 );
xnor \U$26211 ( \26554 , \13664 , \13677 );
not \U$26212 ( \26555 , \26554 );
or \U$26213 ( \26556 , \26553 , \26555 );
or \U$26214 ( \26557 , \26554 , \26552 );
nand \U$26215 ( \26558 , \26556 , \26557 );
not \U$26216 ( \26559 , \26275 );
not \U$26217 ( \26560 , \26270 );
or \U$26218 ( \26561 , \26559 , \26560 );
nand \U$26219 ( \26562 , \26269 , \26264 );
nand \U$26220 ( \26563 , \26561 , \26562 );
xor \U$26221 ( \26564 , \26558 , \26563 );
not \U$26222 ( \26565 , \26564 );
or \U$26223 ( \26566 , \26551 , \26565 );
or \U$26224 ( \26567 , \26564 , \26550 );
nand \U$26225 ( \26568 , \26566 , \26567 );
not \U$26226 ( \26569 , \26568 );
xor \U$26227 ( \26570 , \14003 , \14013 );
xnor \U$26228 ( \26571 , \26570 , \14025 );
not \U$26229 ( \26572 , \26571 );
xor \U$26230 ( \26573 , \14038 , \14048 );
xor \U$26231 ( \26574 , \26573 , \14058 );
not \U$26232 ( \26575 , \26574 );
or \U$26233 ( \26576 , \26572 , \26575 );
or \U$26234 ( \26577 , \26574 , \26571 );
nand \U$26235 ( \26578 , \26576 , \26577 );
not \U$26236 ( \26579 , \26578 );
not \U$26237 ( \26580 , \26198 );
not \U$26238 ( \26581 , \26209 );
or \U$26239 ( \26582 , \26580 , \26581 );
not \U$26240 ( \26583 , \26202 );
not \U$26241 ( \26584 , \26200 );
or \U$26242 ( \26585 , \26583 , \26584 );
nand \U$26243 ( \26586 , \26585 , \26208 );
nand \U$26244 ( \26587 , \26582 , \26586 );
not \U$26245 ( \26588 , \26587 );
not \U$26246 ( \26589 , \26588 );
and \U$26247 ( \26590 , \26579 , \26589 );
and \U$26248 ( \26591 , \26578 , \26588 );
nor \U$26249 ( \26592 , \26590 , \26591 );
not \U$26250 ( \26593 , \26592 );
or \U$26251 ( \26594 , \26569 , \26593 );
or \U$26252 ( \26595 , \26568 , \26592 );
nand \U$26253 ( \26596 , \26594 , \26595 );
xor \U$26254 ( \26597 , \26548 , \26596 );
and \U$26255 ( \26598 , \26541 , \26597 );
not \U$26256 ( \26599 , \26541 );
not \U$26257 ( \26600 , \26597 );
and \U$26258 ( \26601 , \26599 , \26600 );
nor \U$26259 ( \26602 , \26598 , \26601 );
xnor \U$26260 ( \26603 , \26484 , \26602 );
not \U$26261 ( \26604 , \26603 );
and \U$26262 ( \26605 , \26389 , \26604 );
and \U$26263 ( \26606 , \26388 , \26603 );
nor \U$26264 ( \26607 , \26605 , \26606 );
xor \U$26265 ( \26608 , \26338 , \26607 );
xor \U$26266 ( \26609 , \26310 , \26313 );
and \U$26267 ( \26610 , \26609 , \26318 );
and \U$26268 ( \26611 , \26310 , \26313 );
or \U$26269 ( \26612 , \26610 , \26611 );
not \U$26270 ( \26613 , \26612 );
xor \U$26271 ( \26614 , \26608 , \26613 );
nand \U$26272 ( \26615 , \26333 , \26614 );
not \U$26273 ( \26616 , \26401 );
not \U$26274 ( \26617 , \26395 );
or \U$26275 ( \26618 , \26616 , \26617 );
not \U$26276 ( \26619 , \26390 );
nand \U$26277 ( \26620 , \26619 , \26394 );
nand \U$26278 ( \26621 , \26618 , \26620 );
not \U$26279 ( \26622 , \26621 );
xor \U$26280 ( \26623 , \26425 , \26429 );
and \U$26281 ( \26624 , \26623 , \26435 );
and \U$26282 ( \26625 , \26425 , \26429 );
or \U$26283 ( \26626 , \26624 , \26625 );
not \U$26284 ( \26627 , \26626 );
or \U$26285 ( \26628 , \26622 , \26627 );
not \U$26286 ( \26629 , \26626 );
not \U$26287 ( \26630 , \26621 );
nand \U$26288 ( \26631 , \26629 , \26630 );
nand \U$26289 ( \26632 , \26628 , \26631 );
xor \U$26290 ( \26633 , \14027 , \14061 );
xor \U$26291 ( \26634 , \26633 , \14091 );
xnor \U$26292 ( \26635 , \26632 , \26634 );
xnor \U$26293 ( \26636 , \13496 , \13513 );
xor \U$26294 ( \26637 , \13685 , \13593 );
xnor \U$26295 ( \26638 , \26636 , \26637 );
not \U$26296 ( \26639 , \26638 );
not \U$26297 ( \26640 , \26513 );
not \U$26298 ( \26641 , \26640 );
not \U$26299 ( \26642 , \26523 );
or \U$26300 ( \26643 , \26641 , \26642 );
nand \U$26301 ( \26644 , \26508 , \26506 );
nand \U$26302 ( \26645 , \26643 , \26644 );
not \U$26303 ( \26646 , \26645 );
not \U$26304 ( \26647 , \26646 );
or \U$26305 ( \26648 , \26639 , \26647 );
not \U$26306 ( \26649 , \26638 );
nand \U$26307 ( \26650 , \26649 , \26645 );
nand \U$26308 ( \26651 , \26648 , \26650 );
not \U$26309 ( \26652 , \26436 );
not \U$26310 ( \26653 , \26652 );
not \U$26311 ( \26654 , \26456 );
or \U$26312 ( \26655 , \26653 , \26654 );
not \U$26313 ( \26656 , \26450 );
not \U$26314 ( \26657 , \26444 );
or \U$26315 ( \26658 , \26656 , \26657 );
nand \U$26316 ( \26659 , \26658 , \26441 );
nand \U$26317 ( \26660 , \26655 , \26659 );
xor \U$26318 ( \26661 , \26651 , \26660 );
xnor \U$26319 ( \26662 , \26635 , \26661 );
not \U$26320 ( \26663 , \14099 );
not \U$26321 ( \26664 , \14103 );
or \U$26322 ( \26665 , \26663 , \26664 );
or \U$26323 ( \26666 , \14099 , \14103 );
nand \U$26324 ( \26667 , \26665 , \26666 );
xnor \U$26325 ( \26668 , \14140 , \26667 );
not \U$26326 ( \26669 , \26668 );
not \U$26327 ( \26670 , \26669 );
nor \U$26328 ( \26671 , \26357 , \26359 );
or \U$26329 ( \26672 , \26364 , \26671 );
nand \U$26330 ( \26673 , \26672 , \26361 );
not \U$26331 ( \26674 , \26673 );
not \U$26332 ( \26675 , \26674 );
or \U$26333 ( \26676 , \26670 , \26675 );
nand \U$26334 ( \26677 , \26673 , \26668 );
nand \U$26335 ( \26678 , \26676 , \26677 );
not \U$26336 ( \26679 , \26550 );
not \U$26337 ( \26680 , \26679 );
not \U$26338 ( \26681 , \26564 );
or \U$26339 ( \26682 , \26680 , \26681 );
nand \U$26340 ( \26683 , \26563 , \26558 );
nand \U$26341 ( \26684 , \26682 , \26683 );
and \U$26342 ( \26685 , \26678 , \26684 );
not \U$26343 ( \26686 , \26678 );
not \U$26344 ( \26687 , \26684 );
and \U$26345 ( \26688 , \26686 , \26687 );
nor \U$26346 ( \26689 , \26685 , \26688 );
not \U$26347 ( \26690 , \26689 );
xor \U$26348 ( \26691 , \14157 , \14154 );
xor \U$26349 ( \26692 , \26691 , \14152 );
not \U$26350 ( \26693 , \26692 );
not \U$26351 ( \26694 , \26693 );
xor \U$26352 ( \26695 , \13812 , \13818 );
xor \U$26353 ( \26696 , \26695 , \13952 );
not \U$26354 ( \26697 , \26696 );
not \U$26355 ( \26698 , \26697 );
or \U$26356 ( \26699 , \26694 , \26698 );
nand \U$26357 ( \26700 , \26692 , \26696 );
nand \U$26358 ( \26701 , \26699 , \26700 );
not \U$26359 ( \26702 , \26587 );
not \U$26360 ( \26703 , \26578 );
or \U$26361 ( \26704 , \26702 , \26703 );
not \U$26362 ( \26705 , \26571 );
nand \U$26363 ( \26706 , \26705 , \26574 );
nand \U$26364 ( \26707 , \26704 , \26706 );
and \U$26365 ( \26708 , \26701 , \26707 );
not \U$26366 ( \26709 , \26701 );
not \U$26367 ( \26710 , \26707 );
and \U$26368 ( \26711 , \26709 , \26710 );
nor \U$26369 ( \26712 , \26708 , \26711 );
not \U$26370 ( \26713 , \26712 );
not \U$26371 ( \26714 , \26713 );
or \U$26372 ( \26715 , \26690 , \26714 );
not \U$26373 ( \26716 , \26689 );
nand \U$26374 ( \26717 , \26712 , \26716 );
nand \U$26375 ( \26718 , \26715 , \26717 );
not \U$26376 ( \26719 , \26548 );
not \U$26377 ( \26720 , \26596 );
or \U$26378 ( \26721 , \26719 , \26720 );
not \U$26379 ( \26722 , \26592 );
nand \U$26380 ( \26723 , \26722 , \26568 );
nand \U$26381 ( \26724 , \26721 , \26723 );
buf \U$26382 ( \26725 , \26724 );
xor \U$26383 ( \26726 , \26718 , \26725 );
xor \U$26384 ( \26727 , \26662 , \26726 );
not \U$26385 ( \26728 , \26597 );
not \U$26386 ( \26729 , \26541 );
or \U$26387 ( \26730 , \26728 , \26729 );
nand \U$26388 ( \26731 , \26537 , \26492 );
nand \U$26389 ( \26732 , \26730 , \26731 );
xor \U$26390 ( \26733 , \26727 , \26732 );
not \U$26391 ( \26734 , \26733 );
not \U$26392 ( \26735 , \26734 );
not \U$26393 ( \26736 , \26374 );
not \U$26394 ( \26737 , \26355 );
or \U$26395 ( \26738 , \26736 , \26737 );
not \U$26396 ( \26739 , \26365 );
nand \U$26397 ( \26740 , \26739 , \26370 );
nand \U$26398 ( \26741 , \26738 , \26740 );
or \U$26399 ( \26742 , \26525 , \26532 );
nand \U$26400 ( \26743 , \26742 , \26527 );
xor \U$26401 ( \26744 , \14182 , \14236 );
xor \U$26402 ( \26745 , \26744 , \14239 );
not \U$26403 ( \26746 , \26413 );
not \U$26404 ( \26747 , \26409 );
or \U$26405 ( \26748 , \26746 , \26747 );
not \U$26406 ( \26749 , \26408 );
xor \U$26407 ( \26750 , \26401 , \26395 );
nand \U$26408 ( \26751 , \26749 , \26750 );
nand \U$26409 ( \26752 , \26748 , \26751 );
xor \U$26410 ( \26753 , \26745 , \26752 );
xor \U$26411 ( \26754 , \26743 , \26753 );
xor \U$26412 ( \26755 , \26741 , \26754 );
not \U$26413 ( \26756 , \26470 );
not \U$26414 ( \26757 , \26465 );
or \U$26415 ( \26758 , \26756 , \26757 );
nand \U$26416 ( \26759 , \26460 , \26419 );
nand \U$26417 ( \26760 , \26758 , \26759 );
not \U$26418 ( \26761 , \26760 );
xor \U$26419 ( \26762 , \26755 , \26761 );
not \U$26420 ( \26763 , \26762 );
not \U$26421 ( \26764 , \26383 );
not \U$26422 ( \26765 , \26376 );
or \U$26423 ( \26766 , \26764 , \26765 );
not \U$26424 ( \26767 , \26375 );
nand \U$26425 ( \26768 , \26767 , \26349 );
nand \U$26426 ( \26769 , \26766 , \26768 );
not \U$26427 ( \26770 , \26769 );
and \U$26428 ( \26771 , \26763 , \26770 );
and \U$26429 ( \26772 , \26769 , \26762 );
nor \U$26430 ( \26773 , \26771 , \26772 );
not \U$26431 ( \26774 , \26602 );
not \U$26432 ( \26775 , \26484 );
or \U$26433 ( \26776 , \26774 , \26775 );
not \U$26434 ( \26777 , \26475 );
nand \U$26435 ( \26778 , \26777 , \26480 );
nand \U$26436 ( \26779 , \26776 , \26778 );
and \U$26437 ( \26780 , \26773 , \26779 );
not \U$26438 ( \26781 , \26773 );
not \U$26439 ( \26782 , \26779 );
and \U$26440 ( \26783 , \26781 , \26782 );
nor \U$26441 ( \26784 , \26780 , \26783 );
not \U$26442 ( \26785 , \26784 );
or \U$26443 ( \26786 , \26735 , \26785 );
not \U$26444 ( \26787 , \26784 );
nand \U$26445 ( \26788 , \26787 , \26733 );
nand \U$26446 ( \26789 , \26786 , \26788 );
not \U$26447 ( \26790 , \26603 );
not \U$26448 ( \26791 , \26790 );
not \U$26449 ( \26792 , \26388 );
or \U$26450 ( \26793 , \26791 , \26792 );
not \U$26451 ( \26794 , \26384 );
nand \U$26452 ( \26795 , \26794 , \26343 );
nand \U$26453 ( \26796 , \26793 , \26795 );
and \U$26454 ( \26797 , \26789 , \26796 );
not \U$26455 ( \26798 , \26789 );
not \U$26456 ( \26799 , \26796 );
and \U$26457 ( \26800 , \26798 , \26799 );
nor \U$26458 ( \26801 , \26797 , \26800 );
xor \U$26459 ( \26802 , \26338 , \26607 );
and \U$26460 ( \26803 , \26802 , \26613 );
and \U$26461 ( \26804 , \26338 , \26607 );
or \U$26462 ( \26805 , \26803 , \26804 );
nand \U$26463 ( \26806 , \26801 , \26805 );
nand \U$26464 ( \26807 , \26321 , \26615 , \26806 );
xor \U$26465 ( \26808 , \26662 , \26726 );
and \U$26466 ( \26809 , \26808 , \26732 );
and \U$26467 ( \26810 , \26662 , \26726 );
or \U$26468 ( \26811 , \26809 , \26810 );
xor \U$26469 ( \26812 , \14094 , \14096 );
xor \U$26470 ( \26813 , \26812 , \14145 );
not \U$26471 ( \26814 , \26629 );
not \U$26472 ( \26815 , \26621 );
or \U$26473 ( \26816 , \26814 , \26815 );
not \U$26474 ( \26817 , \26630 );
not \U$26475 ( \26818 , \26626 );
or \U$26476 ( \26819 , \26817 , \26818 );
nand \U$26477 ( \26820 , \26819 , \26634 );
nand \U$26478 ( \26821 , \26816 , \26820 );
and \U$26479 ( \26822 , \26813 , \26821 );
not \U$26480 ( \26823 , \26813 );
not \U$26481 ( \26824 , \26821 );
and \U$26482 ( \26825 , \26823 , \26824 );
nor \U$26483 ( \26826 , \26822 , \26825 );
not \U$26484 ( \26827 , \26684 );
not \U$26485 ( \26828 , \26678 );
or \U$26486 ( \26829 , \26827 , \26828 );
nand \U$26487 ( \26830 , \26673 , \26669 );
nand \U$26488 ( \26831 , \26829 , \26830 );
and \U$26489 ( \26832 , \26826 , \26831 );
not \U$26490 ( \26833 , \26826 );
not \U$26491 ( \26834 , \26831 );
and \U$26492 ( \26835 , \26833 , \26834 );
nor \U$26493 ( \26836 , \26832 , \26835 );
not \U$26494 ( \26837 , \26724 );
not \U$26495 ( \26838 , \26689 );
or \U$26496 ( \26839 , \26837 , \26838 );
or \U$26497 ( \26840 , \26724 , \26689 );
nand \U$26498 ( \26841 , \26840 , \26712 );
nand \U$26499 ( \26842 , \26839 , \26841 );
nor \U$26500 ( \26843 , \26836 , \26842 );
not \U$26501 ( \26844 , \26843 );
nand \U$26502 ( \26845 , \26842 , \26836 );
nand \U$26503 ( \26846 , \26844 , \26845 );
not \U$26504 ( \26847 , \26707 );
not \U$26505 ( \26848 , \26693 );
or \U$26506 ( \26849 , \26847 , \26848 );
or \U$26507 ( \26850 , \26693 , \26707 );
nand \U$26508 ( \26851 , \26850 , \26696 );
nand \U$26509 ( \26852 , \26849 , \26851 );
xor \U$26510 ( \26853 , \13955 , \13957 );
xor \U$26511 ( \26854 , \26853 , \13960 );
xor \U$26512 ( \26855 , \26852 , \26854 );
not \U$26513 ( \26856 , \14163 );
nand \U$26514 ( \26857 , \26856 , \14245 );
and \U$26515 ( \26858 , \26857 , \14242 );
not \U$26516 ( \26859 , \26857 );
and \U$26517 ( \26860 , \26859 , \14243 );
nor \U$26518 ( \26861 , \26858 , \26860 );
xor \U$26519 ( \26862 , \26855 , \26861 );
buf \U$26520 ( \26863 , \26862 );
and \U$26521 ( \26864 , \26846 , \26863 );
not \U$26522 ( \26865 , \26846 );
not \U$26523 ( \26866 , \26863 );
and \U$26524 ( \26867 , \26865 , \26866 );
nor \U$26525 ( \26868 , \26864 , \26867 );
xor \U$26526 ( \26869 , \26811 , \26868 );
not \U$26527 ( \26870 , \26635 );
and \U$26528 ( \26871 , \26870 , \26661 );
and \U$26529 ( \26872 , \26651 , \26660 );
nor \U$26530 ( \26873 , \26871 , \26872 );
xnor \U$26531 ( \26874 , \13689 , \13559 );
not \U$26532 ( \26875 , \26874 );
not \U$26533 ( \26876 , \13448 );
not \U$26534 ( \26877 , \13519 );
or \U$26535 ( \26878 , \26876 , \26877 );
or \U$26536 ( \26879 , \13519 , \13448 );
nand \U$26537 ( \26880 , \26878 , \26879 );
not \U$26538 ( \26881 , \26880 );
or \U$26539 ( \26882 , \26875 , \26881 );
or \U$26540 ( \26883 , \26880 , \26874 );
nand \U$26541 ( \26884 , \26882 , \26883 );
not \U$26542 ( \26885 , \26638 );
not \U$26543 ( \26886 , \26645 );
or \U$26544 ( \26887 , \26885 , \26886 );
not \U$26545 ( \26888 , \26636 );
nand \U$26546 ( \26889 , \26888 , \26637 );
nand \U$26547 ( \26890 , \26887 , \26889 );
not \U$26548 ( \26891 , \26890 );
and \U$26549 ( \26892 , \26884 , \26891 );
not \U$26550 ( \26893 , \26884 );
and \U$26551 ( \26894 , \26893 , \26890 );
or \U$26552 ( \26895 , \26892 , \26894 );
not \U$26553 ( \26896 , \26895 );
nand \U$26554 ( \26897 , \26753 , \26743 );
not \U$26555 ( \26898 , \26897 );
and \U$26556 ( \26899 , \26745 , \26752 );
nor \U$26557 ( \26900 , \26898 , \26899 );
not \U$26558 ( \26901 , \26900 );
or \U$26559 ( \26902 , \26896 , \26901 );
not \U$26560 ( \26903 , \26899 );
not \U$26561 ( \26904 , \26903 );
not \U$26562 ( \26905 , \26897 );
or \U$26563 ( \26906 , \26904 , \26905 );
not \U$26564 ( \26907 , \26895 );
nand \U$26565 ( \26908 , \26906 , \26907 );
nand \U$26566 ( \26909 , \26902 , \26908 );
xor \U$26567 ( \26910 , \26873 , \26909 );
not \U$26568 ( \26911 , \26761 );
not \U$26569 ( \26912 , \26911 );
not \U$26570 ( \26913 , \26754 );
or \U$26571 ( \26914 , \26912 , \26913 );
not \U$26572 ( \26915 , \26754 );
not \U$26573 ( \26916 , \26915 );
not \U$26574 ( \26917 , \26761 );
or \U$26575 ( \26918 , \26916 , \26917 );
nand \U$26576 ( \26919 , \26918 , \26741 );
nand \U$26577 ( \26920 , \26914 , \26919 );
xnor \U$26578 ( \26921 , \26910 , \26920 );
xnor \U$26579 ( \26922 , \26869 , \26921 );
not \U$26580 ( \26923 , \26762 );
not \U$26581 ( \26924 , \26782 );
or \U$26582 ( \26925 , \26923 , \26924 );
nand \U$26583 ( \26926 , \26925 , \26769 );
not \U$26584 ( \26927 , \26762 );
nand \U$26585 ( \26928 , \26927 , \26779 );
nand \U$26586 ( \26929 , \26926 , \26928 );
and \U$26587 ( \26930 , \26922 , \26929 );
not \U$26588 ( \26931 , \26922 );
not \U$26589 ( \26932 , \26929 );
and \U$26590 ( \26933 , \26931 , \26932 );
nor \U$26591 ( \26934 , \26930 , \26933 );
not \U$26592 ( \26935 , \26734 );
not \U$26593 ( \26936 , \26784 );
or \U$26594 ( \26937 , \26935 , \26936 );
nand \U$26595 ( \26938 , \26937 , \26796 );
nand \U$26596 ( \26939 , \26938 , \26788 );
not \U$26597 ( \26940 , \26939 );
nand \U$26598 ( \26941 , \26934 , \26940 );
nor \U$26599 ( \26942 , \26854 , \26852 );
or \U$26600 ( \26943 , \26942 , \26861 );
nand \U$26601 ( \26944 , \26854 , \26852 );
nand \U$26602 ( \26945 , \26943 , \26944 );
not \U$26603 ( \26946 , \26945 );
xor \U$26604 ( \26947 , \14148 , \14149 );
xor \U$26605 ( \26948 , \26947 , \14246 );
not \U$26606 ( \26949 , \26948 );
or \U$26607 ( \26950 , \26946 , \26949 );
or \U$26608 ( \26951 , \26948 , \26945 );
and \U$26609 ( \26952 , \13969 , \13809 );
not \U$26610 ( \26953 , \13969 );
not \U$26611 ( \26954 , \13809 );
and \U$26612 ( \26955 , \26953 , \26954 );
nor \U$26613 ( \26956 , \26952 , \26955 );
nand \U$26614 ( \26957 , \26951 , \26956 );
nand \U$26615 ( \26958 , \26950 , \26957 );
not \U$26616 ( \26959 , \26958 );
and \U$26617 ( \26960 , \13542 , \13526 );
not \U$26618 ( \26961 , \13542 );
not \U$26619 ( \26962 , \13526 );
and \U$26620 ( \26963 , \26961 , \26962 );
nor \U$26621 ( \26964 , \26960 , \26963 );
not \U$26622 ( \26965 , \26890 );
not \U$26623 ( \26966 , \26884 );
or \U$26624 ( \26967 , \26965 , \26966 );
not \U$26625 ( \26968 , \26874 );
nand \U$26626 ( \26969 , \26968 , \26880 );
nand \U$26627 ( \26970 , \26967 , \26969 );
xor \U$26628 ( \26971 , \26964 , \26970 );
not \U$26629 ( \26972 , \26821 );
not \U$26630 ( \26973 , \26813 );
or \U$26631 ( \26974 , \26972 , \26973 );
not \U$26632 ( \26975 , \26813 );
nand \U$26633 ( \26976 , \26975 , \26824 );
nand \U$26634 ( \26977 , \26976 , \26831 );
nand \U$26635 ( \26978 , \26974 , \26977 );
and \U$26636 ( \26979 , \26971 , \26978 );
and \U$26637 ( \26980 , \26964 , \26970 );
or \U$26638 ( \26981 , \26979 , \26980 );
not \U$26639 ( \26982 , \26981 );
not \U$26640 ( \26983 , \13997 );
not \U$26641 ( \26984 , \14249 );
and \U$26642 ( \26985 , \26983 , \26984 );
and \U$26643 ( \26986 , \13997 , \14249 );
nor \U$26644 ( \26987 , \26985 , \26986 );
not \U$26645 ( \26988 , \26987 );
or \U$26646 ( \26989 , \26982 , \26988 );
or \U$26647 ( \26990 , \26987 , \26981 );
nand \U$26648 ( \26991 , \26989 , \26990 );
not \U$26649 ( \26992 , \26991 );
or \U$26650 ( \26993 , \26959 , \26992 );
not \U$26651 ( \26994 , \26987 );
nand \U$26652 ( \26995 , \26994 , \26981 );
nand \U$26653 ( \26996 , \26993 , \26995 );
not \U$26654 ( \26997 , \26996 );
and \U$26655 ( \26998 , \13715 , \13744 );
not \U$26656 ( \26999 , \13715 );
and \U$26657 ( \27000 , \26999 , \13717 );
nor \U$26658 ( \27001 , \26998 , \27000 );
xnor \U$26659 ( \27002 , \13741 , \27001 );
and \U$26660 ( \27003 , \26997 , \27002 );
not \U$26661 ( \27004 , \26997 );
not \U$26662 ( \27005 , \27002 );
and \U$26663 ( \27006 , \27004 , \27005 );
nor \U$26664 ( \27007 , \27003 , \27006 );
nand \U$26665 ( \27008 , \14261 , \14256 );
and \U$26666 ( \27009 , \27008 , \13982 );
not \U$26667 ( \27010 , \27008 );
not \U$26668 ( \27011 , \13982 );
and \U$26669 ( \27012 , \27010 , \27011 );
nor \U$26670 ( \27013 , \27009 , \27012 );
nand \U$26671 ( \27014 , \27007 , \27013 );
not \U$26672 ( \27015 , \27014 );
nand \U$26673 ( \27016 , \26997 , \27002 );
not \U$26674 ( \27017 , \27016 );
or \U$26675 ( \27018 , \27015 , \27017 );
not \U$26676 ( \27019 , \13796 );
not \U$26677 ( \27020 , \13794 );
not \U$26678 ( \27021 , \14262 );
not \U$26679 ( \27022 , \27021 );
or \U$26680 ( \27023 , \27020 , \27022 );
nand \U$26681 ( \27024 , \14262 , \13793 );
nand \U$26682 ( \27025 , \27023 , \27024 );
not \U$26683 ( \27026 , \27025 );
or \U$26684 ( \27027 , \27019 , \27026 );
or \U$26685 ( \27028 , \27025 , \13796 );
nand \U$26686 ( \27029 , \27027 , \27028 );
nand \U$26687 ( \27030 , \27018 , \27029 );
and \U$26688 ( \27031 , \26941 , \27030 );
or \U$26689 ( \27032 , \26843 , \26862 );
nand \U$26690 ( \27033 , \27032 , \26845 );
xor \U$26691 ( \27034 , \26964 , \26970 );
xor \U$26692 ( \27035 , \27034 , \26978 );
xor \U$26693 ( \27036 , \27033 , \27035 );
not \U$26694 ( \27037 , \26873 );
not \U$26695 ( \27038 , \27037 );
not \U$26696 ( \27039 , \26909 );
or \U$26697 ( \27040 , \27038 , \27039 );
not \U$26698 ( \27041 , \26903 );
not \U$26699 ( \27042 , \26897 );
or \U$26700 ( \27043 , \27041 , \27042 );
nand \U$26701 ( \27044 , \27043 , \26895 );
nand \U$26702 ( \27045 , \27040 , \27044 );
xor \U$26703 ( \27046 , \27036 , \27045 );
not \U$26704 ( \27047 , \27046 );
xor \U$26705 ( \27048 , \26945 , \26948 );
xor \U$26706 ( \27049 , \27048 , \26956 );
not \U$26707 ( \27050 , \27049 );
not \U$26708 ( \27051 , \27050 );
not \U$26709 ( \27052 , \26811 );
not \U$26710 ( \27053 , \26921 );
or \U$26711 ( \27054 , \27052 , \27053 );
xor \U$26712 ( \27055 , \26909 , \27037 );
buf \U$26713 ( \27056 , \26920 );
nand \U$26714 ( \27057 , \27055 , \27056 );
nand \U$26715 ( \27058 , \27054 , \27057 );
not \U$26716 ( \27059 , \27058 );
or \U$26717 ( \27060 , \27051 , \27059 );
or \U$26718 ( \27061 , \27050 , \27058 );
nand \U$26719 ( \27062 , \27060 , \27061 );
not \U$26720 ( \27063 , \27062 );
or \U$26721 ( \27064 , \27047 , \27063 );
nand \U$26722 ( \27065 , \27058 , \27049 );
nand \U$26723 ( \27066 , \27064 , \27065 );
not \U$26724 ( \27067 , \13800 );
and \U$26725 ( \27068 , \13978 , \27067 );
not \U$26726 ( \27069 , \13978 );
and \U$26727 ( \27070 , \27069 , \13800 );
nor \U$26728 ( \27071 , \27068 , \27070 );
xor \U$26729 ( \27072 , \26981 , \26958 );
xor \U$26730 ( \27073 , \27072 , \26987 );
xor \U$26731 ( \27074 , \27071 , \27073 );
xor \U$26732 ( \27075 , \27035 , \27045 );
buf \U$26733 ( \27076 , \27033 );
and \U$26734 ( \27077 , \27075 , \27076 );
and \U$26735 ( \27078 , \27035 , \27045 );
nor \U$26736 ( \27079 , \27077 , \27078 );
xnor \U$26737 ( \27080 , \27074 , \27079 );
nor \U$26738 ( \27081 , \27066 , \27080 );
not \U$26739 ( \27082 , \27081 );
xor \U$26740 ( \27083 , \27049 , \27046 );
xor \U$26741 ( \27084 , \27083 , \27058 );
not \U$26742 ( \27085 , \27084 );
not \U$26743 ( \27086 , \26811 );
xnor \U$26744 ( \27087 , \26921 , \27086 );
buf \U$26745 ( \27088 , \26868 );
or \U$26746 ( \27089 , \27087 , \27088 );
nand \U$26747 ( \27090 , \27089 , \26929 );
nand \U$26748 ( \27091 , \27087 , \27088 );
nand \U$26749 ( \27092 , \27090 , \27091 );
not \U$26750 ( \27093 , \27092 );
nand \U$26751 ( \27094 , \27085 , \27093 );
xor \U$26752 ( \27095 , \27013 , \27007 );
or \U$26753 ( \27096 , \27073 , \27071 );
not \U$26754 ( \27097 , \27096 );
not \U$26755 ( \27098 , \27079 );
or \U$26756 ( \27099 , \27097 , \27098 );
nand \U$26757 ( \27100 , \27073 , \27071 );
nand \U$26758 ( \27101 , \27099 , \27100 );
nand \U$26759 ( \27102 , \27095 , \27101 );
nand \U$26760 ( \27103 , \27031 , \27082 , \27094 , \27102 );
nor \U$26761 ( \27104 , \26807 , \27103 );
nand \U$26762 ( \27105 , \25956 , \27104 );
not \U$26763 ( \27106 , \25069 );
xor \U$26764 ( \27107 , \25321 , \27106 );
xnor \U$26765 ( \27108 , \27107 , \25550 );
not \U$26766 ( \27109 , \27108 );
not \U$26767 ( \27110 , \25692 );
or \U$26768 ( \27111 , \27109 , \27110 );
or \U$26769 ( \27112 , \25692 , \27108 );
nand \U$26770 ( \27113 , \27111 , \27112 );
buf \U$26771 ( \27114 , \27113 );
xor \U$26772 ( \27115 , \25152 , \25286 );
xor \U$26773 ( \27116 , \27115 , \25149 );
xor \U$26774 ( \27117 , \25541 , \25543 );
xnor \U$26775 ( \27118 , \27117 , \25547 );
nand \U$26776 ( \27119 , \27116 , \27118 );
not \U$26777 ( \27120 , \27119 );
not \U$26778 ( \27121 , \18508 );
and \U$26779 ( \27122 , \1603 , \24305 );
not \U$26780 ( \27123 , \1603 );
and \U$26781 ( \27124 , \27123 , RI9873288_184);
nor \U$26782 ( \27125 , \27122 , \27124 );
not \U$26783 ( \27126 , \27125 );
or \U$26784 ( \27127 , \27121 , \27126 );
nand \U$26785 ( \27128 , \25528 , \17528 );
nand \U$26786 ( \27129 , \27127 , \27128 );
not \U$26787 ( \27130 , \27129 );
not \U$26788 ( \27131 , \18562 );
xor \U$26789 ( \27132 , \9694 , \3568 );
not \U$26790 ( \27133 , \27132 );
or \U$26791 ( \27134 , \27131 , \27133 );
nand \U$26792 ( \27135 , \25504 , \10332 );
nand \U$26793 ( \27136 , \27134 , \27135 );
not \U$26794 ( \27137 , \27136 );
not \U$26795 ( \27138 , \27137 );
not \U$26796 ( \27139 , \13214 );
not \U$26797 ( \27140 , \25577 );
or \U$26798 ( \27141 , \27139 , \27140 );
and \U$26799 ( \27142 , RI9872f40_177, \3859 );
not \U$26800 ( \27143 , RI9872f40_177);
and \U$26801 ( \27144 , \27143 , \3860 );
or \U$26802 ( \27145 , \27142 , \27144 );
nand \U$26803 ( \27146 , \27145 , \9526 );
nand \U$26804 ( \27147 , \27141 , \27146 );
not \U$26805 ( \27148 , \27147 );
or \U$26806 ( \27149 , \27138 , \27148 );
or \U$26807 ( \27150 , \27147 , \27137 );
nand \U$26808 ( \27151 , \27149 , \27150 );
not \U$26809 ( \27152 , \27151 );
or \U$26810 ( \27153 , \27130 , \27152 );
not \U$26811 ( \27154 , \27137 );
nand \U$26812 ( \27155 , \27154 , \27147 );
nand \U$26813 ( \27156 , \27153 , \27155 );
not \U$26814 ( \27157 , \13020 );
not \U$26815 ( \27158 , RI98730a8_180);
not \U$26816 ( \27159 , \5946 );
or \U$26817 ( \27160 , \27158 , \27159 );
or \U$26818 ( \27161 , \1191 , RI98730a8_180);
nand \U$26819 ( \27162 , \27160 , \27161 );
not \U$26820 ( \27163 , \27162 );
or \U$26821 ( \27164 , \27157 , \27163 );
nand \U$26822 ( \27165 , \25649 , \17347 );
nand \U$26823 ( \27166 , \27164 , \27165 );
not \U$26824 ( \27167 , \27166 );
not \U$26825 ( \27168 , \9214 );
not \U$26826 ( \27169 , \25610 );
or \U$26827 ( \27170 , \27168 , \27169 );
not \U$26828 ( \27171 , \9198 );
not \U$26829 ( \27172 , \5393 );
or \U$26830 ( \27173 , \27171 , \27172 );
nand \U$26831 ( \27174 , \5776 , RI9872b80_169);
nand \U$26832 ( \27175 , \27173 , \27174 );
nand \U$26833 ( \27176 , \27175 , \9196 );
nand \U$26834 ( \27177 , \27170 , \27176 );
not \U$26835 ( \27178 , \27177 );
nand \U$26836 ( \27179 , \25835 , \17263 );
not \U$26837 ( \27180 , \27179 );
not \U$26838 ( \27181 , \5720 );
not \U$26839 ( \27182 , RI98733f0_187);
and \U$26840 ( \27183 , \27181 , \27182 );
and \U$26841 ( \27184 , \1253 , RI98733f0_187);
nor \U$26842 ( \27185 , \27183 , \27184 );
not \U$26843 ( \27186 , \17251 );
nor \U$26844 ( \27187 , \27185 , \27186 );
nor \U$26845 ( \27188 , \27180 , \27187 );
not \U$26846 ( \27189 , \27188 );
or \U$26847 ( \27190 , \27178 , \27189 );
not \U$26848 ( \27191 , \27185 );
nand \U$26849 ( \27192 , \27191 , \17252 );
not \U$26850 ( \27193 , \27192 );
not \U$26851 ( \27194 , \27179 );
or \U$26852 ( \27195 , \27193 , \27194 );
not \U$26853 ( \27196 , \27177 );
nand \U$26854 ( \27197 , \27195 , \27196 );
nand \U$26855 ( \27198 , \27190 , \27197 );
not \U$26856 ( \27199 , \27198 );
or \U$26857 ( \27200 , \27167 , \27199 );
not \U$26858 ( \27201 , \27192 );
not \U$26859 ( \27202 , \27179 );
or \U$26860 ( \27203 , \27201 , \27202 );
nand \U$26861 ( \27204 , \27203 , \27177 );
nand \U$26862 ( \27205 , \27200 , \27204 );
xor \U$26863 ( \27206 , \27156 , \27205 );
not \U$26864 ( \27207 , \18615 );
not \U$26865 ( \27208 , RI9873558_190);
not \U$26866 ( \27209 , \1505 );
or \U$26867 ( \27210 , \27208 , \27209 );
not \U$26868 ( \27211 , \892 );
nand \U$26869 ( \27212 , \27211 , \18239 );
nand \U$26870 ( \27213 , \27210 , \27212 );
not \U$26871 ( \27214 , \27213 );
or \U$26872 ( \27215 , \27207 , \27214 );
nand \U$26873 ( \27216 , \25840 , RI9873648_192);
nand \U$26874 ( \27217 , \27215 , \27216 );
not \U$26875 ( \27218 , \9937 );
not \U$26876 ( \27219 , \25662 );
or \U$26877 ( \27220 , \27218 , \27219 );
and \U$26878 ( \27221 , RI9873030_179, \2111 );
not \U$26879 ( \27222 , RI9873030_179);
and \U$26880 ( \27223 , \27222 , \6378 );
nor \U$26881 ( \27224 , \27221 , \27223 );
nand \U$26882 ( \27225 , \27224 , \9952 );
nand \U$26883 ( \27226 , \27220 , \27225 );
xor \U$26884 ( \27227 , \27217 , \27226 );
xnor \U$26885 ( \27228 , \25417 , \25388 );
not \U$26886 ( \27229 , \27228 );
and \U$26887 ( \27230 , \27227 , \27229 );
and \U$26888 ( \27231 , \27217 , \27226 );
or \U$26889 ( \27232 , \27230 , \27231 );
and \U$26890 ( \27233 , \27206 , \27232 );
and \U$26891 ( \27234 , \27156 , \27205 );
or \U$26892 ( \27235 , \27233 , \27234 );
not \U$26893 ( \27236 , \27235 );
not \U$26894 ( \27237 , \5642 );
xnor \U$26895 ( \27238 , \8074 , RI9872568_156);
not \U$26896 ( \27239 , \27238 );
or \U$26897 ( \27240 , \27237 , \27239 );
nand \U$26898 ( \27241 , \25474 , \5653 );
nand \U$26899 ( \27242 , \27240 , \27241 );
not \U$26900 ( \27243 , \7325 );
not \U$26901 ( \27244 , \7333 );
not \U$26902 ( \27245 , \7905 );
or \U$26903 ( \27246 , \27244 , \27245 );
nand \U$26904 ( \27247 , \15875 , RI98729a0_165);
nand \U$26905 ( \27248 , \27246 , \27247 );
not \U$26906 ( \27249 , \27248 );
or \U$26907 ( \27250 , \27243 , \27249 );
nand \U$26908 ( \27251 , \25367 , \7338 );
nand \U$26909 ( \27252 , \27250 , \27251 );
xor \U$26910 ( \27253 , \27242 , \27252 );
not \U$26911 ( \27254 , \8029 );
not \U$26912 ( \27255 , \15389 );
not \U$26913 ( \27256 , \7108 );
or \U$26914 ( \27257 , \27255 , \27256 );
nand \U$26915 ( \27258 , \6308 , RI9872a18_166);
nand \U$26916 ( \27259 , \27257 , \27258 );
not \U$26917 ( \27260 , \27259 );
or \U$26918 ( \27261 , \27254 , \27260 );
or \U$26919 ( \27262 , \25638 , \8040 );
nand \U$26920 ( \27263 , \27261 , \27262 );
and \U$26921 ( \27264 , \27253 , \27263 );
and \U$26922 ( \27265 , \27242 , \27252 );
or \U$26923 ( \27266 , \27264 , \27265 );
not \U$26924 ( \27267 , \27266 );
xor \U$26925 ( \27268 , \25230 , \25236 );
xor \U$26926 ( \27269 , \27268 , \25246 );
xor \U$26927 ( \27270 , \25351 , \27269 );
not \U$26928 ( \27271 , \25373 );
xnor \U$26929 ( \27272 , \27270 , \27271 );
not \U$26930 ( \27273 , \27272 );
or \U$26931 ( \27274 , \27267 , \27273 );
buf \U$26932 ( \27275 , \27271 );
xnor \U$26933 ( \27276 , \27275 , \25351 );
nand \U$26934 ( \27277 , \27276 , \27269 );
nand \U$26935 ( \27278 , \27274 , \27277 );
not \U$26936 ( \27279 , \27278 );
not \U$26937 ( \27280 , \25264 );
not \U$26938 ( \27281 , \25253 );
not \U$26939 ( \27282 , \27281 );
and \U$26940 ( \27283 , \27280 , \27282 );
and \U$26941 ( \27284 , \25264 , \27281 );
nor \U$26942 ( \27285 , \27283 , \27284 );
and \U$26943 ( \27286 , \27279 , \27285 );
not \U$26944 ( \27287 , \27279 );
not \U$26945 ( \27288 , \27285 );
and \U$26946 ( \27289 , \27287 , \27288 );
nor \U$26947 ( \27290 , \27286 , \27289 );
not \U$26948 ( \27291 , \27290 );
or \U$26949 ( \27292 , \27236 , \27291 );
not \U$26950 ( \27293 , \27279 );
nand \U$26951 ( \27294 , \27293 , \27288 );
nand \U$26952 ( \27295 , \27292 , \27294 );
not \U$26953 ( \27296 , \27295 );
xor \U$26954 ( \27297 , \25421 , \25431 );
xor \U$26955 ( \27298 , \27297 , \25442 );
not \U$26956 ( \27299 , \9249 );
not \U$26957 ( \27300 , RI9872bf8_170);
not \U$26958 ( \27301 , \7007 );
or \U$26959 ( \27302 , \27300 , \27301 );
or \U$26960 ( \27303 , \23391 , RI9872bf8_170);
nand \U$26961 ( \27304 , \27302 , \27303 );
not \U$26962 ( \27305 , \27304 );
or \U$26963 ( \27306 , \27299 , \27305 );
nand \U$26964 ( \27307 , \25620 , \9227 );
nand \U$26965 ( \27308 , \27306 , \27307 );
not \U$26966 ( \27309 , \8802 );
not \U$26967 ( \27310 , \25513 );
or \U$26968 ( \27311 , \27309 , \27310 );
not \U$26969 ( \27312 , RI9872d60_173);
not \U$26970 ( \27313 , \5205 );
or \U$26971 ( \27314 , \27312 , \27313 );
or \U$26972 ( \27315 , \4408 , RI9872d60_173);
nand \U$26973 ( \27316 , \27314 , \27315 );
nand \U$26974 ( \27317 , \27316 , \8819 );
nand \U$26975 ( \27318 , \27311 , \27317 );
xor \U$26976 ( \27319 , \27308 , \27318 );
not \U$26977 ( \27320 , \17243 );
and \U$26978 ( \27321 , \6334 , \22675 );
not \U$26979 ( \27322 , \6334 );
and \U$26980 ( \27323 , \27322 , RI9873210_183);
or \U$26981 ( \27324 , \27321 , \27323 );
not \U$26982 ( \27325 , \27324 );
or \U$26983 ( \27326 , \27320 , \27325 );
nand \U$26984 ( \27327 , \25627 , \22670 );
nand \U$26985 ( \27328 , \27326 , \27327 );
and \U$26986 ( \27329 , \27319 , \27328 );
and \U$26987 ( \27330 , \27308 , \27318 );
or \U$26988 ( \27331 , \27329 , \27330 );
xor \U$26989 ( \27332 , \27298 , \27331 );
xor \U$26990 ( \27333 , \25455 , \25476 );
xor \U$26991 ( \27334 , \27333 , \25466 );
and \U$26992 ( \27335 , \27332 , \27334 );
and \U$26993 ( \27336 , \27298 , \27331 );
or \U$26994 ( \27337 , \27335 , \27336 );
not \U$26995 ( \27338 , \27337 );
xor \U$26996 ( \27339 , \25445 , \25378 );
xnor \U$26997 ( \27340 , \27339 , \25485 );
nand \U$26998 ( \27341 , \27338 , \27340 );
not \U$26999 ( \27342 , \27341 );
and \U$27000 ( \27343 , \25564 , \25567 );
not \U$27001 ( \27344 , \25564 );
and \U$27002 ( \27345 , \27344 , \25568 );
nor \U$27003 ( \27346 , \27343 , \27345 );
xor \U$27004 ( \27347 , \27346 , \25597 );
not \U$27005 ( \27348 , \27347 );
or \U$27006 ( \27349 , \27342 , \27348 );
not \U$27007 ( \27350 , \27340 );
nand \U$27008 ( \27351 , \27350 , \27337 );
nand \U$27009 ( \27352 , \27349 , \27351 );
not \U$27010 ( \27353 , \27352 );
or \U$27011 ( \27354 , \27296 , \27353 );
not \U$27012 ( \27355 , \27352 );
not \U$27013 ( \27356 , \27355 );
not \U$27014 ( \27357 , \27295 );
not \U$27015 ( \27358 , \27357 );
or \U$27016 ( \27359 , \27356 , \27358 );
xor \U$27017 ( \27360 , \25496 , \25532 );
xor \U$27018 ( \27361 , \25530 , \25506 );
xor \U$27019 ( \27362 , \27361 , \25517 );
not \U$27020 ( \27363 , \27362 );
xor \U$27021 ( \27364 , \25879 , \25837 );
not \U$27022 ( \27365 , \25183 );
or \U$27023 ( \27366 , \27365 , \1494 );
and \U$27024 ( \27367 , \17862 , RI9871c80_137);
not \U$27025 ( \27368 , \17862 );
and \U$27026 ( \27369 , \27368 , \1584 );
nor \U$27027 ( \27370 , \27367 , \27369 );
not \U$27028 ( \27371 , \27370 );
or \U$27029 ( \27372 , \27371 , \1499 );
nand \U$27030 ( \27373 , \27366 , \27372 );
not \U$27031 ( \27374 , \27373 );
not \U$27032 ( \27375 , \25398 );
not \U$27033 ( \27376 , \25403 );
and \U$27034 ( \27377 , \27375 , \27376 );
and \U$27035 ( \27378 , \25398 , \25403 );
nor \U$27036 ( \27379 , \27377 , \27378 );
not \U$27037 ( \27380 , \27379 );
or \U$27038 ( \27381 , \27374 , \27380 );
or \U$27039 ( \27382 , \27373 , \27379 );
nand \U$27040 ( \27383 , \27381 , \27382 );
not \U$27041 ( \27384 , \25414 );
or \U$27042 ( \27385 , \27384 , \1543 );
xor \U$27043 ( \27386 , \16995 , RI9871b18_134);
not \U$27044 ( \27387 , \27386 );
or \U$27045 ( \27388 , \27387 , \1293 );
nand \U$27046 ( \27389 , \27385 , \27388 );
and \U$27047 ( \27390 , \27383 , \27389 );
not \U$27048 ( \27391 , \27379 );
and \U$27049 ( \27392 , \27391 , \27373 );
nor \U$27050 ( \27393 , \27390 , \27392 );
not \U$27051 ( \27394 , \27393 );
not \U$27052 ( \27395 , \6284 );
not \U$27053 ( \27396 , \7049 );
not \U$27054 ( \27397 , \7467 );
or \U$27055 ( \27398 , \27396 , \27397 );
nand \U$27056 ( \27399 , \17440 , RI98728b0_163);
nand \U$27057 ( \27400 , \27398 , \27399 );
not \U$27058 ( \27401 , \27400 );
or \U$27059 ( \27402 , \27395 , \27401 );
nand \U$27060 ( \27403 , \25464 , \6610 );
nand \U$27061 ( \27404 , \27402 , \27403 );
not \U$27062 ( \27405 , \27404 );
or \U$27063 ( \27406 , \27394 , \27405 );
or \U$27064 ( \27407 , \27404 , \27393 );
nand \U$27065 ( \27408 , \27406 , \27407 );
not \U$27066 ( \27409 , \27408 );
not \U$27067 ( \27410 , \20147 );
not \U$27068 ( \27411 , \25589 );
or \U$27069 ( \27412 , \27410 , \27411 );
not \U$27070 ( \27413 , RI98734e0_189);
not \U$27071 ( \27414 , \6224 );
or \U$27072 ( \27415 , \27413 , \27414 );
or \U$27073 ( \27416 , \18737 , RI98734e0_189);
nand \U$27074 ( \27417 , \27415 , \27416 );
nand \U$27075 ( \27418 , \27417 , \19036 );
nand \U$27076 ( \27419 , \27412 , \27418 );
not \U$27077 ( \27420 , \27419 );
or \U$27078 ( \27421 , \27409 , \27420 );
not \U$27079 ( \27422 , \27393 );
nand \U$27080 ( \27423 , \27422 , \27404 );
nand \U$27081 ( \27424 , \27421 , \27423 );
xor \U$27082 ( \27425 , \27364 , \27424 );
not \U$27083 ( \27426 , \27425 );
or \U$27084 ( \27427 , \27363 , \27426 );
nand \U$27085 ( \27428 , \27424 , \27364 );
nand \U$27086 ( \27429 , \27427 , \27428 );
xor \U$27087 ( \27430 , \27360 , \27429 );
xor \U$27088 ( \27431 , \25612 , \25629 );
xor \U$27089 ( \27432 , \27431 , \25622 );
not \U$27090 ( \27433 , \27432 );
xor \U$27091 ( \27434 , \25641 , \25652 );
xnor \U$27092 ( \27435 , \27434 , \25664 );
xor \U$27093 ( \27436 , \25579 , \25582 );
xnor \U$27094 ( \27437 , \27436 , \25591 );
xnor \U$27095 ( \27438 , \27435 , \27437 );
not \U$27096 ( \27439 , \27438 );
or \U$27097 ( \27440 , \27433 , \27439 );
not \U$27098 ( \27441 , \27435 );
nand \U$27099 ( \27442 , \27437 , \27441 );
nand \U$27100 ( \27443 , \27440 , \27442 );
and \U$27101 ( \27444 , \27430 , \27443 );
and \U$27102 ( \27445 , \27360 , \27429 );
or \U$27103 ( \27446 , \27444 , \27445 );
nand \U$27104 ( \27447 , \27359 , \27446 );
nand \U$27105 ( \27448 , \27354 , \27447 );
not \U$27106 ( \27449 , \27448 );
or \U$27107 ( \27450 , \27120 , \27449 );
not \U$27108 ( \27451 , \27118 );
not \U$27109 ( \27452 , \27116 );
nand \U$27110 ( \27453 , \27451 , \27452 );
nand \U$27111 ( \27454 , \27450 , \27453 );
not \U$27112 ( \27455 , \27454 );
nand \U$27113 ( \27456 , \27114 , \27455 );
not \U$27114 ( \27457 , \27456 );
xor \U$27115 ( \27458 , \25818 , \25913 );
not \U$27116 ( \27459 , \27458 );
xor \U$27117 ( \27460 , \25684 , \25677 );
xnor \U$27118 ( \27461 , \27460 , \25687 );
not \U$27119 ( \27462 , \25491 );
nand \U$27120 ( \27463 , \27462 , \25537 );
not \U$27121 ( \27464 , \27463 );
not \U$27122 ( \27465 , \25535 );
and \U$27123 ( \27466 , \27464 , \27465 );
and \U$27124 ( \27467 , \27463 , \25535 );
nor \U$27125 ( \27468 , \27466 , \27467 );
nor \U$27126 ( \27469 , \27461 , \27468 );
xor \U$27127 ( \27470 , \25902 , \25899 );
xor \U$27128 ( \27471 , \27470 , \25901 );
or \U$27129 ( \27472 , \27469 , \27471 );
nand \U$27130 ( \27473 , \27461 , \27468 );
nand \U$27131 ( \27474 , \27472 , \27473 );
not \U$27132 ( \27475 , \27474 );
xor \U$27133 ( \27476 , \24981 , \25560 );
not \U$27134 ( \27477 , \25065 );
not \U$27135 ( \27478 , \24984 );
and \U$27136 ( \27479 , \27477 , \27478 );
and \U$27137 ( \27480 , \25554 , \24984 );
nor \U$27138 ( \27481 , \27479 , \27480 );
xnor \U$27139 ( \27482 , \27476 , \27481 );
xor \U$27140 ( \27483 , \27482 , \25689 );
nand \U$27141 ( \27484 , \27475 , \27483 );
not \U$27142 ( \27485 , \27484 );
or \U$27143 ( \27486 , \27459 , \27485 );
not \U$27144 ( \27487 , \27483 );
nand \U$27145 ( \27488 , \27487 , \27474 );
nand \U$27146 ( \27489 , \27486 , \27488 );
not \U$27147 ( \27490 , \27489 );
or \U$27148 ( \27491 , \27457 , \27490 );
not \U$27149 ( \27492 , \27114 );
nand \U$27150 ( \27493 , \27492 , \27454 );
nand \U$27151 ( \27494 , \27491 , \27493 );
xor \U$27152 ( \27495 , \25139 , \25146 );
xnor \U$27153 ( \27496 , \27495 , \25311 );
xor \U$27154 ( \27497 , \27494 , \27496 );
xor \U$27155 ( \27498 , \25925 , \25701 );
xor \U$27156 ( \27499 , \27497 , \27498 );
not \U$27157 ( \27500 , \27499 );
xor \U$27158 ( \27501 , \27235 , \27290 );
not \U$27159 ( \27502 , \27501 );
not \U$27160 ( \27503 , \27502 );
xor \U$27161 ( \27504 , \27156 , \27205 );
xor \U$27162 ( \27505 , \27504 , \27232 );
not \U$27163 ( \27506 , \27505 );
not \U$27164 ( \27507 , \27151 );
not \U$27165 ( \27508 , \27129 );
not \U$27166 ( \27509 , \27508 );
and \U$27167 ( \27510 , \27507 , \27509 );
and \U$27168 ( \27511 , \27151 , \27508 );
nor \U$27169 ( \27512 , \27510 , \27511 );
not \U$27170 ( \27513 , \27512 );
not \U$27171 ( \27514 , \27513 );
xor \U$27172 ( \27515 , \27308 , \27318 );
xor \U$27173 ( \27516 , \27515 , \27328 );
not \U$27174 ( \27517 , \27516 );
or \U$27175 ( \27518 , \27514 , \27517 );
not \U$27176 ( \27519 , \27516 );
not \U$27177 ( \27520 , \27519 );
not \U$27178 ( \27521 , \27512 );
or \U$27179 ( \27522 , \27520 , \27521 );
buf \U$27180 ( \27523 , \18704 );
and \U$27181 ( \27524 , \27523 , \924 );
not \U$27182 ( \27525 , \1493 );
not \U$27183 ( \27526 , \27370 );
or \U$27184 ( \27527 , \27525 , \27526 );
and \U$27185 ( \27528 , \18194 , RI9871c80_137);
and \U$27186 ( \27529 , \25166 , \1800 );
nor \U$27187 ( \27530 , \27528 , \27529 );
or \U$27188 ( \27531 , \27530 , \1499 );
nand \U$27189 ( \27532 , \27527 , \27531 );
xor \U$27190 ( \27533 , \27524 , \27532 );
not \U$27191 ( \27534 , \1290 );
not \U$27192 ( \27535 , \27386 );
or \U$27193 ( \27536 , \27534 , \27535 );
not \U$27194 ( \27537 , \1283 );
not \U$27195 ( \27538 , \17702 );
or \U$27196 ( \27539 , \27537 , \27538 );
not \U$27197 ( \27540 , \1283 );
not \U$27198 ( \27541 , \17702 );
nand \U$27199 ( \27542 , \27540 , \27541 );
nand \U$27200 ( \27543 , \27539 , \27542 );
nand \U$27201 ( \27544 , \27543 , \1291 );
nand \U$27202 ( \27545 , \27536 , \27544 );
and \U$27203 ( \27546 , \27533 , \27545 );
and \U$27204 ( \27547 , \27524 , \27532 );
nor \U$27205 ( \27548 , \27546 , \27547 );
not \U$27206 ( \27549 , \1429 );
not \U$27207 ( \27550 , \25384 );
or \U$27208 ( \27551 , \27549 , \27550 );
not \U$27209 ( \27552 , \1850 );
not \U$27210 ( \27553 , \17744 );
or \U$27211 ( \27554 , \27552 , \27553 );
nand \U$27212 ( \27555 , \21529 , RI9871c08_136);
nand \U$27213 ( \27556 , \27554 , \27555 );
nand \U$27214 ( \27557 , \27556 , \1455 );
nand \U$27215 ( \27558 , \27551 , \27557 );
xnor \U$27216 ( \27559 , \27548 , \27558 );
not \U$27217 ( \27560 , \2071 );
and \U$27218 ( \27561 , RI9871aa0_133, \12784 );
not \U$27219 ( \27562 , RI9871aa0_133);
and \U$27220 ( \27563 , \27562 , \13601 );
or \U$27221 ( \27564 , \27561 , \27563 );
not \U$27222 ( \27565 , \27564 );
or \U$27223 ( \27566 , \27560 , \27565 );
nand \U$27224 ( \27567 , \25863 , \2087 );
nand \U$27225 ( \27568 , \27566 , \27567 );
xnor \U$27226 ( \27569 , \27559 , \27568 );
not \U$27227 ( \27570 , \27569 );
not \U$27228 ( \27571 , \2072 );
not \U$27229 ( \27572 , \13268 );
xor \U$27230 ( \27573 , \27572 , RI9871aa0_133);
not \U$27231 ( \27574 , \27573 );
or \U$27232 ( \27575 , \27571 , \27574 );
nand \U$27233 ( \27576 , \27564 , \2087 );
nand \U$27234 ( \27577 , \27575 , \27576 );
not \U$27235 ( \27578 , \27577 );
xor \U$27236 ( \27579 , \27524 , \27532 );
xor \U$27237 ( \27580 , \27579 , \27545 );
not \U$27238 ( \27581 , \27580 );
and \U$27239 ( \27582 , \3154 , \17756 );
not \U$27240 ( \27583 , \3154 );
and \U$27241 ( \27584 , \27583 , \20302 );
nor \U$27242 ( \27585 , \27582 , \27584 );
nand \U$27243 ( \27586 , \27585 , \3170 );
not \U$27244 ( \27587 , \10063 );
not \U$27245 ( \27588 , \27587 );
and \U$27246 ( \27589 , RI9872310_151, \27588 );
not \U$27247 ( \27590 , RI9872310_151);
and \U$27248 ( \27591 , \27590 , \11358 );
or \U$27249 ( \27592 , \27589 , \27591 );
nand \U$27250 ( \27593 , \27592 , \3163 );
and \U$27251 ( \27594 , \27586 , \27593 );
not \U$27252 ( \27595 , \27594 );
or \U$27253 ( \27596 , \27581 , \27595 );
not \U$27254 ( \27597 , \27586 );
not \U$27255 ( \27598 , \27593 );
or \U$27256 ( \27599 , \27597 , \27598 );
not \U$27257 ( \27600 , \27580 );
nand \U$27258 ( \27601 , \27599 , \27600 );
nand \U$27259 ( \27602 , \27596 , \27601 );
not \U$27260 ( \27603 , \27602 );
or \U$27261 ( \27604 , \27578 , \27603 );
not \U$27262 ( \27605 , \27586 );
not \U$27263 ( \27606 , \27593 );
or \U$27264 ( \27607 , \27605 , \27606 );
nand \U$27265 ( \27608 , \27607 , \27580 );
nand \U$27266 ( \27609 , \27604 , \27608 );
not \U$27267 ( \27610 , \27609 );
or \U$27268 ( \27611 , \27570 , \27610 );
or \U$27269 ( \27612 , \27609 , \27569 );
nand \U$27270 ( \27613 , \27611 , \27612 );
not \U$27271 ( \27614 , \27613 );
nand \U$27272 ( \27615 , \27213 , RI9873648_192);
and \U$27273 ( \27616 , RI9873558_190, \820 );
not \U$27274 ( \27617 , RI9873558_190);
and \U$27275 ( \27618 , \27617 , \8005 );
or \U$27276 ( \27619 , \27616 , \27618 );
nand \U$27277 ( \27620 , \27619 , \18615 );
nand \U$27278 ( \27621 , \27615 , \27620 );
not \U$27279 ( \27622 , \27621 );
or \U$27280 ( \27623 , \27614 , \27622 );
not \U$27281 ( \27624 , \27569 );
nand \U$27282 ( \27625 , \27624 , \27609 );
nand \U$27283 ( \27626 , \27623 , \27625 );
nand \U$27284 ( \27627 , \27522 , \27626 );
nand \U$27285 ( \27628 , \27518 , \27627 );
xor \U$27286 ( \27629 , \25775 , \25765 );
xor \U$27287 ( \27630 , \27629 , \25784 );
not \U$27288 ( \27631 , \9214 );
not \U$27289 ( \27632 , \27175 );
or \U$27290 ( \27633 , \27631 , \27632 );
xnor \U$27291 ( \27634 , \6481 , RI9872b80_169);
nand \U$27292 ( \27635 , \27634 , \9196 );
nand \U$27293 ( \27636 , \27633 , \27635 );
not \U$27294 ( \27637 , \9227 );
not \U$27295 ( \27638 , \27304 );
or \U$27296 ( \27639 , \27637 , \27638 );
xor \U$27297 ( \27640 , \5739 , RI9872bf8_170);
nand \U$27298 ( \27641 , \27640 , \9249 );
nand \U$27299 ( \27642 , \27639 , \27641 );
xor \U$27300 ( \27643 , \27636 , \27642 );
not \U$27301 ( \27644 , \13484 );
not \U$27302 ( \27645 , \27324 );
or \U$27303 ( \27646 , \27644 , \27645 );
and \U$27304 ( \27647 , \18012 , \3127 );
not \U$27305 ( \27648 , \18012 );
and \U$27306 ( \27649 , \27648 , \14032 );
nor \U$27307 ( \27650 , \27647 , \27649 );
nand \U$27308 ( \27651 , \27650 , \17243 );
nand \U$27309 ( \27652 , \27646 , \27651 );
and \U$27310 ( \27653 , \27643 , \27652 );
and \U$27311 ( \27654 , \27636 , \27642 );
or \U$27312 ( \27655 , \27653 , \27654 );
xor \U$27313 ( \27656 , \27630 , \27655 );
xor \U$27314 ( \27657 , \27228 , \27226 );
xnor \U$27315 ( \27658 , \27657 , \27217 );
and \U$27316 ( \27659 , \27656 , \27658 );
and \U$27317 ( \27660 , \27630 , \27655 );
or \U$27318 ( \27661 , \27659 , \27660 );
xor \U$27319 ( \27662 , \27628 , \27661 );
not \U$27320 ( \27663 , \27662 );
or \U$27321 ( \27664 , \27506 , \27663 );
nand \U$27322 ( \27665 , \27661 , \27628 );
nand \U$27323 ( \27666 , \27664 , \27665 );
not \U$27324 ( \27667 , \27666 );
not \U$27325 ( \27668 , \27667 );
or \U$27326 ( \27669 , \27503 , \27668 );
xor \U$27327 ( \27670 , \27360 , \27429 );
xor \U$27328 ( \27671 , \27670 , \27443 );
nand \U$27329 ( \27672 , \27669 , \27671 );
not \U$27330 ( \27673 , \27502 );
nand \U$27331 ( \27674 , \27673 , \27666 );
nand \U$27332 ( \27675 , \27672 , \27674 );
not \U$27333 ( \27676 , \27352 );
not \U$27334 ( \27677 , \27357 );
or \U$27335 ( \27678 , \27676 , \27677 );
nand \U$27336 ( \27679 , \27295 , \27355 );
nand \U$27337 ( \27680 , \27678 , \27679 );
and \U$27338 ( \27681 , \27680 , \27446 );
not \U$27339 ( \27682 , \27680 );
not \U$27340 ( \27683 , \27446 );
and \U$27341 ( \27684 , \27682 , \27683 );
nor \U$27342 ( \27685 , \27681 , \27684 );
nor \U$27343 ( \27686 , \27675 , \27685 );
not \U$27344 ( \27687 , \27686 );
xor \U$27345 ( \27688 , \27468 , \27471 );
xnor \U$27346 ( \27689 , \27688 , \27461 );
nand \U$27347 ( \27690 , \27687 , \27689 );
nand \U$27348 ( \27691 , \27675 , \27685 );
nand \U$27349 ( \27692 , \27690 , \27691 );
not \U$27350 ( \27693 , \27692 );
not \U$27351 ( \27694 , \27693 );
xor \U$27352 ( \27695 , \25718 , \25809 );
xnor \U$27353 ( \27696 , \27695 , \25804 );
not \U$27354 ( \27697 , \27696 );
not \U$27355 ( \27698 , \27697 );
not \U$27356 ( \27699 , \25793 );
xor \U$27357 ( \27700 , \25795 , \27699 );
xnor \U$27358 ( \27701 , \27700 , \25797 );
not \U$27359 ( \27702 , \27701 );
not \U$27360 ( \27703 , \27702 );
xor \U$27361 ( \27704 , \25632 , \25666 );
xor \U$27362 ( \27705 , \27704 , \25673 );
not \U$27363 ( \27706 , \27705 );
xor \U$27364 ( \27707 , \25886 , \25826 );
xnor \U$27365 ( \27708 , \27707 , \25889 );
not \U$27366 ( \27709 , \27708 );
or \U$27367 ( \27710 , \27706 , \27709 );
or \U$27368 ( \27711 , \27708 , \27705 );
nand \U$27369 ( \27712 , \27710 , \27711 );
not \U$27370 ( \27713 , \27712 );
or \U$27371 ( \27714 , \27703 , \27713 );
not \U$27372 ( \27715 , \27708 );
nand \U$27373 ( \27716 , \27715 , \27705 );
nand \U$27374 ( \27717 , \27714 , \27716 );
not \U$27375 ( \27718 , \1135 );
not \U$27376 ( \27719 , \25732 );
or \U$27377 ( \27720 , \27718 , \27719 );
and \U$27378 ( \27721 , \17883 , \1111 );
not \U$27379 ( \27722 , \17883 );
and \U$27380 ( \27723 , \27722 , RI98718c0_129);
nor \U$27381 ( \27724 , \27721 , \27723 );
not \U$27382 ( \27725 , \27724 );
nand \U$27383 ( \27726 , \27725 , \1083 );
nand \U$27384 ( \27727 , \27720 , \27726 );
not \U$27385 ( \27728 , \27727 );
not \U$27386 ( \27729 , \3163 );
not \U$27387 ( \27730 , \27585 );
or \U$27388 ( \27731 , \27729 , \27730 );
nand \U$27389 ( \27732 , \25722 , \3169 );
nand \U$27390 ( \27733 , \27731 , \27732 );
not \U$27391 ( \27734 , \796 );
not \U$27392 ( \27735 , \25849 );
or \U$27393 ( \27736 , \27734 , \27735 );
not \U$27394 ( \27737 , \6568 );
not \U$27395 ( \27738 , \19594 );
or \U$27396 ( \27739 , \27737 , \27738 );
not \U$27397 ( \27740 , \19591 );
or \U$27398 ( \27741 , \27740 , \1078 );
nand \U$27399 ( \27742 , \27739 , \27741 );
nand \U$27400 ( \27743 , \27742 , \791 );
nand \U$27401 ( \27744 , \27736 , \27743 );
xor \U$27402 ( \27745 , \27733 , \27744 );
not \U$27403 ( \27746 , \27745 );
or \U$27404 ( \27747 , \27728 , \27746 );
nand \U$27405 ( \27748 , \27744 , \27733 );
nand \U$27406 ( \27749 , \27747 , \27748 );
not \U$27407 ( \27750 , \27749 );
not \U$27408 ( \27751 , \27568 );
not \U$27409 ( \27752 , \27559 );
or \U$27410 ( \27753 , \27751 , \27752 );
not \U$27411 ( \27754 , \27548 );
nand \U$27412 ( \27755 , \27754 , \27558 );
nand \U$27413 ( \27756 , \27753 , \27755 );
not \U$27414 ( \27757 , \27756 );
not \U$27415 ( \27758 , \27757 );
and \U$27416 ( \27759 , \27750 , \27758 );
and \U$27417 ( \27760 , \27749 , \27757 );
nor \U$27418 ( \27761 , \27759 , \27760 );
not \U$27419 ( \27762 , \27761 );
not \U$27420 ( \27763 , \27762 );
not \U$27421 ( \27764 , \17098 );
not \U$27422 ( \27765 , \25761 );
or \U$27423 ( \27766 , \27764 , \27765 );
not \U$27424 ( \27767 , RI98725e0_157);
not \U$27425 ( \27768 , \18498 );
or \U$27426 ( \27769 , \27767 , \27768 );
or \U$27427 ( \27770 , \18498 , RI98725e0_157);
nand \U$27428 ( \27771 , \27769 , \27770 );
nand \U$27429 ( \27772 , \27771 , \18171 );
nand \U$27430 ( \27773 , \27766 , \27772 );
not \U$27431 ( \27774 , \27773 );
not \U$27432 ( \27775 , \4923 );
not \U$27433 ( \27776 , \25782 );
or \U$27434 ( \27777 , \27775 , \27776 );
not \U$27435 ( \27778 , RI9872388_152);
not \U$27436 ( \27779 , \9911 );
or \U$27437 ( \27780 , \27778 , \27779 );
or \U$27438 ( \27781 , \8579 , RI9872388_152);
nand \U$27439 ( \27782 , \27780 , \27781 );
nand \U$27440 ( \27783 , \27782 , \4918 );
nand \U$27441 ( \27784 , \27777 , \27783 );
not \U$27442 ( \27785 , \5034 );
and \U$27443 ( \27786 , RI9872478_154, \9881 );
not \U$27444 ( \27787 , RI9872478_154);
and \U$27445 ( \27788 , \27787 , \9880 );
nor \U$27446 ( \27789 , \27786 , \27788 );
not \U$27447 ( \27790 , \27789 );
or \U$27448 ( \27791 , \27785 , \27790 );
nand \U$27449 ( \27792 , \25747 , \5035 );
nand \U$27450 ( \27793 , \27791 , \27792 );
xor \U$27451 ( \27794 , \27784 , \27793 );
not \U$27452 ( \27795 , \27794 );
or \U$27453 ( \27796 , \27774 , \27795 );
nand \U$27454 ( \27797 , \27784 , \27793 );
nand \U$27455 ( \27798 , \27796 , \27797 );
not \U$27456 ( \27799 , \27798 );
or \U$27457 ( \27800 , \27763 , \27799 );
not \U$27458 ( \27801 , \27757 );
nand \U$27459 ( \27802 , \27801 , \27749 );
nand \U$27460 ( \27803 , \27800 , \27802 );
not \U$27461 ( \27804 , \25737 );
not \U$27462 ( \27805 , \25726 );
or \U$27463 ( \27806 , \27804 , \27805 );
or \U$27464 ( \27807 , \25726 , \25737 );
nand \U$27465 ( \27808 , \27806 , \27807 );
xor \U$27466 ( \27809 , \25749 , \27808 );
not \U$27467 ( \27810 , \3467 );
not \U$27468 ( \27811 , \25771 );
or \U$27469 ( \27812 , \27810 , \27811 );
and \U$27470 ( \27813 , RI98726d0_159, \9849 );
not \U$27471 ( \27814 , RI98726d0_159);
and \U$27472 ( \27815 , \27814 , \8708 );
or \U$27473 ( \27816 , \27813 , \27815 );
nand \U$27474 ( \27817 , \27816 , \3464 );
nand \U$27475 ( \27818 , \27812 , \27817 );
not \U$27476 ( \27819 , \5653 );
not \U$27477 ( \27820 , \27238 );
or \U$27478 ( \27821 , \27819 , \27820 );
not \U$27479 ( \27822 , RI9872568_156);
not \U$27480 ( \27823 , \16946 );
or \U$27481 ( \27824 , \27822 , \27823 );
or \U$27482 ( \27825 , \12717 , RI9872568_156);
nand \U$27483 ( \27826 , \27824 , \27825 );
nand \U$27484 ( \27827 , \27826 , \6063 );
nand \U$27485 ( \27828 , \27821 , \27827 );
xor \U$27486 ( \27829 , \27818 , \27828 );
not \U$27487 ( \27830 , \8041 );
not \U$27488 ( \27831 , \27259 );
or \U$27489 ( \27832 , \27830 , \27831 );
and \U$27490 ( \27833 , RI9872a18_166, \8053 );
not \U$27491 ( \27834 , RI9872a18_166);
and \U$27492 ( \27835 , \27834 , \12802 );
or \U$27493 ( \27836 , \27833 , \27835 );
nand \U$27494 ( \27837 , \27836 , \8029 );
nand \U$27495 ( \27838 , \27832 , \27837 );
and \U$27496 ( \27839 , \27829 , \27838 );
and \U$27497 ( \27840 , \27818 , \27828 );
or \U$27498 ( \27841 , \27839 , \27840 );
xor \U$27499 ( \27842 , \27809 , \27841 );
not \U$27500 ( \27843 , \6610 );
not \U$27501 ( \27844 , \27400 );
or \U$27502 ( \27845 , \27843 , \27844 );
not \U$27503 ( \27846 , \7049 );
not \U$27504 ( \27847 , \9895 );
not \U$27505 ( \27848 , \27847 );
or \U$27506 ( \27849 , \27846 , \27848 );
nand \U$27507 ( \27850 , \8334 , RI98728b0_163);
nand \U$27508 ( \27851 , \27849 , \27850 );
nand \U$27509 ( \27852 , \27851 , \6284 );
nand \U$27510 ( \27853 , \27845 , \27852 );
xor \U$27511 ( \27854 , \27383 , \27389 );
xor \U$27512 ( \27855 , \27853 , \27854 );
not \U$27513 ( \27856 , \7338 );
not \U$27514 ( \27857 , \27248 );
or \U$27515 ( \27858 , \27856 , \27857 );
not \U$27516 ( \27859 , \7333 );
not \U$27517 ( \27860 , \8082 );
or \U$27518 ( \27861 , \27859 , \27860 );
not \U$27519 ( \27862 , \17449 );
nand \U$27520 ( \27863 , \27862 , RI98729a0_165);
nand \U$27521 ( \27864 , \27861 , \27863 );
nand \U$27522 ( \27865 , \27864 , \7325 );
nand \U$27523 ( \27866 , \27858 , \27865 );
not \U$27524 ( \27867 , \27866 );
not \U$27525 ( \27868 , \27867 );
and \U$27526 ( \27869 , \27855 , \27868 );
and \U$27527 ( \27870 , \27853 , \27854 );
or \U$27528 ( \27871 , \27869 , \27870 );
and \U$27529 ( \27872 , \27842 , \27871 );
and \U$27530 ( \27873 , \27809 , \27841 );
or \U$27531 ( \27874 , \27872 , \27873 );
xor \U$27532 ( \27875 , \27803 , \27874 );
not \U$27533 ( \27876 , \8752 );
not \U$27534 ( \27877 , \27145 );
or \U$27535 ( \27878 , \27876 , \27877 );
not \U$27536 ( \27879 , \8732 );
not \U$27537 ( \27880 , \18685 );
or \U$27538 ( \27881 , \27879 , \27880 );
or \U$27539 ( \27882 , \3537 , \8732 );
nand \U$27540 ( \27883 , \27881 , \27882 );
nand \U$27541 ( \27884 , \27883 , \9527 );
nand \U$27542 ( \27885 , \27878 , \27884 );
not \U$27543 ( \27886 , \27885 );
not \U$27544 ( \27887 , \1455 );
not \U$27545 ( \27888 , \17868 );
not \U$27546 ( \27889 , \27888 );
and \U$27547 ( \27890 , \27889 , \3487 );
not \U$27548 ( \27891 , \27889 );
and \U$27549 ( \27892 , \27891 , RI9871c08_136);
nor \U$27550 ( \27893 , \27890 , \27892 );
not \U$27551 ( \27894 , \27893 );
or \U$27552 ( \27895 , \27887 , \27894 );
nand \U$27553 ( \27896 , \27556 , \1428 );
nand \U$27554 ( \27897 , \27895 , \27896 );
or \U$27555 ( \27898 , \27530 , \1494 );
and \U$27556 ( \27899 , \22278 , RI9871c80_137);
and \U$27557 ( \27900 , \21779 , \1584 );
nor \U$27558 ( \27901 , \27899 , \27900 );
or \U$27559 ( \27902 , \27901 , \1499 );
nand \U$27560 ( \27903 , \27898 , \27902 );
not \U$27561 ( \27904 , \27903 );
or \U$27562 ( \27905 , \4044 , \1491 );
or \U$27563 ( \27906 , RI9871b18_134, RI9871cf8_138);
nand \U$27564 ( \27907 , \27906 , \24450 );
nand \U$27565 ( \27908 , \27905 , \27907 , RI9871c80_137);
nor \U$27566 ( \27909 , \27904 , \27908 );
xor \U$27567 ( \27910 , \27897 , \27909 );
or \U$27568 ( \27911 , \27724 , \6671 );
not \U$27569 ( \27912 , RI98718c0_129);
not \U$27570 ( \27913 , \13934 );
or \U$27571 ( \27914 , \27912 , \27913 );
or \U$27572 ( \27915 , \20765 , RI98718c0_129);
nand \U$27573 ( \27916 , \27914 , \27915 );
not \U$27574 ( \27917 , \27916 );
or \U$27575 ( \27918 , \27917 , \1688 );
nand \U$27576 ( \27919 , \27911 , \27918 );
nand \U$27577 ( \27920 , \27910 , \27919 );
nand \U$27578 ( \27921 , \27897 , \27909 );
and \U$27579 ( \27922 , \27920 , \27921 );
not \U$27580 ( \27923 , \27922 );
not \U$27581 ( \27924 , \19046 );
not \U$27582 ( \27925 , \27417 );
or \U$27583 ( \27926 , \27924 , \27925 );
xor \U$27584 ( \27927 , RI98734e0_189, \5908 );
nand \U$27585 ( \27928 , \27927 , \19243 );
nand \U$27586 ( \27929 , \27926 , \27928 );
not \U$27587 ( \27930 , \27929 );
or \U$27588 ( \27931 , \27923 , \27930 );
or \U$27589 ( \27932 , \27929 , \27922 );
nand \U$27590 ( \27933 , \27931 , \27932 );
not \U$27591 ( \27934 , \27933 );
or \U$27592 ( \27935 , \27886 , \27934 );
not \U$27593 ( \27936 , \27922 );
nand \U$27594 ( \27937 , \27936 , \27929 );
nand \U$27595 ( \27938 , \27935 , \27937 );
not \U$27596 ( \27939 , \27938 );
not \U$27597 ( \27940 , \9686 );
not \U$27598 ( \27941 , RI9872e50_175);
not \U$27599 ( \27942 , \18647 );
or \U$27600 ( \27943 , \27941 , \27942 );
or \U$27601 ( \27944 , \4176 , RI9872e50_175);
nand \U$27602 ( \27945 , \27943 , \27944 );
not \U$27603 ( \27946 , \27945 );
or \U$27604 ( \27947 , \27940 , \27946 );
nand \U$27605 ( \27948 , \27132 , \10332 );
nand \U$27606 ( \27949 , \27947 , \27948 );
not \U$27607 ( \27950 , \10624 );
not \U$27608 ( \27951 , \27316 );
or \U$27609 ( \27952 , \27950 , \27951 );
and \U$27610 ( \27953 , RI9872d60_173, \5623 );
not \U$27611 ( \27954 , RI9872d60_173);
and \U$27612 ( \27955 , \27954 , \12971 );
nor \U$27613 ( \27956 , \27953 , \27955 );
nand \U$27614 ( \27957 , \27956 , \10251 );
nand \U$27615 ( \27958 , \27952 , \27957 );
or \U$27616 ( \27959 , \27949 , \27958 );
not \U$27617 ( \27960 , \17528 );
not \U$27618 ( \27961 , \27125 );
or \U$27619 ( \27962 , \27960 , \27961 );
not \U$27620 ( \27963 , \22727 );
not \U$27621 ( \27964 , \1061 );
or \U$27622 ( \27965 , \27963 , \27964 );
not \U$27623 ( \27966 , RI9873288_184);
or \U$27624 ( \27967 , \6573 , \27966 );
nand \U$27625 ( \27968 , \27965 , \27967 );
nand \U$27626 ( \27969 , \27968 , \18508 );
nand \U$27627 ( \27970 , \27962 , \27969 );
nand \U$27628 ( \27971 , \27959 , \27970 );
nand \U$27629 ( \27972 , \27949 , \27958 );
and \U$27630 ( \27973 , \27971 , \27972 );
buf \U$27631 ( \27974 , \25869 );
xor \U$27632 ( \27975 , \25853 , \27974 );
not \U$27633 ( \27976 , \27975 );
and \U$27634 ( \27977 , \27973 , \27976 );
not \U$27635 ( \27978 , \27973 );
and \U$27636 ( \27979 , \27978 , \27975 );
nor \U$27637 ( \27980 , \27977 , \27979 );
not \U$27638 ( \27981 , \27980 );
or \U$27639 ( \27982 , \27939 , \27981 );
not \U$27640 ( \27983 , \27972 );
not \U$27641 ( \27984 , \27971 );
or \U$27642 ( \27985 , \27983 , \27984 );
nand \U$27643 ( \27986 , \27985 , \27975 );
nand \U$27644 ( \27987 , \27982 , \27986 );
and \U$27645 ( \27988 , \27875 , \27987 );
and \U$27646 ( \27989 , \27803 , \27874 );
or \U$27647 ( \27990 , \27988 , \27989 );
not \U$27648 ( \27991 , \27990 );
xor \U$27649 ( \27992 , \27242 , \27252 );
xor \U$27650 ( \27993 , \27992 , \27263 );
xor \U$27651 ( \27994 , \27419 , \27408 );
xor \U$27652 ( \27995 , \27993 , \27994 );
not \U$27653 ( \27996 , \17371 );
not \U$27654 ( \27997 , RI98733f0_187);
not \U$27655 ( \27998 , \17363 );
or \U$27656 ( \27999 , \27997 , \27998 );
or \U$27657 ( \28000 , \1340 , RI98733f0_187);
nand \U$27658 ( \28001 , \27999 , \28000 );
not \U$27659 ( \28002 , \28001 );
or \U$27660 ( \28003 , \27996 , \28002 );
nand \U$27661 ( \28004 , \27191 , \19282 );
nand \U$27662 ( \28005 , \28003 , \28004 );
not \U$27663 ( \28006 , \9952 );
not \U$27664 ( \28007 , \14132 );
not \U$27665 ( \28008 , \5884 );
or \U$27666 ( \28009 , \28007 , \28008 );
nand \U$27667 ( \28010 , \3691 , RI9873030_179);
nand \U$27668 ( \28011 , \28009 , \28010 );
not \U$27669 ( \28012 , \28011 );
or \U$27670 ( \28013 , \28006 , \28012 );
nand \U$27671 ( \28014 , \27224 , \9937 );
nand \U$27672 ( \28015 , \28013 , \28014 );
xor \U$27673 ( \28016 , \28005 , \28015 );
not \U$27674 ( \28017 , \12868 );
not \U$27675 ( \28018 , \27162 );
or \U$27676 ( \28019 , \28017 , \28018 );
and \U$27677 ( \28020 , \1485 , \13022 );
not \U$27678 ( \28021 , \1485 );
and \U$27679 ( \28022 , \28021 , RI98730a8_180);
nor \U$27680 ( \28023 , \28020 , \28022 );
nand \U$27681 ( \28024 , \28023 , \11350 );
nand \U$27682 ( \28025 , \28019 , \28024 );
and \U$27683 ( \28026 , \28016 , \28025 );
and \U$27684 ( \28027 , \28005 , \28015 );
or \U$27685 ( \28028 , \28026 , \28027 );
and \U$27686 ( \28029 , \27995 , \28028 );
and \U$27687 ( \28030 , \27993 , \27994 );
or \U$27688 ( \28031 , \28029 , \28030 );
not \U$27689 ( \28032 , \28031 );
xnor \U$27690 ( \28033 , \25789 , \25755 );
xor \U$27691 ( \28034 , \27266 , \28033 );
xnor \U$27692 ( \28035 , \28034 , \27272 );
not \U$27693 ( \28036 , \28035 );
or \U$27694 ( \28037 , \28032 , \28036 );
not \U$27695 ( \28038 , \28033 );
xor \U$27696 ( \28039 , \27266 , \27272 );
nand \U$27697 ( \28040 , \28038 , \28039 );
nand \U$27698 ( \28041 , \28037 , \28040 );
not \U$27699 ( \28042 , \28041 );
or \U$27700 ( \28043 , \27991 , \28042 );
xor \U$27701 ( \28044 , \27340 , \27337 );
xnor \U$27702 ( \28045 , \28044 , \27347 );
not \U$27703 ( \28046 , \28041 );
not \U$27704 ( \28047 , \27990 );
nand \U$27705 ( \28048 , \28046 , \28047 );
nand \U$27706 ( \28049 , \28045 , \28048 );
nand \U$27707 ( \28050 , \28043 , \28049 );
and \U$27708 ( \28051 , \27717 , \28050 );
not \U$27709 ( \28052 , \27717 );
not \U$27710 ( \28053 , \28050 );
and \U$27711 ( \28054 , \28052 , \28053 );
nor \U$27712 ( \28055 , \28051 , \28054 );
not \U$27713 ( \28056 , \28055 );
or \U$27714 ( \28057 , \27698 , \28056 );
nand \U$27715 ( \28058 , \28050 , \27717 );
nand \U$27716 ( \28059 , \28057 , \28058 );
buf \U$27717 ( \28060 , \27448 );
not \U$27718 ( \28061 , \28060 );
not \U$27719 ( \28062 , \27452 );
not \U$27720 ( \28063 , \27118 );
or \U$27721 ( \28064 , \28062 , \28063 );
or \U$27722 ( \28065 , \27118 , \27452 );
nand \U$27723 ( \28066 , \28064 , \28065 );
not \U$27724 ( \28067 , \28066 );
and \U$27725 ( \28068 , \28061 , \28067 );
and \U$27726 ( \28069 , \28060 , \28066 );
nor \U$27727 ( \28070 , \28068 , \28069 );
and \U$27728 ( \28071 , \28059 , \28070 );
not \U$27729 ( \28072 , \28059 );
not \U$27730 ( \28073 , \28070 );
and \U$27731 ( \28074 , \28072 , \28073 );
nor \U$27732 ( \28075 , \28071 , \28074 );
not \U$27733 ( \28076 , \28075 );
or \U$27734 ( \28077 , \27694 , \28076 );
not \U$27735 ( \28078 , \28055 );
or \U$27736 ( \28079 , \28078 , \27696 );
not \U$27737 ( \28080 , \27717 );
or \U$27738 ( \28081 , \28053 , \28080 );
nand \U$27739 ( \28082 , \28079 , \28081 , \28073 );
nand \U$27740 ( \28083 , \28077 , \28082 );
not \U$27741 ( \28084 , \28083 );
xor \U$27742 ( \28085 , \25708 , \25917 );
xnor \U$27743 ( \28086 , \28085 , \25921 );
not \U$27744 ( \28087 , \28086 );
and \U$27745 ( \28088 , \27113 , \27454 );
not \U$27746 ( \28089 , \27113 );
and \U$27747 ( \28090 , \28089 , \27455 );
nor \U$27748 ( \28091 , \28088 , \28090 );
not \U$27749 ( \28092 , \28091 );
not \U$27750 ( \28093 , \28092 );
not \U$27751 ( \28094 , \27489 );
and \U$27752 ( \28095 , \28093 , \28094 );
and \U$27753 ( \28096 , \27489 , \28092 );
nor \U$27754 ( \28097 , \28095 , \28096 );
not \U$27755 ( \28098 , \28097 );
or \U$27756 ( \28099 , \28087 , \28098 );
or \U$27757 ( \28100 , \28097 , \28086 );
nand \U$27758 ( \28101 , \28099 , \28100 );
not \U$27759 ( \28102 , \28101 );
or \U$27760 ( \28103 , \28084 , \28102 );
not \U$27761 ( \28104 , \28097 );
nand \U$27762 ( \28105 , \28104 , \28086 );
nand \U$27763 ( \28106 , \28103 , \28105 );
nand \U$27764 ( \28107 , \27500 , \28106 );
xor \U$27765 ( \28108 , \27474 , \27483 );
xor \U$27766 ( \28109 , \28108 , \27458 );
not \U$27767 ( \28110 , \28109 );
xnor \U$27768 ( \28111 , \27692 , \28075 );
not \U$27769 ( \28112 , \28111 );
or \U$27770 ( \28113 , \28110 , \28112 );
not \U$27771 ( \28114 , \27712 );
not \U$27772 ( \28115 , \27701 );
and \U$27773 ( \28116 , \28114 , \28115 );
and \U$27774 ( \28117 , \27712 , \27701 );
nor \U$27775 ( \28118 , \28116 , \28117 );
xor \U$27776 ( \28119 , \27362 , \27425 );
xor \U$27777 ( \28120 , \27803 , \27874 );
xor \U$27778 ( \28121 , \28120 , \27987 );
xor \U$27779 ( \28122 , \28119 , \28121 );
xor \U$27780 ( \28123 , \27809 , \27841 );
xor \U$27781 ( \28124 , \28123 , \27871 );
not \U$27782 ( \28125 , \24627 );
not \U$27783 ( \28126 , RI9872f40_177);
not \U$27784 ( \28127 , \14930 );
or \U$27785 ( \28128 , \28126 , \28127 );
or \U$27786 ( \28129 , \14930 , RI9872f40_177);
nand \U$27787 ( \28130 , \28128 , \28129 );
not \U$27788 ( \28131 , \28130 );
or \U$27789 ( \28132 , \28125 , \28131 );
nand \U$27790 ( \28133 , \27883 , \8752 );
nand \U$27791 ( \28134 , \28132 , \28133 );
not \U$27792 ( \28135 , \28134 );
nand \U$27793 ( \28136 , \27945 , \10331 );
not \U$27794 ( \28137 , RI9872e50_175);
not \U$27795 ( \28138 , \5205 );
or \U$27796 ( \28139 , \28137 , \28138 );
or \U$27797 ( \28140 , \12832 , RI9872e50_175);
nand \U$27798 ( \28141 , \28139 , \28140 );
nand \U$27799 ( \28142 , \28141 , \18562 );
nand \U$27800 ( \28143 , \28136 , \28142 );
not \U$27801 ( \28144 , \28143 );
or \U$27802 ( \28145 , \28135 , \28144 );
not \U$27803 ( \28146 , \28134 );
or \U$27804 ( \28147 , \28143 , \28146 );
not \U$27805 ( \28148 , \28142 );
not \U$27806 ( \28149 , \28136 );
or \U$27807 ( \28150 , \28148 , \28149 );
nand \U$27808 ( \28151 , \28150 , \28146 );
nand \U$27809 ( \28152 , \28147 , \28151 );
not \U$27810 ( \28153 , \18508 );
and \U$27811 ( \28154 , RI9873288_184, \17140 );
not \U$27812 ( \28155 , RI9873288_184);
and \U$27813 ( \28156 , \28155 , \1038 );
or \U$27814 ( \28157 , \28154 , \28156 );
not \U$27815 ( \28158 , \28157 );
or \U$27816 ( \28159 , \28153 , \28158 );
nand \U$27817 ( \28160 , \27968 , \17528 );
nand \U$27818 ( \28161 , \28159 , \28160 );
nand \U$27819 ( \28162 , \28152 , \28161 );
nand \U$27820 ( \28163 , \28145 , \28162 );
not \U$27821 ( \28164 , \28163 );
not \U$27822 ( \28165 , \27903 );
not \U$27823 ( \28166 , \27908 );
and \U$27824 ( \28167 , \28165 , \28166 );
and \U$27825 ( \28168 , \27903 , \27908 );
nor \U$27826 ( \28169 , \28167 , \28168 );
not \U$27827 ( \28170 , \28169 );
not \U$27828 ( \28171 , \1290 );
not \U$27829 ( \28172 , \27543 );
or \U$27830 ( \28173 , \28171 , \28172 );
not \U$27831 ( \28174 , \1283 );
not \U$27832 ( \28175 , \24854 );
or \U$27833 ( \28176 , \28174 , \28175 );
or \U$27834 ( \28177 , \24854 , \1283 );
nand \U$27835 ( \28178 , \28176 , \28177 );
nand \U$27836 ( \28179 , \28178 , \1291 );
nand \U$27837 ( \28180 , \28173 , \28179 );
not \U$27838 ( \28181 , \28180 );
and \U$27839 ( \28182 , \28170 , \28181 );
and \U$27840 ( \28183 , \28180 , \28169 );
nor \U$27841 ( \28184 , \28182 , \28183 );
not \U$27842 ( \28185 , \28184 );
not \U$27843 ( \28186 , \28185 );
not \U$27844 ( \28187 , \1134 );
not \U$27845 ( \28188 , \27916 );
or \U$27846 ( \28189 , \28187 , \28188 );
not \U$27847 ( \28190 , \1111 );
not \U$27848 ( \28191 , \17741 );
not \U$27849 ( \28192 , \28191 );
or \U$27850 ( \28193 , \28190 , \28192 );
not \U$27851 ( \28194 , \17912 );
nand \U$27852 ( \28195 , \28194 , RI98718c0_129);
nand \U$27853 ( \28196 , \28193 , \28195 );
nand \U$27854 ( \28197 , \28196 , \1083 );
nand \U$27855 ( \28198 , \28189 , \28197 );
not \U$27856 ( \28199 , \28198 );
or \U$27857 ( \28200 , \28186 , \28199 );
not \U$27858 ( \28201 , \28169 );
nand \U$27859 ( \28202 , \28201 , \28180 );
nand \U$27860 ( \28203 , \28200 , \28202 );
not \U$27861 ( \28204 , \28203 );
not \U$27862 ( \28205 , \28204 );
not \U$27863 ( \28206 , \6286 );
not \U$27864 ( \28207 , \27851 );
or \U$27865 ( \28208 , \28206 , \28207 );
and \U$27866 ( \28209 , RI98728b0_163, \24779 );
not \U$27867 ( \28210 , RI98728b0_163);
and \U$27868 ( \28211 , \28210 , \11627 );
nor \U$27869 ( \28212 , \28209 , \28211 );
nand \U$27870 ( \28213 , \28212 , \6284 );
nand \U$27871 ( \28214 , \28208 , \28213 );
not \U$27872 ( \28215 , \28214 );
or \U$27873 ( \28216 , \28205 , \28215 );
or \U$27874 ( \28217 , \28214 , \28204 );
nand \U$27875 ( \28218 , \28216 , \28217 );
not \U$27876 ( \28219 , \28218 );
not \U$27877 ( \28220 , \20147 );
not \U$27878 ( \28221 , \27927 );
or \U$27879 ( \28222 , \28220 , \28221 );
not \U$27880 ( \28223 , RI98734e0_189);
not \U$27881 ( \28224 , \1252 );
or \U$27882 ( \28225 , \28223 , \28224 );
or \U$27883 ( \28226 , \1252 , RI98734e0_189);
nand \U$27884 ( \28227 , \28225 , \28226 );
nand \U$27885 ( \28228 , \28227 , \19036 );
nand \U$27886 ( \28229 , \28222 , \28228 );
not \U$27887 ( \28230 , \28229 );
or \U$27888 ( \28231 , \28219 , \28230 );
not \U$27889 ( \28232 , \28204 );
nand \U$27890 ( \28233 , \28232 , \28214 );
nand \U$27891 ( \28234 , \28231 , \28233 );
not \U$27892 ( \28235 , \28234 );
not \U$27893 ( \28236 , \7338 );
not \U$27894 ( \28237 , \27864 );
or \U$27895 ( \28238 , \28236 , \28237 );
xor \U$27896 ( \28239 , RI98729a0_165, \8923 );
nand \U$27897 ( \28240 , \28239 , \7325 );
nand \U$27898 ( \28241 , \28238 , \28240 );
not \U$27899 ( \28242 , \8029 );
not \U$27900 ( \28243 , \8031 );
not \U$27901 ( \28244 , \10412 );
or \U$27902 ( \28245 , \28243 , \28244 );
or \U$27903 ( \28246 , \7905 , \8031 );
nand \U$27904 ( \28247 , \28245 , \28246 );
not \U$27905 ( \28248 , \28247 );
or \U$27906 ( \28249 , \28242 , \28248 );
nand \U$27907 ( \28250 , \27836 , \13017 );
nand \U$27908 ( \28251 , \28249 , \28250 );
xor \U$27909 ( \28252 , \28241 , \28251 );
not \U$27910 ( \28253 , \27634 );
not \U$27911 ( \28254 , \9214 );
or \U$27912 ( \28255 , \28253 , \28254 );
not \U$27913 ( \28256 , \11691 );
not \U$27914 ( \28257 , RI9872b80_169);
not \U$27915 ( \28258 , \18809 );
not \U$27916 ( \28259 , \28258 );
or \U$27917 ( \28260 , \28257 , \28259 );
nand \U$27918 ( \28261 , \7108 , \9198 );
nand \U$27919 ( \28262 , \28260 , \28261 );
nand \U$27920 ( \28263 , \28256 , \28262 );
nand \U$27921 ( \28264 , \28255 , \28263 );
nand \U$27922 ( \28265 , \28252 , \28264 );
not \U$27923 ( \28266 , \28265 );
and \U$27924 ( \28267 , \28241 , \28251 );
nor \U$27925 ( \28268 , \28266 , \28267 );
not \U$27926 ( \28269 , \28268 );
or \U$27927 ( \28270 , \28235 , \28269 );
not \U$27928 ( \28271 , \28267 );
not \U$27929 ( \28272 , \28271 );
not \U$27930 ( \28273 , \28265 );
or \U$27931 ( \28274 , \28272 , \28273 );
not \U$27932 ( \28275 , \28234 );
nand \U$27933 ( \28276 , \28274 , \28275 );
nand \U$27934 ( \28277 , \28270 , \28276 );
not \U$27935 ( \28278 , \28277 );
or \U$27936 ( \28279 , \28164 , \28278 );
not \U$27937 ( \28280 , \28271 );
not \U$27938 ( \28281 , \28265 );
or \U$27939 ( \28282 , \28280 , \28281 );
nand \U$27940 ( \28283 , \28282 , \28234 );
nand \U$27941 ( \28284 , \28279 , \28283 );
xor \U$27942 ( \28285 , \28124 , \28284 );
not \U$27943 ( \28286 , \9668 );
not \U$27944 ( \28287 , \27640 );
or \U$27945 ( \28288 , \28286 , \28287 );
not \U$27946 ( \28289 , RI9872bf8_170);
not \U$27947 ( \28290 , \5775 );
or \U$27948 ( \28291 , \28289 , \28290 );
or \U$27949 ( \28292 , \5775 , RI9872bf8_170);
nand \U$27950 ( \28293 , \28291 , \28292 );
nand \U$27951 ( \28294 , \28293 , \9249 );
nand \U$27952 ( \28295 , \28288 , \28294 );
not \U$27953 ( \28296 , \28295 );
not \U$27954 ( \28297 , \13476 );
not \U$27955 ( \28298 , RI9873210_183);
not \U$27956 ( \28299 , \9254 );
or \U$27957 ( \28300 , \28298 , \28299 );
or \U$27958 ( \28301 , \1190 , RI9873210_183);
nand \U$27959 ( \28302 , \28300 , \28301 );
not \U$27960 ( \28303 , \28302 );
or \U$27961 ( \28304 , \28297 , \28303 );
nand \U$27962 ( \28305 , \27650 , \17123 );
nand \U$27963 ( \28306 , \28304 , \28305 );
not \U$27964 ( \28307 , \9312 );
not \U$27965 ( \28308 , RI9872d60_173);
not \U$27966 ( \28309 , \7791 );
or \U$27967 ( \28310 , \28308 , \28309 );
or \U$27968 ( \28311 , \7791 , RI9872d60_173);
nand \U$27969 ( \28312 , \28310 , \28311 );
not \U$27970 ( \28313 , \28312 );
or \U$27971 ( \28314 , \28307 , \28313 );
nand \U$27972 ( \28315 , \27956 , \10624 );
nand \U$27973 ( \28316 , \28314 , \28315 );
and \U$27974 ( \28317 , \28306 , \28316 );
not \U$27975 ( \28318 , \28306 );
not \U$27976 ( \28319 , \28316 );
and \U$27977 ( \28320 , \28318 , \28319 );
nor \U$27978 ( \28321 , \28317 , \28320 );
not \U$27979 ( \28322 , \28321 );
or \U$27980 ( \28323 , \28296 , \28322 );
nand \U$27981 ( \28324 , \28306 , \28316 );
nand \U$27982 ( \28325 , \28323 , \28324 );
xor \U$27983 ( \28326 , \27854 , \27853 );
xor \U$27984 ( \28327 , \28326 , \27867 );
not \U$27985 ( \28328 , \28327 );
nor \U$27986 ( \28329 , \28325 , \28328 );
xnor \U$27987 ( \28330 , \27910 , \27919 );
not \U$27988 ( \28331 , \28330 );
not \U$27989 ( \28332 , RI9873648_192);
not \U$27990 ( \28333 , \27619 );
or \U$27991 ( \28334 , \28332 , \28333 );
xor \U$27992 ( \28335 , RI9873558_190, \846 );
nand \U$27993 ( \28336 , \28335 , \20626 );
nand \U$27994 ( \28337 , \28334 , \28336 );
xor \U$27995 ( \28338 , \28331 , \28337 );
not \U$27996 ( \28339 , \12868 );
not \U$27997 ( \28340 , \28023 );
or \U$27998 ( \28341 , \28339 , \28340 );
xor \U$27999 ( \28342 , RI98730a8_180, \18453 );
nand \U$28000 ( \28343 , \28342 , \13020 );
nand \U$28001 ( \28344 , \28341 , \28343 );
and \U$28002 ( \28345 , \28338 , \28344 );
and \U$28003 ( \28346 , \28331 , \28337 );
nor \U$28004 ( \28347 , \28345 , \28346 );
or \U$28005 ( \28348 , \28329 , \28347 );
nand \U$28006 ( \28349 , \28325 , \28328 );
nand \U$28007 ( \28350 , \28348 , \28349 );
and \U$28008 ( \28351 , \28285 , \28350 );
and \U$28009 ( \28352 , \28124 , \28284 );
or \U$28010 ( \28353 , \28351 , \28352 );
and \U$28011 ( \28354 , \28122 , \28353 );
and \U$28012 ( \28355 , \28119 , \28121 );
nor \U$28013 ( \28356 , \28354 , \28355 );
xor \U$28014 ( \28357 , \28118 , \28356 );
xor \U$28015 ( \28358 , \27432 , \27441 );
xnor \U$28016 ( \28359 , \28358 , \27437 );
not \U$28017 ( \28360 , \28359 );
and \U$28018 ( \28361 , \27745 , \27727 );
not \U$28019 ( \28362 , \27745 );
not \U$28020 ( \28363 , \27727 );
and \U$28021 ( \28364 , \28362 , \28363 );
nor \U$28022 ( \28365 , \28361 , \28364 );
not \U$28023 ( \28366 , \3464 );
not \U$28024 ( \28367 , RI98726d0_159);
not \U$28025 ( \28368 , \9113 );
or \U$28026 ( \28369 , \28367 , \28368 );
or \U$28027 ( \28370 , RI98726d0_159, \9113 );
nand \U$28028 ( \28371 , \28369 , \28370 );
not \U$28029 ( \28372 , \28371 );
or \U$28030 ( \28373 , \28366 , \28372 );
nand \U$28031 ( \28374 , \27816 , \3467 );
nand \U$28032 ( \28375 , \28373 , \28374 );
not \U$28033 ( \28376 , \28375 );
and \U$28034 ( \28377 , \18350 , \13646 );
not \U$28035 ( \28378 , \18350 );
and \U$28036 ( \28379 , \28378 , RI98719b0_131);
nor \U$28037 ( \28380 , \28377 , \28379 );
and \U$28038 ( \28381 , \28380 , \791 );
not \U$28039 ( \28382 , \27742 );
nor \U$28040 ( \28383 , \28382 , \786 );
nor \U$28041 ( \28384 , \28381 , \28383 );
nand \U$28042 ( \28385 , \28376 , \28384 );
not \U$28043 ( \28386 , \28385 );
not \U$28044 ( \28387 , \5034 );
not \U$28045 ( \28388 , RI9872478_154);
not \U$28046 ( \28389 , \8650 );
or \U$28047 ( \28390 , \28388 , \28389 );
or \U$28048 ( \28391 , \11406 , RI9872478_154);
nand \U$28049 ( \28392 , \28390 , \28391 );
not \U$28050 ( \28393 , \28392 );
or \U$28051 ( \28394 , \28387 , \28393 );
nand \U$28052 ( \28395 , \27789 , \5035 );
nand \U$28053 ( \28396 , \28394 , \28395 );
not \U$28054 ( \28397 , \28396 );
or \U$28055 ( \28398 , \28386 , \28397 );
not \U$28056 ( \28399 , \28384 );
nand \U$28057 ( \28400 , \28375 , \28399 );
nand \U$28058 ( \28401 , \28398 , \28400 );
xor \U$28059 ( \28402 , \28365 , \28401 );
not \U$28060 ( \28403 , \4101 );
not \U$28061 ( \28404 , \4092 );
not \U$28062 ( \28405 , \9750 );
or \U$28063 ( \28406 , \28404 , \28405 );
or \U$28064 ( \28407 , \23712 , \6042 );
nand \U$28065 ( \28408 , \28406 , \28407 );
not \U$28066 ( \28409 , \28408 );
or \U$28067 ( \28410 , \28403 , \28409 );
nand \U$28068 ( \28411 , \27771 , \4084 );
nand \U$28069 ( \28412 , \28410 , \28411 );
not \U$28070 ( \28413 , \4918 );
not \U$28071 ( \28414 , RI9872388_152);
not \U$28072 ( \28415 , \10369 );
or \U$28073 ( \28416 , \28414 , \28415 );
or \U$28074 ( \28417 , \8555 , RI9872388_152);
nand \U$28075 ( \28418 , \28416 , \28417 );
not \U$28076 ( \28419 , \28418 );
or \U$28077 ( \28420 , \28413 , \28419 );
nand \U$28078 ( \28421 , \27782 , \4923 );
nand \U$28079 ( \28422 , \28420 , \28421 );
xor \U$28080 ( \28423 , \28412 , \28422 );
not \U$28081 ( \28424 , \5653 );
not \U$28082 ( \28425 , \27826 );
or \U$28083 ( \28426 , \28424 , \28425 );
not \U$28084 ( \28427 , RI9872568_156);
not \U$28085 ( \28428 , \10308 );
or \U$28086 ( \28429 , \28427 , \28428 );
or \U$28087 ( \28430 , \18107 , RI9872568_156);
nand \U$28088 ( \28431 , \28429 , \28430 );
not \U$28089 ( \28432 , \28431 );
not \U$28090 ( \28433 , \9320 );
or \U$28091 ( \28434 , \28432 , \28433 );
nand \U$28092 ( \28435 , \28426 , \28434 );
and \U$28093 ( \28436 , \28423 , \28435 );
and \U$28094 ( \28437 , \28412 , \28422 );
or \U$28095 ( \28438 , \28436 , \28437 );
and \U$28096 ( \28439 , \28402 , \28438 );
and \U$28097 ( \28440 , \28365 , \28401 );
or \U$28098 ( \28441 , \28439 , \28440 );
not \U$28099 ( \28442 , \28441 );
not \U$28100 ( \28443 , \27761 );
not \U$28101 ( \28444 , \27798 );
or \U$28102 ( \28445 , \28443 , \28444 );
or \U$28103 ( \28446 , \27798 , \27761 );
nand \U$28104 ( \28447 , \28445 , \28446 );
not \U$28105 ( \28448 , \28447 );
or \U$28106 ( \28449 , \28442 , \28448 );
or \U$28107 ( \28450 , \28447 , \28441 );
not \U$28108 ( \28451 , \27198 );
not \U$28109 ( \28452 , \27166 );
not \U$28110 ( \28453 , \28452 );
or \U$28111 ( \28454 , \28451 , \28453 );
or \U$28112 ( \28455 , \28452 , \27198 );
nand \U$28113 ( \28456 , \28454 , \28455 );
nand \U$28114 ( \28457 , \28450 , \28456 );
nand \U$28115 ( \28458 , \28449 , \28457 );
xor \U$28116 ( \28459 , \27298 , \27331 );
xor \U$28117 ( \28460 , \28459 , \27334 );
xor \U$28118 ( \28461 , \28458 , \28460 );
not \U$28119 ( \28462 , \28461 );
not \U$28120 ( \28463 , \28462 );
and \U$28121 ( \28464 , \28360 , \28463 );
and \U$28122 ( \28465 , \28458 , \28460 );
nor \U$28123 ( \28466 , \28464 , \28465 );
and \U$28124 ( \28467 , \28357 , \28466 );
and \U$28125 ( \28468 , \28118 , \28356 );
or \U$28126 ( \28469 , \28467 , \28468 );
xor \U$28127 ( \28470 , \27696 , \28080 );
xor \U$28128 ( \28471 , \28470 , \28053 );
xor \U$28129 ( \28472 , \28469 , \28471 );
and \U$28130 ( \28473 , \28041 , \28047 );
not \U$28131 ( \28474 , \28041 );
and \U$28132 ( \28475 , \28474 , \27990 );
nor \U$28133 ( \28476 , \28473 , \28475 );
xor \U$28134 ( \28477 , \28045 , \28476 );
xor \U$28135 ( \28478 , \28031 , \28035 );
xor \U$28136 ( \28479 , \27818 , \27828 );
xor \U$28137 ( \28480 , \28479 , \27838 );
not \U$28138 ( \28481 , \28480 );
xor \U$28139 ( \28482 , \27773 , \27794 );
not \U$28140 ( \28483 , \28482 );
or \U$28141 ( \28484 , \28481 , \28483 );
xor \U$28142 ( \28485 , \27970 , \27958 );
xor \U$28143 ( \28486 , \28485 , \27949 );
not \U$28144 ( \28487 , \28486 );
nand \U$28145 ( \28488 , \28484 , \28487 );
or \U$28146 ( \28489 , \28480 , \28482 );
and \U$28147 ( \28490 , \28488 , \28489 );
not \U$28148 ( \28491 , \28490 );
xor \U$28149 ( \28492 , \27630 , \27655 );
xor \U$28150 ( \28493 , \28492 , \27658 );
not \U$28151 ( \28494 , \28493 );
or \U$28152 ( \28495 , \28491 , \28494 );
or \U$28153 ( \28496 , \28493 , \28490 );
not \U$28154 ( \28497 , \2087 );
not \U$28155 ( \28498 , \27573 );
or \U$28156 ( \28499 , \28497 , \28498 );
not \U$28157 ( \28500 , \2076 );
not \U$28158 ( \28501 , \13281 );
or \U$28159 ( \28502 , \28500 , \28501 );
nand \U$28160 ( \28503 , \24523 , RI9871aa0_133);
nand \U$28161 ( \28504 , \28502 , \28503 );
nand \U$28162 ( \28505 , \28504 , \2071 );
nand \U$28163 ( \28506 , \28499 , \28505 );
not \U$28164 ( \28507 , \28506 );
and \U$28165 ( \28508 , RI98719b0_131, \13860 );
not \U$28166 ( \28509 , RI98719b0_131);
and \U$28167 ( \28510 , \28509 , \20456 );
nor \U$28168 ( \28511 , \28508 , \28510 );
not \U$28169 ( \28512 , \28511 );
not \U$28170 ( \28513 , \792 );
and \U$28171 ( \28514 , \28512 , \28513 );
and \U$28172 ( \28515 , \28380 , \796 );
nor \U$28173 ( \28516 , \28514 , \28515 );
not \U$28174 ( \28517 , \28516 );
not \U$28175 ( \28518 , \3464 );
not \U$28176 ( \28519 , \3593 );
not \U$28177 ( \28520 , \13065 );
or \U$28178 ( \28521 , \28519 , \28520 );
or \U$28179 ( \28522 , \9138 , \4063 );
nand \U$28180 ( \28523 , \28521 , \28522 );
not \U$28181 ( \28524 , \28523 );
or \U$28182 ( \28525 , \28518 , \28524 );
nand \U$28183 ( \28526 , \28371 , \3467 );
nand \U$28184 ( \28527 , \28525 , \28526 );
not \U$28185 ( \28528 , \28527 );
or \U$28186 ( \28529 , \28517 , \28528 );
or \U$28187 ( \28530 , \28527 , \28516 );
nand \U$28188 ( \28531 , \28529 , \28530 );
not \U$28189 ( \28532 , \28531 );
or \U$28190 ( \28533 , \28507 , \28532 );
not \U$28191 ( \28534 , \28516 );
nand \U$28192 ( \28535 , \28534 , \28527 );
nand \U$28193 ( \28536 , \28533 , \28535 );
not \U$28194 ( \28537 , \28536 );
not \U$28195 ( \28538 , \28537 );
not \U$28196 ( \28539 , \9952 );
not \U$28197 ( \28540 , RI9873030_179);
not \U$28198 ( \28541 , \9461 );
or \U$28199 ( \28542 , \28540 , \28541 );
or \U$28200 ( \28543 , \4370 , RI9873030_179);
nand \U$28201 ( \28544 , \28542 , \28543 );
not \U$28202 ( \28545 , \28544 );
or \U$28203 ( \28546 , \28539 , \28545 );
nand \U$28204 ( \28547 , \28011 , \9937 );
nand \U$28205 ( \28548 , \28546 , \28547 );
not \U$28206 ( \28549 , \28548 );
not \U$28207 ( \28550 , \28549 );
or \U$28208 ( \28551 , \28538 , \28550 );
not \U$28209 ( \28552 , \19282 );
not \U$28210 ( \28553 , \28001 );
or \U$28211 ( \28554 , \28552 , \28553 );
and \U$28212 ( \28555 , RI98733f0_187, \4454 );
not \U$28213 ( \28556 , RI98733f0_187);
and \U$28214 ( \28557 , \28556 , \1603 );
nor \U$28215 ( \28558 , \28555 , \28557 );
nand \U$28216 ( \28559 , \28558 , \17371 );
nand \U$28217 ( \28560 , \28554 , \28559 );
nand \U$28218 ( \28561 , \28551 , \28560 );
not \U$28219 ( \28562 , \28537 );
nand \U$28220 ( \28563 , \28562 , \28548 );
nand \U$28221 ( \28564 , \28561 , \28563 );
xor \U$28222 ( \28565 , \27922 , \27885 );
xnor \U$28223 ( \28566 , \28565 , \27929 );
xor \U$28224 ( \28567 , \28564 , \28566 );
xor \U$28225 ( \28568 , \28005 , \28015 );
xor \U$28226 ( \28569 , \28568 , \28025 );
and \U$28227 ( \28570 , \28567 , \28569 );
and \U$28228 ( \28571 , \28564 , \28566 );
or \U$28229 ( \28572 , \28570 , \28571 );
nand \U$28230 ( \28573 , \28496 , \28572 );
nand \U$28231 ( \28574 , \28495 , \28573 );
xor \U$28232 ( \28575 , \28478 , \28574 );
xor \U$28233 ( \28576 , \27662 , \27505 );
and \U$28234 ( \28577 , \28575 , \28576 );
and \U$28235 ( \28578 , \28478 , \28574 );
or \U$28236 ( \28579 , \28577 , \28578 );
not \U$28237 ( \28580 , \28579 );
xor \U$28238 ( \28581 , \28477 , \28580 );
xor \U$28239 ( \28582 , \27501 , \27666 );
xnor \U$28240 ( \28583 , \28582 , \27671 );
and \U$28241 ( \28584 , \28581 , \28583 );
and \U$28242 ( \28585 , \28477 , \28580 );
or \U$28243 ( \28586 , \28584 , \28585 );
and \U$28244 ( \28587 , \28472 , \28586 );
and \U$28245 ( \28588 , \28469 , \28471 );
or \U$28246 ( \28589 , \28587 , \28588 );
not \U$28247 ( \28590 , \28589 );
nand \U$28248 ( \28591 , \28113 , \28590 );
not \U$28249 ( \28592 , \28109 );
not \U$28250 ( \28593 , \28111 );
nand \U$28251 ( \28594 , \28592 , \28593 );
nand \U$28252 ( \28595 , \28591 , \28594 );
not \U$28253 ( \28596 , \28595 );
xor \U$28254 ( \28597 , \28101 , \28083 );
nand \U$28255 ( \28598 , \28596 , \28597 );
nand \U$28256 ( \28599 , \28107 , \28598 );
xor \U$28257 ( \28600 , \25316 , \25318 );
xor \U$28258 ( \28601 , \28600 , \25930 );
xor \U$28259 ( \28602 , \27494 , \27496 );
and \U$28260 ( \28603 , \28602 , \27498 );
and \U$28261 ( \28604 , \27494 , \27496 );
or \U$28262 ( \28605 , \28603 , \28604 );
nor \U$28263 ( \28606 , \28601 , \28605 );
not \U$28264 ( \28607 , \28606 );
xor \U$28265 ( \28608 , \28109 , \28590 );
xnor \U$28266 ( \28609 , \28608 , \28111 );
not \U$28267 ( \28610 , \27686 );
nand \U$28268 ( \28611 , \28610 , \27691 );
not \U$28269 ( \28612 , \28611 );
not \U$28270 ( \28613 , \27689 );
and \U$28271 ( \28614 , \28612 , \28613 );
and \U$28272 ( \28615 , \28611 , \27689 );
nor \U$28273 ( \28616 , \28614 , \28615 );
xor \U$28274 ( \28617 , \28118 , \28356 );
xor \U$28275 ( \28618 , \28617 , \28466 );
not \U$28276 ( \28619 , \28618 );
xor \U$28277 ( \28620 , \28441 , \28447 );
xnor \U$28278 ( \28621 , \28620 , \28456 );
xor \U$28279 ( \28622 , \27516 , \27513 );
xnor \U$28280 ( \28623 , \28622 , \27626 );
xor \U$28281 ( \28624 , \28621 , \28623 );
xor \U$28282 ( \28625 , \28365 , \28401 );
xor \U$28283 ( \28626 , \28625 , \28438 );
not \U$28284 ( \28627 , \3163 );
not \U$28285 ( \28628 , \11455 );
and \U$28286 ( \28629 , RI9872310_151, \28628 );
not \U$28287 ( \28630 , RI9872310_151);
and \U$28288 ( \28631 , \28630 , \12788 );
nor \U$28289 ( \28632 , \28629 , \28631 );
not \U$28290 ( \28633 , \28632 );
or \U$28291 ( \28634 , \28627 , \28633 );
nand \U$28292 ( \28635 , \27592 , \3170 );
nand \U$28293 ( \28636 , \28634 , \28635 );
not \U$28294 ( \28637 , \28636 );
not \U$28295 ( \28638 , \1428 );
not \U$28296 ( \28639 , \27893 );
or \U$28297 ( \28640 , \28638 , \28639 );
and \U$28298 ( \28641 , \24868 , RI9871c08_136);
not \U$28299 ( \28642 , \24868 );
and \U$28300 ( \28643 , \28642 , \3487 );
nor \U$28301 ( \28644 , \28641 , \28643 );
nand \U$28302 ( \28645 , \28644 , \1455 );
nand \U$28303 ( \28646 , \28640 , \28645 );
not \U$28304 ( \28647 , \28646 );
not \U$28305 ( \28648 , \28647 );
not \U$28306 ( \28649 , \1428 );
not \U$28307 ( \28650 , \28644 );
or \U$28308 ( \28651 , \28649 , \28650 );
not \U$28309 ( \28652 , \1850 );
buf \U$28310 ( \28653 , \23933 );
not \U$28311 ( \28654 , \28653 );
or \U$28312 ( \28655 , \28652 , \28654 );
not \U$28313 ( \28656 , \20489 );
not \U$28314 ( \28657 , \28656 );
nand \U$28315 ( \28658 , \28657 , RI9871c08_136);
nand \U$28316 ( \28659 , \28655 , \28658 );
nand \U$28317 ( \28660 , \28659 , \1455 );
nand \U$28318 ( \28661 , \28651 , \28660 );
not \U$28319 ( \28662 , \28661 );
buf \U$28320 ( \28663 , \18704 );
and \U$28321 ( \28664 , \28663 , \1493 );
not \U$28322 ( \28665 , \28664 );
not \U$28323 ( \28666 , \1290 );
not \U$28324 ( \28667 , \28178 );
or \U$28325 ( \28668 , \28666 , \28667 );
and \U$28326 ( \28669 , RI9871b18_134, \18194 );
not \U$28327 ( \28670 , RI9871b18_134);
not \U$28328 ( \28671 , \21773 );
and \U$28329 ( \28672 , \28670 , \28671 );
or \U$28330 ( \28673 , \28669 , \28672 );
nand \U$28331 ( \28674 , \28673 , \1291 );
nand \U$28332 ( \28675 , \28668 , \28674 );
not \U$28333 ( \28676 , \28675 );
not \U$28334 ( \28677 , \28676 );
or \U$28335 ( \28678 , \28665 , \28677 );
not \U$28336 ( \28679 , \28664 );
nand \U$28337 ( \28680 , \28679 , \28675 );
nand \U$28338 ( \28681 , \28678 , \28680 );
not \U$28339 ( \28682 , \28681 );
or \U$28340 ( \28683 , \28662 , \28682 );
nand \U$28341 ( \28684 , \28675 , \28664 );
nand \U$28342 ( \28685 , \28683 , \28684 );
not \U$28343 ( \28686 , \28685 );
or \U$28344 ( \28687 , \28648 , \28686 );
or \U$28345 ( \28688 , \28685 , \28647 );
nand \U$28346 ( \28689 , \28687 , \28688 );
not \U$28347 ( \28690 , \28689 );
or \U$28348 ( \28691 , \28637 , \28690 );
nand \U$28349 ( \28692 , \28685 , \28646 );
nand \U$28350 ( \28693 , \28691 , \28692 );
not \U$28351 ( \28694 , \5847 );
not \U$28352 ( \28695 , \28408 );
or \U$28353 ( \28696 , \28694 , \28695 );
and \U$28354 ( \28697 , RI98725e0_157, \12460 );
not \U$28355 ( \28698 , RI98725e0_157);
and \U$28356 ( \28699 , \28698 , \8708 );
or \U$28357 ( \28700 , \28697 , \28699 );
nand \U$28358 ( \28701 , \28700 , \4101 );
nand \U$28359 ( \28702 , \28696 , \28701 );
not \U$28360 ( \28703 , \4923 );
not \U$28361 ( \28704 , \28418 );
or \U$28362 ( \28705 , \28703 , \28704 );
and \U$28363 ( \28706 , RI9872388_152, \13454 );
not \U$28364 ( \28707 , RI9872388_152);
and \U$28365 ( \28708 , \28707 , \8722 );
or \U$28366 ( \28709 , \28706 , \28708 );
nand \U$28367 ( \28710 , \28709 , \4918 );
nand \U$28368 ( \28711 , \28705 , \28710 );
xor \U$28369 ( \28712 , \28702 , \28711 );
not \U$28370 ( \28713 , \5036 );
not \U$28371 ( \28714 , \28392 );
or \U$28372 ( \28715 , \28713 , \28714 );
not \U$28373 ( \28716 , RI9872478_154);
not \U$28374 ( \28717 , \8840 );
or \U$28375 ( \28718 , \28716 , \28717 );
or \U$28376 ( \28719 , \8840 , RI9872478_154);
nand \U$28377 ( \28720 , \28718 , \28719 );
nand \U$28378 ( \28721 , \28720 , \5034 );
nand \U$28379 ( \28722 , \28715 , \28721 );
and \U$28380 ( \28723 , \28712 , \28722 );
and \U$28381 ( \28724 , \28702 , \28711 );
or \U$28382 ( \28725 , \28723 , \28724 );
xor \U$28383 ( \28726 , \28693 , \28725 );
not \U$28384 ( \28727 , \9320 );
not \U$28385 ( \28728 , RI9872568_156);
not \U$28386 ( \28729 , \8668 );
or \U$28387 ( \28730 , \28728 , \28729 );
or \U$28388 ( \28731 , \8857 , RI9872568_156);
nand \U$28389 ( \28732 , \28730 , \28731 );
not \U$28390 ( \28733 , \28732 );
or \U$28391 ( \28734 , \28727 , \28733 );
nand \U$28392 ( \28735 , \28431 , \5653 );
nand \U$28393 ( \28736 , \28734 , \28735 );
not \U$28394 ( \28737 , \13017 );
not \U$28395 ( \28738 , \28247 );
or \U$28396 ( \28739 , \28737 , \28738 );
not \U$28397 ( \28740 , \15389 );
not \U$28398 ( \28741 , \7003 );
or \U$28399 ( \28742 , \28740 , \28741 );
nand \U$28400 ( \28743 , \8948 , RI9872a18_166);
nand \U$28401 ( \28744 , \28742 , \28743 );
nand \U$28402 ( \28745 , \28744 , \8028 );
nand \U$28403 ( \28746 , \28739 , \28745 );
xor \U$28404 ( \28747 , \28736 , \28746 );
not \U$28405 ( \28748 , \28262 );
not \U$28406 ( \28749 , \9214 );
or \U$28407 ( \28750 , \28748 , \28749 );
and \U$28408 ( \28751 , RI9872b80_169, \8053 );
not \U$28409 ( \28752 , RI9872b80_169);
and \U$28410 ( \28753 , \28752 , \12802 );
or \U$28411 ( \28754 , \28751 , \28753 );
nand \U$28412 ( \28755 , \28754 , \9196 );
nand \U$28413 ( \28756 , \28750 , \28755 );
and \U$28414 ( \28757 , \28747 , \28756 );
and \U$28415 ( \28758 , \28736 , \28746 );
or \U$28416 ( \28759 , \28757 , \28758 );
and \U$28417 ( \28760 , \28726 , \28759 );
and \U$28418 ( \28761 , \28693 , \28725 );
or \U$28419 ( \28762 , \28760 , \28761 );
xor \U$28420 ( \28763 , \28626 , \28762 );
not \U$28421 ( \28764 , \12868 );
not \U$28422 ( \28765 , \28342 );
or \U$28423 ( \28766 , \28764 , \28765 );
and \U$28424 ( \28767 , RI98730a8_180, \8785 );
not \U$28425 ( \28768 , RI98730a8_180);
and \U$28426 ( \28769 , \28768 , \2947 );
nor \U$28427 ( \28770 , \28767 , \28769 );
nand \U$28428 ( \28771 , \28770 , \13020 );
nand \U$28429 ( \28772 , \28766 , \28771 );
not \U$28430 ( \28773 , \28772 );
not \U$28431 ( \28774 , \22167 );
not \U$28432 ( \28775 , \28293 );
or \U$28433 ( \28776 , \28774 , \28775 );
and \U$28434 ( \28777 , RI9872bf8_170, \6481 );
not \U$28435 ( \28778 , RI9872bf8_170);
and \U$28436 ( \28779 , \28778 , \5766 );
or \U$28437 ( \28780 , \28777 , \28779 );
nand \U$28438 ( \28781 , \28780 , \9670 );
nand \U$28439 ( \28782 , \28776 , \28781 );
not \U$28440 ( \28783 , \28782 );
nand \U$28441 ( \28784 , \28773 , \28783 );
not \U$28442 ( \28785 , \28784 );
not \U$28443 ( \28786 , \22670 );
not \U$28444 ( \28787 , \28302 );
or \U$28445 ( \28788 , \28786 , \28787 );
not \U$28446 ( \28789 , RI9873210_183);
and \U$28447 ( \28790 , \1485 , \28789 );
not \U$28448 ( \28791 , \1485 );
and \U$28449 ( \28792 , \28791 , RI9873210_183);
nor \U$28450 ( \28793 , \28790 , \28792 );
nand \U$28451 ( \28794 , \28793 , \18957 );
nand \U$28452 ( \28795 , \28788 , \28794 );
not \U$28453 ( \28796 , \28795 );
or \U$28454 ( \28797 , \28785 , \28796 );
nand \U$28455 ( \28798 , \28772 , \28782 );
nand \U$28456 ( \28799 , \28797 , \28798 );
not \U$28457 ( \28800 , \9527 );
not \U$28458 ( \28801 , RI9872f40_177);
not \U$28459 ( \28802 , \12616 );
or \U$28460 ( \28803 , \28801 , \28802 );
or \U$28461 ( \28804 , \4176 , RI9872f40_177);
nand \U$28462 ( \28805 , \28803 , \28804 );
not \U$28463 ( \28806 , \28805 );
or \U$28464 ( \28807 , \28800 , \28806 );
nand \U$28465 ( \28808 , \28130 , \13214 );
nand \U$28466 ( \28809 , \28807 , \28808 );
not \U$28467 ( \28810 , \28809 );
buf \U$28468 ( \28811 , \19045 );
not \U$28469 ( \28812 , \28811 );
not \U$28470 ( \28813 , \28227 );
or \U$28471 ( \28814 , \28812 , \28813 );
and \U$28472 ( \28815 , RI98734e0_189, \22615 );
not \U$28473 ( \28816 , RI98734e0_189);
and \U$28474 ( \28817 , \28816 , \17363 );
nor \U$28475 ( \28818 , \28815 , \28817 );
nand \U$28476 ( \28819 , \28818 , \19244 );
nand \U$28477 ( \28820 , \28814 , \28819 );
not \U$28478 ( \28821 , \791 );
not \U$28479 ( \28822 , RI98719b0_131);
not \U$28480 ( \28823 , \25380 );
or \U$28481 ( \28824 , \28822 , \28823 );
or \U$28482 ( \28825 , \20765 , RI98719b0_131);
nand \U$28483 ( \28826 , \28824 , \28825 );
not \U$28484 ( \28827 , \28826 );
or \U$28485 ( \28828 , \28821 , \28827 );
not \U$28486 ( \28829 , \28511 );
nand \U$28487 ( \28830 , \28829 , \796 );
nand \U$28488 ( \28831 , \28828 , \28830 );
not \U$28489 ( \28832 , \28831 );
not \U$28490 ( \28833 , \1289 );
and \U$28491 ( \28834 , \21779 , \28833 );
nand \U$28492 ( \28835 , \1287 , RI9871b18_134);
nor \U$28493 ( \28836 , \28834 , \28835 );
not \U$28494 ( \28837 , \1290 );
not \U$28495 ( \28838 , \28673 );
or \U$28496 ( \28839 , \28837 , \28838 );
xor \U$28497 ( \28840 , \18705 , RI9871b18_134);
nand \U$28498 ( \28841 , \28840 , \1291 );
nand \U$28499 ( \28842 , \28839 , \28841 );
and \U$28500 ( \28843 , \28836 , \28842 );
not \U$28501 ( \28844 , \1083 );
and \U$28502 ( \28845 , \22285 , RI98718c0_129);
not \U$28503 ( \28846 , \22285 );
and \U$28504 ( \28847 , \28846 , \1111 );
nor \U$28505 ( \28848 , \28845 , \28847 );
not \U$28506 ( \28849 , \28848 );
or \U$28507 ( \28850 , \28844 , \28849 );
nand \U$28508 ( \28851 , \28196 , \1134 );
nand \U$28509 ( \28852 , \28850 , \28851 );
xor \U$28510 ( \28853 , \28843 , \28852 );
not \U$28511 ( \28854 , \28853 );
or \U$28512 ( \28855 , \28832 , \28854 );
nand \U$28513 ( \28856 , \28852 , \28843 );
nand \U$28514 ( \28857 , \28855 , \28856 );
xor \U$28515 ( \28858 , \28820 , \28857 );
not \U$28516 ( \28859 , \28858 );
or \U$28517 ( \28860 , \28810 , \28859 );
nand \U$28518 ( \28861 , \28820 , \28857 );
nand \U$28519 ( \28862 , \28860 , \28861 );
xor \U$28520 ( \28863 , \28799 , \28862 );
not \U$28521 ( \28864 , \8801 );
not \U$28522 ( \28865 , \28312 );
or \U$28523 ( \28866 , \28864 , \28865 );
and \U$28524 ( \28867 , RI9872d60_173, \4985 );
not \U$28525 ( \28868 , RI9872d60_173);
and \U$28526 ( \28869 , \28868 , \5739 );
or \U$28527 ( \28870 , \28867 , \28869 );
nand \U$28528 ( \28871 , \28870 , \8819 );
nand \U$28529 ( \28872 , \28866 , \28871 );
not \U$28530 ( \28873 , \28872 );
not \U$28531 ( \28874 , \17528 );
not \U$28532 ( \28875 , \28157 );
or \U$28533 ( \28876 , \28874 , \28875 );
not \U$28534 ( \28877 , RI9873288_184);
not \U$28535 ( \28878 , \9263 );
or \U$28536 ( \28879 , \28877 , \28878 );
or \U$28537 ( \28880 , \20638 , RI9873288_184);
nand \U$28538 ( \28881 , \28879 , \28880 );
nand \U$28539 ( \28882 , \28881 , \19641 );
nand \U$28540 ( \28883 , \28876 , \28882 );
not \U$28541 ( \28884 , \10332 );
not \U$28542 ( \28885 , \28141 );
or \U$28543 ( \28886 , \28884 , \28885 );
and \U$28544 ( \28887 , \9694 , \4711 );
not \U$28545 ( \28888 , \9694 );
and \U$28546 ( \28889 , \28888 , \5623 );
nor \U$28547 ( \28890 , \28887 , \28889 );
nand \U$28548 ( \28891 , \28890 , \18562 );
nand \U$28549 ( \28892 , \28886 , \28891 );
and \U$28550 ( \28893 , \28883 , \28892 );
not \U$28551 ( \28894 , \28883 );
not \U$28552 ( \28895 , \28892 );
and \U$28553 ( \28896 , \28894 , \28895 );
nor \U$28554 ( \28897 , \28893 , \28896 );
not \U$28555 ( \28898 , \28897 );
or \U$28556 ( \28899 , \28873 , \28898 );
buf \U$28557 ( \28900 , \28883 );
nand \U$28558 ( \28901 , \28900 , \28892 );
nand \U$28559 ( \28902 , \28899 , \28901 );
and \U$28560 ( \28903 , \28863 , \28902 );
and \U$28561 ( \28904 , \28799 , \28862 );
or \U$28562 ( \28905 , \28903 , \28904 );
and \U$28563 ( \28906 , \28763 , \28905 );
and \U$28564 ( \28907 , \28626 , \28762 );
or \U$28565 ( \28908 , \28906 , \28907 );
not \U$28566 ( \28909 , \28908 );
and \U$28567 ( \28910 , \28624 , \28909 );
and \U$28568 ( \28911 , \28621 , \28623 );
or \U$28569 ( \28912 , \28910 , \28911 );
not \U$28570 ( \28913 , \28912 );
not \U$28571 ( \28914 , \28913 );
xor \U$28572 ( \28915 , \27636 , \27642 );
xor \U$28573 ( \28916 , \28915 , \27652 );
not \U$28574 ( \28917 , \28916 );
and \U$28575 ( \28918 , \28375 , \28399 );
not \U$28576 ( \28919 , \28375 );
and \U$28577 ( \28920 , \28919 , \28384 );
or \U$28578 ( \28921 , \28918 , \28920 );
xnor \U$28579 ( \28922 , \28921 , \28396 );
not \U$28580 ( \28923 , \28922 );
and \U$28581 ( \28924 , RI98729a0_165, \12727 );
not \U$28582 ( \28925 , RI98729a0_165);
and \U$28583 ( \28926 , \28925 , \8333 );
nor \U$28584 ( \28927 , \28924 , \28926 );
not \U$28585 ( \28928 , \28927 );
not \U$28586 ( \28929 , \7326 );
or \U$28587 ( \28930 , \28928 , \28929 );
nand \U$28588 ( \28931 , \28239 , \7338 );
nand \U$28589 ( \28932 , \28930 , \28931 );
not \U$28590 ( \28933 , \28198 );
not \U$28591 ( \28934 , \28184 );
and \U$28592 ( \28935 , \28933 , \28934 );
and \U$28593 ( \28936 , \28198 , \28184 );
nor \U$28594 ( \28937 , \28935 , \28936 );
not \U$28595 ( \28938 , \28937 );
or \U$28596 ( \28939 , \28932 , \28938 );
not \U$28597 ( \28940 , \6610 );
not \U$28598 ( \28941 , \28212 );
or \U$28599 ( \28942 , \28940 , \28941 );
not \U$28600 ( \28943 , \6283 );
and \U$28601 ( \28944 , \5632 , \20430 );
not \U$28602 ( \28945 , \5632 );
and \U$28603 ( \28946 , \28945 , \8877 );
nor \U$28604 ( \28947 , \28944 , \28946 );
nand \U$28605 ( \28948 , \28943 , \28947 );
nand \U$28606 ( \28949 , \28942 , \28948 );
nand \U$28607 ( \28950 , \28939 , \28949 );
nand \U$28608 ( \28951 , \28932 , \28938 );
nand \U$28609 ( \28952 , \28950 , \28951 );
xor \U$28610 ( \28953 , \27577 , \27602 );
xor \U$28611 ( \28954 , \28952 , \28953 );
not \U$28612 ( \28955 , \28954 );
or \U$28613 ( \28956 , \28923 , \28955 );
not \U$28614 ( \28957 , \28951 );
not \U$28615 ( \28958 , \28950 );
or \U$28616 ( \28959 , \28957 , \28958 );
nand \U$28617 ( \28960 , \28959 , \28953 );
nand \U$28618 ( \28961 , \28956 , \28960 );
not \U$28619 ( \28962 , \28961 );
not \U$28620 ( \28963 , \28962 );
nand \U$28621 ( \28964 , \27620 , \27615 );
not \U$28622 ( \28965 , \27613 );
and \U$28623 ( \28966 , \28964 , \28965 );
not \U$28624 ( \28967 , \28964 );
and \U$28625 ( \28968 , \28967 , \27613 );
or \U$28626 ( \28969 , \28966 , \28968 );
not \U$28627 ( \28970 , \28969 );
or \U$28628 ( \28971 , \28963 , \28970 );
or \U$28629 ( \28972 , \28969 , \28962 );
nand \U$28630 ( \28973 , \28971 , \28972 );
not \U$28631 ( \28974 , \28973 );
or \U$28632 ( \28975 , \28917 , \28974 );
nand \U$28633 ( \28976 , \28969 , \28961 );
nand \U$28634 ( \28977 , \28975 , \28976 );
not \U$28635 ( \28978 , \28977 );
xor \U$28636 ( \28979 , \27993 , \27994 );
xor \U$28637 ( \28980 , \28979 , \28028 );
not \U$28638 ( \28981 , \28980 );
or \U$28639 ( \28982 , \28978 , \28981 );
or \U$28640 ( \28983 , \28980 , \28977 );
xor \U$28641 ( \28984 , \27938 , \27980 );
nand \U$28642 ( \28985 , \28983 , \28984 );
nand \U$28643 ( \28986 , \28982 , \28985 );
xor \U$28644 ( \28987 , \28461 , \28986 );
xnor \U$28645 ( \28988 , \28987 , \28359 );
not \U$28646 ( \28989 , \28988 );
or \U$28647 ( \28990 , \28914 , \28989 );
xor \U$28648 ( \28991 , \28462 , \28359 );
nand \U$28649 ( \28992 , \28991 , \28986 );
nand \U$28650 ( \28993 , \28990 , \28992 );
not \U$28651 ( \28994 , \28993 );
not \U$28652 ( \28995 , \28994 );
or \U$28653 ( \28996 , \28619 , \28995 );
xor \U$28654 ( \28997 , \28353 , \28122 );
xor \U$28655 ( \28998 , \28478 , \28574 );
xor \U$28656 ( \28999 , \28998 , \28576 );
xor \U$28657 ( \29000 , \28997 , \28999 );
xor \U$28658 ( \29001 , \28490 , \28572 );
xor \U$28659 ( \29002 , \29001 , \28493 );
not \U$28660 ( \29003 , \29002 );
not \U$28661 ( \29004 , \28482 );
not \U$28662 ( \29005 , \28480 );
or \U$28663 ( \29006 , \29004 , \29005 );
or \U$28664 ( \29007 , \28480 , \28482 );
nand \U$28665 ( \29008 , \29006 , \29007 );
not \U$28666 ( \29009 , \29008 );
not \U$28667 ( \29010 , \29009 );
not \U$28668 ( \29011 , \28487 );
or \U$28669 ( \29012 , \29010 , \29011 );
nand \U$28670 ( \29013 , \28486 , \29008 );
nand \U$28671 ( \29014 , \29012 , \29013 );
not \U$28672 ( \29015 , \29014 );
xor \U$28673 ( \29016 , \28327 , \28325 );
xnor \U$28674 ( \29017 , \29016 , \28347 );
nand \U$28675 ( \29018 , \29015 , \29017 );
xor \U$28676 ( \29019 , \28229 , \28218 );
xor \U$28677 ( \29020 , \28264 , \28252 );
xor \U$28678 ( \29021 , \29019 , \29020 );
not \U$28679 ( \29022 , \9937 );
not \U$28680 ( \29023 , \28544 );
or \U$28681 ( \29024 , \29022 , \29023 );
not \U$28682 ( \29025 , \3537 );
not \U$28683 ( \29026 , RI9873030_179);
and \U$28684 ( \29027 , \29025 , \29026 );
and \U$28685 ( \29028 , \6718 , RI9873030_179);
nor \U$28686 ( \29029 , \29027 , \29028 );
nand \U$28687 ( \29030 , \29029 , \9952 );
nand \U$28688 ( \29031 , \29024 , \29030 );
not \U$28689 ( \29032 , \29031 );
not \U$28690 ( \29033 , RI9873648_192);
not \U$28691 ( \29034 , \28335 );
or \U$28692 ( \29035 , \29033 , \29034 );
not \U$28693 ( \29036 , \18239 );
not \U$28694 ( \29037 , \943 );
or \U$28695 ( \29038 , \29036 , \29037 );
or \U$28696 ( \29039 , \11283 , \18239 );
nand \U$28697 ( \29040 , \29038 , \29039 );
nand \U$28698 ( \29041 , \29040 , \20626 );
nand \U$28699 ( \29042 , \29035 , \29041 );
not \U$28700 ( \29043 , \17263 );
not \U$28701 ( \29044 , \28558 );
or \U$28702 ( \29045 , \29043 , \29044 );
and \U$28703 ( \29046 , RI98733f0_187, \1061 );
not \U$28704 ( \29047 , RI98733f0_187);
and \U$28705 ( \29048 , \29047 , \23043 );
nor \U$28706 ( \29049 , \29046 , \29048 );
nand \U$28707 ( \29050 , \29049 , \17252 );
nand \U$28708 ( \29051 , \29045 , \29050 );
xor \U$28709 ( \29052 , \29042 , \29051 );
not \U$28710 ( \29053 , \29052 );
or \U$28711 ( \29054 , \29032 , \29053 );
nand \U$28712 ( \29055 , \29042 , \29051 );
nand \U$28713 ( \29056 , \29054 , \29055 );
and \U$28714 ( \29057 , \29021 , \29056 );
and \U$28715 ( \29058 , \29019 , \29020 );
or \U$28716 ( \29059 , \29057 , \29058 );
and \U$28717 ( \29060 , \29018 , \29059 );
not \U$28718 ( \29061 , \29014 );
nor \U$28719 ( \29062 , \29017 , \29061 );
nor \U$28720 ( \29063 , \29060 , \29062 );
not \U$28721 ( \29064 , \29063 );
xor \U$28722 ( \29065 , \28124 , \28284 );
xor \U$28723 ( \29066 , \29065 , \28350 );
not \U$28724 ( \29067 , \29066 );
or \U$28725 ( \29068 , \29064 , \29067 );
or \U$28726 ( \29069 , \29063 , \29066 );
nand \U$28727 ( \29070 , \29068 , \29069 );
not \U$28728 ( \29071 , \29070 );
or \U$28729 ( \29072 , \29003 , \29071 );
not \U$28730 ( \29073 , \29063 );
nand \U$28731 ( \29074 , \29073 , \29066 );
nand \U$28732 ( \29075 , \29072 , \29074 );
and \U$28733 ( \29076 , \29000 , \29075 );
and \U$28734 ( \29077 , \28997 , \28999 );
or \U$28735 ( \29078 , \29076 , \29077 );
nand \U$28736 ( \29079 , \28996 , \29078 );
not \U$28737 ( \29080 , \28618 );
nand \U$28738 ( \29081 , \28993 , \29080 );
and \U$28739 ( \29082 , \29079 , \29081 );
xor \U$28740 ( \29083 , \28616 , \29082 );
xor \U$28741 ( \29084 , \28469 , \28471 );
xor \U$28742 ( \29085 , \29084 , \28586 );
and \U$28743 ( \29086 , \29083 , \29085 );
and \U$28744 ( \29087 , \28616 , \29082 );
or \U$28745 ( \29088 , \29086 , \29087 );
nand \U$28746 ( \29089 , \28609 , \29088 );
nand \U$28747 ( \29090 , \28607 , \29089 );
nor \U$28748 ( \29091 , \28599 , \29090 );
xor \U$28749 ( \29092 , \28997 , \28999 );
xor \U$28750 ( \29093 , \29092 , \29075 );
xor \U$28751 ( \29094 , \28412 , \28422 );
xor \U$28752 ( \29095 , \29094 , \28435 );
not \U$28753 ( \29096 , \29095 );
not \U$28754 ( \29097 , \28161 );
and \U$28755 ( \29098 , \28152 , \29097 );
not \U$28756 ( \29099 , \28152 );
and \U$28757 ( \29100 , \29099 , \28161 );
nor \U$28758 ( \29101 , \29098 , \29100 );
nand \U$28759 ( \29102 , \29096 , \29101 );
and \U$28760 ( \29103 , \28560 , \28536 );
not \U$28761 ( \29104 , \28560 );
and \U$28762 ( \29105 , \29104 , \28537 );
nor \U$28763 ( \29106 , \29103 , \29105 );
not \U$28764 ( \29107 , \29106 );
not \U$28765 ( \29108 , \28549 );
and \U$28766 ( \29109 , \29107 , \29108 );
and \U$28767 ( \29110 , \29106 , \28549 );
nor \U$28768 ( \29111 , \29109 , \29110 );
not \U$28769 ( \29112 , \29111 );
and \U$28770 ( \29113 , \29102 , \29112 );
not \U$28771 ( \29114 , \29095 );
nor \U$28772 ( \29115 , \29114 , \29101 );
nor \U$28773 ( \29116 , \29113 , \29115 );
not \U$28774 ( \29117 , \29116 );
not \U$28775 ( \29118 , \29117 );
xor \U$28776 ( \29119 , \28295 , \28319 );
xnor \U$28777 ( \29120 , \29119 , \28306 );
not \U$28778 ( \29121 , \3163 );
not \U$28779 ( \29122 , RI9872310_151);
not \U$28780 ( \29123 , \13268 );
or \U$28781 ( \29124 , \29122 , \29123 );
or \U$28782 ( \29125 , \12773 , RI9872310_151);
nand \U$28783 ( \29126 , \29124 , \29125 );
not \U$28784 ( \29127 , \29126 );
or \U$28785 ( \29128 , \29121 , \29127 );
nand \U$28786 ( \29129 , \28632 , \3170 );
nand \U$28787 ( \29130 , \29128 , \29129 );
not \U$28788 ( \29131 , \2087 );
not \U$28789 ( \29132 , \28504 );
or \U$28790 ( \29133 , \29131 , \29132 );
not \U$28791 ( \29134 , RI9871aa0_133);
not \U$28792 ( \29135 , \18350 );
or \U$28793 ( \29136 , \29134 , \29135 );
not \U$28794 ( \29137 , \13623 );
or \U$28795 ( \29138 , \29137 , RI9871aa0_133);
nand \U$28796 ( \29139 , \29136 , \29138 );
nand \U$28797 ( \29140 , \29139 , \2071 );
nand \U$28798 ( \29141 , \29133 , \29140 );
nor \U$28799 ( \29142 , \29130 , \29141 );
not \U$28800 ( \29143 , \29142 );
not \U$28801 ( \29144 , \29143 );
not \U$28802 ( \29145 , \7188 );
not \U$28803 ( \29146 , \28732 );
or \U$28804 ( \29147 , \29145 , \29146 );
not \U$28805 ( \29148 , RI9872568_156);
not \U$28806 ( \29149 , \8650 );
or \U$28807 ( \29150 , \29148 , \29149 );
or \U$28808 ( \29151 , \11406 , RI9872568_156);
nand \U$28809 ( \29152 , \29150 , \29151 );
nand \U$28810 ( \29153 , \29152 , \9320 );
nand \U$28811 ( \29154 , \29147 , \29153 );
not \U$28812 ( \29155 , \29154 );
or \U$28813 ( \29156 , \29144 , \29155 );
nand \U$28814 ( \29157 , \29130 , \29141 );
nand \U$28815 ( \29158 , \29156 , \29157 );
not \U$28816 ( \29159 , \29158 );
xor \U$28817 ( \29160 , \28689 , \28636 );
not \U$28818 ( \29161 , \8790 );
not \U$28819 ( \29162 , RI98725e0_157);
not \U$28820 ( \29163 , \11371 );
or \U$28821 ( \29164 , \29162 , \29163 );
or \U$28822 ( \29165 , \9114 , RI98725e0_157);
nand \U$28823 ( \29166 , \29164 , \29165 );
not \U$28824 ( \29167 , \29166 );
or \U$28825 ( \29168 , \29161 , \29167 );
nand \U$28826 ( \29169 , \28700 , \4084 );
nand \U$28827 ( \29170 , \29168 , \29169 );
not \U$28828 ( \29171 , \29170 );
not \U$28829 ( \29172 , \3465 );
and \U$28830 ( \29173 , RI98726d0_159, \10064 );
not \U$28831 ( \29174 , RI98726d0_159);
and \U$28832 ( \29175 , \29174 , \27587 );
or \U$28833 ( \29176 , \29173 , \29175 );
not \U$28834 ( \29177 , \29176 );
or \U$28835 ( \29178 , \29172 , \29177 );
nand \U$28836 ( \29179 , \28523 , \3467 );
nand \U$28837 ( \29180 , \29178 , \29179 );
xor \U$28838 ( \29181 , \28661 , \28681 );
xor \U$28839 ( \29182 , \29180 , \29181 );
not \U$28840 ( \29183 , \29182 );
or \U$28841 ( \29184 , \29171 , \29183 );
nand \U$28842 ( \29185 , \29180 , \29181 );
nand \U$28843 ( \29186 , \29184 , \29185 );
xor \U$28844 ( \29187 , \29160 , \29186 );
not \U$28845 ( \29188 , \29187 );
or \U$28846 ( \29189 , \29159 , \29188 );
nand \U$28847 ( \29190 , \29186 , \29160 );
nand \U$28848 ( \29191 , \29189 , \29190 );
or \U$28849 ( \29192 , \29120 , \29191 );
xor \U$28850 ( \29193 , \28330 , \28344 );
xnor \U$28851 ( \29194 , \29193 , \28337 );
nand \U$28852 ( \29195 , \29192 , \29194 );
nand \U$28853 ( \29196 , \29120 , \29191 );
nand \U$28854 ( \29197 , \29195 , \29196 );
not \U$28855 ( \29198 , \29197 );
not \U$28856 ( \29199 , \28163 );
not \U$28857 ( \29200 , \29199 );
not \U$28858 ( \29201 , \28277 );
or \U$28859 ( \29202 , \29200 , \29201 );
or \U$28860 ( \29203 , \28277 , \29199 );
nand \U$28861 ( \29204 , \29202 , \29203 );
not \U$28862 ( \29205 , \29204 );
not \U$28863 ( \29206 , \29205 );
or \U$28864 ( \29207 , \29198 , \29206 );
or \U$28865 ( \29208 , \29205 , \29197 );
nand \U$28866 ( \29209 , \29207 , \29208 );
not \U$28867 ( \29210 , \29209 );
or \U$28868 ( \29211 , \29118 , \29210 );
not \U$28869 ( \29212 , \29205 );
nand \U$28870 ( \29213 , \29212 , \29197 );
nand \U$28871 ( \29214 , \29211 , \29213 );
and \U$28872 ( \29215 , \28949 , \28937 );
not \U$28873 ( \29216 , \28949 );
and \U$28874 ( \29217 , \29216 , \28938 );
nor \U$28875 ( \29218 , \29215 , \29217 );
xnor \U$28876 ( \29219 , \28932 , \29218 );
xor \U$28877 ( \29220 , \28702 , \28711 );
xor \U$28878 ( \29221 , \29220 , \28722 );
xor \U$28879 ( \29222 , \29219 , \29221 );
xor \U$28880 ( \29223 , \28736 , \28746 );
xor \U$28881 ( \29224 , \29223 , \28756 );
and \U$28882 ( \29225 , \29222 , \29224 );
and \U$28883 ( \29226 , \29219 , \29221 );
or \U$28884 ( \29227 , \29225 , \29226 );
not \U$28885 ( \29228 , \29227 );
xor \U$28886 ( \29229 , \28506 , \28531 );
not \U$28887 ( \29230 , \4922 );
not \U$28888 ( \29231 , \28709 );
or \U$28889 ( \29232 , \29230 , \29231 );
not \U$28890 ( \29233 , \7993 );
not \U$28891 ( \29234 , \8694 );
or \U$28892 ( \29235 , \29233 , \29234 );
or \U$28893 ( \29236 , \18329 , \4902 );
nand \U$28894 ( \29237 , \29235 , \29236 );
nand \U$28895 ( \29238 , \29237 , \4918 );
nand \U$28896 ( \29239 , \29232 , \29238 );
not \U$28897 ( \29240 , \29239 );
and \U$28898 ( \29241 , \22459 , \28720 );
not \U$28899 ( \29242 , RI9872478_154);
not \U$28900 ( \29243 , \8554 );
or \U$28901 ( \29244 , \29242 , \29243 );
or \U$28902 ( \29245 , \8554 , RI9872478_154);
nand \U$28903 ( \29246 , \29244 , \29245 );
and \U$28904 ( \29247 , \29246 , \5034 );
nor \U$28905 ( \29248 , \29241 , \29247 );
not \U$28906 ( \29249 , \29248 );
or \U$28907 ( \29250 , \29240 , \29249 );
or \U$28908 ( \29251 , \29248 , \29239 );
nand \U$28909 ( \29252 , \29250 , \29251 );
not \U$28910 ( \29253 , \29252 );
not \U$28911 ( \29254 , \9249 );
and \U$28912 ( \29255 , RI9872bf8_170, \18808 );
not \U$28913 ( \29256 , RI9872bf8_170);
and \U$28914 ( \29257 , \29256 , \7111 );
nor \U$28915 ( \29258 , \29255 , \29257 );
not \U$28916 ( \29259 , \29258 );
or \U$28917 ( \29260 , \29254 , \29259 );
nand \U$28918 ( \29261 , \28780 , \9668 );
nand \U$28919 ( \29262 , \29260 , \29261 );
not \U$28920 ( \29263 , \29262 );
or \U$28921 ( \29264 , \29253 , \29263 );
not \U$28922 ( \29265 , \29248 );
nand \U$28923 ( \29266 , \29265 , \29239 );
nand \U$28924 ( \29267 , \29264 , \29266 );
xor \U$28925 ( \29268 , \29229 , \29267 );
not \U$28926 ( \29269 , \29268 );
not \U$28927 ( \29270 , \9072 );
not \U$28928 ( \29271 , \28744 );
or \U$28929 ( \29272 , \29270 , \29271 );
not \U$28930 ( \29273 , RI9872a18_166);
not \U$28931 ( \29274 , \7466 );
or \U$28932 ( \29275 , \29273 , \29274 );
or \U$28933 ( \29276 , \13824 , RI9872a18_166);
nand \U$28934 ( \29277 , \29275 , \29276 );
nand \U$28935 ( \29278 , \29277 , \8028 );
nand \U$28936 ( \29279 , \29272 , \29278 );
not \U$28937 ( \29280 , \9196 );
not \U$28938 ( \29281 , \11688 );
not \U$28939 ( \29282 , \7905 );
or \U$28940 ( \29283 , \29281 , \29282 );
nand \U$28941 ( \29284 , \6529 , RI9872b80_169);
nand \U$28942 ( \29285 , \29283 , \29284 );
not \U$28943 ( \29286 , \29285 );
or \U$28944 ( \29287 , \29280 , \29286 );
nand \U$28945 ( \29288 , \28754 , \9214 );
nand \U$28946 ( \29289 , \29287 , \29288 );
xor \U$28947 ( \29290 , \29279 , \29289 );
not \U$28948 ( \29291 , \29290 );
not \U$28949 ( \29292 , \7325 );
and \U$28950 ( \29293 , \8074 , \7333 );
not \U$28951 ( \29294 , \8074 );
and \U$28952 ( \29295 , \29294 , RI98729a0_165);
nor \U$28953 ( \29296 , \29293 , \29295 );
not \U$28954 ( \29297 , \29296 );
or \U$28955 ( \29298 , \29292 , \29297 );
nand \U$28956 ( \29299 , \28927 , \7338 );
nand \U$28957 ( \29300 , \29298 , \29299 );
buf \U$28958 ( \29301 , \29300 );
not \U$28959 ( \29302 , \29301 );
or \U$28960 ( \29303 , \29291 , \29302 );
nand \U$28961 ( \29304 , \29289 , \29279 );
nand \U$28962 ( \29305 , \29303 , \29304 );
not \U$28963 ( \29306 , \29305 );
or \U$28964 ( \29307 , \29269 , \29306 );
nand \U$28965 ( \29308 , \29267 , \29229 );
nand \U$28966 ( \29309 , \29307 , \29308 );
xor \U$28967 ( \29310 , \28693 , \28725 );
xor \U$28968 ( \29311 , \29310 , \28759 );
xor \U$28969 ( \29312 , \29309 , \29311 );
not \U$28970 ( \29313 , \29312 );
or \U$28971 ( \29314 , \29228 , \29313 );
nand \U$28972 ( \29315 , \29311 , \29309 );
nand \U$28973 ( \29316 , \29314 , \29315 );
not \U$28974 ( \29317 , \28961 );
xor \U$28975 ( \29318 , \28916 , \29317 );
xnor \U$28976 ( \29319 , \29318 , \28969 );
or \U$28977 ( \29320 , \29316 , \29319 );
xor \U$28978 ( \29321 , \28564 , \28566 );
xor \U$28979 ( \29322 , \29321 , \28569 );
nand \U$28980 ( \29323 , \29320 , \29322 );
nand \U$28981 ( \29324 , \29316 , \29319 );
nand \U$28982 ( \29325 , \29323 , \29324 );
xor \U$28983 ( \29326 , \29214 , \29325 );
xor \U$28984 ( \29327 , \28984 , \28980 );
xor \U$28985 ( \29328 , \29327 , \28977 );
xor \U$28986 ( \29329 , \29326 , \29328 );
and \U$28987 ( \29330 , \29059 , \29014 );
not \U$28988 ( \29331 , \29059 );
and \U$28989 ( \29332 , \29331 , \29061 );
nor \U$28990 ( \29333 , \29330 , \29332 );
not \U$28991 ( \29334 , \29333 );
not \U$28992 ( \29335 , \29017 );
or \U$28993 ( \29336 , \29334 , \29335 );
not \U$28994 ( \29337 , \29017 );
not \U$28995 ( \29338 , \29333 );
nand \U$28996 ( \29339 , \29337 , \29338 );
nand \U$28997 ( \29340 , \29336 , \29339 );
not \U$28998 ( \29341 , \29340 );
xor \U$28999 ( \29342 , \29305 , \29268 );
not \U$29000 ( \29343 , \29342 );
not \U$29001 ( \29344 , \4922 );
not \U$29002 ( \29345 , \29237 );
or \U$29003 ( \29346 , \29344 , \29345 );
not \U$29004 ( \29347 , RI9872388_152);
not \U$29005 ( \29348 , \9849 );
or \U$29006 ( \29349 , \29347 , \29348 );
or \U$29007 ( \29350 , \12460 , RI9872388_152);
nand \U$29008 ( \29351 , \29349 , \29350 );
nand \U$29009 ( \29352 , \29351 , \4918 );
nand \U$29010 ( \29353 , \29346 , \29352 );
not \U$29011 ( \29354 , \22459 );
not \U$29012 ( \29355 , \29246 );
or \U$29013 ( \29356 , \29354 , \29355 );
and \U$29014 ( \29357 , RI9872478_154, \8722 );
not \U$29015 ( \29358 , RI9872478_154);
and \U$29016 ( \29359 , \29358 , \20385 );
nor \U$29017 ( \29360 , \29357 , \29359 );
nand \U$29018 ( \29361 , \29360 , \5034 );
nand \U$29019 ( \29362 , \29356 , \29361 );
xor \U$29020 ( \29363 , \29353 , \29362 );
not \U$29021 ( \29364 , \5653 );
not \U$29022 ( \29365 , \29152 );
or \U$29023 ( \29366 , \29364 , \29365 );
not \U$29024 ( \29367 , \5648 );
not \U$29025 ( \29368 , \12848 );
or \U$29026 ( \29369 , \29367 , \29368 );
or \U$29027 ( \29370 , \18312 , \5648 );
nand \U$29028 ( \29371 , \29369 , \29370 );
nand \U$29029 ( \29372 , \29371 , \6063 );
nand \U$29030 ( \29373 , \29366 , \29372 );
and \U$29031 ( \29374 , \29363 , \29373 );
and \U$29032 ( \29375 , \29353 , \29362 );
or \U$29033 ( \29376 , \29374 , \29375 );
not \U$29034 ( \29377 , \29376 );
not \U$29035 ( \29378 , \796 );
not \U$29036 ( \29379 , \28826 );
or \U$29037 ( \29380 , \29378 , \29379 );
and \U$29038 ( \29381 , RI98719b0_131, \17911 );
not \U$29039 ( \29382 , RI98719b0_131);
and \U$29040 ( \29383 , \29382 , \18841 );
or \U$29041 ( \29384 , \29381 , \29383 );
nand \U$29042 ( \29385 , \29384 , \791 );
nand \U$29043 ( \29386 , \29380 , \29385 );
not \U$29044 ( \29387 , \29386 );
xor \U$29045 ( \29388 , \28836 , \28842 );
not \U$29046 ( \29389 , \1427 );
not \U$29047 ( \29390 , \28659 );
or \U$29048 ( \29391 , \29389 , \29390 );
not \U$29049 ( \29392 , RI9871c08_136);
not \U$29050 ( \29393 , \22466 );
or \U$29051 ( \29394 , \29392 , \29393 );
nand \U$29052 ( \29395 , \24854 , \1850 );
nand \U$29053 ( \29396 , \29394 , \29395 );
nand \U$29054 ( \29397 , \29396 , \1454 );
nand \U$29055 ( \29398 , \29391 , \29397 );
xor \U$29056 ( \29399 , \29388 , \29398 );
not \U$29057 ( \29400 , \29399 );
not \U$29058 ( \29401 , \29400 );
and \U$29059 ( \29402 , \29387 , \29401 );
and \U$29060 ( \29403 , \29386 , \29400 );
nor \U$29061 ( \29404 , \29402 , \29403 );
and \U$29062 ( \29405 , RI9871aa0_133, \13861 );
not \U$29063 ( \29406 , RI9871aa0_133);
and \U$29064 ( \29407 , \29406 , \13860 );
or \U$29065 ( \29408 , \29405 , \29407 );
not \U$29066 ( \29409 , \29408 );
not \U$29067 ( \29410 , \2086 );
and \U$29068 ( \29411 , \29409 , \29410 );
not \U$29069 ( \29412 , \17003 );
and \U$29070 ( \29413 , RI9871aa0_133, \29412 );
not \U$29071 ( \29414 , RI9871aa0_133);
and \U$29072 ( \29415 , \29414 , \13933 );
or \U$29073 ( \29416 , \29413 , \29415 );
and \U$29074 ( \29417 , \29416 , \2071 );
nor \U$29075 ( \29418 , \29411 , \29417 );
not \U$29076 ( \29419 , \29418 );
or \U$29077 ( \29420 , RI98718c0_129, RI98720b8_146);
nand \U$29078 ( \29421 , \29420 , \18704 );
nand \U$29079 ( \29422 , \29421 , \2358 );
not \U$29080 ( \29423 , \29422 );
not \U$29081 ( \29424 , \1427 );
not \U$29082 ( \29425 , \1850 );
not \U$29083 ( \29426 , \28671 );
or \U$29084 ( \29427 , \29425 , \29426 );
nand \U$29085 ( \29428 , \23953 , RI9871c08_136);
nand \U$29086 ( \29429 , \29427 , \29428 );
not \U$29087 ( \29430 , \29429 );
or \U$29088 ( \29431 , \29424 , \29430 );
not \U$29089 ( \29432 , \1850 );
not \U$29090 ( \29433 , \24450 );
or \U$29091 ( \29434 , \29432 , \29433 );
or \U$29092 ( \29435 , \27523 , \1619 );
nand \U$29093 ( \29436 , \29434 , \29435 );
nand \U$29094 ( \29437 , \29436 , \1454 );
nand \U$29095 ( \29438 , \29431 , \29437 );
nand \U$29096 ( \29439 , \29423 , \29438 );
not \U$29097 ( \29440 , \29439 );
not \U$29098 ( \29441 , \791 );
and \U$29099 ( \29442 , RI98719b0_131, \25412 );
not \U$29100 ( \29443 , RI98719b0_131);
and \U$29101 ( \29444 , \29443 , \19412 );
or \U$29102 ( \29445 , \29442 , \29444 );
not \U$29103 ( \29446 , \29445 );
or \U$29104 ( \29447 , \29441 , \29446 );
nand \U$29105 ( \29448 , \29384 , \796 );
nand \U$29106 ( \29449 , \29447 , \29448 );
nand \U$29107 ( \29450 , \29440 , \29449 );
not \U$29108 ( \29451 , \29450 );
or \U$29109 ( \29452 , \29419 , \29451 );
not \U$29110 ( \29453 , \29449 );
nand \U$29111 ( \29454 , \29453 , \29439 );
nand \U$29112 ( \29455 , \29452 , \29454 );
nand \U$29113 ( \29456 , \29404 , \29455 );
not \U$29114 ( \29457 , \29456 );
not \U$29115 ( \29458 , \7338 );
not \U$29116 ( \29459 , \29296 );
or \U$29117 ( \29460 , \29458 , \29459 );
and \U$29118 ( \29461 , RI98729a0_165, \8874 );
not \U$29119 ( \29462 , RI98729a0_165);
not \U$29120 ( \29463 , \8874 );
and \U$29121 ( \29464 , \29462 , \29463 );
or \U$29122 ( \29465 , \29461 , \29464 );
nand \U$29123 ( \29466 , \29465 , \7325 );
nand \U$29124 ( \29467 , \29460 , \29466 );
not \U$29125 ( \29468 , \29467 );
or \U$29126 ( \29469 , \29457 , \29468 );
not \U$29127 ( \29470 , \29404 );
not \U$29128 ( \29471 , \29455 );
nand \U$29129 ( \29472 , \29470 , \29471 );
nand \U$29130 ( \29473 , \29469 , \29472 );
not \U$29131 ( \29474 , \29473 );
nand \U$29132 ( \29475 , \29377 , \29474 );
not \U$29133 ( \29476 , \29475 );
not \U$29134 ( \29477 , \8027 );
and \U$29135 ( \29478 , RI9872a18_166, \9898 );
not \U$29136 ( \29479 , RI9872a18_166);
and \U$29137 ( \29480 , \29479 , \8333 );
nor \U$29138 ( \29481 , \29478 , \29480 );
not \U$29139 ( \29482 , \29481 );
or \U$29140 ( \29483 , \29477 , \29482 );
nand \U$29141 ( \29484 , \29277 , \9071 );
nand \U$29142 ( \29485 , \29483 , \29484 );
not \U$29143 ( \29486 , \29485 );
not \U$29144 ( \29487 , \9668 );
not \U$29145 ( \29488 , \29258 );
or \U$29146 ( \29489 , \29487 , \29488 );
not \U$29147 ( \29490 , RI9872bf8_170);
not \U$29148 ( \29491 , \8053 );
or \U$29149 ( \29492 , \29490 , \29491 );
or \U$29150 ( \29493 , \8053 , RI9872bf8_170);
nand \U$29151 ( \29494 , \29492 , \29493 );
nand \U$29152 ( \29495 , \29494 , \9249 );
nand \U$29153 ( \29496 , \29489 , \29495 );
not \U$29154 ( \29497 , \29496 );
or \U$29155 ( \29498 , \29486 , \29497 );
or \U$29156 ( \29499 , \29496 , \29485 );
not \U$29157 ( \29500 , \9214 );
not \U$29158 ( \29501 , \29285 );
or \U$29159 ( \29502 , \29500 , \29501 );
not \U$29160 ( \29503 , \11688 );
not \U$29161 ( \29504 , \17449 );
or \U$29162 ( \29505 , \29503 , \29504 );
nand \U$29163 ( \29506 , \8948 , RI9872b80_169);
nand \U$29164 ( \29507 , \29505 , \29506 );
nand \U$29165 ( \29508 , \29507 , \9196 );
nand \U$29166 ( \29509 , \29502 , \29508 );
nand \U$29167 ( \29510 , \29499 , \29509 );
nand \U$29168 ( \29511 , \29498 , \29510 );
not \U$29169 ( \29512 , \29511 );
or \U$29170 ( \29513 , \29476 , \29512 );
nand \U$29171 ( \29514 , \29376 , \29473 );
nand \U$29172 ( \29515 , \29513 , \29514 );
not \U$29173 ( \29516 , \29515 );
xor \U$29174 ( \29517 , \29160 , \29186 );
xnor \U$29175 ( \29518 , \29517 , \29158 );
not \U$29176 ( \29519 , \29518 );
or \U$29177 ( \29520 , \29516 , \29519 );
or \U$29178 ( \29521 , \29515 , \29518 );
nand \U$29179 ( \29522 , \29520 , \29521 );
not \U$29180 ( \29523 , \29522 );
or \U$29181 ( \29524 , \29343 , \29523 );
not \U$29182 ( \29525 , \29518 );
nand \U$29183 ( \29526 , \29525 , \29515 );
nand \U$29184 ( \29527 , \29524 , \29526 );
xor \U$29185 ( \29528 , \29095 , \29111 );
not \U$29186 ( \29529 , \29101 );
xnor \U$29187 ( \29530 , \29528 , \29529 );
or \U$29188 ( \29531 , \29527 , \29530 );
xor \U$29189 ( \29532 , \29191 , \29120 );
xor \U$29190 ( \29533 , \29532 , \29194 );
nand \U$29191 ( \29534 , \29531 , \29533 );
nand \U$29192 ( \29535 , \29527 , \29530 );
nand \U$29193 ( \29536 , \29534 , \29535 );
not \U$29194 ( \29537 , \29536 );
not \U$29195 ( \29538 , \29537 );
xor \U$29196 ( \29539 , \29116 , \29205 );
xor \U$29197 ( \29540 , \29539 , \29197 );
not \U$29198 ( \29541 , \29540 );
or \U$29199 ( \29542 , \29538 , \29541 );
or \U$29200 ( \29543 , \29540 , \29537 );
nand \U$29201 ( \29544 , \29542 , \29543 );
not \U$29202 ( \29545 , \29544 );
or \U$29203 ( \29546 , \29341 , \29545 );
nand \U$29204 ( \29547 , \29540 , \29536 );
nand \U$29205 ( \29548 , \29546 , \29547 );
xor \U$29206 ( \29549 , \29329 , \29548 );
xor \U$29207 ( \29550 , \29019 , \29020 );
xor \U$29208 ( \29551 , \29550 , \29056 );
not \U$29209 ( \29552 , \29551 );
not \U$29210 ( \29553 , \28809 );
and \U$29211 ( \29554 , \28858 , \29553 );
not \U$29212 ( \29555 , \28858 );
and \U$29213 ( \29556 , \29555 , \28809 );
nor \U$29214 ( \29557 , \29554 , \29556 );
not \U$29215 ( \29558 , RI9873648_192);
not \U$29216 ( \29559 , \29040 );
or \U$29217 ( \29560 , \29558 , \29559 );
not \U$29218 ( \29561 , \18668 );
xor \U$29219 ( \29562 , RI9873558_190, \29561 );
nand \U$29220 ( \29563 , \29562 , \20626 );
nand \U$29221 ( \29564 , \29560 , \29563 );
not \U$29222 ( \29565 , \29564 );
not \U$29223 ( \29566 , \6284 );
and \U$29224 ( \29567 , RI98728b0_163, \8597 );
not \U$29225 ( \29568 , RI98728b0_163);
not \U$29226 ( \29569 , \8606 );
and \U$29227 ( \29570 , \29568 , \29569 );
nor \U$29228 ( \29571 , \29567 , \29570 );
not \U$29229 ( \29572 , \29571 );
or \U$29230 ( \29573 , \29566 , \29572 );
nand \U$29231 ( \29574 , \28947 , \6286 );
nand \U$29232 ( \29575 , \29573 , \29574 );
not \U$29233 ( \29576 , \29399 );
not \U$29234 ( \29577 , \29386 );
or \U$29235 ( \29578 , \29576 , \29577 );
nand \U$29236 ( \29579 , \29388 , \29398 );
nand \U$29237 ( \29580 , \29578 , \29579 );
and \U$29238 ( \29581 , \29575 , \29580 );
not \U$29239 ( \29582 , \29575 );
not \U$29240 ( \29583 , \29580 );
and \U$29241 ( \29584 , \29582 , \29583 );
nor \U$29242 ( \29585 , \29581 , \29584 );
not \U$29243 ( \29586 , \29585 );
or \U$29244 ( \29587 , \29565 , \29586 );
nand \U$29245 ( \29588 , \29575 , \29580 );
nand \U$29246 ( \29589 , \29587 , \29588 );
not \U$29247 ( \29590 , \29589 );
nand \U$29248 ( \29591 , \29557 , \29590 );
not \U$29249 ( \29592 , \29591 );
xor \U$29250 ( \29593 , \28872 , \28892 );
xor \U$29251 ( \29594 , \29593 , \28900 );
not \U$29252 ( \29595 , \29594 );
or \U$29253 ( \29596 , \29592 , \29595 );
not \U$29254 ( \29597 , \29557 );
nand \U$29255 ( \29598 , \29597 , \29589 );
nand \U$29256 ( \29599 , \29596 , \29598 );
not \U$29257 ( \29600 , \29599 );
not \U$29258 ( \29601 , \29600 );
xor \U$29259 ( \29602 , \28799 , \28862 );
xor \U$29260 ( \29603 , \29602 , \28902 );
not \U$29261 ( \29604 , \29603 );
or \U$29262 ( \29605 , \29601 , \29604 );
or \U$29263 ( \29606 , \29603 , \29600 );
nand \U$29264 ( \29607 , \29605 , \29606 );
not \U$29265 ( \29608 , \29607 );
or \U$29266 ( \29609 , \29552 , \29608 );
not \U$29267 ( \29610 , \29600 );
nand \U$29268 ( \29611 , \29610 , \29603 );
nand \U$29269 ( \29612 , \29609 , \29611 );
not \U$29270 ( \29613 , \29612 );
xor \U$29271 ( \29614 , \28922 , \28954 );
not \U$29272 ( \29615 , \29614 );
not \U$29273 ( \29616 , \17371 );
not \U$29274 ( \29617 , RI98733f0_187);
not \U$29275 ( \29618 , \17140 );
or \U$29276 ( \29619 , \29617 , \29618 );
or \U$29277 ( \29620 , \17143 , RI98733f0_187);
nand \U$29278 ( \29621 , \29619 , \29620 );
not \U$29279 ( \29622 , \29621 );
or \U$29280 ( \29623 , \29616 , \29622 );
nand \U$29281 ( \29624 , \29049 , \17263 );
nand \U$29282 ( \29625 , \29623 , \29624 );
not \U$29283 ( \29626 , \29625 );
xor \U$29284 ( \29627 , \28831 , \28853 );
not \U$29285 ( \29628 , \17347 );
not \U$29286 ( \29629 , \28770 );
or \U$29287 ( \29630 , \29628 , \29629 );
xor \U$29288 ( \29631 , RI98730a8_180, \3239 );
not \U$29289 ( \29632 , \24209 );
not \U$29290 ( \29633 , \29632 );
nand \U$29291 ( \29634 , \29631 , \29633 );
nand \U$29292 ( \29635 , \29630 , \29634 );
xor \U$29293 ( \29636 , \29627 , \29635 );
not \U$29294 ( \29637 , \29636 );
or \U$29295 ( \29638 , \29626 , \29637 );
nand \U$29296 ( \29639 , \29635 , \29627 );
nand \U$29297 ( \29640 , \29638 , \29639 );
not \U$29298 ( \29641 , \29640 );
not \U$29299 ( \29642 , \9294 );
not \U$29300 ( \29643 , RI9872e50_175);
not \U$29301 ( \29644 , \7007 );
or \U$29302 ( \29645 , \29643 , \29644 );
or \U$29303 ( \29646 , \4990 , RI9872e50_175);
nand \U$29304 ( \29647 , \29645 , \29646 );
not \U$29305 ( \29648 , \29647 );
or \U$29306 ( \29649 , \29642 , \29648 );
nand \U$29307 ( \29650 , \28890 , \10331 );
nand \U$29308 ( \29651 , \29649 , \29650 );
not \U$29309 ( \29652 , \29651 );
not \U$29310 ( \29653 , \29652 );
not \U$29311 ( \29654 , \13214 );
not \U$29312 ( \29655 , \28805 );
or \U$29313 ( \29656 , \29654 , \29655 );
not \U$29314 ( \29657 , \14080 );
not \U$29315 ( \29658 , \12832 );
not \U$29316 ( \29659 , \29658 );
or \U$29317 ( \29660 , \29657 , \29659 );
not \U$29318 ( \29661 , \8732 );
nand \U$29319 ( \29662 , \29661 , \5205 );
nand \U$29320 ( \29663 , \29660 , \29662 );
nand \U$29321 ( \29664 , \29663 , \9526 );
nand \U$29322 ( \29665 , \29656 , \29664 );
not \U$29323 ( \29666 , \29665 );
not \U$29324 ( \29667 , \29666 );
or \U$29325 ( \29668 , \29653 , \29667 );
not \U$29326 ( \29669 , \18508 );
not \U$29327 ( \29670 , RI9873288_184);
not \U$29328 ( \29671 , \5946 );
or \U$29329 ( \29672 , \29670 , \29671 );
or \U$29330 ( \29673 , \1190 , RI9873288_184);
nand \U$29331 ( \29674 , \29672 , \29673 );
not \U$29332 ( \29675 , \29674 );
or \U$29333 ( \29676 , \29669 , \29675 );
nand \U$29334 ( \29677 , \28881 , \17528 );
nand \U$29335 ( \29678 , \29676 , \29677 );
nand \U$29336 ( \29679 , \29668 , \29678 );
nand \U$29337 ( \29680 , \29665 , \29651 );
nand \U$29338 ( \29681 , \29679 , \29680 );
not \U$29339 ( \29682 , \29681 );
or \U$29340 ( \29683 , \29641 , \29682 );
or \U$29341 ( \29684 , \29681 , \29640 );
not \U$29342 ( \29685 , \8802 );
not \U$29343 ( \29686 , \28870 );
or \U$29344 ( \29687 , \29685 , \29686 );
and \U$29345 ( \29688 , \5775 , \8807 );
not \U$29346 ( \29689 , \5775 );
and \U$29347 ( \29690 , \29689 , RI9872d60_173);
nor \U$29348 ( \29691 , \29688 , \29690 );
nand \U$29349 ( \29692 , \29691 , \8819 );
nand \U$29350 ( \29693 , \29687 , \29692 );
not \U$29351 ( \29694 , \19243 );
not \U$29352 ( \29695 , \16999 );
not \U$29353 ( \29696 , \1365 );
or \U$29354 ( \29697 , \29695 , \29696 );
or \U$29355 ( \29698 , \1365 , \16999 );
nand \U$29356 ( \29699 , \29697 , \29698 );
not \U$29357 ( \29700 , \29699 );
or \U$29358 ( \29701 , \29694 , \29700 );
nand \U$29359 ( \29702 , \28818 , \19046 );
nand \U$29360 ( \29703 , \29701 , \29702 );
xor \U$29361 ( \29704 , \29693 , \29703 );
not \U$29362 ( \29705 , \13477 );
and \U$29363 ( \29706 , RI9873210_183, \2111 );
not \U$29364 ( \29707 , RI9873210_183);
and \U$29365 ( \29708 , \29707 , \9162 );
nor \U$29366 ( \29709 , \29706 , \29708 );
not \U$29367 ( \29710 , \29709 );
or \U$29368 ( \29711 , \29705 , \29710 );
nand \U$29369 ( \29712 , \28793 , \22670 );
nand \U$29370 ( \29713 , \29711 , \29712 );
and \U$29371 ( \29714 , \29704 , \29713 );
and \U$29372 ( \29715 , \29693 , \29703 );
or \U$29373 ( \29716 , \29714 , \29715 );
nand \U$29374 ( \29717 , \29684 , \29716 );
nand \U$29375 ( \29718 , \29683 , \29717 );
not \U$29376 ( \29719 , \29718 );
not \U$29377 ( \29720 , \29719 );
or \U$29378 ( \29721 , \29615 , \29720 );
or \U$29379 ( \29722 , \29719 , \29614 );
nand \U$29380 ( \29723 , \29721 , \29722 );
not \U$29381 ( \29724 , \29723 );
not \U$29382 ( \29725 , \28772 );
not \U$29383 ( \29726 , \28783 );
and \U$29384 ( \29727 , \29725 , \29726 );
and \U$29385 ( \29728 , \28772 , \28783 );
nor \U$29386 ( \29729 , \29727 , \29728 );
xnor \U$29387 ( \29730 , \28795 , \29729 );
not \U$29388 ( \29731 , \29730 );
and \U$29389 ( \29732 , \1134 , \28848 );
and \U$29390 ( \29733 , RI98718c0_129, \16996 );
not \U$29391 ( \29734 , RI98718c0_129);
and \U$29392 ( \29735 , \29734 , \16995 );
or \U$29393 ( \29736 , \29733 , \29735 );
and \U$29394 ( \29737 , \29736 , \1083 );
nor \U$29395 ( \29738 , \29732 , \29737 );
not \U$29396 ( \29739 , \29738 );
not \U$29397 ( \29740 , \1134 );
not \U$29398 ( \29741 , \29736 );
or \U$29399 ( \29742 , \29740 , \29741 );
not \U$29400 ( \29743 , \1111 );
not \U$29401 ( \29744 , \17703 );
or \U$29402 ( \29745 , \29743 , \29744 );
nand \U$29403 ( \29746 , \27541 , RI98718c0_129);
nand \U$29404 ( \29747 , \29745 , \29746 );
nand \U$29405 ( \29748 , \29747 , \1082 );
nand \U$29406 ( \29749 , \29742 , \29748 );
not \U$29407 ( \29750 , \29749 );
and \U$29408 ( \29751 , \18704 , \1290 );
not \U$29409 ( \29752 , \29751 );
not \U$29410 ( \29753 , \1427 );
not \U$29411 ( \29754 , \29396 );
or \U$29412 ( \29755 , \29753 , \29754 );
nand \U$29413 ( \29756 , \29429 , \1454 );
nand \U$29414 ( \29757 , \29755 , \29756 );
not \U$29415 ( \29758 , \29757 );
not \U$29416 ( \29759 , \29758 );
or \U$29417 ( \29760 , \29752 , \29759 );
not \U$29418 ( \29761 , \29751 );
nand \U$29419 ( \29762 , \29761 , \29757 );
nand \U$29420 ( \29763 , \29760 , \29762 );
not \U$29421 ( \29764 , \29763 );
or \U$29422 ( \29765 , \29750 , \29764 );
nand \U$29423 ( \29766 , \29757 , \29751 );
nand \U$29424 ( \29767 , \29765 , \29766 );
not \U$29425 ( \29768 , \29767 );
or \U$29426 ( \29769 , \29739 , \29768 );
or \U$29427 ( \29770 , \29767 , \29738 );
nand \U$29428 ( \29771 , \29769 , \29770 );
not \U$29429 ( \29772 , \29771 );
not \U$29430 ( \29773 , \4084 );
not \U$29431 ( \29774 , \29166 );
or \U$29432 ( \29775 , \29773 , \29774 );
and \U$29433 ( \29776 , RI98725e0_157, \13067 );
not \U$29434 ( \29777 , RI98725e0_157);
and \U$29435 ( \29778 , \29777 , \24501 );
nor \U$29436 ( \29779 , \29776 , \29778 );
nand \U$29437 ( \29780 , \29779 , \4101 );
nand \U$29438 ( \29781 , \29775 , \29780 );
not \U$29439 ( \29782 , \29781 );
or \U$29440 ( \29783 , \29772 , \29782 );
not \U$29441 ( \29784 , \29738 );
nand \U$29442 ( \29785 , \29784 , \29767 );
nand \U$29443 ( \29786 , \29783 , \29785 );
not \U$29444 ( \29787 , \2087 );
not \U$29445 ( \29788 , \29139 );
or \U$29446 ( \29789 , \29787 , \29788 );
not \U$29447 ( \29790 , \29408 );
nand \U$29448 ( \29791 , \29790 , \2071 );
nand \U$29449 ( \29792 , \29789 , \29791 );
not \U$29450 ( \29793 , \3169 );
not \U$29451 ( \29794 , \29126 );
or \U$29452 ( \29795 , \29793 , \29794 );
not \U$29453 ( \29796 , RI9872310_151);
not \U$29454 ( \29797 , \20928 );
or \U$29455 ( \29798 , \29796 , \29797 );
or \U$29456 ( \29799 , \17090 , RI9872310_151);
nand \U$29457 ( \29800 , \29798 , \29799 );
nand \U$29458 ( \29801 , \29800 , \3163 );
nand \U$29459 ( \29802 , \29795 , \29801 );
xor \U$29460 ( \29803 , \29792 , \29802 );
not \U$29461 ( \29804 , \3467 );
not \U$29462 ( \29805 , \29176 );
or \U$29463 ( \29806 , \29804 , \29805 );
not \U$29464 ( \29807 , RI98726d0_159);
not \U$29465 ( \29808 , \11454 );
not \U$29466 ( \29809 , \29808 );
or \U$29467 ( \29810 , \29807 , \29809 );
or \U$29468 ( \29811 , \12784 , RI98726d0_159);
nand \U$29469 ( \29812 , \29810 , \29811 );
nand \U$29470 ( \29813 , \29812 , \3465 );
nand \U$29471 ( \29814 , \29806 , \29813 );
and \U$29472 ( \29815 , \29803 , \29814 );
and \U$29473 ( \29816 , \29792 , \29802 );
or \U$29474 ( \29817 , \29815 , \29816 );
xor \U$29475 ( \29818 , \29786 , \29817 );
not \U$29476 ( \29819 , \19321 );
not \U$29477 ( \29820 , RI9873030_179);
not \U$29478 ( \29821 , \11672 );
or \U$29479 ( \29822 , \29820 , \29821 );
or \U$29480 ( \29823 , \3568 , RI9873030_179);
nand \U$29481 ( \29824 , \29822 , \29823 );
not \U$29482 ( \29825 , \29824 );
or \U$29483 ( \29826 , \29819 , \29825 );
nand \U$29484 ( \29827 , \29029 , \9937 );
nand \U$29485 ( \29828 , \29826 , \29827 );
and \U$29486 ( \29829 , \29818 , \29828 );
and \U$29487 ( \29830 , \29786 , \29817 );
or \U$29488 ( \29831 , \29829 , \29830 );
not \U$29489 ( \29832 , \29831 );
xor \U$29490 ( \29833 , \29031 , \29832 );
xnor \U$29491 ( \29834 , \29833 , \29052 );
not \U$29492 ( \29835 , \29834 );
or \U$29493 ( \29836 , \29731 , \29835 );
not \U$29494 ( \29837 , \29052 );
not \U$29495 ( \29838 , \29031 );
not \U$29496 ( \29839 , \29838 );
and \U$29497 ( \29840 , \29837 , \29839 );
and \U$29498 ( \29841 , \29052 , \29838 );
nor \U$29499 ( \29842 , \29840 , \29841 );
or \U$29500 ( \29843 , \29832 , \29842 );
nand \U$29501 ( \29844 , \29836 , \29843 );
not \U$29502 ( \29845 , \29844 );
or \U$29503 ( \29846 , \29724 , \29845 );
nand \U$29504 ( \29847 , \29718 , \29614 );
nand \U$29505 ( \29848 , \29846 , \29847 );
xor \U$29506 ( \29849 , \28626 , \28762 );
xor \U$29507 ( \29850 , \29849 , \28905 );
nor \U$29508 ( \29851 , \29848 , \29850 );
or \U$29509 ( \29852 , \29613 , \29851 );
nand \U$29510 ( \29853 , \29848 , \29850 );
nand \U$29511 ( \29854 , \29852 , \29853 );
not \U$29512 ( \29855 , \29854 );
xor \U$29513 ( \29856 , \28621 , \28623 );
xor \U$29514 ( \29857 , \29856 , \28909 );
not \U$29515 ( \29858 , \29857 );
and \U$29516 ( \29859 , \29855 , \29858 );
and \U$29517 ( \29860 , \29854 , \29857 );
nor \U$29518 ( \29861 , \29859 , \29860 );
not \U$29519 ( \29862 , \29002 );
not \U$29520 ( \29863 , \29070 );
not \U$29521 ( \29864 , \29863 );
or \U$29522 ( \29865 , \29862 , \29864 );
not \U$29523 ( \29866 , \29002 );
nand \U$29524 ( \29867 , \29866 , \29070 );
nand \U$29525 ( \29868 , \29865 , \29867 );
xnor \U$29526 ( \29869 , \29861 , \29868 );
and \U$29527 ( \29870 , \29549 , \29869 );
and \U$29528 ( \29871 , \29329 , \29548 );
or \U$29529 ( \29872 , \29870 , \29871 );
not \U$29530 ( \29873 , \29872 );
xor \U$29531 ( \29874 , \29093 , \29873 );
xor \U$29532 ( \29875 , \29214 , \29325 );
and \U$29533 ( \29876 , \29875 , \29328 );
and \U$29534 ( \29877 , \29214 , \29325 );
or \U$29535 ( \29878 , \29876 , \29877 );
xor \U$29536 ( \29879 , \28986 , \28912 );
xnor \U$29537 ( \29880 , \29879 , \28991 );
xor \U$29538 ( \29881 , \29878 , \29880 );
not \U$29539 ( \29882 , \29861 );
not \U$29540 ( \29883 , \29882 );
not \U$29541 ( \29884 , \29868 );
or \U$29542 ( \29885 , \29883 , \29884 );
not \U$29543 ( \29886 , \29857 );
nand \U$29544 ( \29887 , \29886 , \29854 );
nand \U$29545 ( \29888 , \29885 , \29887 );
not \U$29546 ( \29889 , \29888 );
xor \U$29547 ( \29890 , \29881 , \29889 );
xnor \U$29548 ( \29891 , \29874 , \29890 );
xor \U$29549 ( \29892 , \29329 , \29548 );
xor \U$29550 ( \29893 , \29892 , \29869 );
not \U$29551 ( \29894 , \29893 );
not \U$29552 ( \29895 , \29894 );
xor \U$29553 ( \29896 , \29536 , \29340 );
xor \U$29554 ( \29897 , \29896 , \29540 );
not \U$29555 ( \29898 , \29897 );
xor \U$29556 ( \29899 , \29832 , \29730 );
xnor \U$29557 ( \29900 , \29899 , \29842 );
xor \U$29558 ( \29901 , \29590 , \29557 );
xnor \U$29559 ( \29902 , \29901 , \29594 );
nand \U$29560 ( \29903 , \29900 , \29902 );
not \U$29561 ( \29904 , \29511 );
not \U$29562 ( \29905 , \29474 );
not \U$29563 ( \29906 , \29376 );
and \U$29564 ( \29907 , \29905 , \29906 );
and \U$29565 ( \29908 , \29376 , \29474 );
nor \U$29566 ( \29909 , \29907 , \29908 );
not \U$29567 ( \29910 , \29909 );
or \U$29568 ( \29911 , \29904 , \29910 );
or \U$29569 ( \29912 , \29909 , \29511 );
nand \U$29570 ( \29913 , \29911 , \29912 );
buf \U$29571 ( \29914 , \29913 );
not \U$29572 ( \29915 , \24627 );
and \U$29573 ( \29916 , \23391 , \14080 );
not \U$29574 ( \29917 , \23391 );
and \U$29575 ( \29918 , \29917 , RI9872f40_177);
nor \U$29576 ( \29919 , \29916 , \29918 );
not \U$29577 ( \29920 , \29919 );
or \U$29578 ( \29921 , \29915 , \29920 );
not \U$29579 ( \29922 , RI9872f40_177);
not \U$29580 ( \29923 , \4470 );
or \U$29581 ( \29924 , \29922 , \29923 );
or \U$29582 ( \29925 , \4470 , RI9872f40_177);
nand \U$29583 ( \29926 , \29924 , \29925 );
nand \U$29584 ( \29927 , \29926 , \8752 );
nand \U$29585 ( \29928 , \29921 , \29927 );
not \U$29586 ( \29929 , \29928 );
not \U$29587 ( \29930 , \796 );
not \U$29588 ( \29931 , \29445 );
or \U$29589 ( \29932 , \29930 , \29931 );
not \U$29590 ( \29933 , RI98719b0_131);
not \U$29591 ( \29934 , \16996 );
or \U$29592 ( \29935 , \29933 , \29934 );
or \U$29593 ( \29936 , \21553 , RI98719b0_131);
nand \U$29594 ( \29937 , \29935 , \29936 );
nand \U$29595 ( \29938 , \29937 , \791 );
nand \U$29596 ( \29939 , \29932 , \29938 );
not \U$29597 ( \29940 , \29939 );
not \U$29598 ( \29941 , \1134 );
not \U$29599 ( \29942 , \29747 );
or \U$29600 ( \29943 , \29941 , \29942 );
xor \U$29601 ( \29944 , RI98718c0_129, \17862 );
nand \U$29602 ( \29945 , \29944 , \1082 );
nand \U$29603 ( \29946 , \29943 , \29945 );
not \U$29604 ( \29947 , \29946 );
not \U$29605 ( \29948 , \29438 );
not \U$29606 ( \29949 , \29422 );
and \U$29607 ( \29950 , \29948 , \29949 );
and \U$29608 ( \29951 , \29438 , \29422 );
nor \U$29609 ( \29952 , \29950 , \29951 );
not \U$29610 ( \29953 , \29952 );
or \U$29611 ( \29954 , \29947 , \29953 );
or \U$29612 ( \29955 , \29946 , \29952 );
nand \U$29613 ( \29956 , \29954 , \29955 );
not \U$29614 ( \29957 , \29956 );
or \U$29615 ( \29958 , \29940 , \29957 );
not \U$29616 ( \29959 , \29952 );
nand \U$29617 ( \29960 , \29959 , \29946 );
nand \U$29618 ( \29961 , \29958 , \29960 );
not \U$29619 ( \29962 , \29961 );
not \U$29620 ( \29963 , \29962 );
not \U$29621 ( \29964 , \6284 );
not \U$29622 ( \29965 , RI98728b0_163);
not \U$29623 ( \29966 , \8650 );
or \U$29624 ( \29967 , \29965 , \29966 );
or \U$29625 ( \29968 , \11406 , RI98728b0_163);
nand \U$29626 ( \29969 , \29967 , \29968 );
not \U$29627 ( \29970 , \29969 );
or \U$29628 ( \29971 , \29964 , \29970 );
not \U$29629 ( \29972 , RI98728b0_163);
not \U$29630 ( \29973 , \8667 );
or \U$29631 ( \29974 , \29972 , \29973 );
or \U$29632 ( \29975 , \20414 , RI98728b0_163);
nand \U$29633 ( \29976 , \29974 , \29975 );
nand \U$29634 ( \29977 , \29976 , \6286 );
nand \U$29635 ( \29978 , \29971 , \29977 );
not \U$29636 ( \29979 , \29978 );
or \U$29637 ( \29980 , \29963 , \29979 );
or \U$29638 ( \29981 , \29978 , \29962 );
nand \U$29639 ( \29982 , \29980 , \29981 );
not \U$29640 ( \29983 , \29982 );
or \U$29641 ( \29984 , \29929 , \29983 );
not \U$29642 ( \29985 , \29962 );
nand \U$29643 ( \29986 , \29985 , \29978 );
nand \U$29644 ( \29987 , \29984 , \29986 );
not \U$29645 ( \29988 , \29987 );
xor \U$29646 ( \29989 , \29792 , \29802 );
xor \U$29647 ( \29990 , \29989 , \29814 );
not \U$29648 ( \29991 , \3464 );
not \U$29649 ( \29992 , RI98726d0_159);
not \U$29650 ( \29993 , \13268 );
or \U$29651 ( \29994 , \29992 , \29993 );
or \U$29652 ( \29995 , \12773 , RI98726d0_159);
nand \U$29653 ( \29996 , \29994 , \29995 );
not \U$29654 ( \29997 , \29996 );
or \U$29655 ( \29998 , \29991 , \29997 );
nand \U$29656 ( \29999 , \29812 , \3467 );
nand \U$29657 ( \30000 , \29998 , \29999 );
not \U$29658 ( \30001 , \30000 );
not \U$29659 ( \30002 , \4101 );
and \U$29660 ( \30003 , \10064 , \6042 );
not \U$29661 ( \30004 , \10064 );
and \U$29662 ( \30005 , \30004 , RI98725e0_157);
nor \U$29663 ( \30006 , \30003 , \30005 );
not \U$29664 ( \30007 , \30006 );
or \U$29665 ( \30008 , \30002 , \30007 );
nand \U$29666 ( \30009 , \29779 , \4084 );
nand \U$29667 ( \30010 , \30008 , \30009 );
not \U$29668 ( \30011 , \30010 );
nand \U$29669 ( \30012 , \30001 , \30011 );
not \U$29670 ( \30013 , \30012 );
not \U$29671 ( \30014 , \9312 );
and \U$29672 ( \30015 , RI9872d60_173, \5703 );
not \U$29673 ( \30016 , RI9872d60_173);
and \U$29674 ( \30017 , \30016 , \7111 );
nor \U$29675 ( \30018 , \30015 , \30017 );
not \U$29676 ( \30019 , \30018 );
or \U$29677 ( \30020 , \30014 , \30019 );
and \U$29678 ( \30021 , \5761 , \8807 );
not \U$29679 ( \30022 , \5761 );
and \U$29680 ( \30023 , \30022 , RI9872d60_173);
nor \U$29681 ( \30024 , \30021 , \30023 );
nand \U$29682 ( \30025 , \30024 , \10624 );
nand \U$29683 ( \30026 , \30020 , \30025 );
not \U$29684 ( \30027 , \30026 );
or \U$29685 ( \30028 , \30013 , \30027 );
nand \U$29686 ( \30029 , \30010 , \30000 );
nand \U$29687 ( \30030 , \30028 , \30029 );
and \U$29688 ( \30031 , \29990 , \30030 );
not \U$29689 ( \30032 , \29990 );
not \U$29690 ( \30033 , \30030 );
and \U$29691 ( \30034 , \30032 , \30033 );
nor \U$29692 ( \30035 , \30031 , \30034 );
not \U$29693 ( \30036 , \30035 );
or \U$29694 ( \30037 , \29988 , \30036 );
not \U$29695 ( \30038 , \30033 );
nand \U$29696 ( \30039 , \30038 , \29990 );
nand \U$29697 ( \30040 , \30037 , \30039 );
nor \U$29698 ( \30041 , \29914 , \30040 );
and \U$29699 ( \30042 , \29663 , \13214 );
not \U$29700 ( \30043 , \29926 );
nor \U$29701 ( \30044 , \30043 , \18284 );
nor \U$29702 ( \30045 , \30042 , \30044 );
not \U$29703 ( \30046 , \30045 );
not \U$29704 ( \30047 , \30046 );
not \U$29705 ( \30048 , \6285 );
not \U$29706 ( \30049 , \29571 );
or \U$29707 ( \30050 , \30048 , \30049 );
nand \U$29708 ( \30051 , \29976 , \6284 );
nand \U$29709 ( \30052 , \30050 , \30051 );
not \U$29710 ( \30053 , \30052 );
not \U$29711 ( \30054 , \18615 );
and \U$29712 ( \30055 , RI9873558_190, \20612 );
not \U$29713 ( \30056 , RI9873558_190);
and \U$29714 ( \30057 , \30056 , \22615 );
or \U$29715 ( \30058 , \30055 , \30057 );
not \U$29716 ( \30059 , \30058 );
or \U$29717 ( \30060 , \30054 , \30059 );
nand \U$29718 ( \30061 , \29562 , RI9873648_192);
nand \U$29719 ( \30062 , \30060 , \30061 );
not \U$29720 ( \30063 , \30062 );
not \U$29721 ( \30064 , \30063 );
or \U$29722 ( \30065 , \30053 , \30064 );
or \U$29723 ( \30066 , \30063 , \30052 );
nand \U$29724 ( \30067 , \30065 , \30066 );
not \U$29725 ( \30068 , \30067 );
or \U$29726 ( \30069 , \30047 , \30068 );
nand \U$29727 ( \30070 , \30062 , \30052 );
nand \U$29728 ( \30071 , \30069 , \30070 );
not \U$29729 ( \30072 , \29157 );
nor \U$29730 ( \30073 , \30072 , \29142 );
xor \U$29731 ( \30074 , \30073 , \29154 );
not \U$29732 ( \30075 , \30074 );
xnor \U$29733 ( \30076 , \29182 , \29170 );
not \U$29734 ( \30077 , \30076 );
and \U$29735 ( \30078 , \30075 , \30077 );
and \U$29736 ( \30079 , \30074 , \30076 );
nor \U$29737 ( \30080 , \30078 , \30079 );
xor \U$29738 ( \30081 , \30071 , \30080 );
or \U$29739 ( \30082 , \30041 , \30081 );
nand \U$29740 ( \30083 , \30040 , \29914 );
nand \U$29741 ( \30084 , \30082 , \30083 );
nand \U$29742 ( \30085 , \29903 , \30084 );
not \U$29743 ( \30086 , \29900 );
not \U$29744 ( \30087 , \29902 );
nand \U$29745 ( \30088 , \30086 , \30087 );
and \U$29746 ( \30089 , \30085 , \30088 );
not \U$29747 ( \30090 , \30089 );
not \U$29748 ( \30091 , \30090 );
and \U$29749 ( \30092 , \29844 , \29723 );
not \U$29750 ( \30093 , \29844 );
not \U$29751 ( \30094 , \29723 );
and \U$29752 ( \30095 , \30093 , \30094 );
nor \U$29753 ( \30096 , \30092 , \30095 );
not \U$29754 ( \30097 , \30096 );
not \U$29755 ( \30098 , \30097 );
not \U$29756 ( \30099 , \29551 );
not \U$29757 ( \30100 , \29607 );
not \U$29758 ( \30101 , \30100 );
or \U$29759 ( \30102 , \30099 , \30101 );
not \U$29760 ( \30103 , \29551 );
nand \U$29761 ( \30104 , \30103 , \29607 );
nand \U$29762 ( \30105 , \30102 , \30104 );
not \U$29763 ( \30106 , \30105 );
or \U$29764 ( \30107 , \30098 , \30106 );
or \U$29765 ( \30108 , \30105 , \30097 );
nand \U$29766 ( \30109 , \30107 , \30108 );
not \U$29767 ( \30110 , \30109 );
or \U$29768 ( \30111 , \30091 , \30110 );
not \U$29769 ( \30112 , \30097 );
nand \U$29770 ( \30113 , \30112 , \30105 );
nand \U$29771 ( \30114 , \30111 , \30113 );
not \U$29772 ( \30115 , \30114 );
nand \U$29773 ( \30116 , \29898 , \30115 );
xor \U$29774 ( \30117 , \29530 , \29527 );
xor \U$29775 ( \30118 , \30117 , \29533 );
xor \U$29776 ( \30119 , \30052 , \30063 );
xnor \U$29777 ( \30120 , \30119 , \30045 );
not \U$29778 ( \30121 , \30120 );
not \U$29779 ( \30122 , \8801 );
not \U$29780 ( \30123 , \29691 );
or \U$29781 ( \30124 , \30122 , \30123 );
nand \U$29782 ( \30125 , \30024 , \8819 );
nand \U$29783 ( \30126 , \30124 , \30125 );
not \U$29784 ( \30127 , \10332 );
not \U$29785 ( \30128 , \29647 );
or \U$29786 ( \30129 , \30127 , \30128 );
and \U$29787 ( \30130 , RI9872e50_175, \24185 );
not \U$29788 ( \30131 , RI9872e50_175);
and \U$29789 ( \30132 , \30131 , \22314 );
nor \U$29790 ( \30133 , \30130 , \30132 );
nand \U$29791 ( \30134 , \30133 , \9686 );
nand \U$29792 ( \30135 , \30129 , \30134 );
not \U$29793 ( \30136 , \30135 );
xor \U$29794 ( \30137 , \30126 , \30136 );
not \U$29795 ( \30138 , \17528 );
not \U$29796 ( \30139 , \29674 );
or \U$29797 ( \30140 , \30138 , \30139 );
not \U$29798 ( \30141 , \22715 );
not \U$29799 ( \30142 , \18004 );
not \U$29800 ( \30143 , \30142 );
or \U$29801 ( \30144 , \30141 , \30143 );
or \U$29802 ( \30145 , \30142 , \27966 );
nand \U$29803 ( \30146 , \30144 , \30145 );
nand \U$29804 ( \30147 , \30146 , \18508 );
nand \U$29805 ( \30148 , \30140 , \30147 );
xnor \U$29806 ( \30149 , \30137 , \30148 );
not \U$29807 ( \30150 , \30149 );
not \U$29808 ( \30151 , \30150 );
or \U$29809 ( \30152 , \30121 , \30151 );
not \U$29810 ( \30153 , \13477 );
not \U$29811 ( \30154 , RI9873210_183);
not \U$29812 ( \30155 , \2947 );
or \U$29813 ( \30156 , \30154 , \30155 );
or \U$29814 ( \30157 , \2947 , RI9873210_183);
nand \U$29815 ( \30158 , \30156 , \30157 );
not \U$29816 ( \30159 , \30158 );
or \U$29817 ( \30160 , \30153 , \30159 );
nand \U$29818 ( \30161 , \29709 , \17234 );
nand \U$29819 ( \30162 , \30160 , \30161 );
not \U$29820 ( \30163 , \20147 );
not \U$29821 ( \30164 , \29699 );
or \U$29822 ( \30165 , \30163 , \30164 );
and \U$29823 ( \30166 , RI98734e0_189, \1061 );
not \U$29824 ( \30167 , RI98734e0_189);
and \U$29825 ( \30168 , \30167 , \6572 );
nor \U$29826 ( \30169 , \30166 , \30168 );
nand \U$29827 ( \30170 , \30169 , \24076 );
nand \U$29828 ( \30171 , \30165 , \30170 );
not \U$29829 ( \30172 , \30171 );
not \U$29830 ( \30173 , \12867 );
not \U$29831 ( \30174 , \29631 );
or \U$29832 ( \30175 , \30173 , \30174 );
xor \U$29833 ( \30176 , RI98730a8_180, \3536 );
nand \U$29834 ( \30177 , \30176 , \13020 );
nand \U$29835 ( \30178 , \30175 , \30177 );
not \U$29836 ( \30179 , \30178 );
not \U$29837 ( \30180 , \30179 );
or \U$29838 ( \30181 , \30172 , \30180 );
or \U$29839 ( \30182 , \30179 , \30171 );
nand \U$29840 ( \30183 , \30181 , \30182 );
xor \U$29841 ( \30184 , \30162 , \30183 );
nand \U$29842 ( \30185 , \30152 , \30184 );
not \U$29843 ( \30186 , \30120 );
nand \U$29844 ( \30187 , \30186 , \30149 );
nand \U$29845 ( \30188 , \30185 , \30187 );
not \U$29846 ( \30189 , \30188 );
not \U$29847 ( \30190 , \9272 );
not \U$29848 ( \30191 , \30133 );
or \U$29849 ( \30192 , \30190 , \30191 );
xor \U$29850 ( \30193 , RI9872e50_175, \5392 );
nand \U$29851 ( \30194 , \30193 , \18562 );
nand \U$29852 ( \30195 , \30192 , \30194 );
not \U$29853 ( \30196 , \24209 );
not \U$29854 ( \30197 , RI98730a8_180);
not \U$29855 ( \30198 , \3567 );
or \U$29856 ( \30199 , \30197 , \30198 );
or \U$29857 ( \30200 , \3567 , RI98730a8_180);
nand \U$29858 ( \30201 , \30199 , \30200 );
not \U$29859 ( \30202 , \30201 );
or \U$29860 ( \30203 , \30196 , \30202 );
nand \U$29861 ( \30204 , \30176 , \22618 );
nand \U$29862 ( \30205 , \30203 , \30204 );
xor \U$29863 ( \30206 , \30195 , \30205 );
not \U$29864 ( \30207 , \18508 );
xor \U$29865 ( \30208 , RI9873288_184, \18453 );
not \U$29866 ( \30209 , \30208 );
or \U$29867 ( \30210 , \30207 , \30209 );
nand \U$29868 ( \30211 , \30146 , \17528 );
nand \U$29869 ( \30212 , \30210 , \30211 );
and \U$29870 ( \30213 , \30206 , \30212 );
and \U$29871 ( \30214 , \30195 , \30205 );
or \U$29872 ( \30215 , \30213 , \30214 );
xor \U$29873 ( \30216 , \29353 , \29362 );
xor \U$29874 ( \30217 , \30216 , \29373 );
xor \U$29875 ( \30218 , \30215 , \30217 );
xor \U$29876 ( \30219 , \29485 , \29496 );
xor \U$29877 ( \30220 , \30219 , \29509 );
and \U$29878 ( \30221 , \30218 , \30220 );
and \U$29879 ( \30222 , \30215 , \30217 );
or \U$29880 ( \30223 , \30221 , \30222 );
not \U$29881 ( \30224 , \30223 );
not \U$29882 ( \30225 , \29252 );
and \U$29883 ( \30226 , \29262 , \30225 );
not \U$29884 ( \30227 , \29262 );
and \U$29885 ( \30228 , \30227 , \29252 );
nor \U$29886 ( \30229 , \30226 , \30228 );
xor \U$29887 ( \30230 , \29301 , \30229 );
xor \U$29888 ( \30231 , \30230 , \29290 );
xor \U$29889 ( \30232 , \29781 , \29771 );
not \U$29890 ( \30233 , \30232 );
not \U$29891 ( \30234 , \19282 );
not \U$29892 ( \30235 , \29621 );
or \U$29893 ( \30236 , \30234 , \30235 );
and \U$29894 ( \30237 , RI98733f0_187, \20637 );
not \U$29895 ( \30238 , RI98733f0_187);
and \U$29896 ( \30239 , \30238 , \1209 );
nor \U$29897 ( \30240 , \30237 , \30239 );
nand \U$29898 ( \30241 , \30240 , \17371 );
nand \U$29899 ( \30242 , \30236 , \30241 );
not \U$29900 ( \30243 , \30242 );
or \U$29901 ( \30244 , \30233 , \30243 );
or \U$29902 ( \30245 , \30242 , \30232 );
not \U$29903 ( \30246 , \13109 );
and \U$29904 ( \30247 , RI9873030_179, \4176 );
not \U$29905 ( \30248 , RI9873030_179);
and \U$29906 ( \30249 , \30248 , \5594 );
or \U$29907 ( \30250 , \30247 , \30249 );
not \U$29908 ( \30251 , \30250 );
or \U$29909 ( \30252 , \30246 , \30251 );
nand \U$29910 ( \30253 , \29824 , \9937 );
nand \U$29911 ( \30254 , \30252 , \30253 );
nand \U$29912 ( \30255 , \30245 , \30254 );
nand \U$29913 ( \30256 , \30244 , \30255 );
and \U$29914 ( \30257 , \30231 , \30256 );
not \U$29915 ( \30258 , \30231 );
not \U$29916 ( \30259 , \30256 );
and \U$29917 ( \30260 , \30258 , \30259 );
nor \U$29918 ( \30261 , \30257 , \30260 );
nand \U$29919 ( \30262 , \30224 , \30261 );
not \U$29920 ( \30263 , \30262 );
or \U$29921 ( \30264 , \30189 , \30263 );
not \U$29922 ( \30265 , \30261 );
nand \U$29923 ( \30266 , \30265 , \30223 );
nand \U$29924 ( \30267 , \30264 , \30266 );
not \U$29925 ( \30268 , \30126 );
nand \U$29926 ( \30269 , \30268 , \30136 );
nand \U$29927 ( \30270 , \30148 , \30269 );
nand \U$29928 ( \30271 , \30135 , \30126 );
nand \U$29929 ( \30272 , \30270 , \30271 );
xor \U$29930 ( \30273 , \29564 , \29585 );
xor \U$29931 ( \30274 , \30272 , \30273 );
not \U$29932 ( \30275 , \30162 );
not \U$29933 ( \30276 , \30183 );
or \U$29934 ( \30277 , \30275 , \30276 );
nand \U$29935 ( \30278 , \30178 , \30171 );
nand \U$29936 ( \30279 , \30277 , \30278 );
and \U$29937 ( \30280 , \30274 , \30279 );
not \U$29938 ( \30281 , \30274 );
not \U$29939 ( \30282 , \30279 );
and \U$29940 ( \30283 , \30281 , \30282 );
nor \U$29941 ( \30284 , \30280 , \30283 );
not \U$29942 ( \30285 , \30284 );
not \U$29943 ( \30286 , \7338 );
not \U$29944 ( \30287 , RI98729a0_165);
not \U$29945 ( \30288 , \18110 );
or \U$29946 ( \30289 , \30287 , \30288 );
or \U$29947 ( \30290 , \8607 , RI98729a0_165);
nand \U$29948 ( \30291 , \30289 , \30290 );
not \U$29949 ( \30292 , \30291 );
or \U$29950 ( \30293 , \30286 , \30292 );
and \U$29951 ( \30294 , \9882 , \7333 );
not \U$29952 ( \30295 , \9882 );
and \U$29953 ( \30296 , \30295 , RI98729a0_165);
nor \U$29954 ( \30297 , \30294 , \30296 );
nand \U$29955 ( \30298 , \30297 , \7325 );
nand \U$29956 ( \30299 , \30293 , \30298 );
not \U$29957 ( \30300 , \30299 );
not \U$29958 ( \30301 , \9072 );
and \U$29959 ( \30302 , RI9872a18_166, \9598 );
not \U$29960 ( \30303 , RI9872a18_166);
and \U$29961 ( \30304 , \30303 , \9599 );
nor \U$29962 ( \30305 , \30302 , \30304 );
not \U$29963 ( \30306 , \30305 );
or \U$29964 ( \30307 , \30301 , \30306 );
not \U$29965 ( \30308 , RI9872a18_166);
not \U$29966 ( \30309 , \16942 );
or \U$29967 ( \30310 , \30308 , \30309 );
or \U$29968 ( \30311 , \8620 , RI9872a18_166);
nand \U$29969 ( \30312 , \30310 , \30311 );
nand \U$29970 ( \30313 , \30312 , \8028 );
nand \U$29971 ( \30314 , \30307 , \30313 );
not \U$29972 ( \30315 , \30314 );
not \U$29973 ( \30316 , \3163 );
not \U$29974 ( \30317 , RI9872310_151);
not \U$29975 ( \30318 , \13934 );
or \U$29976 ( \30319 , \30317 , \30318 );
not \U$29977 ( \30320 , \17005 );
or \U$29978 ( \30321 , \30320 , RI9872310_151);
nand \U$29979 ( \30322 , \30319 , \30321 );
not \U$29980 ( \30323 , \30322 );
or \U$29981 ( \30324 , \30316 , \30323 );
and \U$29982 ( \30325 , RI9872310_151, \25224 );
not \U$29983 ( \30326 , RI9872310_151);
and \U$29984 ( \30327 , \30326 , \17883 );
or \U$29985 ( \30328 , \30325 , \30327 );
nand \U$29986 ( \30329 , \30328 , \3169 );
nand \U$29987 ( \30330 , \30324 , \30329 );
not \U$29988 ( \30331 , \30330 );
and \U$29989 ( \30332 , RI98718c0_129, \23949 );
not \U$29990 ( \30333 , RI98718c0_129);
and \U$29991 ( \30334 , \30333 , \23952 );
or \U$29992 ( \30335 , \30332 , \30334 );
not \U$29993 ( \30336 , \30335 );
or \U$29994 ( \30337 , \30336 , \6671 );
and \U$29995 ( \30338 , RI98718c0_129, \24449 );
not \U$29996 ( \30339 , RI98718c0_129);
and \U$29997 ( \30340 , \30339 , \18704 );
nor \U$29998 ( \30341 , \30338 , \30340 );
not \U$29999 ( \30342 , \1082 );
or \U$30000 ( \30343 , \30341 , \30342 );
nand \U$30001 ( \30344 , \30337 , \30343 );
nand \U$30002 ( \30345 , \24450 , \1079 );
nand \U$30003 ( \30346 , \30345 , \1080 , RI98718c0_129);
not \U$30004 ( \30347 , \30346 );
and \U$30005 ( \30348 , \30344 , \30347 );
not \U$30006 ( \30349 , \2071 );
not \U$30007 ( \30350 , \17869 );
and \U$30008 ( \30351 , RI9871aa0_133, \30350 );
not \U$30009 ( \30352 , RI9871aa0_133);
and \U$30010 ( \30353 , \30352 , \25409 );
or \U$30011 ( \30354 , \30351 , \30353 );
not \U$30012 ( \30355 , \30354 );
or \U$30013 ( \30356 , \30349 , \30355 );
not \U$30014 ( \30357 , RI9871aa0_133);
not \U$30015 ( \30358 , \17911 );
or \U$30016 ( \30359 , \30357 , \30358 );
or \U$30017 ( \30360 , \17908 , RI9871aa0_133);
nand \U$30018 ( \30361 , \30359 , \30360 );
nand \U$30019 ( \30362 , \30361 , \2087 );
nand \U$30020 ( \30363 , \30356 , \30362 );
xor \U$30021 ( \30364 , \30348 , \30363 );
not \U$30022 ( \30365 , \30364 );
or \U$30023 ( \30366 , \30331 , \30365 );
nand \U$30024 ( \30367 , \30363 , \30348 );
nand \U$30025 ( \30368 , \30366 , \30367 );
not \U$30026 ( \30369 , \30368 );
and \U$30027 ( \30370 , \30315 , \30369 );
not \U$30028 ( \30371 , \30315 );
and \U$30029 ( \30372 , \30371 , \30368 );
nor \U$30030 ( \30373 , \30370 , \30372 );
not \U$30031 ( \30374 , \30373 );
or \U$30032 ( \30375 , \30300 , \30374 );
nand \U$30033 ( \30376 , \30314 , \30368 );
nand \U$30034 ( \30377 , \30375 , \30376 );
not \U$30035 ( \30378 , \30377 );
not \U$30036 ( \30379 , \30000 );
not \U$30037 ( \30380 , \30011 );
or \U$30038 ( \30381 , \30379 , \30380 );
not \U$30039 ( \30382 , \30000 );
nand \U$30040 ( \30383 , \30382 , \30010 );
nand \U$30041 ( \30384 , \30381 , \30383 );
not \U$30042 ( \30385 , \3163 );
and \U$30043 ( \30386 , RI9872310_151, \20787 );
not \U$30044 ( \30387 , RI9872310_151);
and \U$30045 ( \30388 , \30387 , \22391 );
or \U$30046 ( \30389 , \30386 , \30388 );
not \U$30047 ( \30390 , \30389 );
or \U$30048 ( \30391 , \30385 , \30390 );
nand \U$30049 ( \30392 , \29800 , \3170 );
nand \U$30050 ( \30393 , \30391 , \30392 );
not \U$30051 ( \30394 , \30393 );
xnor \U$30052 ( \30395 , \29763 , \29749 );
not \U$30053 ( \30396 , \30395 );
and \U$30054 ( \30397 , \30394 , \30396 );
and \U$30055 ( \30398 , \30393 , \30395 );
nor \U$30056 ( \30399 , \30397 , \30398 );
not \U$30057 ( \30400 , \30399 );
not \U$30058 ( \30401 , \4918 );
and \U$30059 ( \30402 , RI9872388_152, \18344 );
not \U$30060 ( \30403 , RI9872388_152);
and \U$30061 ( \30404 , \30403 , \9113 );
nor \U$30062 ( \30405 , \30402 , \30404 );
not \U$30063 ( \30406 , \30405 );
or \U$30064 ( \30407 , \30401 , \30406 );
nand \U$30065 ( \30408 , \29351 , \4923 );
nand \U$30066 ( \30409 , \30407 , \30408 );
not \U$30067 ( \30410 , \30409 );
and \U$30068 ( \30411 , \30400 , \30410 );
and \U$30069 ( \30412 , \30399 , \30409 );
nor \U$30070 ( \30413 , \30411 , \30412 );
xor \U$30071 ( \30414 , \30384 , \30413 );
buf \U$30072 ( \30415 , \30026 );
xnor \U$30073 ( \30416 , \30414 , \30415 );
not \U$30074 ( \30417 , \30416 );
or \U$30075 ( \30418 , \30378 , \30417 );
not \U$30076 ( \30419 , \30413 );
xor \U$30077 ( \30420 , \30384 , \30415 );
nand \U$30078 ( \30421 , \30419 , \30420 );
nand \U$30079 ( \30422 , \30418 , \30421 );
not \U$30080 ( \30423 , \30422 );
and \U$30081 ( \30424 , \18704 , \1427 );
not \U$30082 ( \30425 , \1134 );
not \U$30083 ( \30426 , \29944 );
or \U$30084 ( \30427 , \30425 , \30426 );
nand \U$30085 ( \30428 , \30335 , \1082 );
nand \U$30086 ( \30429 , \30427 , \30428 );
xor \U$30087 ( \30430 , \30424 , \30429 );
not \U$30088 ( \30431 , \796 );
not \U$30089 ( \30432 , \29937 );
or \U$30090 ( \30433 , \30431 , \30432 );
not \U$30091 ( \30434 , RI98719b0_131);
not \U$30092 ( \30435 , \28657 );
or \U$30093 ( \30436 , \30434 , \30435 );
or \U$30094 ( \30437 , \20490 , RI98719b0_131);
nand \U$30095 ( \30438 , \30436 , \30437 );
nand \U$30096 ( \30439 , \30438 , \791 );
nand \U$30097 ( \30440 , \30433 , \30439 );
and \U$30098 ( \30441 , \30430 , \30440 );
and \U$30099 ( \30442 , \30424 , \30429 );
nor \U$30100 ( \30443 , \30441 , \30442 );
not \U$30101 ( \30444 , \30443 );
not \U$30102 ( \30445 , \2085 );
not \U$30103 ( \30446 , \29416 );
or \U$30104 ( \30447 , \30445 , \30446 );
nand \U$30105 ( \30448 , \30361 , \2071 );
nand \U$30106 ( \30449 , \30447 , \30448 );
nand \U$30107 ( \30450 , \30444 , \30449 );
not \U$30108 ( \30451 , \30450 );
not \U$30109 ( \30452 , \4918 );
not \U$30110 ( \30453 , \4902 );
not \U$30111 ( \30454 , \9138 );
or \U$30112 ( \30455 , \30453 , \30454 );
nand \U$30113 ( \30456 , \20303 , RI9872388_152);
nand \U$30114 ( \30457 , \30455 , \30456 );
not \U$30115 ( \30458 , \30457 );
or \U$30116 ( \30459 , \30452 , \30458 );
nand \U$30117 ( \30460 , \30405 , \4922 );
nand \U$30118 ( \30461 , \30459 , \30460 );
not \U$30119 ( \30462 , \30461 );
not \U$30120 ( \30463 , \30462 );
or \U$30121 ( \30464 , \30451 , \30463 );
not \U$30122 ( \30465 , \30449 );
nand \U$30123 ( \30466 , \30465 , \30443 );
nand \U$30124 ( \30467 , \30464 , \30466 );
not \U$30125 ( \30468 , \4084 );
not \U$30126 ( \30469 , \30006 );
or \U$30127 ( \30470 , \30468 , \30469 );
not \U$30128 ( \30471 , RI98725e0_157);
not \U$30129 ( \30472 , \11453 );
or \U$30130 ( \30473 , \30471 , \30472 );
or \U$30131 ( \30474 , \11453 , RI98725e0_157);
nand \U$30132 ( \30475 , \30473 , \30474 );
nand \U$30133 ( \30476 , \30475 , \4101 );
nand \U$30134 ( \30477 , \30470 , \30476 );
not \U$30135 ( \30478 , \3170 );
not \U$30136 ( \30479 , \30389 );
or \U$30137 ( \30480 , \30478 , \30479 );
nand \U$30138 ( \30481 , \30328 , \3163 );
nand \U$30139 ( \30482 , \30480 , \30481 );
or \U$30140 ( \30483 , \30477 , \30482 );
and \U$30141 ( \30484 , \29996 , \3467 );
and \U$30142 ( \30485 , RI98726d0_159, \17090 );
not \U$30143 ( \30486 , RI98726d0_159);
and \U$30144 ( \30487 , \30486 , \13281 );
or \U$30145 ( \30488 , \30485 , \30487 );
and \U$30146 ( \30489 , \30488 , \3464 );
nor \U$30147 ( \30490 , \30484 , \30489 );
not \U$30148 ( \30491 , \30490 );
nand \U$30149 ( \30492 , \30483 , \30491 );
nand \U$30150 ( \30493 , \30477 , \30482 );
nand \U$30151 ( \30494 , \30467 , \30492 , \30493 );
not \U$30152 ( \30495 , \30494 );
not \U$30153 ( \30496 , \7188 );
and \U$30154 ( \30497 , RI9872568_156, \8555 );
not \U$30155 ( \30498 , RI9872568_156);
and \U$30156 ( \30499 , \30498 , \10372 );
or \U$30157 ( \30500 , \30497 , \30499 );
not \U$30158 ( \30501 , \30500 );
or \U$30159 ( \30502 , \30496 , \30501 );
xor \U$30160 ( \30503 , \20386 , RI9872568_156);
nand \U$30161 ( \30504 , \30503 , \9320 );
nand \U$30162 ( \30505 , \30502 , \30504 );
not \U$30163 ( \30506 , \30505 );
xor \U$30164 ( \30507 , \29956 , \29939 );
not \U$30165 ( \30508 , \9214 );
not \U$30166 ( \30509 , \21642 );
and \U$30167 ( \30510 , RI9872b80_169, \30509 );
not \U$30168 ( \30511 , RI9872b80_169);
and \U$30169 ( \30512 , \30511 , \18128 );
nor \U$30170 ( \30513 , \30510 , \30512 );
not \U$30171 ( \30514 , \30513 );
or \U$30172 ( \30515 , \30508 , \30514 );
not \U$30173 ( \30516 , RI9872b80_169);
not \U$30174 ( \30517 , \8334 );
or \U$30175 ( \30518 , \30516 , \30517 );
or \U$30176 ( \30519 , \8334 , RI9872b80_169);
nand \U$30177 ( \30520 , \30518 , \30519 );
nand \U$30178 ( \30521 , \30520 , \9196 );
nand \U$30179 ( \30522 , \30515 , \30521 );
xor \U$30180 ( \30523 , \30507 , \30522 );
not \U$30181 ( \30524 , \30523 );
or \U$30182 ( \30525 , \30506 , \30524 );
nand \U$30183 ( \30526 , \30522 , \30507 );
nand \U$30184 ( \30527 , \30525 , \30526 );
not \U$30185 ( \30528 , \30527 );
or \U$30186 ( \30529 , \30495 , \30528 );
not \U$30187 ( \30530 , \30467 );
nand \U$30188 ( \30531 , \30492 , \30493 );
nand \U$30189 ( \30532 , \30530 , \30531 );
nand \U$30190 ( \30533 , \30529 , \30532 );
not \U$30191 ( \30534 , \30533 );
xor \U$30192 ( \30535 , \30232 , \30242 );
xnor \U$30193 ( \30536 , \30535 , \30254 );
nand \U$30194 ( \30537 , \30534 , \30536 );
not \U$30195 ( \30538 , \30537 );
or \U$30196 ( \30539 , \30423 , \30538 );
not \U$30197 ( \30540 , \30536 );
nand \U$30198 ( \30541 , \30540 , \30533 );
nand \U$30199 ( \30542 , \30539 , \30541 );
not \U$30200 ( \30543 , \30542 );
or \U$30201 ( \30544 , \30285 , \30543 );
or \U$30202 ( \30545 , \30542 , \30284 );
xor \U$30203 ( \30546 , \29693 , \29703 );
xor \U$30204 ( \30547 , \30546 , \29713 );
xor \U$30205 ( \30548 , \29636 , \29625 );
xor \U$30206 ( \30549 , \30547 , \30548 );
xor \U$30207 ( \30550 , \29651 , \29666 );
xnor \U$30208 ( \30551 , \30550 , \29678 );
xor \U$30209 ( \30552 , \30549 , \30551 );
nand \U$30210 ( \30553 , \30545 , \30552 );
nand \U$30211 ( \30554 , \30544 , \30553 );
xor \U$30212 ( \30555 , \30267 , \30554 );
xor \U$30213 ( \30556 , \29219 , \29221 );
xor \U$30214 ( \30557 , \30556 , \29224 );
buf \U$30215 ( \30558 , \30229 );
not \U$30216 ( \30559 , \30558 );
xor \U$30217 ( \30560 , \29300 , \29279 );
xnor \U$30218 ( \30561 , \30560 , \29289 );
not \U$30219 ( \30562 , \30561 );
or \U$30220 ( \30563 , \30559 , \30562 );
nand \U$30221 ( \30564 , \30563 , \30256 );
or \U$30222 ( \30565 , \30561 , \30558 );
nand \U$30223 ( \30566 , \30564 , \30565 );
xor \U$30224 ( \30567 , \30557 , \30566 );
xor \U$30225 ( \30568 , \30547 , \30548 );
and \U$30226 ( \30569 , \30568 , \30551 );
and \U$30227 ( \30570 , \30547 , \30548 );
or \U$30228 ( \30571 , \30569 , \30570 );
xor \U$30229 ( \30572 , \30567 , \30571 );
and \U$30230 ( \30573 , \30555 , \30572 );
and \U$30231 ( \30574 , \30267 , \30554 );
or \U$30232 ( \30575 , \30573 , \30574 );
xor \U$30233 ( \30576 , \30118 , \30575 );
xor \U$30234 ( \30577 , \29786 , \29817 );
xor \U$30235 ( \30578 , \30577 , \29828 );
not \U$30236 ( \30579 , \30578 );
not \U$30237 ( \30580 , \5035 );
not \U$30238 ( \30581 , \29360 );
or \U$30239 ( \30582 , \30580 , \30581 );
and \U$30240 ( \30583 , RI9872478_154, \8696 );
not \U$30241 ( \30584 , RI9872478_154);
and \U$30242 ( \30585 , \30584 , \9750 );
or \U$30243 ( \30586 , \30583 , \30585 );
nand \U$30244 ( \30587 , \30586 , \5034 );
nand \U$30245 ( \30588 , \30582 , \30587 );
not \U$30246 ( \30589 , \30588 );
not \U$30247 ( \30590 , \9249 );
not \U$30248 ( \30591 , \9244 );
not \U$30249 ( \30592 , \7905 );
or \U$30250 ( \30593 , \30591 , \30592 );
nand \U$30251 ( \30594 , \15875 , RI9872bf8_170);
nand \U$30252 ( \30595 , \30593 , \30594 );
not \U$30253 ( \30596 , \30595 );
or \U$30254 ( \30597 , \30590 , \30596 );
nand \U$30255 ( \30598 , \29494 , \22167 );
nand \U$30256 ( \30599 , \30597 , \30598 );
not \U$30257 ( \30600 , \30599 );
or \U$30258 ( \30601 , \30589 , \30600 );
or \U$30259 ( \30602 , \30599 , \30588 );
not \U$30260 ( \30603 , \5642 );
not \U$30261 ( \30604 , \30500 );
or \U$30262 ( \30605 , \30603 , \30604 );
nand \U$30263 ( \30606 , \29371 , \5653 );
nand \U$30264 ( \30607 , \30605 , \30606 );
nand \U$30265 ( \30608 , \30602 , \30607 );
nand \U$30266 ( \30609 , \30601 , \30608 );
not \U$30267 ( \30610 , \30609 );
not \U$30268 ( \30611 , \30409 );
not \U$30269 ( \30612 , \30399 );
not \U$30270 ( \30613 , \30612 );
or \U$30271 ( \30614 , \30611 , \30613 );
not \U$30272 ( \30615 , \30395 );
nand \U$30273 ( \30616 , \30615 , \30393 );
nand \U$30274 ( \30617 , \30614 , \30616 );
not \U$30275 ( \30618 , \30617 );
not \U$30276 ( \30619 , \8027 );
not \U$30277 ( \30620 , \30305 );
or \U$30278 ( \30621 , \30619 , \30620 );
nand \U$30279 ( \30622 , \29481 , \8039 );
nand \U$30280 ( \30623 , \30621 , \30622 );
not \U$30281 ( \30624 , \30623 );
not \U$30282 ( \30625 , \30624 );
not \U$30283 ( \30626 , \7326 );
not \U$30284 ( \30627 , \30291 );
or \U$30285 ( \30628 , \30626 , \30627 );
nand \U$30286 ( \30629 , \29465 , \7338 );
nand \U$30287 ( \30630 , \30628 , \30629 );
not \U$30288 ( \30631 , \30630 );
not \U$30289 ( \30632 , \30631 );
or \U$30290 ( \30633 , \30625 , \30632 );
not \U$30291 ( \30634 , \9196 );
not \U$30292 ( \30635 , \30513 );
or \U$30293 ( \30636 , \30634 , \30635 );
nand \U$30294 ( \30637 , \29507 , \9214 );
nand \U$30295 ( \30638 , \30636 , \30637 );
nand \U$30296 ( \30639 , \30633 , \30638 );
not \U$30297 ( \30640 , \30624 );
nand \U$30298 ( \30641 , \30640 , \30630 );
and \U$30299 ( \30642 , \30639 , \30641 );
not \U$30300 ( \30643 , \30642 );
or \U$30301 ( \30644 , \30618 , \30643 );
not \U$30302 ( \30645 , \30641 );
not \U$30303 ( \30646 , \30639 );
or \U$30304 ( \30647 , \30645 , \30646 );
not \U$30305 ( \30648 , \30617 );
nand \U$30306 ( \30649 , \30647 , \30648 );
nand \U$30307 ( \30650 , \30644 , \30649 );
not \U$30308 ( \30651 , \30650 );
or \U$30309 ( \30652 , \30610 , \30651 );
not \U$30310 ( \30653 , \30641 );
not \U$30311 ( \30654 , \30639 );
or \U$30312 ( \30655 , \30653 , \30654 );
nand \U$30313 ( \30656 , \30655 , \30617 );
nand \U$30314 ( \30657 , \30652 , \30656 );
not \U$30315 ( \30658 , \30657 );
nand \U$30316 ( \30659 , \30579 , \30658 );
not \U$30317 ( \30660 , \30659 );
not \U$30318 ( \30661 , \9937 );
not \U$30319 ( \30662 , \30250 );
or \U$30320 ( \30663 , \30661 , \30662 );
and \U$30321 ( \30664 , RI9873030_179, \5205 );
not \U$30322 ( \30665 , RI9873030_179);
and \U$30323 ( \30666 , \30665 , \5611 );
or \U$30324 ( \30667 , \30664 , \30666 );
nand \U$30325 ( \30668 , \30667 , \19321 );
nand \U$30326 ( \30669 , \30663 , \30668 );
not \U$30327 ( \30670 , \30669 );
not \U$30328 ( \30671 , \30240 );
not \U$30329 ( \30672 , \19282 );
or \U$30330 ( \30673 , \30671 , \30672 );
xor \U$30331 ( \30674 , \1168 , RI98733f0_187);
buf \U$30332 ( \30675 , \1183 );
xnor \U$30333 ( \30676 , \30674 , \30675 );
or \U$30334 ( \30677 , \30676 , \18079 );
nand \U$30335 ( \30678 , \30673 , \30677 );
not \U$30336 ( \30679 , \30678 );
xor \U$30337 ( \30680 , \29439 , \29449 );
xnor \U$30338 ( \30681 , \30680 , \29418 );
not \U$30339 ( \30682 , \30681 );
and \U$30340 ( \30683 , \30679 , \30682 );
and \U$30341 ( \30684 , \30678 , \30681 );
nor \U$30342 ( \30685 , \30683 , \30684 );
not \U$30343 ( \30686 , \30685 );
not \U$30344 ( \30687 , \30686 );
or \U$30345 ( \30688 , \30670 , \30687 );
not \U$30346 ( \30689 , \30681 );
nand \U$30347 ( \30690 , \30689 , \30678 );
nand \U$30348 ( \30691 , \30688 , \30690 );
not \U$30349 ( \30692 , \30691 );
not \U$30350 ( \30693 , \18615 );
xor \U$30351 ( \30694 , RI9873558_190, \1365 );
not \U$30352 ( \30695 , \30694 );
or \U$30353 ( \30696 , \30693 , \30695 );
nand \U$30354 ( \30697 , \30058 , RI9873648_192);
nand \U$30355 ( \30698 , \30696 , \30697 );
not \U$30356 ( \30699 , \19243 );
xor \U$30357 ( \30700 , RI98734e0_189, \18571 );
not \U$30358 ( \30701 , \30700 );
or \U$30359 ( \30702 , \30699 , \30701 );
nand \U$30360 ( \30703 , \30169 , \20147 );
nand \U$30361 ( \30704 , \30702 , \30703 );
and \U$30362 ( \30705 , \30698 , \30704 );
not \U$30363 ( \30706 , \30705 );
xor \U$30364 ( \30707 , \30698 , \30704 );
not \U$30365 ( \30708 , \17123 );
not \U$30366 ( \30709 , \30158 );
or \U$30367 ( \30710 , \30708 , \30709 );
xor \U$30368 ( \30711 , RI9873210_183, \3239 );
nand \U$30369 ( \30712 , \30711 , \13477 );
nand \U$30370 ( \30713 , \30710 , \30712 );
nand \U$30371 ( \30714 , \30707 , \30713 );
nand \U$30372 ( \30715 , \30706 , \30714 );
nand \U$30373 ( \30716 , \29472 , \29456 );
xnor \U$30374 ( \30717 , \30716 , \29467 );
xor \U$30375 ( \30718 , \30715 , \30717 );
not \U$30376 ( \30719 , \30718 );
or \U$30377 ( \30720 , \30692 , \30719 );
not \U$30378 ( \30721 , \30705 );
not \U$30379 ( \30722 , \30721 );
not \U$30380 ( \30723 , \30714 );
or \U$30381 ( \30724 , \30722 , \30723 );
nand \U$30382 ( \30725 , \30724 , \30717 );
nand \U$30383 ( \30726 , \30720 , \30725 );
not \U$30384 ( \30727 , \30726 );
or \U$30385 ( \30728 , \30660 , \30727 );
nand \U$30386 ( \30729 , \30657 , \30578 );
nand \U$30387 ( \30730 , \30728 , \30729 );
not \U$30388 ( \30731 , \30730 );
xnor \U$30389 ( \30732 , \29522 , \29342 );
not \U$30390 ( \30733 , \30732 );
and \U$30391 ( \30734 , \30731 , \30733 );
and \U$30392 ( \30735 , \30730 , \30732 );
nor \U$30393 ( \30736 , \30734 , \30735 );
not \U$30394 ( \30737 , \30074 );
nand \U$30395 ( \30738 , \30737 , \30076 );
not \U$30396 ( \30739 , \30738 );
not \U$30397 ( \30740 , \30071 );
or \U$30398 ( \30741 , \30739 , \30740 );
not \U$30399 ( \30742 , \30076 );
nand \U$30400 ( \30743 , \30742 , \30074 );
nand \U$30401 ( \30744 , \30741 , \30743 );
not \U$30402 ( \30745 , \30744 );
not \U$30403 ( \30746 , \29681 );
not \U$30404 ( \30747 , \29716 );
and \U$30405 ( \30748 , \29640 , \30747 );
not \U$30406 ( \30749 , \29640 );
and \U$30407 ( \30750 , \30749 , \29716 );
nor \U$30408 ( \30751 , \30748 , \30750 );
not \U$30409 ( \30752 , \30751 );
or \U$30410 ( \30753 , \30746 , \30752 );
not \U$30411 ( \30754 , \30751 );
not \U$30412 ( \30755 , \29681 );
nand \U$30413 ( \30756 , \30754 , \30755 );
nand \U$30414 ( \30757 , \30753 , \30756 );
xor \U$30415 ( \30758 , \30745 , \30757 );
not \U$30416 ( \30759 , \30279 );
not \U$30417 ( \30760 , \30274 );
or \U$30418 ( \30761 , \30759 , \30760 );
not \U$30419 ( \30762 , \30271 );
not \U$30420 ( \30763 , \30270 );
or \U$30421 ( \30764 , \30762 , \30763 );
nand \U$30422 ( \30765 , \30764 , \30273 );
nand \U$30423 ( \30766 , \30761 , \30765 );
not \U$30424 ( \30767 , \30766 );
xnor \U$30425 ( \30768 , \30758 , \30767 );
or \U$30426 ( \30769 , \30736 , \30768 );
not \U$30427 ( \30770 , \30732 );
nand \U$30428 ( \30771 , \30770 , \30730 );
nand \U$30429 ( \30772 , \30769 , \30771 );
and \U$30430 ( \30773 , \30576 , \30772 );
and \U$30431 ( \30774 , \30118 , \30575 );
or \U$30432 ( \30775 , \30773 , \30774 );
nand \U$30433 ( \30776 , \30116 , \30775 );
buf \U$30434 ( \30777 , \29897 );
nand \U$30435 ( \30778 , \30777 , \30114 );
nand \U$30436 ( \30779 , \30776 , \30778 );
xor \U$30437 ( \30780 , \29322 , \29319 );
xnor \U$30438 ( \30781 , \30780 , \29316 );
not \U$30439 ( \30782 , \30757 );
and \U$30440 ( \30783 , \30766 , \30744 );
not \U$30441 ( \30784 , \30766 );
and \U$30442 ( \30785 , \30784 , \30745 );
nor \U$30443 ( \30786 , \30783 , \30785 );
not \U$30444 ( \30787 , \30786 );
or \U$30445 ( \30788 , \30782 , \30787 );
not \U$30446 ( \30789 , \30767 );
nand \U$30447 ( \30790 , \30789 , \30744 );
nand \U$30448 ( \30791 , \30788 , \30790 );
not \U$30449 ( \30792 , \30791 );
or \U$30450 ( \30793 , \30566 , \30557 );
and \U$30451 ( \30794 , \30793 , \30571 );
and \U$30452 ( \30795 , \30566 , \30557 );
nor \U$30453 ( \30796 , \30794 , \30795 );
not \U$30454 ( \30797 , \30796 );
and \U$30455 ( \30798 , \29312 , \29227 );
not \U$30456 ( \30799 , \29312 );
not \U$30457 ( \30800 , \29227 );
and \U$30458 ( \30801 , \30799 , \30800 );
nor \U$30459 ( \30802 , \30798 , \30801 );
not \U$30460 ( \30803 , \30802 );
or \U$30461 ( \30804 , \30797 , \30803 );
or \U$30462 ( \30805 , \30802 , \30796 );
nand \U$30463 ( \30806 , \30804 , \30805 );
not \U$30464 ( \30807 , \30806 );
or \U$30465 ( \30808 , \30792 , \30807 );
not \U$30466 ( \30809 , \30796 );
nand \U$30467 ( \30810 , \30809 , \30802 );
nand \U$30468 ( \30811 , \30808 , \30810 );
not \U$30469 ( \30812 , \30811 );
xor \U$30470 ( \30813 , \30781 , \30812 );
not \U$30471 ( \30814 , \29851 );
nand \U$30472 ( \30815 , \30814 , \29853 );
and \U$30473 ( \30816 , \30815 , \29612 );
not \U$30474 ( \30817 , \30815 );
and \U$30475 ( \30818 , \30817 , \29613 );
nor \U$30476 ( \30819 , \30816 , \30818 );
and \U$30477 ( \30820 , \30813 , \30819 );
and \U$30478 ( \30821 , \30781 , \30812 );
or \U$30479 ( \30822 , \30820 , \30821 );
xnor \U$30480 ( \30823 , \30779 , \30822 );
not \U$30481 ( \30824 , \30823 );
or \U$30482 ( \30825 , \29895 , \30824 );
nand \U$30483 ( \30826 , \30776 , \30778 , \30822 );
nand \U$30484 ( \30827 , \30825 , \30826 );
nand \U$30485 ( \30828 , \29891 , \30827 );
not \U$30486 ( \30829 , \29893 );
not \U$30487 ( \30830 , \30823 );
or \U$30488 ( \30831 , \30829 , \30830 );
or \U$30489 ( \30832 , \30823 , \29893 );
nand \U$30490 ( \30833 , \30831 , \30832 );
xor \U$30491 ( \30834 , \30114 , \30777 );
not \U$30492 ( \30835 , \30775 );
xnor \U$30493 ( \30836 , \30834 , \30835 );
not \U$30494 ( \30837 , \30836 );
not \U$30495 ( \30838 , \30837 );
xor \U$30496 ( \30839 , \30781 , \30812 );
xor \U$30497 ( \30840 , \30839 , \30819 );
not \U$30498 ( \30841 , \30840 );
or \U$30499 ( \30842 , \30838 , \30841 );
not \U$30500 ( \30843 , \30840 );
not \U$30501 ( \30844 , \30843 );
not \U$30502 ( \30845 , \30836 );
or \U$30503 ( \30846 , \30844 , \30845 );
and \U$30504 ( \30847 , \30736 , \30768 );
not \U$30505 ( \30848 , \30736 );
not \U$30506 ( \30849 , \30768 );
and \U$30507 ( \30850 , \30848 , \30849 );
nor \U$30508 ( \30851 , \30847 , \30850 );
not \U$30509 ( \30852 , \30851 );
xor \U$30510 ( \30853 , \29913 , \30040 );
xor \U$30511 ( \30854 , \30853 , \30081 );
not \U$30512 ( \30855 , \30854 );
xor \U$30513 ( \30856 , \30578 , \30658 );
xor \U$30514 ( \30857 , \30856 , \30726 );
not \U$30515 ( \30858 , \30857 );
or \U$30516 ( \30859 , \30855 , \30858 );
not \U$30517 ( \30860 , \13020 );
and \U$30518 ( \30861 , RI98730a8_180, \5596 );
not \U$30519 ( \30862 , RI98730a8_180);
and \U$30520 ( \30863 , \30862 , \4177 );
or \U$30521 ( \30864 , \30861 , \30863 );
not \U$30522 ( \30865 , \30864 );
or \U$30523 ( \30866 , \30860 , \30865 );
nand \U$30524 ( \30867 , \30201 , \12868 );
nand \U$30525 ( \30868 , \30866 , \30867 );
not \U$30526 ( \30869 , \30868 );
not \U$30527 ( \30870 , \19046 );
not \U$30528 ( \30871 , \30700 );
or \U$30529 ( \30872 , \30870 , \30871 );
xor \U$30530 ( \30873 , RI98734e0_189, \20637 );
nand \U$30531 ( \30874 , \30873 , \19244 );
nand \U$30532 ( \30875 , \30872 , \30874 );
not \U$30533 ( \30876 , \30875 );
not \U$30534 ( \30877 , \30676 );
not \U$30535 ( \30878 , \17620 );
and \U$30536 ( \30879 , \30877 , \30878 );
not \U$30537 ( \30880 , \17539 );
not \U$30538 ( \30881 , \30142 );
or \U$30539 ( \30882 , \30880 , \30881 );
or \U$30540 ( \30883 , \30142 , \17539 );
nand \U$30541 ( \30884 , \30882 , \30883 );
not \U$30542 ( \30885 , \30884 );
not \U$30543 ( \30886 , \17251 );
nor \U$30544 ( \30887 , \30885 , \30886 );
nor \U$30545 ( \30888 , \30879 , \30887 );
not \U$30546 ( \30889 , \30888 );
or \U$30547 ( \30890 , \30876 , \30889 );
or \U$30548 ( \30891 , \30888 , \30875 );
nand \U$30549 ( \30892 , \30890 , \30891 );
not \U$30550 ( \30893 , \30892 );
or \U$30551 ( \30894 , \30869 , \30893 );
not \U$30552 ( \30895 , \30888 );
nand \U$30553 ( \30896 , \30895 , \30875 );
nand \U$30554 ( \30897 , \30894 , \30896 );
not \U$30555 ( \30898 , \30897 );
xor \U$30556 ( \30899 , \29982 , \29928 );
not \U$30557 ( \30900 , \30899 );
not \U$30558 ( \30901 , \22167 );
not \U$30559 ( \30902 , \30595 );
or \U$30560 ( \30903 , \30901 , \30902 );
xor \U$30561 ( \30904 , \17072 , RI9872bf8_170);
not \U$30562 ( \30905 , \30904 );
nand \U$30563 ( \30906 , \30905 , \9249 );
nand \U$30564 ( \30907 , \30903 , \30906 );
not \U$30565 ( \30908 , \30907 );
not \U$30566 ( \30909 , \8801 );
not \U$30567 ( \30910 , \30018 );
or \U$30568 ( \30911 , \30909 , \30910 );
and \U$30569 ( \30912 , RI9872d60_173, \6296 );
not \U$30570 ( \30913 , RI9872d60_173);
and \U$30571 ( \30914 , \30913 , \8052 );
nor \U$30572 ( \30915 , \30912 , \30914 );
nand \U$30573 ( \30916 , \30915 , \22664 );
nand \U$30574 ( \30917 , \30911 , \30916 );
not \U$30575 ( \30918 , \5035 );
not \U$30576 ( \30919 , \30586 );
or \U$30577 ( \30920 , \30918 , \30919 );
and \U$30578 ( \30921 , \5025 , \9849 );
not \U$30579 ( \30922 , \5025 );
and \U$30580 ( \30923 , \30922 , \8707 );
nor \U$30581 ( \30924 , \30921 , \30923 );
nand \U$30582 ( \30925 , \30924 , \5034 );
nand \U$30583 ( \30926 , \30920 , \30925 );
and \U$30584 ( \30927 , \30917 , \30926 );
not \U$30585 ( \30928 , \30917 );
not \U$30586 ( \30929 , \30926 );
and \U$30587 ( \30930 , \30928 , \30929 );
nor \U$30588 ( \30931 , \30927 , \30930 );
not \U$30589 ( \30932 , \30931 );
or \U$30590 ( \30933 , \30908 , \30932 );
nand \U$30591 ( \30934 , \30917 , \30926 );
nand \U$30592 ( \30935 , \30933 , \30934 );
not \U$30593 ( \30936 , \30935 );
not \U$30594 ( \30937 , \30936 );
or \U$30595 ( \30938 , \30900 , \30937 );
or \U$30596 ( \30939 , \30936 , \30899 );
nand \U$30597 ( \30940 , \30938 , \30939 );
not \U$30598 ( \30941 , \30940 );
or \U$30599 ( \30942 , \30898 , \30941 );
not \U$30600 ( \30943 , \30936 );
nand \U$30601 ( \30944 , \30943 , \30899 );
nand \U$30602 ( \30945 , \30942 , \30944 );
not \U$30603 ( \30946 , \30945 );
and \U$30604 ( \30947 , \30630 , \30623 );
not \U$30605 ( \30948 , \30630 );
and \U$30606 ( \30949 , \30948 , \30624 );
nor \U$30607 ( \30950 , \30947 , \30949 );
xor \U$30608 ( \30951 , \30950 , \30638 );
not \U$30609 ( \30952 , \9272 );
not \U$30610 ( \30953 , \30193 );
or \U$30611 ( \30954 , \30952 , \30953 );
not \U$30612 ( \30955 , RI9872e50_175);
not \U$30613 ( \30956 , \5761 );
or \U$30614 ( \30957 , \30955 , \30956 );
or \U$30615 ( \30958 , \5761 , RI9872e50_175);
nand \U$30616 ( \30959 , \30957 , \30958 );
nand \U$30617 ( \30960 , \30959 , \18562 );
nand \U$30618 ( \30961 , \30954 , \30960 );
not \U$30619 ( \30962 , \30961 );
buf \U$30620 ( \30963 , \13483 );
not \U$30621 ( \30964 , \30963 );
not \U$30622 ( \30965 , \30711 );
or \U$30623 ( \30966 , \30964 , \30965 );
and \U$30624 ( \30967 , RI9873210_183, \3536 );
not \U$30625 ( \30968 , RI9873210_183);
and \U$30626 ( \30969 , \30968 , \3541 );
nor \U$30627 ( \30970 , \30967 , \30969 );
nand \U$30628 ( \30971 , \30970 , \13476 );
nand \U$30629 ( \30972 , \30966 , \30971 );
not \U$30630 ( \30973 , \30972 );
or \U$30631 ( \30974 , \30962 , \30973 );
or \U$30632 ( \30975 , \30972 , \30961 );
not \U$30633 ( \30976 , RI9873648_192);
not \U$30634 ( \30977 , \30694 );
or \U$30635 ( \30978 , \30976 , \30977 );
and \U$30636 ( \30979 , RI9873558_190, \1061 );
not \U$30637 ( \30980 , RI9873558_190);
and \U$30638 ( \30981 , \30980 , \23043 );
nor \U$30639 ( \30982 , \30979 , \30981 );
nand \U$30640 ( \30983 , \30982 , \18615 );
nand \U$30641 ( \30984 , \30978 , \30983 );
nand \U$30642 ( \30985 , \30975 , \30984 );
nand \U$30643 ( \30986 , \30974 , \30985 );
nor \U$30644 ( \30987 , \30951 , \30986 );
xnor \U$30645 ( \30988 , \30607 , \30588 );
xor \U$30646 ( \30989 , \30599 , \30988 );
or \U$30647 ( \30990 , \30987 , \30989 );
nand \U$30648 ( \30991 , \30951 , \30986 );
nand \U$30649 ( \30992 , \30990 , \30991 );
not \U$30650 ( \30993 , \30992 );
xnor \U$30651 ( \30994 , \30035 , \29987 );
not \U$30652 ( \30995 , \30994 );
or \U$30653 ( \30996 , \30993 , \30995 );
or \U$30654 ( \30997 , \30994 , \30992 );
nand \U$30655 ( \30998 , \30996 , \30997 );
not \U$30656 ( \30999 , \30998 );
or \U$30657 ( \31000 , \30946 , \30999 );
not \U$30658 ( \31001 , \30994 );
nand \U$30659 ( \31002 , \31001 , \30992 );
nand \U$30660 ( \31003 , \31000 , \31002 );
nand \U$30661 ( \31004 , \30859 , \31003 );
not \U$30662 ( \31005 , \30854 );
not \U$30663 ( \31006 , \30857 );
nand \U$30664 ( \31007 , \31005 , \31006 );
and \U$30665 ( \31008 , \31004 , \31007 );
nand \U$30666 ( \31009 , \30088 , \29903 );
and \U$30667 ( \31010 , \31009 , \30084 );
not \U$30668 ( \31011 , \31009 );
not \U$30669 ( \31012 , \30084 );
and \U$30670 ( \31013 , \31011 , \31012 );
nor \U$30671 ( \31014 , \31010 , \31013 );
and \U$30672 ( \31015 , \31008 , \31014 );
not \U$30673 ( \31016 , \31008 );
not \U$30674 ( \31017 , \31014 );
and \U$30675 ( \31018 , \31016 , \31017 );
nor \U$30676 ( \31019 , \31015 , \31018 );
not \U$30677 ( \31020 , \31019 );
or \U$30678 ( \31021 , \30852 , \31020 );
not \U$30679 ( \31022 , \31007 );
not \U$30680 ( \31023 , \31004 );
or \U$30681 ( \31024 , \31022 , \31023 );
nand \U$30682 ( \31025 , \31024 , \31017 );
nand \U$30683 ( \31026 , \31021 , \31025 );
not \U$30684 ( \31027 , \31026 );
not \U$30685 ( \31028 , \30791 );
not \U$30686 ( \31029 , \31028 );
not \U$30687 ( \31030 , \30806 );
and \U$30688 ( \31031 , \31029 , \31030 );
and \U$30689 ( \31032 , \30806 , \31028 );
nor \U$30690 ( \31033 , \31031 , \31032 );
not \U$30691 ( \31034 , \31033 );
xor \U$30692 ( \31035 , \30096 , \30089 );
xnor \U$30693 ( \31036 , \31035 , \30105 );
not \U$30694 ( \31037 , \31036 );
or \U$30695 ( \31038 , \31034 , \31037 );
or \U$30696 ( \31039 , \31036 , \31033 );
nand \U$30697 ( \31040 , \31038 , \31039 );
not \U$30698 ( \31041 , \31040 );
or \U$30699 ( \31042 , \31027 , \31041 );
not \U$30700 ( \31043 , \31033 );
nand \U$30701 ( \31044 , \31043 , \31036 );
nand \U$30702 ( \31045 , \31042 , \31044 );
not \U$30703 ( \31046 , \31045 );
nand \U$30704 ( \31047 , \30846 , \31046 );
nand \U$30705 ( \31048 , \30842 , \31047 );
nand \U$30706 ( \31049 , \30833 , \31048 );
and \U$30707 ( \31050 , \30828 , \31049 );
xor \U$30708 ( \31051 , \28616 , \29082 );
xor \U$30709 ( \31052 , \31051 , \29085 );
xor \U$30710 ( \31053 , \28477 , \28580 );
xor \U$30711 ( \31054 , \31053 , \28583 );
nand \U$30712 ( \31055 , \29880 , \29878 );
not \U$30713 ( \31056 , \31055 );
not \U$30714 ( \31057 , \29880 );
not \U$30715 ( \31058 , \29878 );
and \U$30716 ( \31059 , \31057 , \31058 );
nor \U$30717 ( \31060 , \31059 , \29889 );
nor \U$30718 ( \31061 , \31056 , \31060 );
xor \U$30719 ( \31062 , \31054 , \31061 );
and \U$30720 ( \31063 , \28994 , \28618 );
not \U$30721 ( \31064 , \28994 );
and \U$30722 ( \31065 , \31064 , \29080 );
nor \U$30723 ( \31066 , \31063 , \31065 );
xnor \U$30724 ( \31067 , \29078 , \31066 );
and \U$30725 ( \31068 , \31062 , \31067 );
and \U$30726 ( \31069 , \31054 , \31061 );
or \U$30727 ( \31070 , \31068 , \31069 );
nand \U$30728 ( \31071 , \31052 , \31070 );
xor \U$30729 ( \31072 , \31054 , \31061 );
xor \U$30730 ( \31073 , \31072 , \31067 );
not \U$30731 ( \31074 , \29093 );
not \U$30732 ( \31075 , \31074 );
not \U$30733 ( \31076 , \29890 );
or \U$30734 ( \31077 , \31075 , \31076 );
not \U$30735 ( \31078 , \29873 );
nand \U$30736 ( \31079 , \31077 , \31078 );
not \U$30737 ( \31080 , \29890 );
nand \U$30738 ( \31081 , \31080 , \29093 );
nand \U$30739 ( \31082 , \31079 , \31081 );
not \U$30740 ( \31083 , \31082 );
nand \U$30741 ( \31084 , \31073 , \31083 );
and \U$30742 ( \31085 , \31050 , \31071 , \31084 );
xor \U$30743 ( \31086 , \30223 , \30265 );
xnor \U$30744 ( \31087 , \31086 , \30188 );
not \U$30745 ( \31088 , \31087 );
not \U$30746 ( \31089 , \31088 );
not \U$30747 ( \31090 , \30184 );
not \U$30748 ( \31091 , \30120 );
or \U$30749 ( \31092 , \31090 , \31091 );
or \U$30750 ( \31093 , \30120 , \30184 );
nand \U$30751 ( \31094 , \31092 , \31093 );
and \U$30752 ( \31095 , \31094 , \30150 );
not \U$30753 ( \31096 , \31094 );
and \U$30754 ( \31097 , \31096 , \30149 );
nor \U$30755 ( \31098 , \31095 , \31097 );
not \U$30756 ( \31099 , \11198 );
not \U$30757 ( \31100 , \29919 );
or \U$30758 ( \31101 , \31099 , \31100 );
not \U$30759 ( \31102 , RI9872f40_177);
not \U$30760 ( \31103 , \5736 );
or \U$30761 ( \31104 , \31102 , \31103 );
or \U$30762 ( \31105 , \5736 , RI9872f40_177);
nand \U$30763 ( \31106 , \31104 , \31105 );
nand \U$30764 ( \31107 , \31106 , \8743 );
nand \U$30765 ( \31108 , \31101 , \31107 );
not \U$30766 ( \31109 , \31108 );
not \U$30767 ( \31110 , \17528 );
not \U$30768 ( \31111 , \30208 );
or \U$30769 ( \31112 , \31110 , \31111 );
not \U$30770 ( \31113 , RI9873288_184);
not \U$30771 ( \31114 , \2947 );
or \U$30772 ( \31115 , \31113 , \31114 );
or \U$30773 ( \31116 , \2947 , RI9873288_184);
nand \U$30774 ( \31117 , \31115 , \31116 );
nand \U$30775 ( \31118 , \31117 , \18508 );
nand \U$30776 ( \31119 , \31112 , \31118 );
not \U$30777 ( \31120 , \6286 );
not \U$30778 ( \31121 , \29969 );
or \U$30779 ( \31122 , \31120 , \31121 );
not \U$30780 ( \31123 , RI98728b0_163);
not \U$30781 ( \31124 , \18309 );
or \U$30782 ( \31125 , \31123 , \31124 );
nand \U$30783 ( \31126 , \8580 , \7049 );
nand \U$30784 ( \31127 , \31125 , \31126 );
nand \U$30785 ( \31128 , \31127 , \6284 );
nand \U$30786 ( \31129 , \31122 , \31128 );
and \U$30787 ( \31130 , \31119 , \31129 );
not \U$30788 ( \31131 , \31119 );
not \U$30789 ( \31132 , \31129 );
and \U$30790 ( \31133 , \31131 , \31132 );
nor \U$30791 ( \31134 , \31130 , \31133 );
not \U$30792 ( \31135 , \31134 );
or \U$30793 ( \31136 , \31109 , \31135 );
nand \U$30794 ( \31137 , \31119 , \31129 );
nand \U$30795 ( \31138 , \31136 , \31137 );
not \U$30796 ( \31139 , \31138 );
not \U$30797 ( \31140 , \9937 );
not \U$30798 ( \31141 , \30667 );
or \U$30799 ( \31142 , \31140 , \31141 );
and \U$30800 ( \31143 , RI9873030_179, \12971 );
not \U$30801 ( \31144 , RI9873030_179);
and \U$30802 ( \31145 , \31144 , \5623 );
or \U$30803 ( \31146 , \31143 , \31145 );
nand \U$30804 ( \31147 , \31146 , \19321 );
nand \U$30805 ( \31148 , \31142 , \31147 );
not \U$30806 ( \31149 , \31148 );
xor \U$30807 ( \31150 , \30449 , \30443 );
and \U$30808 ( \31151 , \31150 , \30461 );
not \U$30809 ( \31152 , \31150 );
and \U$30810 ( \31153 , \31152 , \30462 );
or \U$30811 ( \31154 , \31151 , \31153 );
not \U$30812 ( \31155 , \3467 );
not \U$30813 ( \31156 , \30488 );
or \U$30814 ( \31157 , \31155 , \31156 );
not \U$30815 ( \31158 , RI98726d0_159);
not \U$30816 ( \31159 , \24758 );
or \U$30817 ( \31160 , \31158 , \31159 );
or \U$30818 ( \31161 , \22392 , RI98726d0_159);
nand \U$30819 ( \31162 , \31160 , \31161 );
nand \U$30820 ( \31163 , \31162 , \3465 );
nand \U$30821 ( \31164 , \31157 , \31163 );
not \U$30822 ( \31165 , \31164 );
xnor \U$30823 ( \31166 , \30440 , \30430 );
not \U$30824 ( \31167 , \31166 );
not \U$30825 ( \31168 , \4101 );
not \U$30826 ( \31169 , RI98725e0_157);
not \U$30827 ( \31170 , \12772 );
or \U$30828 ( \31171 , \31169 , \31170 );
or \U$30829 ( \31172 , \12772 , RI98725e0_157);
nand \U$30830 ( \31173 , \31171 , \31172 );
not \U$30831 ( \31174 , \31173 );
or \U$30832 ( \31175 , \31168 , \31174 );
not \U$30833 ( \31176 , \4084 );
not \U$30834 ( \31177 , \31176 );
nand \U$30835 ( \31178 , \31177 , \30475 );
nand \U$30836 ( \31179 , \31175 , \31178 );
not \U$30837 ( \31180 , \31179 );
or \U$30838 ( \31181 , \31167 , \31180 );
or \U$30839 ( \31182 , \31179 , \31166 );
nand \U$30840 ( \31183 , \31181 , \31182 );
not \U$30841 ( \31184 , \31183 );
or \U$30842 ( \31185 , \31165 , \31184 );
not \U$30843 ( \31186 , \31166 );
nand \U$30844 ( \31187 , \31186 , \31179 );
nand \U$30845 ( \31188 , \31185 , \31187 );
and \U$30846 ( \31189 , \31154 , \31188 );
not \U$30847 ( \31190 , \31154 );
not \U$30848 ( \31191 , \31188 );
and \U$30849 ( \31192 , \31190 , \31191 );
nor \U$30850 ( \31193 , \31189 , \31192 );
not \U$30851 ( \31194 , \31193 );
or \U$30852 ( \31195 , \31149 , \31194 );
nand \U$30853 ( \31196 , \31188 , \31154 );
nand \U$30854 ( \31197 , \31195 , \31196 );
not \U$30855 ( \31198 , \31197 );
nand \U$30856 ( \31199 , \31139 , \31198 );
xor \U$30857 ( \31200 , \30707 , \30713 );
and \U$30858 ( \31201 , \31199 , \31200 );
nor \U$30859 ( \31202 , \31139 , \31198 );
nor \U$30860 ( \31203 , \31201 , \31202 );
nand \U$30861 ( \31204 , \31098 , \31203 );
not \U$30862 ( \31205 , \31204 );
not \U$30863 ( \31206 , \796 );
not \U$30864 ( \31207 , \30438 );
or \U$30865 ( \31208 , \31206 , \31207 );
and \U$30866 ( \31209 , \1078 , \19542 );
not \U$30867 ( \31210 , \1078 );
and \U$30868 ( \31211 , \31210 , \17862 );
nor \U$30869 ( \31212 , \31209 , \31211 );
nand \U$30870 ( \31213 , \31212 , \791 );
nand \U$30871 ( \31214 , \31208 , \31213 );
not \U$30872 ( \31215 , \30344 );
not \U$30873 ( \31216 , \30346 );
and \U$30874 ( \31217 , \31215 , \31216 );
and \U$30875 ( \31218 , \30344 , \30346 );
nor \U$30876 ( \31219 , \31217 , \31218 );
xnor \U$30877 ( \31220 , \31214 , \31219 );
not \U$30878 ( \31221 , \31220 );
not \U$30879 ( \31222 , \3169 );
not \U$30880 ( \31223 , \30322 );
or \U$30881 ( \31224 , \31222 , \31223 );
not \U$30882 ( \31225 , \3154 );
not \U$30883 ( \31226 , \21529 );
not \U$30884 ( \31227 , \31226 );
or \U$30885 ( \31228 , \31225 , \31227 );
nand \U$30886 ( \31229 , \17908 , RI9872310_151);
nand \U$30887 ( \31230 , \31228 , \31229 );
nand \U$30888 ( \31231 , \31230 , \3163 );
nand \U$30889 ( \31232 , \31224 , \31231 );
not \U$30890 ( \31233 , \31232 );
or \U$30891 ( \31234 , \31221 , \31233 );
not \U$30892 ( \31235 , \31219 );
nand \U$30893 ( \31236 , \31235 , \31214 );
nand \U$30894 ( \31237 , \31234 , \31236 );
not \U$30895 ( \31238 , \31237 );
not \U$30896 ( \31239 , \8028 );
and \U$30897 ( \31240 , RI9872a18_166, \8597 );
not \U$30898 ( \31241 , RI9872a18_166);
and \U$30899 ( \31242 , \31241 , \18110 );
nor \U$30900 ( \31243 , \31240 , \31242 );
not \U$30901 ( \31244 , \31243 );
or \U$30902 ( \31245 , \31239 , \31244 );
nand \U$30903 ( \31246 , \30312 , \9071 );
nand \U$30904 ( \31247 , \31245 , \31246 );
not \U$30905 ( \31248 , \31247 );
xor \U$30906 ( \31249 , \31238 , \31248 );
and \U$30907 ( \31250 , RI9872b80_169, \9599 );
not \U$30908 ( \31251 , RI9872b80_169);
and \U$30909 ( \31252 , \31251 , \13358 );
or \U$30910 ( \31253 , \31250 , \31252 );
and \U$30911 ( \31254 , \9196 , \31253 );
and \U$30912 ( \31255 , \30520 , \9214 );
nor \U$30913 ( \31256 , \31254 , \31255 );
and \U$30914 ( \31257 , \31249 , \31256 );
and \U$30915 ( \31258 , \31238 , \31248 );
or \U$30916 ( \31259 , \31257 , \31258 );
not \U$30917 ( \31260 , \31259 );
not \U$30918 ( \31261 , \31260 );
xor \U$30919 ( \31262 , \30477 , \30482 );
xnor \U$30920 ( \31263 , \31262 , \30490 );
not \U$30921 ( \31264 , \31263 );
not \U$30922 ( \31265 , \31264 );
not \U$30923 ( \31266 , \18562 );
and \U$30924 ( \31267 , \7111 , \18862 );
not \U$30925 ( \31268 , \7111 );
and \U$30926 ( \31269 , \31268 , RI9872e50_175);
nor \U$30927 ( \31270 , \31267 , \31269 );
not \U$30928 ( \31271 , \31270 );
or \U$30929 ( \31272 , \31266 , \31271 );
nand \U$30930 ( \31273 , \30959 , \9273 );
nand \U$30931 ( \31274 , \31272 , \31273 );
not \U$30932 ( \31275 , \31274 );
not \U$30933 ( \31276 , \30904 );
not \U$30934 ( \31277 , \9227 );
not \U$30935 ( \31278 , \31277 );
and \U$30936 ( \31279 , \31276 , \31278 );
not \U$30937 ( \31280 , \9185 );
not \U$30938 ( \31281 , \21641 );
or \U$30939 ( \31282 , \31280 , \31281 );
or \U$30940 ( \31283 , \21641 , \9244 );
nand \U$30941 ( \31284 , \31282 , \31283 );
and \U$30942 ( \31285 , \9249 , \31284 );
nor \U$30943 ( \31286 , \31279 , \31285 );
not \U$30944 ( \31287 , \31286 );
not \U$30945 ( \31288 , \8818 );
xor \U$30946 ( \31289 , RI9872d60_173, \10411 );
not \U$30947 ( \31290 , \31289 );
or \U$30948 ( \31291 , \31288 , \31290 );
nand \U$30949 ( \31292 , \30915 , \8800 );
nand \U$30950 ( \31293 , \31291 , \31292 );
not \U$30951 ( \31294 , \31293 );
or \U$30952 ( \31295 , \31287 , \31294 );
or \U$30953 ( \31296 , \31293 , \31286 );
nand \U$30954 ( \31297 , \31295 , \31296 );
not \U$30955 ( \31298 , \31297 );
or \U$30956 ( \31299 , \31275 , \31298 );
not \U$30957 ( \31300 , \31286 );
nand \U$30958 ( \31301 , \31300 , \31293 );
nand \U$30959 ( \31302 , \31299 , \31301 );
not \U$30960 ( \31303 , \31302 );
or \U$30961 ( \31304 , \31265 , \31303 );
or \U$30962 ( \31305 , \31302 , \31264 );
nand \U$30963 ( \31306 , \31304 , \31305 );
not \U$30964 ( \31307 , \31306 );
or \U$30965 ( \31308 , \31261 , \31307 );
nand \U$30966 ( \31309 , \31302 , \31263 );
nand \U$30967 ( \31310 , \31308 , \31309 );
not \U$30968 ( \31311 , \31310 );
xor \U$30969 ( \31312 , \30195 , \30205 );
xor \U$30970 ( \31313 , \31312 , \30212 );
xor \U$30971 ( \31314 , \30669 , \31313 );
xnor \U$30972 ( \31315 , \31314 , \30685 );
not \U$30973 ( \31316 , \31315 );
or \U$30974 ( \31317 , \31311 , \31316 );
buf \U$30975 ( \31318 , \30685 );
nand \U$30976 ( \31319 , \31318 , \30669 );
not \U$30977 ( \31320 , \31319 );
not \U$30978 ( \31321 , \31318 );
not \U$30979 ( \31322 , \30669 );
nand \U$30980 ( \31323 , \31321 , \31322 );
not \U$30981 ( \31324 , \31323 );
or \U$30982 ( \31325 , \31320 , \31324 );
nand \U$30983 ( \31326 , \31325 , \31313 );
nand \U$30984 ( \31327 , \31317 , \31326 );
not \U$30985 ( \31328 , \31327 );
or \U$30986 ( \31329 , \31205 , \31328 );
not \U$30987 ( \31330 , \31098 );
not \U$30988 ( \31331 , \31203 );
nand \U$30989 ( \31332 , \31330 , \31331 );
nand \U$30990 ( \31333 , \31329 , \31332 );
and \U$30991 ( \31334 , \30650 , \30609 );
not \U$30992 ( \31335 , \30650 );
not \U$30993 ( \31336 , \30609 );
and \U$30994 ( \31337 , \31335 , \31336 );
nor \U$30995 ( \31338 , \31334 , \31337 );
xor \U$30996 ( \31339 , \30215 , \30217 );
xor \U$30997 ( \31340 , \31339 , \30220 );
xor \U$30998 ( \31341 , \31338 , \31340 );
not \U$30999 ( \31342 , \30691 );
not \U$31000 ( \31343 , \31342 );
not \U$31001 ( \31344 , \30718 );
or \U$31002 ( \31345 , \31343 , \31344 );
or \U$31003 ( \31346 , \30718 , \31342 );
nand \U$31004 ( \31347 , \31345 , \31346 );
and \U$31005 ( \31348 , \31341 , \31347 );
and \U$31006 ( \31349 , \31338 , \31340 );
or \U$31007 ( \31350 , \31348 , \31349 );
xor \U$31008 ( \31351 , \31333 , \31350 );
not \U$31009 ( \31352 , \31351 );
or \U$31010 ( \31353 , \31089 , \31352 );
nand \U$31011 ( \31354 , \31333 , \31350 );
nand \U$31012 ( \31355 , \31353 , \31354 );
xor \U$31013 ( \31356 , \30267 , \30554 );
xor \U$31014 ( \31357 , \31356 , \30572 );
or \U$31015 ( \31358 , \31355 , \31357 );
not \U$31016 ( \31359 , \31358 );
not \U$31017 ( \31360 , \30284 );
and \U$31018 ( \31361 , \30552 , \31360 );
not \U$31019 ( \31362 , \30552 );
and \U$31020 ( \31363 , \31362 , \30284 );
nor \U$31021 ( \31364 , \31361 , \31363 );
not \U$31022 ( \31365 , \31364 );
xor \U$31023 ( \31366 , \30542 , \31365 );
not \U$31024 ( \31367 , \31003 );
not \U$31025 ( \31368 , \30854 );
and \U$31026 ( \31369 , \31367 , \31368 );
and \U$31027 ( \31370 , \31003 , \30854 );
nor \U$31028 ( \31371 , \31369 , \31370 );
and \U$31029 ( \31372 , \31371 , \30857 );
not \U$31030 ( \31373 , \31371 );
and \U$31031 ( \31374 , \31373 , \31006 );
nor \U$31032 ( \31375 , \31372 , \31374 );
xor \U$31033 ( \31376 , \31366 , \31375 );
nand \U$31034 ( \31377 , \30537 , \30541 );
and \U$31035 ( \31378 , \31377 , \30422 );
not \U$31036 ( \31379 , \31377 );
not \U$31037 ( \31380 , \30422 );
and \U$31038 ( \31381 , \31379 , \31380 );
nor \U$31039 ( \31382 , \31378 , \31381 );
not \U$31040 ( \31383 , \19036 );
not \U$31041 ( \31384 , \16999 );
not \U$31042 ( \31385 , \5947 );
or \U$31043 ( \31386 , \31384 , \31385 );
or \U$31044 ( \31387 , \18937 , \16999 );
nand \U$31045 ( \31388 , \31386 , \31387 );
not \U$31046 ( \31389 , \31388 );
or \U$31047 ( \31390 , \31383 , \31389 );
nand \U$31048 ( \31391 , \30873 , \20147 );
nand \U$31049 ( \31392 , \31390 , \31391 );
not \U$31050 ( \31393 , \31392 );
and \U$31051 ( \31394 , \30970 , \22670 );
not \U$31052 ( \31395 , RI9873210_183);
not \U$31053 ( \31396 , \11672 );
or \U$31054 ( \31397 , \31395 , \31396 );
or \U$31055 ( \31398 , \3568 , RI9873210_183);
nand \U$31056 ( \31399 , \31397 , \31398 );
and \U$31057 ( \31400 , \31399 , \18957 );
nor \U$31058 ( \31401 , \31394 , \31400 );
nand \U$31059 ( \31402 , \31393 , \31401 );
not \U$31060 ( \31403 , \31402 );
xor \U$31061 ( \31404 , RI9873288_184, \3239 );
not \U$31062 ( \31405 , \31404 );
not \U$31063 ( \31406 , \18508 );
or \U$31064 ( \31407 , \31405 , \31406 );
nand \U$31065 ( \31408 , \31117 , \17528 );
nand \U$31066 ( \31409 , \31407 , \31408 );
not \U$31067 ( \31410 , \31409 );
or \U$31068 ( \31411 , \31403 , \31410 );
not \U$31069 ( \31412 , \31401 );
nand \U$31070 ( \31413 , \31412 , \31392 );
nand \U$31071 ( \31414 , \31411 , \31413 );
not \U$31072 ( \31415 , \31414 );
not \U$31073 ( \31416 , \30299 );
not \U$31074 ( \31417 , \31416 );
not \U$31075 ( \31418 , \30373 );
or \U$31076 ( \31419 , \31417 , \31418 );
or \U$31077 ( \31420 , \30373 , \31416 );
nand \U$31078 ( \31421 , \31419 , \31420 );
not \U$31079 ( \31422 , \30523 );
not \U$31080 ( \31423 , \30505 );
not \U$31081 ( \31424 , \31423 );
and \U$31082 ( \31425 , \31422 , \31424 );
and \U$31083 ( \31426 , \30523 , \31423 );
nor \U$31084 ( \31427 , \31425 , \31426 );
xnor \U$31085 ( \31428 , \31421 , \31427 );
not \U$31086 ( \31429 , \31428 );
or \U$31087 ( \31430 , \31415 , \31429 );
not \U$31088 ( \31431 , \31427 );
nand \U$31089 ( \31432 , \31431 , \31421 );
nand \U$31090 ( \31433 , \31430 , \31432 );
not \U$31091 ( \31434 , \31433 );
nand \U$31092 ( \31435 , \30494 , \30532 );
not \U$31093 ( \31436 , \31435 );
not \U$31094 ( \31437 , \30527 );
and \U$31095 ( \31438 , \31436 , \31437 );
and \U$31096 ( \31439 , \30527 , \31435 );
nor \U$31097 ( \31440 , \31438 , \31439 );
not \U$31098 ( \31441 , \31440 );
not \U$31099 ( \31442 , \30377 );
not \U$31100 ( \31443 , \30416 );
not \U$31101 ( \31444 , \31443 );
or \U$31102 ( \31445 , \31442 , \31444 );
not \U$31103 ( \31446 , \30377 );
nand \U$31104 ( \31447 , \31446 , \30416 );
nand \U$31105 ( \31448 , \31445 , \31447 );
not \U$31106 ( \31449 , \31448 );
or \U$31107 ( \31450 , \31441 , \31449 );
or \U$31108 ( \31451 , \31448 , \31440 );
nand \U$31109 ( \31452 , \31450 , \31451 );
not \U$31110 ( \31453 , \31452 );
or \U$31111 ( \31454 , \31434 , \31453 );
not \U$31112 ( \31455 , \31440 );
nand \U$31113 ( \31456 , \31455 , \31448 );
nand \U$31114 ( \31457 , \31454 , \31456 );
not \U$31115 ( \31458 , \31457 );
xor \U$31116 ( \31459 , \31382 , \31458 );
not \U$31117 ( \31460 , \17347 );
not \U$31118 ( \31461 , \30864 );
or \U$31119 ( \31462 , \31460 , \31461 );
xnor \U$31120 ( \31463 , RI98730a8_180, \5205 );
nand \U$31121 ( \31464 , \31463 , \13020 );
nand \U$31122 ( \31465 , \31462 , \31464 );
not \U$31123 ( \31466 , \31465 );
xor \U$31124 ( \31467 , \30364 , \30330 );
not \U$31125 ( \31468 , \31467 );
not \U$31126 ( \31469 , \18615 );
not \U$31127 ( \31470 , RI9873558_190);
not \U$31128 ( \31471 , \18572 );
or \U$31129 ( \31472 , \31470 , \31471 );
or \U$31130 ( \31473 , \18572 , RI9873558_190);
nand \U$31131 ( \31474 , \31472 , \31473 );
not \U$31132 ( \31475 , \31474 );
or \U$31133 ( \31476 , \31469 , \31475 );
nand \U$31134 ( \31477 , \30982 , RI9873648_192);
nand \U$31135 ( \31478 , \31476 , \31477 );
not \U$31136 ( \31479 , \31478 );
not \U$31137 ( \31480 , \31479 );
or \U$31138 ( \31481 , \31468 , \31480 );
not \U$31139 ( \31482 , \31467 );
nand \U$31140 ( \31483 , \31482 , \31478 );
nand \U$31141 ( \31484 , \31481 , \31483 );
not \U$31142 ( \31485 , \31484 );
or \U$31143 ( \31486 , \31466 , \31485 );
nand \U$31144 ( \31487 , \31478 , \31467 );
nand \U$31145 ( \31488 , \31486 , \31487 );
not \U$31146 ( \31489 , \5653 );
not \U$31147 ( \31490 , \30503 );
or \U$31148 ( \31491 , \31489 , \31490 );
and \U$31149 ( \31492 , \9750 , RI9872568_156);
not \U$31150 ( \31493 , \9750 );
and \U$31151 ( \31494 , \31493 , \5648 );
nor \U$31152 ( \31495 , \31492 , \31494 );
nand \U$31153 ( \31496 , \31495 , \5642 );
nand \U$31154 ( \31497 , \31491 , \31496 );
not \U$31155 ( \31498 , \31497 );
not \U$31156 ( \31499 , \4918 );
and \U$31157 ( \31500 , RI9872388_152, \13391 );
not \U$31158 ( \31501 , RI9872388_152);
and \U$31159 ( \31502 , \31501 , \13876 );
or \U$31160 ( \31503 , \31500 , \31502 );
not \U$31161 ( \31504 , \31503 );
or \U$31162 ( \31505 , \31499 , \31504 );
nand \U$31163 ( \31506 , \30457 , \4922 );
nand \U$31164 ( \31507 , \31505 , \31506 );
not \U$31165 ( \31508 , \5034 );
and \U$31166 ( \31509 , RI9872478_154, \17897 );
not \U$31167 ( \31510 , RI9872478_154);
not \U$31168 ( \31511 , \11370 );
and \U$31169 ( \31512 , \31510 , \31511 );
nor \U$31170 ( \31513 , \31509 , \31512 );
not \U$31171 ( \31514 , \31513 );
or \U$31172 ( \31515 , \31508 , \31514 );
nand \U$31173 ( \31516 , \30924 , \22459 );
nand \U$31174 ( \31517 , \31515 , \31516 );
and \U$31175 ( \31518 , \31507 , \31517 );
not \U$31176 ( \31519 , \31507 );
not \U$31177 ( \31520 , \31517 );
and \U$31178 ( \31521 , \31519 , \31520 );
nor \U$31179 ( \31522 , \31518 , \31521 );
not \U$31180 ( \31523 , \31522 );
or \U$31181 ( \31524 , \31498 , \31523 );
nand \U$31182 ( \31525 , \31507 , \31517 );
nand \U$31183 ( \31526 , \31524 , \31525 );
not \U$31184 ( \31527 , \6284 );
not \U$31185 ( \31528 , RI98728b0_163);
not \U$31186 ( \31529 , \8555 );
or \U$31187 ( \31530 , \31528 , \31529 );
or \U$31188 ( \31531 , \10369 , RI98728b0_163);
nand \U$31189 ( \31532 , \31530 , \31531 );
not \U$31190 ( \31533 , \31532 );
or \U$31191 ( \31534 , \31527 , \31533 );
nand \U$31192 ( \31535 , \31127 , \6610 );
nand \U$31193 ( \31536 , \31534 , \31535 );
not \U$31194 ( \31537 , \8752 );
not \U$31195 ( \31538 , \31106 );
or \U$31196 ( \31539 , \31537 , \31538 );
and \U$31197 ( \31540 , \8732 , \5775 );
not \U$31198 ( \31541 , \8732 );
and \U$31199 ( \31542 , \31541 , \6185 );
nor \U$31200 ( \31543 , \31540 , \31542 );
nand \U$31201 ( \31544 , \31543 , \24627 );
nand \U$31202 ( \31545 , \31539 , \31544 );
xor \U$31203 ( \31546 , \31536 , \31545 );
not \U$31204 ( \31547 , \7325 );
not \U$31205 ( \31548 , RI98729a0_165);
not \U$31206 ( \31549 , \11406 );
or \U$31207 ( \31550 , \31548 , \31549 );
or \U$31208 ( \31551 , \11406 , RI98729a0_165);
nand \U$31209 ( \31552 , \31550 , \31551 );
not \U$31210 ( \31553 , \31552 );
or \U$31211 ( \31554 , \31547 , \31553 );
nand \U$31212 ( \31555 , \30297 , \7338 );
nand \U$31213 ( \31556 , \31554 , \31555 );
and \U$31214 ( \31557 , \31546 , \31556 );
and \U$31215 ( \31558 , \31536 , \31545 );
or \U$31216 ( \31559 , \31557 , \31558 );
and \U$31217 ( \31560 , \31526 , \31559 );
or \U$31218 ( \31561 , \31488 , \31560 );
or \U$31219 ( \31562 , \31559 , \31526 );
nand \U$31220 ( \31563 , \31561 , \31562 );
not \U$31221 ( \31564 , \31563 );
not \U$31222 ( \31565 , \31564 );
not \U$31223 ( \31566 , \30868 );
not \U$31224 ( \31567 , \30892 );
not \U$31225 ( \31568 , \31567 );
or \U$31226 ( \31569 , \31566 , \31568 );
not \U$31227 ( \31570 , \30868 );
nand \U$31228 ( \31571 , \31570 , \30892 );
nand \U$31229 ( \31572 , \31569 , \31571 );
buf \U$31230 ( \31573 , \30931 );
and \U$31231 ( \31574 , \31573 , \30907 );
not \U$31232 ( \31575 , \31573 );
not \U$31233 ( \31576 , \30907 );
and \U$31234 ( \31577 , \31575 , \31576 );
nor \U$31235 ( \31578 , \31574 , \31577 );
buf \U$31236 ( \31579 , \31578 );
nor \U$31237 ( \31580 , \31572 , \31579 );
not \U$31238 ( \31581 , \9937 );
not \U$31239 ( \31582 , \31146 );
or \U$31240 ( \31583 , \31581 , \31582 );
and \U$31241 ( \31584 , RI9873030_179, \4989 );
not \U$31242 ( \31585 , RI9873030_179);
and \U$31243 ( \31586 , \31585 , \23391 );
nor \U$31244 ( \31587 , \31584 , \31586 );
nand \U$31245 ( \31588 , \31587 , \9952 );
nand \U$31246 ( \31589 , \31583 , \31588 );
not \U$31247 ( \31590 , \31589 );
not \U$31248 ( \31591 , \4084 );
not \U$31249 ( \31592 , \31173 );
or \U$31250 ( \31593 , \31591 , \31592 );
not \U$31251 ( \31594 , \4088 );
not \U$31252 ( \31595 , \13281 );
or \U$31253 ( \31596 , \31594 , \31595 );
nand \U$31254 ( \31597 , \17090 , RI98725e0_157);
nand \U$31255 ( \31598 , \31596 , \31597 );
nand \U$31256 ( \31599 , \31598 , \4101 );
nand \U$31257 ( \31600 , \31593 , \31599 );
not \U$31258 ( \31601 , \31600 );
not \U$31259 ( \31602 , \2087 );
not \U$31260 ( \31603 , \30354 );
or \U$31261 ( \31604 , \31602 , \31603 );
and \U$31262 ( \31605 , RI9871aa0_133, \19519 );
not \U$31263 ( \31606 , RI9871aa0_133);
and \U$31264 ( \31607 , \31606 , \24867 );
nor \U$31265 ( \31608 , \31605 , \31607 );
nand \U$31266 ( \31609 , \31608 , \2071 );
nand \U$31267 ( \31610 , \31604 , \31609 );
not \U$31268 ( \31611 , \2085 );
not \U$31269 ( \31612 , \31608 );
or \U$31270 ( \31613 , \31611 , \31612 );
and \U$31271 ( \31614 , \2076 , \28657 );
not \U$31272 ( \31615 , \2076 );
and \U$31273 ( \31616 , \31615 , \17702 );
nor \U$31274 ( \31617 , \31614 , \31616 );
nand \U$31275 ( \31618 , \31617 , \2070 );
nand \U$31276 ( \31619 , \31613 , \31618 );
not \U$31277 ( \31620 , \31619 );
nand \U$31278 ( \31621 , \21779 , \1134 );
not \U$31279 ( \31622 , \31621 );
not \U$31280 ( \31623 , \796 );
not \U$31281 ( \31624 , \31212 );
or \U$31282 ( \31625 , \31623 , \31624 );
and \U$31283 ( \31626 , RI98719b0_131, \23952 );
not \U$31284 ( \31627 , RI98719b0_131);
and \U$31285 ( \31628 , \31627 , \21773 );
nor \U$31286 ( \31629 , \31626 , \31628 );
nand \U$31287 ( \31630 , \31629 , \791 );
nand \U$31288 ( \31631 , \31625 , \31630 );
not \U$31289 ( \31632 , \31631 );
or \U$31290 ( \31633 , \31622 , \31632 );
or \U$31291 ( \31634 , \31631 , \31621 );
nand \U$31292 ( \31635 , \31633 , \31634 );
not \U$31293 ( \31636 , \31635 );
or \U$31294 ( \31637 , \31620 , \31636 );
not \U$31295 ( \31638 , \31621 );
nand \U$31296 ( \31639 , \31638 , \31631 );
nand \U$31297 ( \31640 , \31637 , \31639 );
and \U$31298 ( \31641 , \31610 , \31640 );
not \U$31299 ( \31642 , \31610 );
not \U$31300 ( \31643 , \31640 );
and \U$31301 ( \31644 , \31642 , \31643 );
nor \U$31302 ( \31645 , \31641 , \31644 );
not \U$31303 ( \31646 , \31645 );
or \U$31304 ( \31647 , \31601 , \31646 );
nand \U$31305 ( \31648 , \31640 , \31610 );
nand \U$31306 ( \31649 , \31647 , \31648 );
not \U$31307 ( \31650 , \31649 );
not \U$31308 ( \31651 , \17252 );
not \U$31309 ( \31652 , \2110 );
and \U$31310 ( \31653 , RI98733f0_187, \31652 );
not \U$31311 ( \31654 , RI98733f0_187);
and \U$31312 ( \31655 , \31654 , \2110 );
or \U$31313 ( \31656 , \31653 , \31655 );
not \U$31314 ( \31657 , \31656 );
or \U$31315 ( \31658 , \31651 , \31657 );
nand \U$31316 ( \31659 , \30884 , \19282 );
nand \U$31317 ( \31660 , \31658 , \31659 );
xnor \U$31318 ( \31661 , \31650 , \31660 );
not \U$31319 ( \31662 , \31661 );
or \U$31320 ( \31663 , \31590 , \31662 );
not \U$31321 ( \31664 , \31650 );
nand \U$31322 ( \31665 , \31664 , \31660 );
nand \U$31323 ( \31666 , \31663 , \31665 );
not \U$31324 ( \31667 , \31666 );
or \U$31325 ( \31668 , \31580 , \31667 );
nand \U$31326 ( \31669 , \31572 , \31579 );
nand \U$31327 ( \31670 , \31668 , \31669 );
buf \U$31328 ( \31671 , \31670 );
not \U$31329 ( \31672 , \31671 );
or \U$31330 ( \31673 , \31565 , \31672 );
xor \U$31331 ( \31674 , \30986 , \30951 );
xnor \U$31332 ( \31675 , \31674 , \30989 );
not \U$31333 ( \31676 , \31675 );
nand \U$31334 ( \31677 , \31673 , \31676 );
or \U$31335 ( \31678 , \31671 , \31564 );
nand \U$31336 ( \31679 , \31677 , \31678 );
and \U$31337 ( \31680 , \31459 , \31679 );
and \U$31338 ( \31681 , \31382 , \31458 );
nor \U$31339 ( \31682 , \31680 , \31681 );
and \U$31340 ( \31683 , \31376 , \31682 );
and \U$31341 ( \31684 , \31366 , \31375 );
or \U$31342 ( \31685 , \31683 , \31684 );
not \U$31343 ( \31686 , \31685 );
or \U$31344 ( \31687 , \31359 , \31686 );
nand \U$31345 ( \31688 , \31355 , \31357 );
nand \U$31346 ( \31689 , \31687 , \31688 );
not \U$31347 ( \31690 , \31689 );
xor \U$31348 ( \31691 , \30118 , \30575 );
xor \U$31349 ( \31692 , \31691 , \30772 );
not \U$31350 ( \31693 , \31692 );
not \U$31351 ( \31694 , \31693 );
xor \U$31352 ( \31695 , \31033 , \31036 );
xnor \U$31353 ( \31696 , \31695 , \31026 );
not \U$31354 ( \31697 , \31696 );
or \U$31355 ( \31698 , \31694 , \31697 );
or \U$31356 ( \31699 , \31696 , \31693 );
nand \U$31357 ( \31700 , \31698 , \31699 );
not \U$31358 ( \31701 , \31700 );
or \U$31359 ( \31702 , \31690 , \31701 );
nand \U$31360 ( \31703 , \31696 , \31692 );
nand \U$31361 ( \31704 , \31702 , \31703 );
xor \U$31362 ( \31705 , \30840 , \31045 );
xnor \U$31363 ( \31706 , \31705 , \30836 );
nor \U$31364 ( \31707 , \31704 , \31706 );
xor \U$31365 ( \31708 , \31692 , \31689 );
xor \U$31366 ( \31709 , \31708 , \31696 );
not \U$31367 ( \31710 , \31357 );
not \U$31368 ( \31711 , \31355 );
or \U$31369 ( \31712 , \31710 , \31711 );
or \U$31370 ( \31713 , \31355 , \31357 );
nand \U$31371 ( \31714 , \31712 , \31713 );
xor \U$31372 ( \31715 , \31685 , \31714 );
not \U$31373 ( \31716 , \31715 );
not \U$31374 ( \31717 , \31716 );
and \U$31375 ( \31718 , \31019 , \30851 );
not \U$31376 ( \31719 , \31019 );
not \U$31377 ( \31720 , \30851 );
and \U$31378 ( \31721 , \31719 , \31720 );
nor \U$31379 ( \31722 , \31718 , \31721 );
not \U$31380 ( \31723 , \31722 );
xor \U$31381 ( \31724 , \31338 , \31340 );
xor \U$31382 ( \31725 , \31724 , \31347 );
not \U$31383 ( \31726 , \31725 );
xor \U$31384 ( \31727 , \31310 , \31315 );
not \U$31385 ( \31728 , \31727 );
xor \U$31386 ( \31729 , \31148 , \31193 );
not \U$31387 ( \31730 , \31108 );
not \U$31388 ( \31731 , \31134 );
not \U$31389 ( \31732 , \31731 );
or \U$31390 ( \31733 , \31730 , \31732 );
not \U$31391 ( \31734 , \31108 );
nand \U$31392 ( \31735 , \31734 , \31134 );
nand \U$31393 ( \31736 , \31733 , \31735 );
or \U$31394 ( \31737 , \31729 , \31736 );
xor \U$31395 ( \31738 , \30961 , \30984 );
xnor \U$31396 ( \31739 , \31738 , \30972 );
not \U$31397 ( \31740 , \31739 );
nand \U$31398 ( \31741 , \31737 , \31740 );
nand \U$31399 ( \31742 , \31736 , \31729 );
nand \U$31400 ( \31743 , \31741 , \31742 );
not \U$31401 ( \31744 , \31743 );
not \U$31402 ( \31745 , \30940 );
not \U$31403 ( \31746 , \30897 );
not \U$31404 ( \31747 , \31746 );
and \U$31405 ( \31748 , \31745 , \31747 );
and \U$31406 ( \31749 , \30940 , \31746 );
nor \U$31407 ( \31750 , \31748 , \31749 );
nand \U$31408 ( \31751 , \31744 , \31750 );
not \U$31409 ( \31752 , \31751 );
or \U$31410 ( \31753 , \31728 , \31752 );
not \U$31411 ( \31754 , \31750 );
nand \U$31412 ( \31755 , \31754 , \31743 );
nand \U$31413 ( \31756 , \31753 , \31755 );
not \U$31414 ( \31757 , \31756 );
xor \U$31415 ( \31758 , \30998 , \30945 );
not \U$31416 ( \31759 , \31758 );
nand \U$31417 ( \31760 , \31757 , \31759 );
not \U$31418 ( \31761 , \31760 );
or \U$31419 ( \31762 , \31726 , \31761 );
not \U$31420 ( \31763 , \31759 );
nand \U$31421 ( \31764 , \31763 , \31756 );
nand \U$31422 ( \31765 , \31762 , \31764 );
not \U$31423 ( \31766 , \31087 );
not \U$31424 ( \31767 , \31351 );
or \U$31425 ( \31768 , \31766 , \31767 );
or \U$31426 ( \31769 , \31351 , \31087 );
nand \U$31427 ( \31770 , \31768 , \31769 );
xor \U$31428 ( \31771 , \31765 , \31770 );
and \U$31429 ( \31772 , \31200 , \31198 );
not \U$31430 ( \31773 , \31200 );
not \U$31431 ( \31774 , \31148 );
not \U$31432 ( \31775 , \31193 );
or \U$31433 ( \31776 , \31774 , \31775 );
nand \U$31434 ( \31777 , \31776 , \31196 );
and \U$31435 ( \31778 , \31773 , \31777 );
or \U$31436 ( \31779 , \31772 , \31778 );
xor \U$31437 ( \31780 , \31779 , \31139 );
not \U$31438 ( \31781 , \5653 );
not \U$31439 ( \31782 , \31495 );
or \U$31440 ( \31783 , \31781 , \31782 );
not \U$31441 ( \31784 , RI9872568_156);
not \U$31442 ( \31785 , \12460 );
or \U$31443 ( \31786 , \31784 , \31785 );
or \U$31444 ( \31787 , \12460 , RI9872568_156);
nand \U$31445 ( \31788 , \31786 , \31787 );
nand \U$31446 ( \31789 , \31788 , \5642 );
nand \U$31447 ( \31790 , \31783 , \31789 );
not \U$31448 ( \31791 , \8801 );
not \U$31449 ( \31792 , \31289 );
or \U$31450 ( \31793 , \31791 , \31792 );
not \U$31451 ( \31794 , RI9872d60_173);
not \U$31452 ( \31795 , \10582 );
or \U$31453 ( \31796 , \31794 , \31795 );
or \U$31454 ( \31797 , \20583 , RI9872d60_173);
nand \U$31455 ( \31798 , \31796 , \31797 );
nand \U$31456 ( \31799 , \31798 , \8819 );
nand \U$31457 ( \31800 , \31793 , \31799 );
xor \U$31458 ( \31801 , \31790 , \31800 );
not \U$31459 ( \31802 , \10331 );
not \U$31460 ( \31803 , \31270 );
or \U$31461 ( \31804 , \31802 , \31803 );
and \U$31462 ( \31805 , \9694 , \8903 );
not \U$31463 ( \31806 , \9694 );
and \U$31464 ( \31807 , \31806 , \6296 );
nor \U$31465 ( \31808 , \31805 , \31807 );
nand \U$31466 ( \31809 , \31808 , \18562 );
nand \U$31467 ( \31810 , \31804 , \31809 );
and \U$31468 ( \31811 , \31801 , \31810 );
and \U$31469 ( \31812 , \31790 , \31800 );
or \U$31470 ( \31813 , \31811 , \31812 );
not \U$31471 ( \31814 , \31813 );
xor \U$31472 ( \31815 , \31183 , \31164 );
not \U$31473 ( \31816 , \31815 );
nand \U$31474 ( \31817 , \31284 , \9227 );
not \U$31475 ( \31818 , \9244 );
not \U$31476 ( \31819 , \8916 );
or \U$31477 ( \31820 , \31818 , \31819 );
or \U$31478 ( \31821 , \9898 , \9185 );
nand \U$31479 ( \31822 , \31820 , \31821 );
nand \U$31480 ( \31823 , \31822 , \9249 );
nand \U$31481 ( \31824 , \31817 , \31823 );
xor \U$31482 ( \31825 , \31232 , \31220 );
xor \U$31483 ( \31826 , \31824 , \31825 );
not \U$31484 ( \31827 , \9214 );
not \U$31485 ( \31828 , \31253 );
or \U$31486 ( \31829 , \31827 , \31828 );
and \U$31487 ( \31830 , RI9872b80_169, \8878 );
not \U$31488 ( \31831 , RI9872b80_169);
and \U$31489 ( \31832 , \31831 , \29463 );
or \U$31490 ( \31833 , \31830 , \31832 );
nand \U$31491 ( \31834 , \31833 , \9196 );
nand \U$31492 ( \31835 , \31829 , \31834 );
nand \U$31493 ( \31836 , \31826 , \31835 );
not \U$31494 ( \31837 , \31817 );
not \U$31495 ( \31838 , \31823 );
or \U$31496 ( \31839 , \31837 , \31838 );
nand \U$31497 ( \31840 , \31839 , \31825 );
and \U$31498 ( \31841 , \31836 , \31840 );
not \U$31499 ( \31842 , \31841 );
or \U$31500 ( \31843 , \31816 , \31842 );
not \U$31501 ( \31844 , \31840 );
not \U$31502 ( \31845 , \31836 );
or \U$31503 ( \31846 , \31844 , \31845 );
not \U$31504 ( \31847 , \31815 );
nand \U$31505 ( \31848 , \31846 , \31847 );
nand \U$31506 ( \31849 , \31843 , \31848 );
not \U$31507 ( \31850 , \31849 );
or \U$31508 ( \31851 , \31814 , \31850 );
not \U$31509 ( \31852 , \31840 );
not \U$31510 ( \31853 , \31836 );
or \U$31511 ( \31854 , \31852 , \31853 );
nand \U$31512 ( \31855 , \31854 , \31815 );
nand \U$31513 ( \31856 , \31851 , \31855 );
or \U$31514 ( \31857 , RI9871a28_132, RI9871aa0_133);
nand \U$31515 ( \31858 , \31857 , \18704 );
and \U$31516 ( \31859 , \31858 , \1687 );
not \U$31517 ( \31860 , \796 );
not \U$31518 ( \31861 , \31629 );
or \U$31519 ( \31862 , \31860 , \31861 );
not \U$31520 ( \31863 , \1078 );
not \U$31521 ( \31864 , \18704 );
or \U$31522 ( \31865 , \31863 , \31864 );
or \U$31523 ( \31866 , \27523 , \1078 );
nand \U$31524 ( \31867 , \31865 , \31866 );
nand \U$31525 ( \31868 , \31867 , \791 );
nand \U$31526 ( \31869 , \31862 , \31868 );
and \U$31527 ( \31870 , \31859 , \31869 );
not \U$31528 ( \31871 , \3163 );
not \U$31529 ( \31872 , RI9872310_151);
not \U$31530 ( \31873 , \30350 );
or \U$31531 ( \31874 , \31872 , \31873 );
not \U$31532 ( \31875 , \17725 );
or \U$31533 ( \31876 , \31875 , RI9872310_151);
nand \U$31534 ( \31877 , \31874 , \31876 );
not \U$31535 ( \31878 , \31877 );
or \U$31536 ( \31879 , \31871 , \31878 );
nand \U$31537 ( \31880 , \31230 , \3169 );
nand \U$31538 ( \31881 , \31879 , \31880 );
xor \U$31539 ( \31882 , \31870 , \31881 );
not \U$31540 ( \31883 , \3467 );
not \U$31541 ( \31884 , \3593 );
not \U$31542 ( \31885 , \17014 );
or \U$31543 ( \31886 , \31884 , \31885 );
or \U$31544 ( \31887 , \17014 , \3593 );
nand \U$31545 ( \31888 , \31886 , \31887 );
not \U$31546 ( \31889 , \31888 );
or \U$31547 ( \31890 , \31883 , \31889 );
not \U$31548 ( \31891 , RI98726d0_159);
not \U$31549 ( \31892 , \20449 );
or \U$31550 ( \31893 , \31891 , \31892 );
or \U$31551 ( \31894 , \20764 , RI98726d0_159);
nand \U$31552 ( \31895 , \31893 , \31894 );
nand \U$31553 ( \31896 , \31895 , \3464 );
nand \U$31554 ( \31897 , \31890 , \31896 );
and \U$31555 ( \31898 , \31882 , \31897 );
and \U$31556 ( \31899 , \31870 , \31881 );
or \U$31557 ( \31900 , \31898 , \31899 );
not \U$31558 ( \31901 , \9072 );
not \U$31559 ( \31902 , \31243 );
or \U$31560 ( \31903 , \31901 , \31902 );
not \U$31561 ( \31904 , \20414 );
xor \U$31562 ( \31905 , RI9872a18_166, \31904 );
nand \U$31563 ( \31906 , \31905 , \8027 );
nand \U$31564 ( \31907 , \31903 , \31906 );
xor \U$31565 ( \31908 , \31900 , \31907 );
not \U$31566 ( \31909 , \7338 );
not \U$31567 ( \31910 , \31552 );
or \U$31568 ( \31911 , \31909 , \31910 );
and \U$31569 ( \31912 , RI98729a0_165, \8575 );
not \U$31570 ( \31913 , RI98729a0_165);
and \U$31571 ( \31914 , \31913 , \8576 );
nor \U$31572 ( \31915 , \31912 , \31914 );
nand \U$31573 ( \31916 , \31915 , \7325 );
nand \U$31574 ( \31917 , \31911 , \31916 );
and \U$31575 ( \31918 , \31908 , \31917 );
and \U$31576 ( \31919 , \31900 , \31907 );
or \U$31577 ( \31920 , \31918 , \31919 );
not \U$31578 ( \31921 , \31920 );
not \U$31579 ( \31922 , RI9872478_154);
not \U$31580 ( \31923 , \13066 );
or \U$31581 ( \31924 , \31922 , \31923 );
or \U$31582 ( \31925 , \12597 , RI9872478_154);
nand \U$31583 ( \31926 , \31924 , \31925 );
not \U$31584 ( \31927 , \31926 );
not \U$31585 ( \31928 , \5034 );
or \U$31586 ( \31929 , \31927 , \31928 );
not \U$31587 ( \31930 , \31513 );
or \U$31588 ( \31931 , \31930 , \5795 );
nand \U$31589 ( \31932 , \31929 , \31931 );
not \U$31590 ( \31933 , \31932 );
not \U$31591 ( \31934 , \31162 );
nor \U$31592 ( \31935 , \31934 , \3591 );
and \U$31593 ( \31936 , \31888 , \3464 );
nor \U$31594 ( \31937 , \31935 , \31936 );
not \U$31595 ( \31938 , \31937 );
not \U$31596 ( \31939 , \4923 );
not \U$31597 ( \31940 , \31503 );
or \U$31598 ( \31941 , \31939 , \31940 );
and \U$31599 ( \31942 , RI9872388_152, \12783 );
not \U$31600 ( \31943 , RI9872388_152);
and \U$31601 ( \31944 , \31943 , \18151 );
nor \U$31602 ( \31945 , \31942 , \31944 );
nand \U$31603 ( \31946 , \31945 , \4918 );
nand \U$31604 ( \31947 , \31941 , \31946 );
not \U$31605 ( \31948 , \31947 );
or \U$31606 ( \31949 , \31938 , \31948 );
or \U$31607 ( \31950 , \31947 , \31937 );
nand \U$31608 ( \31951 , \31949 , \31950 );
not \U$31609 ( \31952 , \31951 );
or \U$31610 ( \31953 , \31933 , \31952 );
not \U$31611 ( \31954 , \31937 );
nand \U$31612 ( \31955 , \31954 , \31947 );
nand \U$31613 ( \31956 , \31953 , \31955 );
xor \U$31614 ( \31957 , \31497 , \31522 );
xor \U$31615 ( \31958 , \31956 , \31957 );
not \U$31616 ( \31959 , \31958 );
or \U$31617 ( \31960 , \31921 , \31959 );
nand \U$31618 ( \31961 , \31957 , \31956 );
nand \U$31619 ( \31962 , \31960 , \31961 );
nand \U$31620 ( \31963 , \31856 , \31962 );
not \U$31621 ( \31964 , \31963 );
not \U$31622 ( \31965 , \6285 );
not \U$31623 ( \31966 , \31532 );
or \U$31624 ( \31967 , \31965 , \31966 );
not \U$31625 ( \31968 , RI98728b0_163);
not \U$31626 ( \31969 , \13454 );
or \U$31627 ( \31970 , \31968 , \31969 );
or \U$31628 ( \31971 , \9924 , RI98728b0_163);
nand \U$31629 ( \31972 , \31970 , \31971 );
nand \U$31630 ( \31973 , \31972 , \6282 );
nand \U$31631 ( \31974 , \31967 , \31973 );
not \U$31632 ( \31975 , \11198 );
not \U$31633 ( \31976 , \31543 );
or \U$31634 ( \31977 , \31975 , \31976 );
and \U$31635 ( \31978 , \5760 , \8732 );
not \U$31636 ( \31979 , \5760 );
and \U$31637 ( \31980 , \31979 , RI9872f40_177);
nor \U$31638 ( \31981 , \31978 , \31980 );
nand \U$31639 ( \31982 , \8742 , \31981 );
nand \U$31640 ( \31983 , \31977 , \31982 );
xor \U$31641 ( \31984 , \31974 , \31983 );
not \U$31642 ( \31985 , \31984 );
not \U$31643 ( \31986 , \20147 );
not \U$31644 ( \31987 , \31388 );
or \U$31645 ( \31988 , \31986 , \31987 );
and \U$31646 ( \31989 , RI98734e0_189, \1485 );
not \U$31647 ( \31990 , RI98734e0_189);
and \U$31648 ( \31991 , \31990 , \1486 );
or \U$31649 ( \31992 , \31989 , \31991 );
nand \U$31650 ( \31993 , \31992 , \19243 );
nand \U$31651 ( \31994 , \31988 , \31993 );
not \U$31652 ( \31995 , \31994 );
or \U$31653 ( \31996 , \31985 , \31995 );
nand \U$31654 ( \31997 , \31974 , \31983 );
nand \U$31655 ( \31998 , \31996 , \31997 );
not \U$31656 ( \31999 , \31998 );
not \U$31657 ( \32000 , \17347 );
not \U$31658 ( \32001 , \31463 );
or \U$31659 ( \32002 , \32000 , \32001 );
not \U$31660 ( \32003 , RI98730a8_180);
not \U$31661 ( \32004 , \4470 );
or \U$31662 ( \32005 , \32003 , \32004 );
or \U$31663 ( \32006 , \4470 , RI98730a8_180);
nand \U$31664 ( \32007 , \32005 , \32006 );
nand \U$31665 ( \32008 , \32007 , \13020 );
nand \U$31666 ( \32009 , \32002 , \32008 );
not \U$31667 ( \32010 , \9937 );
not \U$31668 ( \32011 , \31587 );
or \U$31669 ( \32012 , \32010 , \32011 );
and \U$31670 ( \32013 , \5736 , \9946 );
not \U$31671 ( \32014 , \5736 );
and \U$31672 ( \32015 , \32014 , RI9873030_179);
nor \U$31673 ( \32016 , \32013 , \32015 );
nand \U$31674 ( \32017 , \32016 , \12507 );
nand \U$31675 ( \32018 , \32012 , \32017 );
nor \U$31676 ( \32019 , \32009 , \32018 );
and \U$31677 ( \32020 , \17539 , \8785 );
not \U$31678 ( \32021 , \17539 );
and \U$31679 ( \32022 , \32021 , \2947 );
nor \U$31680 ( \32023 , \32020 , \32022 );
not \U$31681 ( \32024 , \32023 );
not \U$31682 ( \32025 , \30886 );
and \U$31683 ( \32026 , \32024 , \32025 );
and \U$31684 ( \32027 , \31656 , \19282 );
nor \U$31685 ( \32028 , \32026 , \32027 );
or \U$31686 ( \32029 , \32019 , \32028 );
nand \U$31687 ( \32030 , \32009 , \32018 );
nand \U$31688 ( \32031 , \32029 , \32030 );
not \U$31689 ( \32032 , \32031 );
not \U$31690 ( \32033 , RI9873648_192);
not \U$31691 ( \32034 , \31474 );
or \U$31692 ( \32035 , \32033 , \32034 );
not \U$31693 ( \32036 , \18239 );
not \U$31694 ( \32037 , \11113 );
or \U$31695 ( \32038 , \32036 , \32037 );
or \U$31696 ( \32039 , \9262 , \18239 );
nand \U$31697 ( \32040 , \32038 , \32039 );
nand \U$31698 ( \32041 , \32040 , \18615 );
nand \U$31699 ( \32042 , \32035 , \32041 );
not \U$31700 ( \32043 , \17528 );
not \U$31701 ( \32044 , \31404 );
or \U$31702 ( \32045 , \32043 , \32044 );
not \U$31703 ( \32046 , \22727 );
not \U$31704 ( \32047 , \3536 );
or \U$31705 ( \32048 , \32046 , \32047 );
or \U$31706 ( \32049 , \6718 , \22715 );
nand \U$31707 ( \32050 , \32048 , \32049 );
nand \U$31708 ( \32051 , \32050 , \19641 );
nand \U$31709 ( \32052 , \32045 , \32051 );
or \U$31710 ( \32053 , \32042 , \32052 );
not \U$31711 ( \32054 , \18957 );
and \U$31712 ( \32055 , \18012 , \5595 );
not \U$31713 ( \32056 , \18012 );
and \U$31714 ( \32057 , \32056 , \5594 );
nor \U$31715 ( \32058 , \32055 , \32057 );
not \U$31716 ( \32059 , \32058 );
or \U$31717 ( \32060 , \32054 , \32059 );
nand \U$31718 ( \32061 , \31399 , \22670 );
nand \U$31719 ( \32062 , \32060 , \32061 );
nand \U$31720 ( \32063 , \32053 , \32062 );
nand \U$31721 ( \32064 , \32042 , \32052 );
nand \U$31722 ( \32065 , \32063 , \32064 );
not \U$31723 ( \32066 , \32065 );
not \U$31724 ( \32067 , \32066 );
or \U$31725 ( \32068 , \32032 , \32067 );
or \U$31726 ( \32069 , \32066 , \32031 );
nand \U$31727 ( \32070 , \32068 , \32069 );
not \U$31728 ( \32071 , \32070 );
or \U$31729 ( \32072 , \31999 , \32071 );
not \U$31730 ( \32073 , \32066 );
nand \U$31731 ( \32074 , \32073 , \32031 );
nand \U$31732 ( \32075 , \32072 , \32074 );
not \U$31733 ( \32076 , \32075 );
not \U$31734 ( \32077 , \32076 );
or \U$31735 ( \32078 , \31964 , \32077 );
or \U$31736 ( \32079 , \31856 , \31962 );
nand \U$31737 ( \32080 , \32078 , \32079 );
xor \U$31738 ( \32081 , \31780 , \32080 );
xor \U$31739 ( \32082 , \31440 , \31448 );
xor \U$31740 ( \32083 , \32082 , \31433 );
and \U$31741 ( \32084 , \32081 , \32083 );
and \U$31742 ( \32085 , \31780 , \32080 );
or \U$31743 ( \32086 , \32084 , \32085 );
xor \U$31744 ( \32087 , \31331 , \31330 );
xnor \U$31745 ( \32088 , \32087 , \31327 );
nand \U$31746 ( \32089 , \32086 , \32088 );
not \U$31747 ( \32090 , \32089 );
not \U$31748 ( \32091 , \31459 );
and \U$31749 ( \32092 , \31679 , \32091 );
not \U$31750 ( \32093 , \31679 );
and \U$31751 ( \32094 , \32093 , \31459 );
nor \U$31752 ( \32095 , \32092 , \32094 );
not \U$31753 ( \32096 , \32095 );
or \U$31754 ( \32097 , \32090 , \32096 );
or \U$31755 ( \32098 , \32086 , \32088 );
nand \U$31756 ( \32099 , \32097 , \32098 );
nand \U$31757 ( \32100 , \31771 , \32099 );
not \U$31758 ( \32101 , \32100 );
and \U$31759 ( \32102 , \31765 , \31770 );
nor \U$31760 ( \32103 , \32101 , \32102 );
not \U$31761 ( \32104 , \32103 );
or \U$31762 ( \32105 , \31723 , \32104 );
not \U$31763 ( \32106 , \32102 );
not \U$31764 ( \32107 , \32106 );
not \U$31765 ( \32108 , \32100 );
or \U$31766 ( \32109 , \32107 , \32108 );
not \U$31767 ( \32110 , \31722 );
nand \U$31768 ( \32111 , \32109 , \32110 );
nand \U$31769 ( \32112 , \32105 , \32111 );
not \U$31770 ( \32113 , \32112 );
or \U$31771 ( \32114 , \31717 , \32113 );
not \U$31772 ( \32115 , \32106 );
not \U$31773 ( \32116 , \32100 );
or \U$31774 ( \32117 , \32115 , \32116 );
nand \U$31775 ( \32118 , \32117 , \31722 );
nand \U$31776 ( \32119 , \32114 , \32118 );
nor \U$31777 ( \32120 , \31709 , \32119 );
nor \U$31778 ( \32121 , \31707 , \32120 );
nand \U$31779 ( \32122 , \32098 , \32089 );
not \U$31780 ( \32123 , \32122 );
buf \U$31781 ( \32124 , \32095 );
not \U$31782 ( \32125 , \32124 );
and \U$31783 ( \32126 , \32123 , \32125 );
and \U$31784 ( \32127 , \32122 , \32124 );
nor \U$31785 ( \32128 , \32126 , \32127 );
not \U$31786 ( \32129 , \31750 );
xor \U$31787 ( \32130 , \31743 , \32129 );
not \U$31788 ( \32131 , \31727 );
xnor \U$31789 ( \32132 , \32130 , \32131 );
not \U$31790 ( \32133 , \32132 );
xnor \U$31791 ( \32134 , \31962 , \31856 );
and \U$31792 ( \32135 , \32134 , \32076 );
not \U$31793 ( \32136 , \32134 );
and \U$31794 ( \32137 , \32136 , \32075 );
nor \U$31795 ( \32138 , \32135 , \32137 );
not \U$31796 ( \32139 , \32138 );
and \U$31797 ( \32140 , \31826 , \31835 );
not \U$31798 ( \32141 , \31826 );
not \U$31799 ( \32142 , \31835 );
and \U$31800 ( \32143 , \32141 , \32142 );
nor \U$31801 ( \32144 , \32140 , \32143 );
xor \U$31802 ( \32145 , \31900 , \31907 );
xor \U$31803 ( \32146 , \32145 , \31917 );
xor \U$31804 ( \32147 , \32144 , \32146 );
xor \U$31805 ( \32148 , \31790 , \31800 );
xor \U$31806 ( \32149 , \32148 , \31810 );
and \U$31807 ( \32150 , \32147 , \32149 );
and \U$31808 ( \32151 , \32144 , \32146 );
or \U$31809 ( \32152 , \32150 , \32151 );
not \U$31810 ( \32153 , \32152 );
xor \U$31811 ( \32154 , \31600 , \31645 );
not \U$31812 ( \32155 , \31598 );
or \U$31813 ( \32156 , \32155 , \6048 );
not \U$31814 ( \32157 , RI98725e0_157);
not \U$31815 ( \32158 , \17783 );
or \U$31816 ( \32159 , \32157 , \32158 );
or \U$31817 ( \32160 , \17783 , RI98725e0_157);
nand \U$31818 ( \32161 , \32159 , \32160 );
not \U$31819 ( \32162 , \32161 );
or \U$31820 ( \32163 , \32162 , \4100 );
nand \U$31821 ( \32164 , \32156 , \32163 );
not \U$31822 ( \32165 , \32164 );
not \U$31823 ( \32166 , \31635 );
xor \U$31824 ( \32167 , \31619 , \32166 );
not \U$31825 ( \32168 , \32167 );
not \U$31826 ( \32169 , \4918 );
not \U$31827 ( \32170 , \4902 );
not \U$31828 ( \32171 , \14193 );
or \U$31829 ( \32172 , \32170 , \32171 );
not \U$31830 ( \32173 , \12773 );
or \U$31831 ( \32174 , \32173 , \4902 );
nand \U$31832 ( \32175 , \32172 , \32174 );
not \U$31833 ( \32176 , \32175 );
or \U$31834 ( \32177 , \32169 , \32176 );
not \U$31835 ( \32178 , \4922 );
not \U$31836 ( \32179 , \32178 );
nand \U$31837 ( \32180 , \32179 , \31945 );
nand \U$31838 ( \32181 , \32177 , \32180 );
not \U$31839 ( \32182 , \32181 );
or \U$31840 ( \32183 , \32168 , \32182 );
or \U$31841 ( \32184 , \32181 , \32167 );
nand \U$31842 ( \32185 , \32183 , \32184 );
not \U$31843 ( \32186 , \32185 );
or \U$31844 ( \32187 , \32165 , \32186 );
not \U$31845 ( \32188 , \32167 );
nand \U$31846 ( \32189 , \32188 , \32181 );
nand \U$31847 ( \32190 , \32187 , \32189 );
xor \U$31848 ( \32191 , \32154 , \32190 );
xor \U$31849 ( \32192 , \31932 , \31951 );
and \U$31850 ( \32193 , \32191 , \32192 );
and \U$31851 ( \32194 , \32154 , \32190 );
nor \U$31852 ( \32195 , \32193 , \32194 );
not \U$31853 ( \32196 , \32195 );
not \U$31854 ( \32197 , \9196 );
xor \U$31855 ( \32198 , RI9872b80_169, \8596 );
not \U$31856 ( \32199 , \32198 );
or \U$31857 ( \32200 , \32197 , \32199 );
nand \U$31858 ( \32201 , \31833 , \9214 );
nand \U$31859 ( \32202 , \32200 , \32201 );
not \U$31860 ( \32203 , \32202 );
not \U$31861 ( \32204 , \31895 );
not \U$31862 ( \32205 , \3467 );
or \U$31863 ( \32206 , \32204 , \32205 );
not \U$31864 ( \32207 , \4063 );
not \U$31865 ( \32208 , \17741 );
not \U$31866 ( \32209 , \32208 );
or \U$31867 ( \32210 , \32207 , \32209 );
nand \U$31868 ( \32211 , \17911 , RI98726d0_159);
nand \U$31869 ( \32212 , \32210 , \32211 );
nand \U$31870 ( \32213 , \32212 , \3464 );
nand \U$31871 ( \32214 , \32206 , \32213 );
xor \U$31872 ( \32215 , \31859 , \31869 );
not \U$31873 ( \32216 , \2085 );
not \U$31874 ( \32217 , \31617 );
or \U$31875 ( \32218 , \32216 , \32217 );
not \U$31876 ( \32219 , \2076 );
not \U$31877 ( \32220 , \17862 );
or \U$31878 ( \32221 , \32219 , \32220 );
or \U$31879 ( \32222 , \17862 , \2080 );
nand \U$31880 ( \32223 , \32221 , \32222 );
nand \U$31881 ( \32224 , \32223 , \2070 );
nand \U$31882 ( \32225 , \32218 , \32224 );
xor \U$31883 ( \32226 , \32215 , \32225 );
and \U$31884 ( \32227 , \32214 , \32226 );
and \U$31885 ( \32228 , \32215 , \32225 );
nor \U$31886 ( \32229 , \32227 , \32228 );
not \U$31887 ( \32230 , \32229 );
not \U$31888 ( \32231 , \9071 );
not \U$31889 ( \32232 , \31905 );
or \U$31890 ( \32233 , \32231 , \32232 );
xor \U$31891 ( \32234 , RI9872a18_166, \8640 );
nand \U$31892 ( \32235 , \32234 , \8027 );
nand \U$31893 ( \32236 , \32233 , \32235 );
not \U$31894 ( \32237 , \32236 );
or \U$31895 ( \32238 , \32230 , \32237 );
or \U$31896 ( \32239 , \32236 , \32229 );
nand \U$31897 ( \32240 , \32238 , \32239 );
not \U$31898 ( \32241 , \32240 );
or \U$31899 ( \32242 , \32203 , \32241 );
not \U$31900 ( \32243 , \32229 );
nand \U$31901 ( \32244 , \32243 , \32236 );
nand \U$31902 ( \32245 , \32242 , \32244 );
not \U$31903 ( \32246 , \32245 );
not \U$31904 ( \32247 , \6063 );
not \U$31905 ( \32248 , \5644 );
not \U$31906 ( \32249 , \11370 );
or \U$31907 ( \32250 , \32248 , \32249 );
or \U$31908 ( \32251 , \17897 , \5648 );
nand \U$31909 ( \32252 , \32250 , \32251 );
not \U$31910 ( \32253 , \32252 );
or \U$31911 ( \32254 , \32247 , \32253 );
nand \U$31912 ( \32255 , \31788 , \5653 );
nand \U$31913 ( \32256 , \32254 , \32255 );
not \U$31914 ( \32257 , \32256 );
and \U$31915 ( \32258 , \5035 , \31926 );
xor \U$31916 ( \32259 , RI9872478_154, \27587 );
and \U$31917 ( \32260 , \32259 , \5034 );
nor \U$31918 ( \32261 , \32258 , \32260 );
not \U$31919 ( \32262 , \32261 );
or \U$31920 ( \32263 , \32257 , \32262 );
or \U$31921 ( \32264 , \32261 , \32256 );
nand \U$31922 ( \32265 , \32263 , \32264 );
not \U$31923 ( \32266 , \32265 );
not \U$31924 ( \32267 , \9293 );
xor \U$31925 ( \32268 , RI9872e50_175, \6528 );
not \U$31926 ( \32269 , \32268 );
or \U$31927 ( \32270 , \32267 , \32269 );
nand \U$31928 ( \32271 , \31808 , \10331 );
nand \U$31929 ( \32272 , \32270 , \32271 );
not \U$31930 ( \32273 , \32272 );
or \U$31931 ( \32274 , \32266 , \32273 );
not \U$31932 ( \32275 , \32261 );
nand \U$31933 ( \32276 , \32275 , \32256 );
nand \U$31934 ( \32277 , \32274 , \32276 );
not \U$31935 ( \32278 , \32277 );
nand \U$31936 ( \32279 , \32246 , \32278 );
not \U$31937 ( \32280 , \32279 );
not \U$31938 ( \32281 , \8801 );
not \U$31939 ( \32282 , \31798 );
or \U$31940 ( \32283 , \32281 , \32282 );
not \U$31941 ( \32284 , \8807 );
not \U$31942 ( \32285 , \21641 );
or \U$31943 ( \32286 , \32284 , \32285 );
or \U$31944 ( \32287 , \21641 , \8811 );
nand \U$31945 ( \32288 , \32286 , \32287 );
nand \U$31946 ( \32289 , \32288 , \22664 );
nand \U$31947 ( \32290 , \32283 , \32289 );
not \U$31948 ( \32291 , \32290 );
buf \U$31949 ( \32292 , \9249 );
not \U$31950 ( \32293 , \32292 );
not \U$31951 ( \32294 , \9244 );
not \U$31952 ( \32295 , \9598 );
or \U$31953 ( \32296 , \32294 , \32295 );
or \U$31954 ( \32297 , \10391 , \9244 );
nand \U$31955 ( \32298 , \32296 , \32297 );
not \U$31956 ( \32299 , \32298 );
or \U$31957 ( \32300 , \32293 , \32299 );
nand \U$31958 ( \32301 , \31822 , \9227 );
nand \U$31959 ( \32302 , \32300 , \32301 );
not \U$31960 ( \32303 , \8742 );
not \U$31961 ( \32304 , \8732 );
not \U$31962 ( \32305 , \5703 );
or \U$31963 ( \32306 , \32304 , \32305 );
or \U$31964 ( \32307 , \8732 , \5703 );
nand \U$31965 ( \32308 , \32306 , \32307 );
not \U$31966 ( \32309 , \32308 );
or \U$31967 ( \32310 , \32303 , \32309 );
nand \U$31968 ( \32311 , \31981 , \11198 );
nand \U$31969 ( \32312 , \32310 , \32311 );
xor \U$31970 ( \32313 , \32302 , \32312 );
not \U$31971 ( \32314 , \32313 );
or \U$31972 ( \32315 , \32291 , \32314 );
nand \U$31973 ( \32316 , \32312 , \32302 );
nand \U$31974 ( \32317 , \32315 , \32316 );
not \U$31975 ( \32318 , \32317 );
or \U$31976 ( \32319 , \32280 , \32318 );
nand \U$31977 ( \32320 , \32277 , \32245 );
nand \U$31978 ( \32321 , \32319 , \32320 );
not \U$31979 ( \32322 , \32321 );
or \U$31980 ( \32323 , \32196 , \32322 );
or \U$31981 ( \32324 , \32321 , \32195 );
nand \U$31982 ( \32325 , \32323 , \32324 );
not \U$31983 ( \32326 , \32325 );
or \U$31984 ( \32327 , \32153 , \32326 );
not \U$31985 ( \32328 , \32195 );
nand \U$31986 ( \32329 , \32328 , \32321 );
nand \U$31987 ( \32330 , \32327 , \32329 );
not \U$31988 ( \32331 , \32330 );
xor \U$31989 ( \32332 , \31666 , \31578 );
xnor \U$31990 ( \32333 , \32332 , \31572 );
not \U$31991 ( \32334 , \32333 );
or \U$31992 ( \32335 , \32331 , \32334 );
or \U$31993 ( \32336 , \32333 , \32330 );
nand \U$31994 ( \32337 , \32335 , \32336 );
not \U$31995 ( \32338 , \32337 );
or \U$31996 ( \32339 , \32139 , \32338 );
not \U$31997 ( \32340 , \32333 );
nand \U$31998 ( \32341 , \32340 , \32330 );
nand \U$31999 ( \32342 , \32339 , \32341 );
not \U$32000 ( \32343 , \32342 );
not \U$32001 ( \32344 , \32343 );
or \U$32002 ( \32345 , \32133 , \32344 );
or \U$32003 ( \32346 , \32343 , \32132 );
nand \U$32004 ( \32347 , \32345 , \32346 );
xnor \U$32005 ( \32348 , \31297 , \31274 );
not \U$32006 ( \32349 , \32348 );
not \U$32007 ( \32350 , \32349 );
xor \U$32008 ( \32351 , \31238 , \31248 );
xor \U$32009 ( \32352 , \32351 , \31256 );
not \U$32010 ( \32353 , \32352 );
not \U$32011 ( \32354 , \32353 );
or \U$32012 ( \32355 , \32350 , \32354 );
not \U$32013 ( \32356 , \32352 );
not \U$32014 ( \32357 , \32348 );
or \U$32015 ( \32358 , \32356 , \32357 );
xor \U$32016 ( \32359 , \31536 , \31545 );
xor \U$32017 ( \32360 , \32359 , \31556 );
nand \U$32018 ( \32361 , \32358 , \32360 );
nand \U$32019 ( \32362 , \32355 , \32361 );
not \U$32020 ( \32363 , \31488 );
xor \U$32021 ( \32364 , \31526 , \31559 );
not \U$32022 ( \32365 , \32364 );
and \U$32023 ( \32366 , \32363 , \32365 );
and \U$32024 ( \32367 , \31488 , \32364 );
nor \U$32025 ( \32368 , \32366 , \32367 );
xor \U$32026 ( \32369 , \32362 , \32368 );
xor \U$32027 ( \32370 , \31263 , \31259 );
xnor \U$32028 ( \32371 , \32370 , \31302 );
xor \U$32029 ( \32372 , \32369 , \32371 );
not \U$32030 ( \32373 , \32028 );
xor \U$32031 ( \32374 , \32018 , \32373 );
xnor \U$32032 ( \32375 , \32374 , \32009 );
not \U$32033 ( \32376 , \32375 );
not \U$32034 ( \32377 , \32376 );
not \U$32035 ( \32378 , \4922 );
not \U$32036 ( \32379 , \32175 );
or \U$32037 ( \32380 , \32378 , \32379 );
not \U$32038 ( \32381 , RI9872388_152);
not \U$32039 ( \32382 , \19591 );
or \U$32040 ( \32383 , \32381 , \32382 );
or \U$32041 ( \32384 , \20928 , RI9872388_152);
nand \U$32042 ( \32385 , \32383 , \32384 );
nand \U$32043 ( \32386 , \32385 , \4918 );
nand \U$32044 ( \32387 , \32380 , \32386 );
not \U$32045 ( \32388 , \32387 );
not \U$32046 ( \32389 , \3169 );
not \U$32047 ( \32390 , \31877 );
or \U$32048 ( \32391 , \32389 , \32390 );
and \U$32049 ( \32392 , RI9872310_151, \16996 );
not \U$32050 ( \32393 , RI9872310_151);
and \U$32051 ( \32394 , \32393 , \16995 );
or \U$32052 ( \32395 , \32392 , \32394 );
nand \U$32053 ( \32396 , \32395 , \3163 );
nand \U$32054 ( \32397 , \32391 , \32396 );
not \U$32055 ( \32398 , \3169 );
not \U$32056 ( \32399 , \32395 );
or \U$32057 ( \32400 , \32398 , \32399 );
not \U$32058 ( \32401 , RI9872310_151);
not \U$32059 ( \32402 , \20490 );
or \U$32060 ( \32403 , \32401 , \32402 );
or \U$32061 ( \32404 , \20490 , RI9872310_151);
nand \U$32062 ( \32405 , \32403 , \32404 );
nand \U$32063 ( \32406 , \32405 , \3163 );
nand \U$32064 ( \32407 , \32400 , \32406 );
not \U$32065 ( \32408 , \32407 );
not \U$32066 ( \32409 , \2085 );
not \U$32067 ( \32410 , \32223 );
or \U$32068 ( \32411 , \32409 , \32410 );
not \U$32069 ( \32412 , \23947 );
not \U$32070 ( \32413 , RI9871aa0_133);
or \U$32071 ( \32414 , \32412 , \32413 );
or \U$32072 ( \32415 , \21773 , RI9871aa0_133);
nand \U$32073 ( \32416 , \32414 , \32415 );
nand \U$32074 ( \32417 , \32416 , \2070 );
nand \U$32075 ( \32418 , \32411 , \32417 );
and \U$32076 ( \32419 , \18704 , \796 );
xor \U$32077 ( \32420 , \32418 , \32419 );
not \U$32078 ( \32421 , \32420 );
or \U$32079 ( \32422 , \32408 , \32421 );
nand \U$32080 ( \32423 , \32418 , \32419 );
nand \U$32081 ( \32424 , \32422 , \32423 );
and \U$32082 ( \32425 , \32397 , \32424 );
not \U$32083 ( \32426 , \32397 );
not \U$32084 ( \32427 , \32424 );
and \U$32085 ( \32428 , \32426 , \32427 );
nor \U$32086 ( \32429 , \32425 , \32428 );
not \U$32087 ( \32430 , \32429 );
or \U$32088 ( \32431 , \32388 , \32430 );
nand \U$32089 ( \32432 , \32424 , \32397 );
nand \U$32090 ( \32433 , \32431 , \32432 );
not \U$32091 ( \32434 , \13109 );
and \U$32092 ( \32435 , \5775 , \14132 );
not \U$32093 ( \32436 , \5775 );
and \U$32094 ( \32437 , \32436 , RI9873030_179);
nor \U$32095 ( \32438 , \32435 , \32437 );
not \U$32096 ( \32439 , \32438 );
or \U$32097 ( \32440 , \32434 , \32439 );
nand \U$32098 ( \32441 , \32016 , \9937 );
nand \U$32099 ( \32442 , \32440 , \32441 );
xor \U$32100 ( \32443 , \32433 , \32442 );
not \U$32101 ( \32444 , \4084 );
not \U$32102 ( \32445 , \32161 );
or \U$32103 ( \32446 , \32444 , \32445 );
xor \U$32104 ( \32447 , \24439 , RI98725e0_157);
nand \U$32105 ( \32448 , \32447 , \4101 );
nand \U$32106 ( \32449 , \32446 , \32448 );
not \U$32107 ( \32450 , \5035 );
not \U$32108 ( \32451 , \32259 );
or \U$32109 ( \32452 , \32450 , \32451 );
xor \U$32110 ( \32453 , RI9872478_154, \21392 );
nand \U$32111 ( \32454 , \32453 , \5034 );
nand \U$32112 ( \32455 , \32452 , \32454 );
xor \U$32113 ( \32456 , \32449 , \32455 );
not \U$32114 ( \32457 , \5641 );
and \U$32115 ( \32458 , RI9872568_156, \13066 );
not \U$32116 ( \32459 , RI9872568_156);
and \U$32117 ( \32460 , \32459 , \13067 );
or \U$32118 ( \32461 , \32458 , \32460 );
not \U$32119 ( \32462 , \32461 );
or \U$32120 ( \32463 , \32457 , \32462 );
nand \U$32121 ( \32464 , \32252 , \5653 );
nand \U$32122 ( \32465 , \32463 , \32464 );
and \U$32123 ( \32466 , \32456 , \32465 );
and \U$32124 ( \32467 , \32449 , \32455 );
or \U$32125 ( \32468 , \32466 , \32467 );
and \U$32126 ( \32469 , \32443 , \32468 );
and \U$32127 ( \32470 , \32433 , \32442 );
or \U$32128 ( \32471 , \32469 , \32470 );
not \U$32129 ( \32472 , \32471 );
xor \U$32130 ( \32473 , \31984 , \32472 );
xnor \U$32131 ( \32474 , \32473 , \31994 );
not \U$32132 ( \32475 , \32474 );
or \U$32133 ( \32476 , \32377 , \32475 );
not \U$32134 ( \32477 , \32472 );
xor \U$32135 ( \32478 , \31994 , \31984 );
nand \U$32136 ( \32479 , \32477 , \32478 );
nand \U$32137 ( \32480 , \32476 , \32479 );
not \U$32138 ( \32481 , \32480 );
not \U$32139 ( \32482 , \32070 );
not \U$32140 ( \32483 , \31998 );
not \U$32141 ( \32484 , \32483 );
or \U$32142 ( \32485 , \32482 , \32484 );
or \U$32143 ( \32486 , \32070 , \32483 );
nand \U$32144 ( \32487 , \32485 , \32486 );
not \U$32145 ( \32488 , \32487 );
xor \U$32146 ( \32489 , \32352 , \32360 );
xnor \U$32147 ( \32490 , \32348 , \32489 );
nand \U$32148 ( \32491 , \32488 , \32490 );
not \U$32149 ( \32492 , \32491 );
or \U$32150 ( \32493 , \32481 , \32492 );
not \U$32151 ( \32494 , \32490 );
nand \U$32152 ( \32495 , \32494 , \32487 );
nand \U$32153 ( \32496 , \32493 , \32495 );
xor \U$32154 ( \32497 , \32372 , \32496 );
xor \U$32155 ( \32498 , \31870 , \31881 );
xor \U$32156 ( \32499 , \32498 , \31897 );
not \U$32157 ( \32500 , \29633 );
and \U$32158 ( \32501 , RI98730a8_180, \4960 );
not \U$32159 ( \32502 , RI98730a8_180);
and \U$32160 ( \32503 , \32502 , \23391 );
nor \U$32161 ( \32504 , \32501 , \32503 );
not \U$32162 ( \32505 , \32504 );
or \U$32163 ( \32506 , \32500 , \32505 );
nand \U$32164 ( \32507 , \32007 , \12867 );
nand \U$32165 ( \32508 , \32506 , \32507 );
xor \U$32166 ( \32509 , \32499 , \32508 );
and \U$32167 ( \32510 , RI98733f0_187, \3240 );
not \U$32168 ( \32511 , RI98733f0_187);
and \U$32169 ( \32512 , \32511 , \3859 );
nor \U$32170 ( \32513 , \32510 , \32512 );
not \U$32171 ( \32514 , \32513 );
or \U$32172 ( \32515 , \32514 , \27186 );
not \U$32173 ( \32516 , \32023 );
nand \U$32174 ( \32517 , \32516 , \17263 );
nand \U$32175 ( \32518 , \32515 , \32517 );
and \U$32176 ( \32519 , \32509 , \32518 );
and \U$32177 ( \32520 , \32499 , \32508 );
or \U$32178 ( \32521 , \32519 , \32520 );
not \U$32179 ( \32522 , \32521 );
not \U$32180 ( \32523 , \17544 );
not \U$32181 ( \32524 , RI9873288_184);
not \U$32182 ( \32525 , \14930 );
or \U$32183 ( \32526 , \32524 , \32525 );
or \U$32184 ( \32527 , \14930 , RI9873288_184);
nand \U$32185 ( \32528 , \32526 , \32527 );
not \U$32186 ( \32529 , \32528 );
or \U$32187 ( \32530 , \32523 , \32529 );
nand \U$32188 ( \32531 , \32050 , \17528 );
nand \U$32189 ( \32532 , \32530 , \32531 );
not \U$32190 ( \32533 , \6610 );
not \U$32191 ( \32534 , \31972 );
or \U$32192 ( \32535 , \32533 , \32534 );
and \U$32193 ( \32536 , \8695 , RI98728b0_163);
not \U$32194 ( \32537 , \8695 );
and \U$32195 ( \32538 , \32537 , \7049 );
nor \U$32196 ( \32539 , \32536 , \32538 );
nand \U$32197 ( \32540 , \32539 , \6284 );
nand \U$32198 ( \32541 , \32535 , \32540 );
xor \U$32199 ( \32542 , \32532 , \32541 );
not \U$32200 ( \32543 , \7325 );
not \U$32201 ( \32544 , \7333 );
not \U$32202 ( \32545 , \10372 );
or \U$32203 ( \32546 , \32544 , \32545 );
nand \U$32204 ( \32547 , \8555 , RI98729a0_165);
nand \U$32205 ( \32548 , \32546 , \32547 );
not \U$32206 ( \32549 , \32548 );
or \U$32207 ( \32550 , \32543 , \32549 );
nand \U$32208 ( \32551 , \31915 , \7338 );
nand \U$32209 ( \32552 , \32550 , \32551 );
and \U$32210 ( \32553 , \32542 , \32552 );
and \U$32211 ( \32554 , \32532 , \32541 );
nor \U$32212 ( \32555 , \32553 , \32554 );
not \U$32213 ( \32556 , \32555 );
and \U$32214 ( \32557 , \32522 , \32556 );
and \U$32215 ( \32558 , \32521 , \32555 );
nor \U$32216 ( \32559 , \32557 , \32558 );
not \U$32217 ( \32560 , \32559 );
not \U$32218 ( \32561 , \32560 );
not \U$32219 ( \32562 , \19046 );
not \U$32220 ( \32563 , \31992 );
or \U$32221 ( \32564 , \32562 , \32563 );
not \U$32222 ( \32565 , RI98734e0_189);
not \U$32223 ( \32566 , \31652 );
or \U$32224 ( \32567 , \32565 , \32566 );
nand \U$32225 ( \32568 , \18453 , \16999 );
nand \U$32226 ( \32569 , \32567 , \32568 );
nand \U$32227 ( \32570 , \32569 , \19244 );
nand \U$32228 ( \32571 , \32564 , \32570 );
not \U$32229 ( \32572 , \32571 );
not \U$32230 ( \32573 , \22670 );
not \U$32231 ( \32574 , \32058 );
or \U$32232 ( \32575 , \32573 , \32574 );
and \U$32233 ( \32576 , RI9873210_183, \4408 );
not \U$32234 ( \32577 , RI9873210_183);
not \U$32235 ( \32578 , \5205 );
and \U$32236 ( \32579 , \32577 , \32578 );
or \U$32237 ( \32580 , \32576 , \32579 );
nand \U$32238 ( \32581 , \32580 , \18957 );
nand \U$32239 ( \32582 , \32575 , \32581 );
not \U$32240 ( \32583 , \32582 );
not \U$32241 ( \32584 , \32583 );
not \U$32242 ( \32585 , \20626 );
not \U$32243 ( \32586 , \18239 );
not \U$32244 ( \32587 , \11755 );
or \U$32245 ( \32588 , \32586 , \32587 );
or \U$32246 ( \32589 , \3395 , \18239 );
nand \U$32247 ( \32590 , \32588 , \32589 );
not \U$32248 ( \32591 , \32590 );
or \U$32249 ( \32592 , \32585 , \32591 );
nand \U$32250 ( \32593 , \32040 , RI9873648_192);
nand \U$32251 ( \32594 , \32592 , \32593 );
not \U$32252 ( \32595 , \32594 );
or \U$32253 ( \32596 , \32584 , \32595 );
or \U$32254 ( \32597 , \32594 , \32583 );
nand \U$32255 ( \32598 , \32596 , \32597 );
not \U$32256 ( \32599 , \32598 );
or \U$32257 ( \32600 , \32572 , \32599 );
nand \U$32258 ( \32601 , \32594 , \32582 );
nand \U$32259 ( \32602 , \32600 , \32601 );
not \U$32260 ( \32603 , \32602 );
or \U$32261 ( \32604 , \32561 , \32603 );
not \U$32262 ( \32605 , \32555 );
nand \U$32263 ( \32606 , \32605 , \32521 );
nand \U$32264 ( \32607 , \32604 , \32606 );
not \U$32265 ( \32608 , \32607 );
not \U$32266 ( \32609 , \31813 );
not \U$32267 ( \32610 , \32609 );
not \U$32268 ( \32611 , \31849 );
and \U$32269 ( \32612 , \32610 , \32611 );
and \U$32270 ( \32613 , \31849 , \32609 );
nor \U$32271 ( \32614 , \32612 , \32613 );
not \U$32272 ( \32615 , \31958 );
not \U$32273 ( \32616 , \31920 );
not \U$32274 ( \32617 , \32616 );
and \U$32275 ( \32618 , \32615 , \32617 );
and \U$32276 ( \32619 , \31958 , \32616 );
nor \U$32277 ( \32620 , \32618 , \32619 );
xor \U$32278 ( \32621 , \32614 , \32620 );
not \U$32279 ( \32622 , \32621 );
or \U$32280 ( \32623 , \32608 , \32622 );
or \U$32281 ( \32624 , \32614 , \32620 );
nand \U$32282 ( \32625 , \32623 , \32624 );
and \U$32283 ( \32626 , \32497 , \32625 );
and \U$32284 ( \32627 , \32372 , \32496 );
or \U$32285 ( \32628 , \32626 , \32627 );
and \U$32286 ( \32629 , \32347 , \32628 );
not \U$32287 ( \32630 , \32347 );
not \U$32288 ( \32631 , \32628 );
and \U$32289 ( \32632 , \32630 , \32631 );
nor \U$32290 ( \32633 , \32629 , \32632 );
xor \U$32291 ( \32634 , \32362 , \32368 );
and \U$32292 ( \32635 , \32634 , \32371 );
and \U$32293 ( \32636 , \32362 , \32368 );
or \U$32294 ( \32637 , \32635 , \32636 );
xor \U$32295 ( \32638 , \31563 , \31675 );
xnor \U$32296 ( \32639 , \32638 , \31670 );
not \U$32297 ( \32640 , \32639 );
xor \U$32298 ( \32641 , \32637 , \32640 );
not \U$32299 ( \32642 , \31736 );
not \U$32300 ( \32643 , \32642 );
not \U$32301 ( \32644 , \31740 );
not \U$32302 ( \32645 , \31729 );
not \U$32303 ( \32646 , \32645 );
or \U$32304 ( \32647 , \32644 , \32646 );
nand \U$32305 ( \32648 , \31729 , \31739 );
nand \U$32306 ( \32649 , \32647 , \32648 );
not \U$32307 ( \32650 , \32649 );
or \U$32308 ( \32651 , \32643 , \32650 );
or \U$32309 ( \32652 , \32649 , \32642 );
nand \U$32310 ( \32653 , \32651 , \32652 );
xor \U$32311 ( \32654 , \31428 , \31414 );
xor \U$32312 ( \32655 , \32653 , \32654 );
xor \U$32313 ( \32656 , \31409 , \31401 );
xor \U$32314 ( \32657 , \31392 , \32656 );
not \U$32315 ( \32658 , \32657 );
not \U$32316 ( \32659 , \32658 );
xor \U$32317 ( \32660 , \31650 , \31589 );
xnor \U$32318 ( \32661 , \32660 , \31660 );
not \U$32319 ( \32662 , \32661 );
not \U$32320 ( \32663 , \32662 );
xnor \U$32321 ( \32664 , \31484 , \31465 );
not \U$32322 ( \32665 , \32664 );
not \U$32323 ( \32666 , \32665 );
or \U$32324 ( \32667 , \32663 , \32666 );
nand \U$32325 ( \32668 , \32664 , \32661 );
nand \U$32326 ( \32669 , \32667 , \32668 );
not \U$32327 ( \32670 , \32669 );
or \U$32328 ( \32671 , \32659 , \32670 );
not \U$32329 ( \32672 , \32662 );
nand \U$32330 ( \32673 , \32672 , \32665 );
nand \U$32331 ( \32674 , \32671 , \32673 );
and \U$32332 ( \32675 , \32655 , \32674 );
and \U$32333 ( \32676 , \32653 , \32654 );
or \U$32334 ( \32677 , \32675 , \32676 );
not \U$32335 ( \32678 , \32677 );
xnor \U$32336 ( \32679 , \32641 , \32678 );
xor \U$32337 ( \32680 , \31780 , \32080 );
xor \U$32338 ( \32681 , \32680 , \32083 );
nand \U$32339 ( \32682 , \32679 , \32681 );
nand \U$32340 ( \32683 , \32633 , \32682 );
not \U$32341 ( \32684 , \32679 );
not \U$32342 ( \32685 , \32681 );
nand \U$32343 ( \32686 , \32684 , \32685 );
nand \U$32344 ( \32687 , \32683 , \32686 );
not \U$32345 ( \32688 , \32687 );
xor \U$32346 ( \32689 , \32128 , \32688 );
not \U$32347 ( \32690 , \32628 );
not \U$32348 ( \32691 , \32347 );
or \U$32349 ( \32692 , \32690 , \32691 );
not \U$32350 ( \32693 , \32343 );
nand \U$32351 ( \32694 , \32693 , \32132 );
nand \U$32352 ( \32695 , \32692 , \32694 );
not \U$32353 ( \32696 , \32695 );
nand \U$32354 ( \32697 , \32677 , \32639 );
nand \U$32355 ( \32698 , \32639 , \32637 );
nand \U$32356 ( \32699 , \32677 , \32637 );
nand \U$32357 ( \32700 , \32697 , \32698 , \32699 );
not \U$32358 ( \32701 , \32700 );
not \U$32359 ( \32702 , \32701 );
not \U$32360 ( \32703 , \31758 );
not \U$32361 ( \32704 , \31756 );
or \U$32362 ( \32705 , \32703 , \32704 );
or \U$32363 ( \32706 , \31756 , \31758 );
nand \U$32364 ( \32707 , \32705 , \32706 );
not \U$32365 ( \32708 , \32707 );
not \U$32366 ( \32709 , \31725 );
and \U$32367 ( \32710 , \32708 , \32709 );
and \U$32368 ( \32711 , \32707 , \31725 );
nor \U$32369 ( \32712 , \32710 , \32711 );
not \U$32370 ( \32713 , \32712 );
not \U$32371 ( \32714 , \32713 );
or \U$32372 ( \32715 , \32702 , \32714 );
nand \U$32373 ( \32716 , \32712 , \32700 );
nand \U$32374 ( \32717 , \32715 , \32716 );
not \U$32375 ( \32718 , \32717 );
not \U$32376 ( \32719 , \32718 );
or \U$32377 ( \32720 , \32696 , \32719 );
not \U$32378 ( \32721 , \32695 );
nand \U$32379 ( \32722 , \32717 , \32721 );
nand \U$32380 ( \32723 , \32720 , \32722 );
buf \U$32381 ( \32724 , \32723 );
xnor \U$32382 ( \32725 , \32689 , \32724 );
nand \U$32383 ( \32726 , \32686 , \32682 );
and \U$32384 ( \32727 , \32726 , \32633 );
not \U$32385 ( \32728 , \32726 );
not \U$32386 ( \32729 , \32633 );
and \U$32387 ( \32730 , \32728 , \32729 );
nor \U$32388 ( \32731 , \32727 , \32730 );
not \U$32389 ( \32732 , \32731 );
not \U$32390 ( \32733 , \32732 );
xor \U$32391 ( \32734 , \32062 , \32042 );
xnor \U$32392 ( \32735 , \32734 , \32052 );
not \U$32393 ( \32736 , \32192 );
and \U$32394 ( \32737 , \32191 , \32736 );
not \U$32395 ( \32738 , \32191 );
and \U$32396 ( \32739 , \32738 , \32192 );
nor \U$32397 ( \32740 , \32737 , \32739 );
nand \U$32398 ( \32741 , \32735 , \32740 );
not \U$32399 ( \32742 , \32741 );
not \U$32400 ( \32743 , \7338 );
not \U$32401 ( \32744 , \32548 );
or \U$32402 ( \32745 , \32743 , \32744 );
not \U$32403 ( \32746 , RI98729a0_165);
not \U$32404 ( \32747 , \18498 );
or \U$32405 ( \32748 , \32746 , \32747 );
or \U$32406 ( \32749 , \13454 , RI98729a0_165);
nand \U$32407 ( \32750 , \32748 , \32749 );
nand \U$32408 ( \32751 , \32750 , \7325 );
nand \U$32409 ( \32752 , \32745 , \32751 );
not \U$32410 ( \32753 , \32752 );
not \U$32411 ( \32754 , \8039 );
not \U$32412 ( \32755 , \32234 );
or \U$32413 ( \32756 , \32754 , \32755 );
xor \U$32414 ( \32757 , RI9872a18_166, \8574 );
nand \U$32415 ( \32758 , \32757 , \8027 );
nand \U$32416 ( \32759 , \32756 , \32758 );
not \U$32417 ( \32760 , \32759 );
not \U$32418 ( \32761 , \4101 );
and \U$32419 ( \32762 , RI98725e0_157, \18709 );
not \U$32420 ( \32763 , RI98725e0_157);
and \U$32421 ( \32764 , \32763 , \25380 );
nor \U$32422 ( \32765 , \32762 , \32764 );
not \U$32423 ( \32766 , \32765 );
or \U$32424 ( \32767 , \32761 , \32766 );
nand \U$32425 ( \32768 , \32447 , \4084 );
nand \U$32426 ( \32769 , \32767 , \32768 );
not \U$32427 ( \32770 , \32769 );
or \U$32428 ( \32771 , RI9872298_150, RI9872310_151);
nand \U$32429 ( \32772 , \32771 , \24450 );
nand \U$32430 ( \32773 , \32772 , \1390 );
not \U$32431 ( \32774 , \32773 );
not \U$32432 ( \32775 , \2085 );
not \U$32433 ( \32776 , \32416 );
or \U$32434 ( \32777 , \32775 , \32776 );
and \U$32435 ( \32778 , RI9871aa0_133, \21779 );
not \U$32436 ( \32779 , RI9871aa0_133);
and \U$32437 ( \32780 , \32779 , \22278 );
nor \U$32438 ( \32781 , \32778 , \32780 );
nand \U$32439 ( \32782 , \32781 , \2070 );
nand \U$32440 ( \32783 , \32777 , \32782 );
nand \U$32441 ( \32784 , \32774 , \32783 );
not \U$32442 ( \32785 , \32784 );
not \U$32443 ( \32786 , \3467 );
not \U$32444 ( \32787 , \32212 );
or \U$32445 ( \32788 , \32786 , \32787 );
and \U$32446 ( \32789 , \17726 , \4063 );
not \U$32447 ( \32790 , \17726 );
and \U$32448 ( \32791 , \32790 , RI98726d0_159);
nor \U$32449 ( \32792 , \32789 , \32791 );
nand \U$32450 ( \32793 , \32792 , \3464 );
nand \U$32451 ( \32794 , \32788 , \32793 );
not \U$32452 ( \32795 , \32794 );
or \U$32453 ( \32796 , \32785 , \32795 );
or \U$32454 ( \32797 , \32794 , \32784 );
nand \U$32455 ( \32798 , \32796 , \32797 );
not \U$32456 ( \32799 , \32798 );
or \U$32457 ( \32800 , \32770 , \32799 );
not \U$32458 ( \32801 , \32784 );
nand \U$32459 ( \32802 , \32801 , \32794 );
nand \U$32460 ( \32803 , \32800 , \32802 );
xnor \U$32461 ( \32804 , \32760 , \32803 );
not \U$32462 ( \32805 , \32804 );
or \U$32463 ( \32806 , \32753 , \32805 );
nand \U$32464 ( \32807 , \32759 , \32803 );
nand \U$32465 ( \32808 , \32806 , \32807 );
not \U$32466 ( \32809 , \32808 );
xnor \U$32467 ( \32810 , \32185 , \32164 );
not \U$32468 ( \32811 , \32810 );
and \U$32469 ( \32812 , \32272 , \32265 );
not \U$32470 ( \32813 , \32272 );
not \U$32471 ( \32814 , \32265 );
and \U$32472 ( \32815 , \32813 , \32814 );
nor \U$32473 ( \32816 , \32812 , \32815 );
not \U$32474 ( \32817 , \32816 );
or \U$32475 ( \32818 , \32811 , \32817 );
or \U$32476 ( \32819 , \32816 , \32810 );
nand \U$32477 ( \32820 , \32818 , \32819 );
not \U$32478 ( \32821 , \32820 );
or \U$32479 ( \32822 , \32809 , \32821 );
not \U$32480 ( \32823 , \32810 );
nand \U$32481 ( \32824 , \32823 , \32816 );
nand \U$32482 ( \32825 , \32822 , \32824 );
not \U$32483 ( \32826 , \32825 );
or \U$32484 ( \32827 , \32742 , \32826 );
not \U$32485 ( \32828 , \32735 );
not \U$32486 ( \32829 , \32740 );
nand \U$32487 ( \32830 , \32828 , \32829 );
nand \U$32488 ( \32831 , \32827 , \32830 );
not \U$32489 ( \32832 , \32831 );
not \U$32490 ( \32833 , \32669 );
not \U$32491 ( \32834 , \32657 );
and \U$32492 ( \32835 , \32833 , \32834 );
and \U$32493 ( \32836 , \32669 , \32657 );
nor \U$32494 ( \32837 , \32835 , \32836 );
not \U$32495 ( \32838 , \32837 );
or \U$32496 ( \32839 , \32832 , \32838 );
or \U$32497 ( \32840 , \32837 , \32831 );
nand \U$32498 ( \32841 , \32839 , \32840 );
not \U$32499 ( \32842 , \12867 );
not \U$32500 ( \32843 , \32504 );
or \U$32501 ( \32844 , \32842 , \32843 );
not \U$32502 ( \32845 , RI98730a8_180);
not \U$32503 ( \32846 , \4985 );
or \U$32504 ( \32847 , \32845 , \32846 );
or \U$32505 ( \32848 , \4985 , RI98730a8_180);
nand \U$32506 ( \32849 , \32847 , \32848 );
nand \U$32507 ( \32850 , \32849 , \24209 );
nand \U$32508 ( \32851 , \32844 , \32850 );
not \U$32509 ( \32852 , \32851 );
not \U$32510 ( \32853 , \32852 );
not \U$32511 ( \32854 , \19243 );
not \U$32512 ( \32855 , RI98734e0_189);
not \U$32513 ( \32856 , \2947 );
or \U$32514 ( \32857 , \32855 , \32856 );
or \U$32515 ( \32858 , \2947 , RI98734e0_189);
nand \U$32516 ( \32859 , \32857 , \32858 );
not \U$32517 ( \32860 , \32859 );
or \U$32518 ( \32861 , \32854 , \32860 );
nand \U$32519 ( \32862 , \32569 , \20147 );
nand \U$32520 ( \32863 , \32861 , \32862 );
not \U$32521 ( \32864 , \32863 );
not \U$32522 ( \32865 , \32864 );
or \U$32523 ( \32866 , \32853 , \32865 );
not \U$32524 ( \32867 , \17234 );
not \U$32525 ( \32868 , \32580 );
or \U$32526 ( \32869 , \32867 , \32868 );
and \U$32527 ( \32870 , RI9873210_183, \12971 );
not \U$32528 ( \32871 , RI9873210_183);
and \U$32529 ( \32872 , \32871 , \5623 );
or \U$32530 ( \32873 , \32870 , \32872 );
nand \U$32531 ( \32874 , \32873 , \17243 );
nand \U$32532 ( \32875 , \32869 , \32874 );
nand \U$32533 ( \32876 , \32866 , \32875 );
nand \U$32534 ( \32877 , \32851 , \32863 );
nand \U$32535 ( \32878 , \32876 , \32877 );
not \U$32536 ( \32879 , \32878 );
xnor \U$32537 ( \32880 , \32240 , \32202 );
not \U$32538 ( \32881 , \32880 );
xor \U$32539 ( \32882 , \32302 , \32290 );
xor \U$32540 ( \32883 , \32882 , \32312 );
not \U$32541 ( \32884 , \32883 );
or \U$32542 ( \32885 , \32881 , \32884 );
or \U$32543 ( \32886 , \32883 , \32880 );
nand \U$32544 ( \32887 , \32885 , \32886 );
not \U$32545 ( \32888 , \32887 );
or \U$32546 ( \32889 , \32879 , \32888 );
not \U$32547 ( \32890 , \32880 );
nand \U$32548 ( \32891 , \32890 , \32883 );
nand \U$32549 ( \32892 , \32889 , \32891 );
not \U$32550 ( \32893 , \32892 );
not \U$32551 ( \32894 , \9668 );
not \U$32552 ( \32895 , \32298 );
or \U$32553 ( \32896 , \32894 , \32895 );
and \U$32554 ( \32897 , RI9872bf8_170, \22347 );
not \U$32555 ( \32898 , RI9872bf8_170);
and \U$32556 ( \32899 , \32898 , \8873 );
or \U$32557 ( \32900 , \32897 , \32899 );
nand \U$32558 ( \32901 , \32900 , \32292 );
nand \U$32559 ( \32902 , \32896 , \32901 );
not \U$32560 ( \32903 , \32902 );
not \U$32561 ( \32904 , \32226 );
not \U$32562 ( \32905 , \32904 );
not \U$32563 ( \32906 , \32214 );
or \U$32564 ( \32907 , \32905 , \32906 );
or \U$32565 ( \32908 , \32214 , \32904 );
nand \U$32566 ( \32909 , \32907 , \32908 );
not \U$32567 ( \32910 , \9214 );
not \U$32568 ( \32911 , \32198 );
or \U$32569 ( \32912 , \32910 , \32911 );
not \U$32570 ( \32913 , RI9872b80_169);
not \U$32571 ( \32914 , \20414 );
or \U$32572 ( \32915 , \32913 , \32914 );
or \U$32573 ( \32916 , \20414 , RI9872b80_169);
nand \U$32574 ( \32917 , \32915 , \32916 );
nand \U$32575 ( \32918 , \32917 , \9195 );
nand \U$32576 ( \32919 , \32912 , \32918 );
xor \U$32577 ( \32920 , \32909 , \32919 );
not \U$32578 ( \32921 , \32920 );
or \U$32579 ( \32922 , \32903 , \32921 );
nand \U$32580 ( \32923 , \32919 , \32909 );
nand \U$32581 ( \32924 , \32922 , \32923 );
not \U$32582 ( \32925 , \32924 );
not \U$32583 ( \32926 , \8800 );
not \U$32584 ( \32927 , \32288 );
or \U$32585 ( \32928 , \32926 , \32927 );
not \U$32586 ( \32929 , RI9872d60_173);
not \U$32587 ( \32930 , \8915 );
or \U$32588 ( \32931 , \32929 , \32930 );
or \U$32589 ( \32932 , \8333 , RI9872d60_173);
nand \U$32590 ( \32933 , \32931 , \32932 );
nand \U$32591 ( \32934 , \32933 , \8818 );
nand \U$32592 ( \32935 , \32928 , \32934 );
not \U$32593 ( \32936 , \32935 );
not \U$32594 ( \32937 , \32936 );
not \U$32595 ( \32938 , \11198 );
not \U$32596 ( \32939 , \32308 );
or \U$32597 ( \32940 , \32938 , \32939 );
and \U$32598 ( \32941 , \8732 , \8052 );
not \U$32599 ( \32942 , \8732 );
and \U$32600 ( \32943 , \32942 , \6296 );
nor \U$32601 ( \32944 , \32941 , \32943 );
nand \U$32602 ( \32945 , \32944 , \9525 );
nand \U$32603 ( \32946 , \32940 , \32945 );
not \U$32604 ( \32947 , \32946 );
not \U$32605 ( \32948 , \32947 );
or \U$32606 ( \32949 , \32937 , \32948 );
not \U$32607 ( \32950 , \10331 );
not \U$32608 ( \32951 , \32268 );
or \U$32609 ( \32952 , \32950 , \32951 );
not \U$32610 ( \32953 , RI9872e50_175);
not \U$32611 ( \32954 , \32953 );
not \U$32612 ( \32955 , \8942 );
or \U$32613 ( \32956 , \32954 , \32955 );
nand \U$32614 ( \32957 , \8943 , RI9872e50_175);
nand \U$32615 ( \32958 , \32956 , \32957 );
nand \U$32616 ( \32959 , \32958 , \9294 );
nand \U$32617 ( \32960 , \32952 , \32959 );
nand \U$32618 ( \32961 , \32949 , \32960 );
nand \U$32619 ( \32962 , \32946 , \32935 );
nand \U$32620 ( \32963 , \32925 , \32961 , \32962 );
not \U$32621 ( \32964 , \32963 );
buf \U$32622 ( \32965 , \18508 );
not \U$32623 ( \32966 , \32965 );
not \U$32624 ( \32967 , RI9873288_184);
and \U$32625 ( \32968 , \32967 , \12616 );
not \U$32626 ( \32969 , \32967 );
and \U$32627 ( \32970 , \32969 , \5594 );
nor \U$32628 ( \32971 , \32968 , \32970 );
not \U$32629 ( \32972 , \32971 );
or \U$32630 ( \32973 , \32966 , \32972 );
nand \U$32631 ( \32974 , \32528 , \17528 );
nand \U$32632 ( \32975 , \32973 , \32974 );
not \U$32633 ( \32976 , \32975 );
not \U$32634 ( \32977 , \6610 );
not \U$32635 ( \32978 , \32539 );
or \U$32636 ( \32979 , \32977 , \32978 );
and \U$32637 ( \32980 , RI98728b0_163, \12460 );
not \U$32638 ( \32981 , RI98728b0_163);
and \U$32639 ( \32982 , \32981 , \8708 );
or \U$32640 ( \32983 , \32980 , \32982 );
nand \U$32641 ( \32984 , \32983 , \6282 );
nand \U$32642 ( \32985 , \32979 , \32984 );
not \U$32643 ( \32986 , \32985 );
or \U$32644 ( \32987 , \32976 , \32986 );
not \U$32645 ( \32988 , \32985 );
not \U$32646 ( \32989 , \32988 );
not \U$32647 ( \32990 , \32975 );
not \U$32648 ( \32991 , \32990 );
or \U$32649 ( \32992 , \32989 , \32991 );
not \U$32650 ( \32993 , RI9873648_192);
not \U$32651 ( \32994 , \32590 );
or \U$32652 ( \32995 , \32993 , \32994 );
and \U$32653 ( \32996 , RI9873558_190, \6382 );
not \U$32654 ( \32997 , RI9873558_190);
and \U$32655 ( \32998 , \32997 , \1485 );
nor \U$32656 ( \32999 , \32996 , \32998 );
nand \U$32657 ( \33000 , \32999 , \20626 );
nand \U$32658 ( \33001 , \32995 , \33000 );
nand \U$32659 ( \33002 , \32992 , \33001 );
nand \U$32660 ( \33003 , \32987 , \33002 );
not \U$32661 ( \33004 , \33003 );
or \U$32662 ( \33005 , \32964 , \33004 );
nand \U$32663 ( \33006 , \32961 , \32962 );
nand \U$32664 ( \33007 , \33006 , \32924 );
nand \U$32665 ( \33008 , \33005 , \33007 );
not \U$32666 ( \33009 , \32245 );
not \U$32667 ( \33010 , \32278 );
or \U$32668 ( \33011 , \33009 , \33010 );
or \U$32669 ( \33012 , \32278 , \32245 );
nand \U$32670 ( \33013 , \33011 , \33012 );
xnor \U$32671 ( \33014 , \32317 , \33013 );
xnor \U$32672 ( \33015 , \33008 , \33014 );
not \U$32673 ( \33016 , \33015 );
or \U$32674 ( \33017 , \32893 , \33016 );
not \U$32675 ( \33018 , \33014 );
nand \U$32676 ( \33019 , \33018 , \33008 );
nand \U$32677 ( \33020 , \33017 , \33019 );
xor \U$32678 ( \33021 , \32841 , \33020 );
not \U$32679 ( \33022 , \33021 );
nand \U$32680 ( \33023 , \32491 , \32495 );
buf \U$32681 ( \33024 , \32480 );
and \U$32682 ( \33025 , \33023 , \33024 );
not \U$32683 ( \33026 , \33023 );
not \U$32684 ( \33027 , \33024 );
and \U$32685 ( \33028 , \33026 , \33027 );
nor \U$32686 ( \33029 , \33025 , \33028 );
not \U$32687 ( \33030 , \33029 );
not \U$32688 ( \33031 , \17234 );
not \U$32689 ( \33032 , \32873 );
or \U$32690 ( \33033 , \33031 , \33032 );
xnor \U$32691 ( \33034 , \4988 , RI9873210_183);
nand \U$32692 ( \33035 , \33034 , \13477 );
nand \U$32693 ( \33036 , \33033 , \33035 );
not \U$32694 ( \33037 , \33036 );
xnor \U$32695 ( \33038 , \32798 , \32769 );
not \U$32696 ( \33039 , \33038 );
not \U$32697 ( \33040 , \20147 );
not \U$32698 ( \33041 , \32859 );
or \U$32699 ( \33042 , \33040 , \33041 );
not \U$32700 ( \33043 , \19304 );
and \U$32701 ( \33044 , \16999 , \33043 );
not \U$32702 ( \33045 , \16999 );
and \U$32703 ( \33046 , \33045 , \3239 );
nor \U$32704 ( \33047 , \33044 , \33046 );
nand \U$32705 ( \33048 , \33047 , \19035 );
nand \U$32706 ( \33049 , \33042 , \33048 );
not \U$32707 ( \33050 , \33049 );
or \U$32708 ( \33051 , \33039 , \33050 );
or \U$32709 ( \33052 , \33049 , \33038 );
nand \U$32710 ( \33053 , \33051 , \33052 );
not \U$32711 ( \33054 , \33053 );
or \U$32712 ( \33055 , \33037 , \33054 );
not \U$32713 ( \33056 , \33038 );
nand \U$32714 ( \33057 , \33056 , \33049 );
nand \U$32715 ( \33058 , \33055 , \33057 );
not \U$32716 ( \33059 , \33058 );
not \U$32717 ( \33060 , \8027 );
not \U$32718 ( \33061 , RI9872a18_166);
not \U$32719 ( \33062 , \8554 );
or \U$32720 ( \33063 , \33061 , \33062 );
or \U$32721 ( \33064 , \8554 , RI9872a18_166);
nand \U$32722 ( \33065 , \33063 , \33064 );
not \U$32723 ( \33066 , \33065 );
or \U$32724 ( \33067 , \33060 , \33066 );
nand \U$32725 ( \33068 , \32757 , \9071 );
nand \U$32726 ( \33069 , \33067 , \33068 );
not \U$32727 ( \33070 , \3169 );
not \U$32728 ( \33071 , \32405 );
or \U$32729 ( \33072 , \33070 , \33071 );
not \U$32730 ( \33073 , RI9872310_151);
not \U$32731 ( \33074 , \19542 );
or \U$32732 ( \33075 , \33073 , \33074 );
nand \U$32733 ( \33076 , \24854 , \3154 );
nand \U$32734 ( \33077 , \33075 , \33076 );
nand \U$32735 ( \33078 , \33077 , \3163 );
nand \U$32736 ( \33079 , \33072 , \33078 );
not \U$32737 ( \33080 , \33079 );
xor \U$32738 ( \33081 , \32783 , \32773 );
not \U$32739 ( \33082 , \33081 );
or \U$32740 ( \33083 , \33080 , \33082 );
or \U$32741 ( \33084 , \33079 , \33081 );
nand \U$32742 ( \33085 , \33083 , \33084 );
not \U$32743 ( \33086 , \33085 );
not \U$32744 ( \33087 , \4084 );
not \U$32745 ( \33088 , \32765 );
or \U$32746 ( \33089 , \33087 , \33088 );
not \U$32747 ( \33090 , \4088 );
not \U$32748 ( \33091 , \28191 );
or \U$32749 ( \33092 , \33090 , \33091 );
nand \U$32750 ( \33093 , \17911 , RI98725e0_157);
nand \U$32751 ( \33094 , \33092 , \33093 );
nand \U$32752 ( \33095 , \33094 , \4101 );
nand \U$32753 ( \33096 , \33089 , \33095 );
not \U$32754 ( \33097 , \33096 );
or \U$32755 ( \33098 , \33086 , \33097 );
not \U$32756 ( \33099 , \33081 );
nand \U$32757 ( \33100 , \33099 , \33079 );
nand \U$32758 ( \33101 , \33098 , \33100 );
and \U$32759 ( \33102 , \33069 , \33101 );
not \U$32760 ( \33103 , \33069 );
not \U$32761 ( \33104 , \33101 );
and \U$32762 ( \33105 , \33103 , \33104 );
nor \U$32763 ( \33106 , \33102 , \33105 );
not \U$32764 ( \33107 , \33106 );
not \U$32765 ( \33108 , \18672 );
not \U$32766 ( \33109 , \14132 );
not \U$32767 ( \33110 , \6303 );
or \U$32768 ( \33111 , \33109 , \33110 );
nand \U$32769 ( \33112 , \21955 , RI9873030_179);
nand \U$32770 ( \33113 , \33111 , \33112 );
not \U$32771 ( \33114 , \33113 );
or \U$32772 ( \33115 , \33108 , \33114 );
and \U$32773 ( \33116 , RI9873030_179, \5761 );
not \U$32774 ( \33117 , RI9873030_179);
and \U$32775 ( \33118 , \33117 , \6058 );
or \U$32776 ( \33119 , \33116 , \33118 );
nand \U$32777 ( \33120 , \33119 , \9937 );
nand \U$32778 ( \33121 , \33115 , \33120 );
not \U$32779 ( \33122 , \33121 );
or \U$32780 ( \33123 , \33107 , \33122 );
nand \U$32781 ( \33124 , \33069 , \33101 );
nand \U$32782 ( \33125 , \33123 , \33124 );
not \U$32783 ( \33126 , \33125 );
and \U$32784 ( \33127 , RI98728b0_163, \11371 );
not \U$32785 ( \33128 , RI98728b0_163);
and \U$32786 ( \33129 , \33128 , \18344 );
or \U$32787 ( \33130 , \33127 , \33129 );
nand \U$32788 ( \33131 , \33130 , \6282 );
not \U$32789 ( \33132 , \32385 );
not \U$32790 ( \33133 , \33132 );
not \U$32791 ( \33134 , \32178 );
and \U$32792 ( \33135 , \33133 , \33134 );
and \U$32793 ( \33136 , RI9872388_152, \29137 );
not \U$32794 ( \33137 , RI9872388_152);
and \U$32795 ( \33138 , \33137 , \22395 );
or \U$32796 ( \33139 , \33136 , \33138 );
and \U$32797 ( \33140 , \33139 , \4918 );
nor \U$32798 ( \33141 , \33135 , \33140 );
nand \U$32799 ( \33142 , \32983 , \6286 );
nand \U$32800 ( \33143 , \33131 , \33141 , \33142 );
not \U$32801 ( \33144 , \33143 );
not \U$32802 ( \33145 , \9526 );
not \U$32803 ( \33146 , \8732 );
not \U$32804 ( \33147 , \6528 );
or \U$32805 ( \33148 , \33146 , \33147 );
or \U$32806 ( \33149 , \10412 , \8732 );
nand \U$32807 ( \33150 , \33148 , \33149 );
not \U$32808 ( \33151 , \33150 );
or \U$32809 ( \33152 , \33145 , \33151 );
nand \U$32810 ( \33153 , \32944 , \11198 );
nand \U$32811 ( \33154 , \33152 , \33153 );
not \U$32812 ( \33155 , \33154 );
or \U$32813 ( \33156 , \33144 , \33155 );
not \U$32814 ( \33157 , \33141 );
nand \U$32815 ( \33158 , \33131 , \33142 );
nand \U$32816 ( \33159 , \33157 , \33158 );
nand \U$32817 ( \33160 , \33156 , \33159 );
not \U$32818 ( \33161 , \33160 );
not \U$32819 ( \33162 , \33161 );
or \U$32820 ( \33163 , \33126 , \33162 );
not \U$32821 ( \33164 , \33125 );
nand \U$32822 ( \33165 , \33164 , \33160 );
nand \U$32823 ( \33166 , \33163 , \33165 );
not \U$32824 ( \33167 , \33166 );
or \U$32825 ( \33168 , \33059 , \33167 );
nand \U$32826 ( \33169 , \33160 , \33125 );
nand \U$32827 ( \33170 , \33168 , \33169 );
xor \U$32828 ( \33171 , \32902 , \32920 );
not \U$32829 ( \33172 , \7326 );
not \U$32830 ( \33173 , \7333 );
not \U$32831 ( \33174 , \9750 );
or \U$32832 ( \33175 , \33173 , \33174 );
or \U$32833 ( \33176 , \24808 , \7333 );
nand \U$32834 ( \33177 , \33175 , \33176 );
not \U$32835 ( \33178 , \33177 );
or \U$32836 ( \33179 , \33172 , \33178 );
nand \U$32837 ( \33180 , \32750 , \7338 );
nand \U$32838 ( \33181 , \33179 , \33180 );
not \U$32839 ( \33182 , \33181 );
not \U$32840 ( \33183 , \9195 );
xor \U$32841 ( \33184 , RI9872b80_169, \8640 );
not \U$32842 ( \33185 , \33184 );
or \U$32843 ( \33186 , \33183 , \33185 );
nand \U$32844 ( \33187 , \32917 , \9214 );
nand \U$32845 ( \33188 , \33186 , \33187 );
not \U$32846 ( \33189 , \33188 );
nand \U$32847 ( \33190 , \33182 , \33189 );
not \U$32848 ( \33191 , \33190 );
not \U$32849 ( \33192 , \17528 );
not \U$32850 ( \33193 , \32971 );
or \U$32851 ( \33194 , \33192 , \33193 );
and \U$32852 ( \33195 , RI9873288_184, \4408 );
not \U$32853 ( \33196 , RI9873288_184);
and \U$32854 ( \33197 , \33196 , \22043 );
or \U$32855 ( \33198 , \33195 , \33197 );
nand \U$32856 ( \33199 , \33198 , \17544 );
nand \U$32857 ( \33200 , \33194 , \33199 );
not \U$32858 ( \33201 , \33200 );
or \U$32859 ( \33202 , \33191 , \33201 );
nand \U$32860 ( \33203 , \33188 , \33181 );
nand \U$32861 ( \33204 , \33202 , \33203 );
xor \U$32862 ( \33205 , \33171 , \33204 );
not \U$32863 ( \33206 , \22618 );
not \U$32864 ( \33207 , \32849 );
or \U$32865 ( \33208 , \33206 , \33207 );
not \U$32866 ( \33209 , \5775 );
xor \U$32867 ( \33210 , RI98730a8_180, \33209 );
nand \U$32868 ( \33211 , \33210 , \24209 );
nand \U$32869 ( \33212 , \33208 , \33211 );
not \U$32870 ( \33213 , \17251 );
not \U$32871 ( \33214 , \17539 );
not \U$32872 ( \33215 , \16906 );
or \U$32873 ( \33216 , \33214 , \33215 );
not \U$32874 ( \33217 , \17522 );
nand \U$32875 ( \33218 , \33217 , \14930 );
nand \U$32876 ( \33219 , \33216 , \33218 );
not \U$32877 ( \33220 , \33219 );
or \U$32878 ( \33221 , \33213 , \33220 );
not \U$32879 ( \33222 , \17539 );
not \U$32880 ( \33223 , \3536 );
or \U$32881 ( \33224 , \33222 , \33223 );
or \U$32882 ( \33225 , \3537 , \17539 );
nand \U$32883 ( \33226 , \33224 , \33225 );
nand \U$32884 ( \33227 , \33226 , \17263 );
nand \U$32885 ( \33228 , \33221 , \33227 );
xor \U$32886 ( \33229 , \33212 , \33228 );
not \U$32887 ( \33230 , \18545 );
not \U$32888 ( \33231 , RI9873558_190);
not \U$32889 ( \33232 , \6378 );
or \U$32890 ( \33233 , \33231 , \33232 );
or \U$32891 ( \33234 , \7164 , RI9873558_190);
nand \U$32892 ( \33235 , \33233 , \33234 );
not \U$32893 ( \33236 , \33235 );
or \U$32894 ( \33237 , \33230 , \33236 );
nand \U$32895 ( \33238 , \32999 , RI9873648_192);
nand \U$32896 ( \33239 , \33237 , \33238 );
and \U$32897 ( \33240 , \33229 , \33239 );
and \U$32898 ( \33241 , \33212 , \33228 );
or \U$32899 ( \33242 , \33240 , \33241 );
and \U$32900 ( \33243 , \33205 , \33242 );
and \U$32901 ( \33244 , \33171 , \33204 );
or \U$32902 ( \33245 , \33243 , \33244 );
xor \U$32903 ( \33246 , \33170 , \33245 );
not \U$32904 ( \33247 , \33003 );
and \U$32905 ( \33248 , \33006 , \32924 );
not \U$32906 ( \33249 , \33006 );
and \U$32907 ( \33250 , \33249 , \32925 );
nor \U$32908 ( \33251 , \33248 , \33250 );
not \U$32909 ( \33252 , \33251 );
and \U$32910 ( \33253 , \33247 , \33252 );
and \U$32911 ( \33254 , \33003 , \33251 );
nor \U$32912 ( \33255 , \33253 , \33254 );
and \U$32913 ( \33256 , \33246 , \33255 );
and \U$32914 ( \33257 , \33170 , \33245 );
or \U$32915 ( \33258 , \33256 , \33257 );
not \U$32916 ( \33259 , \33258 );
xor \U$32917 ( \33260 , \32433 , \32442 );
xor \U$32918 ( \33261 , \33260 , \32468 );
not \U$32919 ( \33262 , \8818 );
not \U$32920 ( \33263 , \11627 );
xor \U$32921 ( \33264 , RI9872d60_173, \33263 );
not \U$32922 ( \33265 , \33264 );
or \U$32923 ( \33266 , \33262 , \33265 );
nand \U$32924 ( \33267 , \32933 , \8800 );
nand \U$32925 ( \33268 , \33266 , \33267 );
not \U$32926 ( \33269 , \33268 );
not \U$32927 ( \33270 , \9249 );
and \U$32928 ( \33271 , RI9872bf8_170, \8596 );
not \U$32929 ( \33272 , RI9872bf8_170);
and \U$32930 ( \33273 , \33272 , \18110 );
nor \U$32931 ( \33274 , \33271 , \33273 );
not \U$32932 ( \33275 , \33274 );
or \U$32933 ( \33276 , \33270 , \33275 );
nand \U$32934 ( \33277 , \32900 , \22167 );
nand \U$32935 ( \33278 , \33276 , \33277 );
not \U$32936 ( \33279 , \33278 );
or \U$32937 ( \33280 , \33269 , \33279 );
not \U$32938 ( \33281 , \33278 );
not \U$32939 ( \33282 , \33281 );
not \U$32940 ( \33283 , \33268 );
not \U$32941 ( \33284 , \33283 );
or \U$32942 ( \33285 , \33282 , \33284 );
not \U$32943 ( \33286 , \9273 );
not \U$32944 ( \33287 , \32958 );
or \U$32945 ( \33288 , \33286 , \33287 );
not \U$32946 ( \33289 , RI9872e50_175);
not \U$32947 ( \33290 , \7466 );
or \U$32948 ( \33291 , \33289 , \33290 );
or \U$32949 ( \33292 , \8924 , RI9872e50_175);
nand \U$32950 ( \33293 , \33291 , \33292 );
nand \U$32951 ( \33294 , \33293 , \9294 );
nand \U$32952 ( \33295 , \33288 , \33294 );
nand \U$32953 ( \33296 , \33285 , \33295 );
nand \U$32954 ( \33297 , \33280 , \33296 );
not \U$32955 ( \33298 , \33297 );
xor \U$32956 ( \33299 , \32449 , \32455 );
xor \U$32957 ( \33300 , \33299 , \32465 );
not \U$32958 ( \33301 , \33300 );
not \U$32959 ( \33302 , \5653 );
not \U$32960 ( \33303 , \32461 );
or \U$32961 ( \33304 , \33302 , \33303 );
and \U$32962 ( \33305 , RI9872568_156, \13391 );
not \U$32963 ( \33306 , RI9872568_156);
not \U$32964 ( \33307 , \13391 );
and \U$32965 ( \33308 , \33306 , \33307 );
or \U$32966 ( \33309 , \33305 , \33308 );
nand \U$32967 ( \33310 , \33309 , \6063 );
nand \U$32968 ( \33311 , \33304 , \33310 );
xor \U$32969 ( \33312 , \32407 , \32420 );
not \U$32970 ( \33313 , \33312 );
not \U$32971 ( \33314 , \5034 );
and \U$32972 ( \33315 , RI9872478_154, \17081 );
not \U$32973 ( \33316 , RI9872478_154);
and \U$32974 ( \33317 , \33316 , \12773 );
nor \U$32975 ( \33318 , \33315 , \33317 );
not \U$32976 ( \33319 , \33318 );
or \U$32977 ( \33320 , \33314 , \33319 );
nand \U$32978 ( \33321 , \32453 , \5035 );
nand \U$32979 ( \33322 , \33320 , \33321 );
not \U$32980 ( \33323 , \33322 );
not \U$32981 ( \33324 , \33323 );
or \U$32982 ( \33325 , \33313 , \33324 );
or \U$32983 ( \33326 , \33323 , \33312 );
nand \U$32984 ( \33327 , \33325 , \33326 );
and \U$32985 ( \33328 , \33311 , \33327 );
not \U$32986 ( \33329 , \33312 );
nor \U$32987 ( \33330 , \33329 , \33323 );
nor \U$32988 ( \33331 , \33328 , \33330 );
not \U$32989 ( \33332 , \33331 );
or \U$32990 ( \33333 , \33301 , \33332 );
or \U$32991 ( \33334 , \33331 , \33300 );
nand \U$32992 ( \33335 , \33333 , \33334 );
not \U$32993 ( \33336 , \33335 );
or \U$32994 ( \33337 , \33298 , \33336 );
not \U$32995 ( \33338 , \33331 );
nand \U$32996 ( \33339 , \33338 , \33300 );
nand \U$32997 ( \33340 , \33337 , \33339 );
xor \U$32998 ( \33341 , \33261 , \33340 );
xor \U$32999 ( \33342 , \32499 , \32508 );
xor \U$33000 ( \33343 , \33342 , \32518 );
and \U$33001 ( \33344 , \33341 , \33343 );
and \U$33002 ( \33345 , \33261 , \33340 );
or \U$33003 ( \33346 , \33344 , \33345 );
xor \U$33004 ( \33347 , \32375 , \33346 );
xnor \U$33005 ( \33348 , \33347 , \32474 );
not \U$33006 ( \33349 , \33348 );
or \U$33007 ( \33350 , \33259 , \33349 );
and \U$33008 ( \33351 , \32474 , \32375 );
not \U$33009 ( \33352 , \32474 );
and \U$33010 ( \33353 , \33352 , \32376 );
or \U$33011 ( \33354 , \33351 , \33353 );
nand \U$33012 ( \33355 , \33354 , \33346 );
nand \U$33013 ( \33356 , \33350 , \33355 );
not \U$33014 ( \33357 , \33356 );
or \U$33015 ( \33358 , \33030 , \33357 );
or \U$33016 ( \33359 , \33356 , \33029 );
nand \U$33017 ( \33360 , \33358 , \33359 );
not \U$33018 ( \33361 , \33360 );
or \U$33019 ( \33362 , \33022 , \33361 );
not \U$33020 ( \33363 , \33029 );
nand \U$33021 ( \33364 , \33363 , \33356 );
nand \U$33022 ( \33365 , \33362 , \33364 );
xnor \U$33023 ( \33366 , \32337 , \32138 );
xor \U$33024 ( \33367 , \32372 , \32496 );
xor \U$33025 ( \33368 , \33367 , \32625 );
xnor \U$33026 ( \33369 , \33366 , \33368 );
nand \U$33027 ( \33370 , \33365 , \33369 );
not \U$33028 ( \33371 , \33366 );
nand \U$33029 ( \33372 , \33371 , \33368 );
nand \U$33030 ( \33373 , \33370 , \33372 );
xor \U$33031 ( \33374 , \32653 , \32654 );
xor \U$33032 ( \33375 , \33374 , \32674 );
not \U$33033 ( \33376 , \33020 );
not \U$33034 ( \33377 , \32841 );
or \U$33035 ( \33378 , \33376 , \33377 );
not \U$33036 ( \33379 , \32837 );
nand \U$33037 ( \33380 , \33379 , \32831 );
nand \U$33038 ( \33381 , \33378 , \33380 );
xor \U$33039 ( \33382 , \33375 , \33381 );
not \U$33040 ( \33383 , \33382 );
xor \U$33041 ( \33384 , \32144 , \32146 );
xor \U$33042 ( \33385 , \33384 , \32149 );
not \U$33043 ( \33386 , \33385 );
xnor \U$33044 ( \33387 , \32602 , \32560 );
not \U$33045 ( \33388 , \33387 );
not \U$33046 ( \33389 , \33388 );
or \U$33047 ( \33390 , \33386 , \33389 );
not \U$33048 ( \33391 , \33385 );
not \U$33049 ( \33392 , \33391 );
not \U$33050 ( \33393 , \33387 );
or \U$33051 ( \33394 , \33392 , \33393 );
not \U$33052 ( \33395 , \32552 );
not \U$33053 ( \33396 , \33395 );
not \U$33054 ( \33397 , \32542 );
or \U$33055 ( \33398 , \33396 , \33397 );
or \U$33056 ( \33399 , \32542 , \33395 );
nand \U$33057 ( \33400 , \33398 , \33399 );
not \U$33058 ( \33401 , \33400 );
xor \U$33059 ( \33402 , \32571 , \32583 );
xnor \U$33060 ( \33403 , \33402 , \32594 );
not \U$33061 ( \33404 , \33403 );
or \U$33062 ( \33405 , \33401 , \33404 );
or \U$33063 ( \33406 , \33403 , \33400 );
not \U$33064 ( \33407 , \9937 );
not \U$33065 ( \33408 , \32438 );
or \U$33066 ( \33409 , \33407 , \33408 );
nand \U$33067 ( \33410 , \33119 , \18672 );
nand \U$33068 ( \33411 , \33409 , \33410 );
not \U$33069 ( \33412 , \33411 );
not \U$33070 ( \33413 , \19282 );
not \U$33071 ( \33414 , \32513 );
or \U$33072 ( \33415 , \33413 , \33414 );
nand \U$33073 ( \33416 , \33226 , \17252 );
nand \U$33074 ( \33417 , \33415 , \33416 );
xor \U$33075 ( \33418 , \32387 , \32429 );
xor \U$33076 ( \33419 , \33417 , \33418 );
not \U$33077 ( \33420 , \33419 );
or \U$33078 ( \33421 , \33412 , \33420 );
nand \U$33079 ( \33422 , \33417 , \33418 );
nand \U$33080 ( \33423 , \33421 , \33422 );
nand \U$33081 ( \33424 , \33406 , \33423 );
nand \U$33082 ( \33425 , \33405 , \33424 );
nand \U$33083 ( \33426 , \33394 , \33425 );
nand \U$33084 ( \33427 , \33390 , \33426 );
not \U$33085 ( \33428 , \33427 );
xnor \U$33086 ( \33429 , \32325 , \32152 );
not \U$33087 ( \33430 , \33429 );
not \U$33088 ( \33431 , \33430 );
xor \U$33089 ( \33432 , \32607 , \32621 );
not \U$33090 ( \33433 , \33432 );
not \U$33091 ( \33434 , \33433 );
or \U$33092 ( \33435 , \33431 , \33434 );
nand \U$33093 ( \33436 , \33432 , \33429 );
nand \U$33094 ( \33437 , \33435 , \33436 );
not \U$33095 ( \33438 , \33437 );
or \U$33096 ( \33439 , \33428 , \33438 );
nand \U$33097 ( \33440 , \33432 , \33430 );
nand \U$33098 ( \33441 , \33439 , \33440 );
not \U$33099 ( \33442 , \33441 );
or \U$33100 ( \33443 , \33383 , \33442 );
nand \U$33101 ( \33444 , \33375 , \33381 );
nand \U$33102 ( \33445 , \33443 , \33444 );
xor \U$33103 ( \33446 , \33373 , \33445 );
not \U$33104 ( \33447 , \33446 );
or \U$33105 ( \33448 , \32733 , \33447 );
not \U$33106 ( \33449 , \33372 );
not \U$33107 ( \33450 , \33370 );
or \U$33108 ( \33451 , \33449 , \33450 );
nand \U$33109 ( \33452 , \33451 , \33445 );
nand \U$33110 ( \33453 , \33448 , \33452 );
not \U$33111 ( \33454 , \33453 );
nand \U$33112 ( \33455 , \32725 , \33454 );
and \U$33113 ( \33456 , \33365 , \33369 );
not \U$33114 ( \33457 , \33365 );
not \U$33115 ( \33458 , \33369 );
and \U$33116 ( \33459 , \33457 , \33458 );
nor \U$33117 ( \33460 , \33456 , \33459 );
not \U$33118 ( \33461 , \33460 );
xor \U$33119 ( \33462 , \33441 , \33382 );
not \U$33120 ( \33463 , \33462 );
not \U$33121 ( \33464 , \33463 );
xor \U$33122 ( \33465 , \33348 , \33258 );
not \U$33123 ( \33466 , \33465 );
xor \U$33124 ( \33467 , \33261 , \33340 );
xor \U$33125 ( \33468 , \33467 , \33343 );
xor \U$33126 ( \33469 , \33400 , \33423 );
xor \U$33127 ( \33470 , \33469 , \33403 );
xor \U$33128 ( \33471 , \33468 , \33470 );
not \U$33129 ( \33472 , \3467 );
and \U$33130 ( \33473 , RI98726d0_159, \21553 );
not \U$33131 ( \33474 , RI98726d0_159);
and \U$33132 ( \33475 , \33474 , \24868 );
or \U$33133 ( \33476 , \33473 , \33475 );
not \U$33134 ( \33477 , \33476 );
or \U$33135 ( \33478 , \33472 , \33477 );
not \U$33136 ( \33479 , \27541 );
and \U$33137 ( \33480 , RI98726d0_159, \33479 );
not \U$33138 ( \33481 , RI98726d0_159);
not \U$33139 ( \33482 , \28653 );
and \U$33140 ( \33483 , \33481 , \33482 );
nor \U$33141 ( \33484 , \33480 , \33483 );
nand \U$33142 ( \33485 , \33484 , \3464 );
nand \U$33143 ( \33486 , \33478 , \33485 );
not \U$33144 ( \33487 , \33486 );
and \U$33145 ( \33488 , \21779 , \2085 );
not \U$33146 ( \33489 , \33488 );
not \U$33147 ( \33490 , \3169 );
not \U$33148 ( \33491 , \33077 );
or \U$33149 ( \33492 , \33490 , \33491 );
not \U$33150 ( \33493 , RI9872310_151);
not \U$33151 ( \33494 , \21773 );
or \U$33152 ( \33495 , \33493 , \33494 );
nand \U$33153 ( \33496 , \23948 , \3154 );
nand \U$33154 ( \33497 , \33495 , \33496 );
nand \U$33155 ( \33498 , \33497 , \3162 );
nand \U$33156 ( \33499 , \33492 , \33498 );
not \U$33157 ( \33500 , \33499 );
not \U$33158 ( \33501 , \33500 );
or \U$33159 ( \33502 , \33489 , \33501 );
not \U$33160 ( \33503 , \33488 );
nand \U$33161 ( \33504 , \33503 , \33499 );
nand \U$33162 ( \33505 , \33502 , \33504 );
not \U$33163 ( \33506 , \33505 );
or \U$33164 ( \33507 , \33487 , \33506 );
nand \U$33165 ( \33508 , \33499 , \33488 );
nand \U$33166 ( \33509 , \33507 , \33508 );
not \U$33167 ( \33510 , \33509 );
not \U$33168 ( \33511 , \3467 );
not \U$33169 ( \33512 , \32792 );
or \U$33170 ( \33513 , \33511 , \33512 );
nand \U$33171 ( \33514 , \33476 , \3464 );
nand \U$33172 ( \33515 , \33513 , \33514 );
not \U$33173 ( \33516 , \33515 );
not \U$33174 ( \33517 , \33516 );
and \U$33175 ( \33518 , \33510 , \33517 );
and \U$33176 ( \33519 , \33509 , \33516 );
nor \U$33177 ( \33520 , \33518 , \33519 );
not \U$33178 ( \33521 , \33520 );
not \U$33179 ( \33522 , \33521 );
not \U$33180 ( \33523 , \5653 );
not \U$33181 ( \33524 , \33309 );
or \U$33182 ( \33525 , \33523 , \33524 );
and \U$33183 ( \33526 , RI9872568_156, \18155 );
not \U$33184 ( \33527 , RI9872568_156);
and \U$33185 ( \33528 , \33527 , \18152 );
nor \U$33186 ( \33529 , \33526 , \33528 );
not \U$33187 ( \33530 , \33529 );
nand \U$33188 ( \33531 , \33530 , \6063 );
nand \U$33189 ( \33532 , \33525 , \33531 );
not \U$33190 ( \33533 , \33532 );
or \U$33191 ( \33534 , \33522 , \33533 );
nand \U$33192 ( \33535 , \33509 , \33515 );
nand \U$33193 ( \33536 , \33534 , \33535 );
not \U$33194 ( \33537 , \6284 );
not \U$33195 ( \33538 , \5632 );
not \U$33196 ( \33539 , \17757 );
not \U$33197 ( \33540 , \33539 );
or \U$33198 ( \33541 , \33538 , \33540 );
nand \U$33199 ( \33542 , \13066 , RI98728b0_163);
nand \U$33200 ( \33543 , \33541 , \33542 );
not \U$33201 ( \33544 , \33543 );
or \U$33202 ( \33545 , \33537 , \33544 );
nand \U$33203 ( \33546 , \33130 , \6286 );
nand \U$33204 ( \33547 , \33545 , \33546 );
not \U$33205 ( \33548 , \33547 );
not \U$33206 ( \33549 , \4922 );
not \U$33207 ( \33550 , \33139 );
or \U$33208 ( \33551 , \33549 , \33550 );
not \U$33209 ( \33552 , \4902 );
not \U$33210 ( \33553 , \13861 );
or \U$33211 ( \33554 , \33552 , \33553 );
or \U$33212 ( \33555 , \17883 , \4902 );
nand \U$33213 ( \33556 , \33554 , \33555 );
nand \U$33214 ( \33557 , \33556 , \4918 );
nand \U$33215 ( \33558 , \33551 , \33557 );
not \U$33216 ( \33559 , \33558 );
not \U$33217 ( \33560 , \5035 );
not \U$33218 ( \33561 , \33318 );
or \U$33219 ( \33562 , \33560 , \33561 );
and \U$33220 ( \33563 , RI9872478_154, \13281 );
not \U$33221 ( \33564 , RI9872478_154);
and \U$33222 ( \33565 , \33564 , \19591 );
nor \U$33223 ( \33566 , \33563 , \33565 );
nand \U$33224 ( \33567 , \33566 , \5034 );
nand \U$33225 ( \33568 , \33562 , \33567 );
not \U$33226 ( \33569 , \33568 );
not \U$33227 ( \33570 , \33569 );
or \U$33228 ( \33571 , \33559 , \33570 );
or \U$33229 ( \33572 , \33569 , \33558 );
nand \U$33230 ( \33573 , \33571 , \33572 );
not \U$33231 ( \33574 , \33573 );
or \U$33232 ( \33575 , \33548 , \33574 );
nand \U$33233 ( \33576 , \33568 , \33558 );
nand \U$33234 ( \33577 , \33575 , \33576 );
xor \U$33235 ( \33578 , \33536 , \33577 );
not \U$33236 ( \33579 , \9249 );
not \U$33237 ( \33580 , RI9872bf8_170);
not \U$33238 ( \33581 , \8857 );
or \U$33239 ( \33582 , \33580 , \33581 );
nand \U$33240 ( \33583 , \9881 , \9185 );
nand \U$33241 ( \33584 , \33582 , \33583 );
not \U$33242 ( \33585 , \33584 );
or \U$33243 ( \33586 , \33579 , \33585 );
nand \U$33244 ( \33587 , \33274 , \22167 );
nand \U$33245 ( \33588 , \33586 , \33587 );
not \U$33246 ( \33589 , \33588 );
and \U$33247 ( \33590 , RI9873030_179, \8053 );
not \U$33248 ( \33591 , RI9873030_179);
and \U$33249 ( \33592 , \33591 , \22516 );
nor \U$33250 ( \33593 , \33590 , \33592 );
not \U$33251 ( \33594 , \33593 );
not \U$33252 ( \33595 , \19320 );
and \U$33253 ( \33596 , \33594 , \33595 );
and \U$33254 ( \33597 , \33113 , \9937 );
nor \U$33255 ( \33598 , \33596 , \33597 );
xor \U$33256 ( \33599 , \33085 , \33096 );
not \U$33257 ( \33600 , \33599 );
and \U$33258 ( \33601 , \33598 , \33600 );
not \U$33259 ( \33602 , \33598 );
and \U$33260 ( \33603 , \33602 , \33599 );
nor \U$33261 ( \33604 , \33601 , \33603 );
not \U$33262 ( \33605 , \33604 );
or \U$33263 ( \33606 , \33589 , \33605 );
not \U$33264 ( \33607 , \33598 );
nand \U$33265 ( \33608 , \33607 , \33599 );
nand \U$33266 ( \33609 , \33606 , \33608 );
and \U$33267 ( \33610 , \33578 , \33609 );
and \U$33268 ( \33611 , \33536 , \33577 );
or \U$33269 ( \33612 , \33610 , \33611 );
not \U$33270 ( \33613 , \33612 );
xor \U$33271 ( \33614 , \32863 , \32852 );
xor \U$33272 ( \33615 , \33614 , \32875 );
not \U$33273 ( \33616 , \33615 );
xor \U$33274 ( \33617 , \33418 , \33411 );
xor \U$33275 ( \33618 , \33617 , \33417 );
not \U$33276 ( \33619 , \33618 );
or \U$33277 ( \33620 , \33616 , \33619 );
or \U$33278 ( \33621 , \33618 , \33615 );
nand \U$33279 ( \33622 , \33620 , \33621 );
not \U$33280 ( \33623 , \33622 );
or \U$33281 ( \33624 , \33613 , \33623 );
not \U$33282 ( \33625 , \33615 );
nand \U$33283 ( \33626 , \33625 , \33618 );
nand \U$33284 ( \33627 , \33624 , \33626 );
and \U$33285 ( \33628 , \33471 , \33627 );
and \U$33286 ( \33629 , \33468 , \33470 );
or \U$33287 ( \33630 , \33628 , \33629 );
not \U$33288 ( \33631 , \33630 );
not \U$33289 ( \33632 , \33631 );
xor \U$33290 ( \33633 , \32559 , \33385 );
xnor \U$33291 ( \33634 , \33633 , \32602 );
not \U$33292 ( \33635 , \33425 );
and \U$33293 ( \33636 , \33634 , \33635 );
not \U$33294 ( \33637 , \33634 );
and \U$33295 ( \33638 , \33637 , \33425 );
nor \U$33296 ( \33639 , \33636 , \33638 );
not \U$33297 ( \33640 , \33639 );
not \U$33298 ( \33641 , \33640 );
or \U$33299 ( \33642 , \33632 , \33641 );
nand \U$33300 ( \33643 , \33639 , \33630 );
nand \U$33301 ( \33644 , \33642 , \33643 );
not \U$33302 ( \33645 , \33644 );
or \U$33303 ( \33646 , \33466 , \33645 );
nand \U$33304 ( \33647 , \33640 , \33630 );
nand \U$33305 ( \33648 , \33646 , \33647 );
not \U$33306 ( \33649 , \33648 );
not \U$33307 ( \33650 , \32808 );
and \U$33308 ( \33651 , \32820 , \33650 );
not \U$33309 ( \33652 , \32820 );
and \U$33310 ( \33653 , \33652 , \32808 );
or \U$33311 ( \33654 , \33651 , \33653 );
not \U$33312 ( \33655 , \33654 );
not \U$33313 ( \33656 , \32878 );
not \U$33314 ( \33657 , \32887 );
not \U$33315 ( \33658 , \33657 );
or \U$33316 ( \33659 , \33656 , \33658 );
not \U$33317 ( \33660 , \32878 );
nand \U$33318 ( \33661 , \33660 , \32887 );
nand \U$33319 ( \33662 , \33659 , \33661 );
not \U$33320 ( \33663 , \33662 );
or \U$33321 ( \33664 , \33655 , \33663 );
or \U$33322 ( \33665 , \33662 , \33654 );
xor \U$33323 ( \33666 , \32985 , \32990 );
xor \U$33324 ( \33667 , \33666 , \33001 );
not \U$33325 ( \33668 , \33667 );
not \U$33326 ( \33669 , \33668 );
xor \U$33327 ( \33670 , \32803 , \32760 );
xor \U$33328 ( \33671 , \33670 , \32752 );
not \U$33329 ( \33672 , \33671 );
and \U$33330 ( \33673 , \32935 , \32946 );
not \U$33331 ( \33674 , \32935 );
and \U$33332 ( \33675 , \33674 , \32947 );
nor \U$33333 ( \33676 , \33673 , \33675 );
xor \U$33334 ( \33677 , \33676 , \32960 );
not \U$33335 ( \33678 , \33677 );
or \U$33336 ( \33679 , \33672 , \33678 );
or \U$33337 ( \33680 , \33677 , \33671 );
nand \U$33338 ( \33681 , \33679 , \33680 );
not \U$33339 ( \33682 , \33681 );
or \U$33340 ( \33683 , \33669 , \33682 );
not \U$33341 ( \33684 , \33671 );
nand \U$33342 ( \33685 , \33684 , \33677 );
nand \U$33343 ( \33686 , \33683 , \33685 );
nand \U$33344 ( \33687 , \33665 , \33686 );
nand \U$33345 ( \33688 , \33664 , \33687 );
nand \U$33346 ( \33689 , \32830 , \32741 );
and \U$33347 ( \33690 , \33689 , \32825 );
not \U$33348 ( \33691 , \33689 );
not \U$33349 ( \33692 , \32825 );
and \U$33350 ( \33693 , \33691 , \33692 );
nor \U$33351 ( \33694 , \33690 , \33693 );
not \U$33352 ( \33695 , \33694 );
or \U$33353 ( \33696 , \33688 , \33695 );
not \U$33354 ( \33697 , \32892 );
not \U$33355 ( \33698 , \33697 );
not \U$33356 ( \33699 , \33015 );
or \U$33357 ( \33700 , \33698 , \33699 );
or \U$33358 ( \33701 , \33015 , \33697 );
nand \U$33359 ( \33702 , \33700 , \33701 );
nand \U$33360 ( \33703 , \33696 , \33702 );
nand \U$33361 ( \33704 , \33688 , \33695 );
and \U$33362 ( \33705 , \33703 , \33704 );
xor \U$33363 ( \33706 , \33427 , \33705 );
xnor \U$33364 ( \33707 , \33706 , \33437 );
not \U$33365 ( \33708 , \33707 );
or \U$33366 ( \33709 , \33649 , \33708 );
not \U$33367 ( \33710 , \33705 );
xor \U$33368 ( \33711 , \33437 , \33427 );
nand \U$33369 ( \33712 , \33710 , \33711 );
nand \U$33370 ( \33713 , \33709 , \33712 );
not \U$33371 ( \33714 , \33713 );
or \U$33372 ( \33715 , \33464 , \33714 );
or \U$33373 ( \33716 , \33713 , \33463 );
nand \U$33374 ( \33717 , \33715 , \33716 );
not \U$33375 ( \33718 , \33717 );
or \U$33376 ( \33719 , \33461 , \33718 );
nand \U$33377 ( \33720 , \33713 , \33462 );
nand \U$33378 ( \33721 , \33719 , \33720 );
not \U$33379 ( \33722 , \32731 );
not \U$33380 ( \33723 , \33446 );
or \U$33381 ( \33724 , \33722 , \33723 );
or \U$33382 ( \33725 , \33446 , \32731 );
nand \U$33383 ( \33726 , \33724 , \33725 );
nor \U$33384 ( \33727 , \33721 , \33726 );
not \U$33385 ( \33728 , \33727 );
xor \U$33386 ( \33729 , \33463 , \33460 );
xnor \U$33387 ( \33730 , \33729 , \33713 );
not \U$33388 ( \33731 , \33654 );
not \U$33389 ( \33732 , \33731 );
not \U$33390 ( \33733 , \33662 );
or \U$33391 ( \33734 , \33732 , \33733 );
or \U$33392 ( \33735 , \33662 , \33731 );
nand \U$33393 ( \33736 , \33734 , \33735 );
not \U$33394 ( \33737 , \33736 );
xor \U$33395 ( \33738 , \33686 , \33737 );
not \U$33396 ( \33739 , \33738 );
not \U$33397 ( \33740 , \33612 );
and \U$33398 ( \33741 , \33622 , \33740 );
not \U$33399 ( \33742 , \33622 );
and \U$33400 ( \33743 , \33742 , \33612 );
nor \U$33401 ( \33744 , \33741 , \33743 );
not \U$33402 ( \33745 , \33744 );
not \U$33403 ( \33746 , \33745 );
not \U$33404 ( \33747 , \33667 );
not \U$33405 ( \33748 , \33681 );
or \U$33406 ( \33749 , \33747 , \33748 );
or \U$33407 ( \33750 , \33681 , \33667 );
nand \U$33408 ( \33751 , \33749 , \33750 );
xor \U$33409 ( \33752 , \33171 , \33204 );
xor \U$33410 ( \33753 , \33752 , \33242 );
xor \U$33411 ( \33754 , \33751 , \33753 );
not \U$33412 ( \33755 , \33754 );
or \U$33413 ( \33756 , \33746 , \33755 );
nand \U$33414 ( \33757 , \33751 , \33753 );
nand \U$33415 ( \33758 , \33756 , \33757 );
not \U$33416 ( \33759 , \33758 );
not \U$33417 ( \33760 , \33759 );
or \U$33418 ( \33761 , \33739 , \33760 );
xor \U$33419 ( \33762 , \33468 , \33470 );
xor \U$33420 ( \33763 , \33762 , \33627 );
nand \U$33421 ( \33764 , \33761 , \33763 );
not \U$33422 ( \33765 , \33738 );
nand \U$33423 ( \33766 , \33765 , \33758 );
nand \U$33424 ( \33767 , \33764 , \33766 );
not \U$33425 ( \33768 , \33767 );
xor \U$33426 ( \33769 , \33170 , \33245 );
xor \U$33427 ( \33770 , \33769 , \33255 );
buf \U$33428 ( \33771 , \33770 );
not \U$33429 ( \33772 , \33771 );
not \U$33430 ( \33773 , \33772 );
xor \U$33431 ( \33774 , \33038 , \33036 );
xnor \U$33432 ( \33775 , \33774 , \33049 );
xor \U$33433 ( \33776 , \33212 , \33228 );
xor \U$33434 ( \33777 , \33776 , \33239 );
xor \U$33435 ( \33778 , \33775 , \33777 );
not \U$33436 ( \33779 , \7326 );
and \U$33437 ( \33780 , \9114 , \7333 );
not \U$33438 ( \33781 , \9114 );
and \U$33439 ( \33782 , \33781 , RI98729a0_165);
nor \U$33440 ( \33783 , \33780 , \33782 );
not \U$33441 ( \33784 , \33783 );
or \U$33442 ( \33785 , \33779 , \33784 );
and \U$33443 ( \33786 , \9850 , \7333 );
not \U$33444 ( \33787 , \9850 );
and \U$33445 ( \33788 , \33787 , RI98729a0_165);
nor \U$33446 ( \33789 , \33786 , \33788 );
nand \U$33447 ( \33790 , \33789 , \7338 );
nand \U$33448 ( \33791 , \33785 , \33790 );
not \U$33449 ( \33792 , \33791 );
not \U$33450 ( \33793 , \33529 );
not \U$33451 ( \33794 , \5653 );
not \U$33452 ( \33795 , \33794 );
and \U$33453 ( \33796 , \33793 , \33795 );
not \U$33454 ( \33797 , RI9872568_156);
not \U$33455 ( \33798 , \13268 );
or \U$33456 ( \33799 , \33797 , \33798 );
or \U$33457 ( \33800 , \25847 , RI9872568_156);
nand \U$33458 ( \33801 , \33799 , \33800 );
and \U$33459 ( \33802 , \33801 , \6063 );
nor \U$33460 ( \33803 , \33796 , \33802 );
xor \U$33461 ( \33804 , \33505 , \33486 );
xnor \U$33462 ( \33805 , \33803 , \33804 );
not \U$33463 ( \33806 , \33805 );
or \U$33464 ( \33807 , \33792 , \33806 );
not \U$33465 ( \33808 , \33803 );
nand \U$33466 ( \33809 , \33808 , \33804 );
nand \U$33467 ( \33810 , \33807 , \33809 );
not \U$33468 ( \33811 , \33810 );
xor \U$33469 ( \33812 , \33520 , \33532 );
buf \U$33470 ( \33813 , \33812 );
not \U$33471 ( \33814 , \33813 );
not \U$33472 ( \33815 , \17371 );
and \U$33473 ( \33816 , RI98733f0_187, \11028 );
not \U$33474 ( \33817 , RI98733f0_187);
and \U$33475 ( \33818 , \33817 , \5599 );
or \U$33476 ( \33819 , \33816 , \33818 );
not \U$33477 ( \33820 , \33819 );
or \U$33478 ( \33821 , \33815 , \33820 );
nand \U$33479 ( \33822 , \33219 , \19282 );
nand \U$33480 ( \33823 , \33821 , \33822 );
not \U$33481 ( \33824 , \33823 );
or \U$33482 ( \33825 , \33814 , \33824 );
or \U$33483 ( \33826 , \33823 , \33813 );
nand \U$33484 ( \33827 , \33825 , \33826 );
not \U$33485 ( \33828 , \33827 );
or \U$33486 ( \33829 , \33811 , \33828 );
not \U$33487 ( \33830 , \33813 );
nand \U$33488 ( \33831 , \33830 , \33823 );
nand \U$33489 ( \33832 , \33829 , \33831 );
and \U$33490 ( \33833 , \33778 , \33832 );
and \U$33491 ( \33834 , \33775 , \33777 );
or \U$33492 ( \33835 , \33833 , \33834 );
not \U$33493 ( \33836 , \33835 );
xnor \U$33494 ( \33837 , \33335 , \33297 );
and \U$33495 ( \33838 , \33283 , \33281 );
not \U$33496 ( \33839 , \33283 );
and \U$33497 ( \33840 , \33839 , \33278 );
nor \U$33498 ( \33841 , \33838 , \33840 );
not \U$33499 ( \33842 , \33295 );
and \U$33500 ( \33843 , \33841 , \33842 );
not \U$33501 ( \33844 , \33841 );
and \U$33502 ( \33845 , \33844 , \33295 );
nor \U$33503 ( \33846 , \33843 , \33845 );
not \U$33504 ( \33847 , \33846 );
not \U$33505 ( \33848 , \33847 );
xor \U$33506 ( \33849 , \33181 , \33189 );
xnor \U$33507 ( \33850 , \33849 , \33200 );
not \U$33508 ( \33851 , \33850 );
or \U$33509 ( \33852 , \33848 , \33851 );
not \U$33510 ( \33853 , \33846 );
not \U$33511 ( \33854 , \33850 );
not \U$33512 ( \33855 , \33854 );
or \U$33513 ( \33856 , \33853 , \33855 );
not \U$33514 ( \33857 , \19046 );
not \U$33515 ( \33858 , \33047 );
or \U$33516 ( \33859 , \33857 , \33858 );
not \U$33517 ( \33860 , \16999 );
not \U$33518 ( \33861 , \3537 );
or \U$33519 ( \33862 , \33860 , \33861 );
or \U$33520 ( \33863 , \16891 , \16999 );
nand \U$33521 ( \33864 , \33862 , \33863 );
nand \U$33522 ( \33865 , \33864 , \24076 );
nand \U$33523 ( \33866 , \33859 , \33865 );
not \U$33524 ( \33867 , \33866 );
nand \U$33525 ( \33868 , \33198 , \17528 );
not \U$33526 ( \33869 , RI9873288_184);
not \U$33527 ( \33870 , \4470 );
or \U$33528 ( \33871 , \33869 , \33870 );
or \U$33529 ( \33872 , \4470 , RI9873288_184);
nand \U$33530 ( \33873 , \33871 , \33872 );
nand \U$33531 ( \33874 , \33873 , \17544 );
nand \U$33532 ( \33875 , \33868 , \33874 );
not \U$33533 ( \33876 , \7338 );
not \U$33534 ( \33877 , \33177 );
or \U$33535 ( \33878 , \33876 , \33877 );
nand \U$33536 ( \33879 , \33789 , \7325 );
nand \U$33537 ( \33880 , \33878 , \33879 );
xor \U$33538 ( \33881 , \33875 , \33880 );
not \U$33539 ( \33882 , \33881 );
or \U$33540 ( \33883 , \33867 , \33882 );
not \U$33541 ( \33884 , \33874 );
not \U$33542 ( \33885 , \33868 );
or \U$33543 ( \33886 , \33884 , \33885 );
nand \U$33544 ( \33887 , \33886 , \33880 );
nand \U$33545 ( \33888 , \33883 , \33887 );
nand \U$33546 ( \33889 , \33856 , \33888 );
nand \U$33547 ( \33890 , \33852 , \33889 );
xnor \U$33548 ( \33891 , \33837 , \33890 );
not \U$33549 ( \33892 , \33891 );
or \U$33550 ( \33893 , \33836 , \33892 );
not \U$33551 ( \33894 , \33837 );
nand \U$33552 ( \33895 , \33894 , \33890 );
nand \U$33553 ( \33896 , \33893 , \33895 );
not \U$33554 ( \33897 , \33896 );
not \U$33555 ( \33898 , \33897 );
or \U$33556 ( \33899 , \33773 , \33898 );
not \U$33557 ( \33900 , \20626 );
not \U$33558 ( \33901 , RI9873558_190);
not \U$33559 ( \33902 , \2947 );
or \U$33560 ( \33903 , \33901 , \33902 );
or \U$33561 ( \33904 , \2947 , RI9873558_190);
nand \U$33562 ( \33905 , \33903 , \33904 );
not \U$33563 ( \33906 , \33905 );
or \U$33564 ( \33907 , \33900 , \33906 );
nand \U$33565 ( \33908 , \33235 , RI9873648_192);
nand \U$33566 ( \33909 , \33907 , \33908 );
not \U$33567 ( \33910 , \33909 );
not \U$33568 ( \33911 , \22618 );
not \U$33569 ( \33912 , \33210 );
or \U$33570 ( \33913 , \33911 , \33912 );
not \U$33571 ( \33914 , \13022 );
not \U$33572 ( \33915 , \6058 );
or \U$33573 ( \33916 , \33914 , \33915 );
or \U$33574 ( \33917 , \6480 , \13022 );
nand \U$33575 ( \33918 , \33916 , \33917 );
nand \U$33576 ( \33919 , \33918 , \24209 );
nand \U$33577 ( \33920 , \33913 , \33919 );
not \U$33578 ( \33921 , \33920 );
buf \U$33579 ( \33922 , \30963 );
nand \U$33580 ( \33923 , \33034 , \33922 );
not \U$33581 ( \33924 , \33923 );
not \U$33582 ( \33925 , RI9873210_183);
not \U$33583 ( \33926 , \24185 );
not \U$33584 ( \33927 , \33926 );
or \U$33585 ( \33928 , \33925 , \33927 );
or \U$33586 ( \33929 , \33926 , RI9873210_183);
nand \U$33587 ( \33930 , \33928 , \33929 );
and \U$33588 ( \33931 , \33930 , \13476 );
nor \U$33589 ( \33932 , \33924 , \33931 );
not \U$33590 ( \33933 , \33932 );
or \U$33591 ( \33934 , \33921 , \33933 );
not \U$33592 ( \33935 , \33931 );
not \U$33593 ( \33936 , \33935 );
not \U$33594 ( \33937 , \33923 );
or \U$33595 ( \33938 , \33936 , \33937 );
not \U$33596 ( \33939 , \33920 );
nand \U$33597 ( \33940 , \33938 , \33939 );
nand \U$33598 ( \33941 , \33934 , \33940 );
not \U$33599 ( \33942 , \33941 );
or \U$33600 ( \33943 , \33910 , \33942 );
not \U$33601 ( \33944 , \33935 );
not \U$33602 ( \33945 , \33923 );
or \U$33603 ( \33946 , \33944 , \33945 );
nand \U$33604 ( \33947 , \33946 , \33920 );
nand \U$33605 ( \33948 , \33943 , \33947 );
not \U$33606 ( \33949 , \33948 );
not \U$33607 ( \33950 , \8028 );
not \U$33608 ( \33951 , RI9872a18_166);
not \U$33609 ( \33952 , \18498 );
or \U$33610 ( \33953 , \33951 , \33952 );
or \U$33611 ( \33954 , \9924 , RI9872a18_166);
nand \U$33612 ( \33955 , \33953 , \33954 );
not \U$33613 ( \33956 , \33955 );
or \U$33614 ( \33957 , \33950 , \33956 );
nand \U$33615 ( \33958 , \33065 , \8041 );
nand \U$33616 ( \33959 , \33957 , \33958 );
not \U$33617 ( \33960 , \33959 );
not \U$33618 ( \33961 , \9214 );
not \U$33619 ( \33962 , \33184 );
or \U$33620 ( \33963 , \33961 , \33962 );
not \U$33621 ( \33964 , \18308 );
not \U$33622 ( \33965 , RI9872b80_169);
and \U$33623 ( \33966 , \33964 , \33965 );
and \U$33624 ( \33967 , \24368 , RI9872b80_169);
nor \U$33625 ( \33968 , \33966 , \33967 );
nand \U$33626 ( \33969 , \33968 , \9196 );
nand \U$33627 ( \33970 , \33963 , \33969 );
not \U$33628 ( \33971 , \4918 );
not \U$33629 ( \33972 , RI9872388_152);
not \U$33630 ( \33973 , \25380 );
or \U$33631 ( \33974 , \33972 , \33973 );
or \U$33632 ( \33975 , \20765 , RI9872388_152);
nand \U$33633 ( \33976 , \33974 , \33975 );
not \U$33634 ( \33977 , \33976 );
or \U$33635 ( \33978 , \33971 , \33977 );
nand \U$33636 ( \33979 , \33556 , \4922 );
nand \U$33637 ( \33980 , \33978 , \33979 );
not \U$33638 ( \33981 , \33980 );
not \U$33639 ( \33982 , \4084 );
not \U$33640 ( \33983 , \33094 );
or \U$33641 ( \33984 , \33982 , \33983 );
not \U$33642 ( \33985 , RI98725e0_157);
buf \U$33643 ( \33986 , \19411 );
not \U$33644 ( \33987 , \33986 );
or \U$33645 ( \33988 , \33985 , \33987 );
or \U$33646 ( \33989 , \33986 , RI98725e0_157);
nand \U$33647 ( \33990 , \33988 , \33989 );
nand \U$33648 ( \33991 , \33990 , \4101 );
nand \U$33649 ( \33992 , \33984 , \33991 );
not \U$33650 ( \33993 , \3169 );
not \U$33651 ( \33994 , \33497 );
or \U$33652 ( \33995 , \33993 , \33994 );
xor \U$33653 ( \33996 , \21779 , RI9872310_151);
nand \U$33654 ( \33997 , \33996 , \3162 );
nand \U$33655 ( \33998 , \33995 , \33997 );
or \U$33656 ( \33999 , RI98726d0_159, RI9872748_160);
nand \U$33657 ( \34000 , \33999 , \24450 );
nand \U$33658 ( \34001 , \34000 , \2975 );
not \U$33659 ( \34002 , \34001 );
and \U$33660 ( \34003 , \33998 , \34002 );
xor \U$33661 ( \34004 , \33992 , \34003 );
not \U$33662 ( \34005 , \34004 );
or \U$33663 ( \34006 , \33981 , \34005 );
nand \U$33664 ( \34007 , \33992 , \34003 );
nand \U$33665 ( \34008 , \34006 , \34007 );
and \U$33666 ( \34009 , \33970 , \34008 );
not \U$33667 ( \34010 , \33970 );
not \U$33668 ( \34011 , \34008 );
and \U$33669 ( \34012 , \34010 , \34011 );
nor \U$33670 ( \34013 , \34009 , \34012 );
not \U$33671 ( \34014 , \34013 );
or \U$33672 ( \34015 , \33960 , \34014 );
nand \U$33673 ( \34016 , \33970 , \34008 );
nand \U$33674 ( \34017 , \34015 , \34016 );
not \U$33675 ( \34018 , \33121 );
not \U$33676 ( \34019 , \33106 );
not \U$33677 ( \34020 , \34019 );
and \U$33678 ( \34021 , \34018 , \34020 );
and \U$33679 ( \34022 , \33121 , \34019 );
nor \U$33680 ( \34023 , \34021 , \34022 );
and \U$33681 ( \34024 , \34017 , \34023 );
not \U$33682 ( \34025 , \34017 );
not \U$33683 ( \34026 , \34023 );
and \U$33684 ( \34027 , \34025 , \34026 );
or \U$33685 ( \34028 , \34024 , \34027 );
not \U$33686 ( \34029 , \34028 );
or \U$33687 ( \34030 , \33949 , \34029 );
nand \U$33688 ( \34031 , \34017 , \34026 );
nand \U$33689 ( \34032 , \34030 , \34031 );
not \U$33690 ( \34033 , \34032 );
not \U$33691 ( \34034 , \33311 );
not \U$33692 ( \34035 , \34034 );
not \U$33693 ( \34036 , \33327 );
or \U$33694 ( \34037 , \34035 , \34036 );
or \U$33695 ( \34038 , \33327 , \34034 );
nand \U$33696 ( \34039 , \34037 , \34038 );
not \U$33697 ( \34040 , \33154 );
xnor \U$33698 ( \34041 , \33158 , \33141 );
not \U$33699 ( \34042 , \34041 );
and \U$33700 ( \34043 , \34040 , \34042 );
buf \U$33701 ( \34044 , \33154 );
and \U$33702 ( \34045 , \34044 , \34041 );
nor \U$33703 ( \34046 , \34043 , \34045 );
xor \U$33704 ( \34047 , \34039 , \34046 );
not \U$33705 ( \34048 , \8752 );
not \U$33706 ( \34049 , \33150 );
or \U$33707 ( \34050 , \34048 , \34049 );
not \U$33708 ( \34051 , RI9872f40_177);
not \U$33709 ( \34052 , \20583 );
or \U$33710 ( \34053 , \34051 , \34052 );
or \U$33711 ( \34054 , \8943 , RI9872f40_177);
nand \U$33712 ( \34055 , \34053 , \34054 );
nand \U$33713 ( \34056 , \34055 , \8743 );
nand \U$33714 ( \34057 , \34050 , \34056 );
not \U$33715 ( \34058 , \34057 );
and \U$33716 ( \34059 , \33293 , \10331 );
xnor \U$33717 ( \34060 , \8333 , RI9872e50_175);
and \U$33718 ( \34061 , \34060 , \9294 );
nor \U$33719 ( \34062 , \34059 , \34061 );
not \U$33720 ( \34063 , \34062 );
not \U$33721 ( \34064 , \33264 );
not \U$33722 ( \34065 , \10624 );
or \U$33723 ( \34066 , \34064 , \34065 );
not \U$33724 ( \34067 , RI9872d60_173);
not \U$33725 ( \34068 , \12712 );
or \U$33726 ( \34069 , \34067 , \34068 );
nand \U$33727 ( \34070 , \29463 , \8807 );
nand \U$33728 ( \34071 , \34069 , \34070 );
nand \U$33729 ( \34072 , \34071 , \8818 );
nand \U$33730 ( \34073 , \34066 , \34072 );
not \U$33731 ( \34074 , \34073 );
or \U$33732 ( \34075 , \34063 , \34074 );
or \U$33733 ( \34076 , \34062 , \34073 );
nand \U$33734 ( \34077 , \34075 , \34076 );
not \U$33735 ( \34078 , \34077 );
or \U$33736 ( \34079 , \34058 , \34078 );
not \U$33737 ( \34080 , \34062 );
nand \U$33738 ( \34081 , \34080 , \34073 );
nand \U$33739 ( \34082 , \34079 , \34081 );
and \U$33740 ( \34083 , \34047 , \34082 );
and \U$33741 ( \34084 , \34039 , \34046 );
or \U$33742 ( \34085 , \34083 , \34084 );
not \U$33743 ( \34086 , \33058 );
not \U$33744 ( \34087 , \34086 );
not \U$33745 ( \34088 , \33166 );
or \U$33746 ( \34089 , \34087 , \34088 );
or \U$33747 ( \34090 , \33166 , \34086 );
nand \U$33748 ( \34091 , \34089 , \34090 );
xor \U$33749 ( \34092 , \34085 , \34091 );
not \U$33750 ( \34093 , \34092 );
or \U$33751 ( \34094 , \34033 , \34093 );
nand \U$33752 ( \34095 , \34091 , \34085 );
nand \U$33753 ( \34096 , \34094 , \34095 );
nand \U$33754 ( \34097 , \33899 , \34096 );
nand \U$33755 ( \34098 , \33896 , \33771 );
nand \U$33756 ( \34099 , \34097 , \34098 );
not \U$33757 ( \34100 , \34099 );
xor \U$33758 ( \34101 , \33694 , \33688 );
xor \U$33759 ( \34102 , \34101 , \33702 );
nand \U$33760 ( \34103 , \34100 , \34102 );
not \U$33761 ( \34104 , \34103 );
or \U$33762 ( \34105 , \33768 , \34104 );
not \U$33763 ( \34106 , \34102 );
nand \U$33764 ( \34107 , \34106 , \34099 );
nand \U$33765 ( \34108 , \34105 , \34107 );
not \U$33766 ( \34109 , \34108 );
not \U$33767 ( \34110 , \33021 );
and \U$33768 ( \34111 , \33360 , \34110 );
not \U$33769 ( \34112 , \33360 );
and \U$33770 ( \34113 , \34112 , \33021 );
nor \U$33771 ( \34114 , \34111 , \34113 );
not \U$33772 ( \34115 , \34114 );
or \U$33773 ( \34116 , \34109 , \34115 );
or \U$33774 ( \34117 , \34108 , \34114 );
nand \U$33775 ( \34118 , \34116 , \34117 );
not \U$33776 ( \34119 , \34118 );
xnor \U$33777 ( \34120 , \33707 , \33648 );
not \U$33778 ( \34121 , \34120 );
not \U$33779 ( \34122 , \34121 );
or \U$33780 ( \34123 , \34119 , \34122 );
not \U$33781 ( \34124 , \34114 );
nand \U$33782 ( \34125 , \34124 , \34108 );
nand \U$33783 ( \34126 , \34123 , \34125 );
nor \U$33784 ( \34127 , \33730 , \34126 );
not \U$33785 ( \34128 , \34127 );
not \U$33786 ( \34129 , \34121 );
not \U$33787 ( \34130 , \34118 );
not \U$33788 ( \34131 , \34130 );
or \U$33789 ( \34132 , \34129 , \34131 );
nand \U$33790 ( \34133 , \34120 , \34118 );
nand \U$33791 ( \34134 , \34132 , \34133 );
not \U$33792 ( \34135 , \9227 );
not \U$33793 ( \34136 , RI9872bf8_170);
not \U$33794 ( \34137 , \8650 );
or \U$33795 ( \34138 , \34136 , \34137 );
or \U$33796 ( \34139 , \11406 , RI9872bf8_170);
nand \U$33797 ( \34140 , \34138 , \34139 );
not \U$33798 ( \34141 , \34140 );
or \U$33799 ( \34142 , \34135 , \34141 );
and \U$33800 ( \34143 , RI9872bf8_170, \8841 );
not \U$33801 ( \34144 , RI9872bf8_170);
and \U$33802 ( \34145 , \34144 , \12848 );
or \U$33803 ( \34146 , \34143 , \34145 );
nand \U$33804 ( \34147 , \34146 , \32292 );
nand \U$33805 ( \34148 , \34142 , \34147 );
not \U$33806 ( \34149 , \34148 );
not \U$33807 ( \34150 , \8801 );
not \U$33808 ( \34151 , RI9872d60_173);
not \U$33809 ( \34152 , \18110 );
or \U$33810 ( \34153 , \34151 , \34152 );
or \U$33811 ( \34154 , \8607 , RI9872d60_173);
nand \U$33812 ( \34155 , \34153 , \34154 );
not \U$33813 ( \34156 , \34155 );
or \U$33814 ( \34157 , \34150 , \34156 );
not \U$33815 ( \34158 , RI9872d60_173);
not \U$33816 ( \34159 , \9880 );
or \U$33817 ( \34160 , \34158 , \34159 );
or \U$33818 ( \34161 , \9880 , RI9872d60_173);
nand \U$33819 ( \34162 , \34160 , \34161 );
nand \U$33820 ( \34163 , \34162 , \22664 );
nand \U$33821 ( \34164 , \34157 , \34163 );
not \U$33822 ( \34165 , \34164 );
or \U$33823 ( \34166 , \34149 , \34165 );
or \U$33824 ( \34167 , \34164 , \34148 );
not \U$33825 ( \34168 , \9214 );
and \U$33826 ( \34169 , \13298 , \11688 );
not \U$33827 ( \34170 , \13298 );
and \U$33828 ( \34171 , \34170 , RI9872b80_169);
nor \U$33829 ( \34172 , \34169 , \34171 );
not \U$33830 ( \34173 , \34172 );
or \U$33831 ( \34174 , \34168 , \34173 );
not \U$33832 ( \34175 , RI9872b80_169);
not \U$33833 ( \34176 , \18498 );
or \U$33834 ( \34177 , \34175 , \34176 );
or \U$33835 ( \34178 , \9924 , RI9872b80_169);
nand \U$33836 ( \34179 , \34177 , \34178 );
nand \U$33837 ( \34180 , \34179 , \9196 );
nand \U$33838 ( \34181 , \34174 , \34180 );
nand \U$33839 ( \34182 , \34167 , \34181 );
nand \U$33840 ( \34183 , \34166 , \34182 );
not \U$33841 ( \34184 , \34183 );
not \U$33842 ( \34185 , \33791 );
not \U$33843 ( \34186 , \34185 );
not \U$33844 ( \34187 , \33805 );
or \U$33845 ( \34188 , \34186 , \34187 );
not \U$33846 ( \34189 , \33805 );
nand \U$33847 ( \34190 , \34189 , \33791 );
nand \U$33848 ( \34191 , \34188 , \34190 );
not \U$33849 ( \34192 , \34191 );
or \U$33850 ( \34193 , \34184 , \34192 );
not \U$33851 ( \34194 , \34191 );
not \U$33852 ( \34195 , \34194 );
not \U$33853 ( \34196 , \34183 );
not \U$33854 ( \34197 , \34196 );
or \U$33855 ( \34198 , \34195 , \34197 );
not \U$33856 ( \34199 , \8039 );
not \U$33857 ( \34200 , \8031 );
not \U$33858 ( \34201 , \18329 );
or \U$33859 ( \34202 , \34200 , \34201 );
or \U$33860 ( \34203 , \9750 , \8031 );
nand \U$33861 ( \34204 , \34202 , \34203 );
not \U$33862 ( \34205 , \34204 );
or \U$33863 ( \34206 , \34199 , \34205 );
xnor \U$33864 ( \34207 , RI9872a18_166, \12460 );
nand \U$33865 ( \34208 , \34207 , \8027 );
nand \U$33866 ( \34209 , \34206 , \34208 );
not \U$33867 ( \34210 , \34209 );
not \U$33868 ( \34211 , \3467 );
and \U$33869 ( \34212 , RI98726d0_159, \18195 );
not \U$33870 ( \34213 , RI98726d0_159);
and \U$33871 ( \34214 , \34213 , \18194 );
nor \U$33872 ( \34215 , \34212 , \34214 );
not \U$33873 ( \34216 , \34215 );
or \U$33874 ( \34217 , \34211 , \34216 );
and \U$33875 ( \34218 , RI98726d0_159, \24450 );
not \U$33876 ( \34219 , RI98726d0_159);
and \U$33877 ( \34220 , \34219 , \24449 );
nor \U$33878 ( \34221 , \34218 , \34220 );
nand \U$33879 ( \34222 , \34221 , \3464 );
nand \U$33880 ( \34223 , \34217 , \34222 );
not \U$33881 ( \34224 , \34223 );
nand \U$33882 ( \34225 , \18704 , \3456 );
nand \U$33883 ( \34226 , \34225 , \3457 , RI98726d0_159);
nor \U$33884 ( \34227 , \34224 , \34226 );
not \U$33885 ( \34228 , \4918 );
not \U$33886 ( \34229 , RI9872388_152);
not \U$33887 ( \34230 , \24470 );
or \U$33888 ( \34231 , \34229 , \34230 );
or \U$33889 ( \34232 , \31875 , RI9872388_152);
nand \U$33890 ( \34233 , \34231 , \34232 );
not \U$33891 ( \34234 , \34233 );
or \U$33892 ( \34235 , \34228 , \34234 );
and \U$33893 ( \34236 , RI9872388_152, \17908 );
not \U$33894 ( \34237 , RI9872388_152);
and \U$33895 ( \34238 , \34237 , \17912 );
or \U$33896 ( \34239 , \34236 , \34238 );
nand \U$33897 ( \34240 , \34239 , \4922 );
nand \U$33898 ( \34241 , \34235 , \34240 );
xor \U$33899 ( \34242 , \34227 , \34241 );
not \U$33900 ( \34243 , \5034 );
not \U$33901 ( \34244 , \5025 );
not \U$33902 ( \34245 , \18713 );
or \U$33903 ( \34246 , \34244 , \34245 );
nand \U$33904 ( \34247 , \25380 , RI9872478_154);
nand \U$33905 ( \34248 , \34246 , \34247 );
not \U$33906 ( \34249 , \34248 );
or \U$33907 ( \34250 , \34243 , \34249 );
and \U$33908 ( \34251 , RI9872478_154, \13860 );
not \U$33909 ( \34252 , RI9872478_154);
and \U$33910 ( \34253 , \34252 , \17883 );
or \U$33911 ( \34254 , \34251 , \34253 );
nand \U$33912 ( \34255 , \34254 , \5035 );
nand \U$33913 ( \34256 , \34250 , \34255 );
and \U$33914 ( \34257 , \34242 , \34256 );
and \U$33915 ( \34258 , \34227 , \34241 );
nor \U$33916 ( \34259 , \34257 , \34258 );
not \U$33917 ( \34260 , \34259 );
or \U$33918 ( \34261 , \34210 , \34260 );
or \U$33919 ( \34262 , \34209 , \34259 );
nand \U$33920 ( \34263 , \34261 , \34262 );
not \U$33921 ( \34264 , \34263 );
not \U$33922 ( \34265 , \12867 );
not \U$33923 ( \34266 , RI98730a8_180);
not \U$33924 ( \34267 , \9556 );
or \U$33925 ( \34268 , \34266 , \34267 );
or \U$33926 ( \34269 , \6308 , RI98730a8_180);
nand \U$33927 ( \34270 , \34268 , \34269 );
not \U$33928 ( \34271 , \34270 );
or \U$33929 ( \34272 , \34265 , \34271 );
not \U$33930 ( \34273 , \13022 );
not \U$33931 ( \34274 , \12802 );
or \U$33932 ( \34275 , \34273 , \34274 );
nand \U$33933 ( \34276 , \8904 , RI98730a8_180);
nand \U$33934 ( \34277 , \34275 , \34276 );
nand \U$33935 ( \34278 , \34277 , \13020 );
nand \U$33936 ( \34279 , \34272 , \34278 );
not \U$33937 ( \34280 , \34279 );
or \U$33938 ( \34281 , \34264 , \34280 );
not \U$33939 ( \34282 , \34259 );
nand \U$33940 ( \34283 , \34282 , \34209 );
nand \U$33941 ( \34284 , \34281 , \34283 );
nand \U$33942 ( \34285 , \34198 , \34284 );
nand \U$33943 ( \34286 , \34193 , \34285 );
not \U$33944 ( \34287 , \34286 );
xor \U$33945 ( \34288 , \33812 , \33810 );
xor \U$33946 ( \34289 , \34288 , \33823 );
not \U$33947 ( \34290 , \34289 );
not \U$33948 ( \34291 , \34290 );
or \U$33949 ( \34292 , \34287 , \34291 );
not \U$33950 ( \34293 , \34286 );
not \U$33951 ( \34294 , \34293 );
not \U$33952 ( \34295 , \34289 );
or \U$33953 ( \34296 , \34294 , \34295 );
not \U$33954 ( \34297 , \11198 );
not \U$33955 ( \34298 , \34055 );
or \U$33956 ( \34299 , \34297 , \34298 );
not \U$33957 ( \34300 , RI9872f40_177);
not \U$33958 ( \34301 , \13824 );
or \U$33959 ( \34302 , \34300 , \34301 );
or \U$33960 ( \34303 , \21642 , RI9872f40_177);
nand \U$33961 ( \34304 , \34302 , \34303 );
nand \U$33962 ( \34305 , \34304 , \9526 );
nand \U$33963 ( \34306 , \34299 , \34305 );
not \U$33964 ( \34307 , \34306 );
not \U$33965 ( \34308 , \5632 );
not \U$33966 ( \34309 , \13876 );
or \U$33967 ( \34310 , \34308 , \34309 );
not \U$33968 ( \34311 , \13387 );
nand \U$33969 ( \34312 , \34311 , RI98728b0_163);
nand \U$33970 ( \34313 , \34310 , \34312 );
nand \U$33971 ( \34314 , \34313 , \6282 );
nand \U$33972 ( \34315 , \33543 , \6285 );
nand \U$33973 ( \34316 , \34314 , \34315 );
not \U$33974 ( \34317 , \5035 );
not \U$33975 ( \34318 , \33566 );
or \U$33976 ( \34319 , \34317 , \34318 );
not \U$33977 ( \34320 , \17783 );
xor \U$33978 ( \34321 , RI9872478_154, \34320 );
nand \U$33979 ( \34322 , \34321 , \5034 );
nand \U$33980 ( \34323 , \34319 , \34322 );
xor \U$33981 ( \34324 , \34316 , \34323 );
not \U$33982 ( \34325 , \34324 );
and \U$33983 ( \34326 , \34307 , \34325 );
and \U$33984 ( \34327 , \34306 , \34324 );
nor \U$33985 ( \34328 , \34326 , \34327 );
not \U$33986 ( \34329 , \34328 );
not \U$33987 ( \34330 , \5653 );
not \U$33988 ( \34331 , \33801 );
or \U$33989 ( \34332 , \34330 , \34331 );
and \U$33990 ( \34333 , RI9872568_156, \19591 );
not \U$33991 ( \34334 , RI9872568_156);
and \U$33992 ( \34335 , \34334 , \13281 );
or \U$33993 ( \34336 , \34333 , \34335 );
nand \U$33994 ( \34337 , \34336 , \5641 );
nand \U$33995 ( \34338 , \34332 , \34337 );
not \U$33996 ( \34339 , \34338 );
not \U$33997 ( \34340 , \5035 );
not \U$33998 ( \34341 , \34321 );
or \U$33999 ( \34342 , \34340 , \34341 );
nand \U$34000 ( \34343 , \34254 , \5034 );
nand \U$34001 ( \34344 , \34342 , \34343 );
not \U$34002 ( \34345 , \34344 );
or \U$34003 ( \34346 , \34339 , \34345 );
not \U$34004 ( \34347 , \6285 );
not \U$34005 ( \34348 , \34313 );
or \U$34006 ( \34349 , \34347 , \34348 );
and \U$34007 ( \34350 , RI98728b0_163, \21393 );
not \U$34008 ( \34351 , RI98728b0_163);
and \U$34009 ( \34352 , \34351 , \11454 );
or \U$34010 ( \34353 , \34350 , \34352 );
nand \U$34011 ( \34354 , \34353 , \6282 );
nand \U$34012 ( \34355 , \34349 , \34354 );
not \U$34013 ( \34356 , \34355 );
not \U$34014 ( \34357 , \34344 );
and \U$34015 ( \34358 , \34338 , \34357 );
not \U$34016 ( \34359 , \34338 );
and \U$34017 ( \34360 , \34359 , \34344 );
nor \U$34018 ( \34361 , \34358 , \34360 );
or \U$34019 ( \34362 , \34356 , \34361 );
nand \U$34020 ( \34363 , \34346 , \34362 );
not \U$34021 ( \34364 , \34363 );
or \U$34022 ( \34365 , \34329 , \34364 );
not \U$34023 ( \34366 , \34363 );
not \U$34024 ( \34367 , \34366 );
not \U$34025 ( \34368 , \34328 );
not \U$34026 ( \34369 , \34368 );
or \U$34027 ( \34370 , \34367 , \34369 );
not \U$34028 ( \34371 , \24627 );
and \U$34029 ( \34372 , RI9872f40_177, \12727 );
not \U$34030 ( \34373 , RI9872f40_177);
and \U$34031 ( \34374 , \34373 , \8334 );
nor \U$34032 ( \34375 , \34372 , \34374 );
not \U$34033 ( \34376 , \34375 );
or \U$34034 ( \34377 , \34371 , \34376 );
nand \U$34035 ( \34378 , \34304 , \11198 );
nand \U$34036 ( \34379 , \34377 , \34378 );
not \U$34037 ( \34380 , \34379 );
not \U$34038 ( \34381 , \9272 );
not \U$34039 ( \34382 , RI9872e50_175);
not \U$34040 ( \34383 , \21518 );
or \U$34041 ( \34384 , \34382 , \34383 );
or \U$34042 ( \34385 , \8074 , RI9872e50_175);
nand \U$34043 ( \34386 , \34384 , \34385 );
not \U$34044 ( \34387 , \34386 );
or \U$34045 ( \34388 , \34381 , \34387 );
and \U$34046 ( \34389 , RI9872e50_175, \8877 );
not \U$34047 ( \34390 , RI9872e50_175);
and \U$34048 ( \34391 , \34390 , \8620 );
nor \U$34049 ( \34392 , \34389 , \34391 );
nand \U$34050 ( \34393 , \34392 , \9293 );
nand \U$34051 ( \34394 , \34388 , \34393 );
and \U$34052 ( \34395 , \33998 , \34001 );
not \U$34053 ( \34396 , \33998 );
and \U$34054 ( \34397 , \34396 , \34002 );
nor \U$34055 ( \34398 , \34395 , \34397 );
not \U$34056 ( \34399 , \34398 );
not \U$34057 ( \34400 , \34399 );
not \U$34058 ( \34401 , \3467 );
not \U$34059 ( \34402 , \33484 );
or \U$34060 ( \34403 , \34401 , \34402 );
not \U$34061 ( \34404 , \4063 );
not \U$34062 ( \34405 , \17862 );
or \U$34063 ( \34406 , \34404 , \34405 );
not \U$34064 ( \34407 , \17862 );
not \U$34065 ( \34408 , \34407 );
or \U$34066 ( \34409 , \34408 , \4063 );
nand \U$34067 ( \34410 , \34406 , \34409 );
nand \U$34068 ( \34411 , \34410 , \3464 );
nand \U$34069 ( \34412 , \34403 , \34411 );
not \U$34070 ( \34413 , \34412 );
not \U$34071 ( \34414 , \34413 );
or \U$34072 ( \34415 , \34400 , \34414 );
nand \U$34073 ( \34416 , \34398 , \34412 );
nand \U$34074 ( \34417 , \34415 , \34416 );
not \U$34075 ( \34418 , \33990 );
or \U$34076 ( \34419 , \34418 , \31176 );
and \U$34077 ( \34420 , RI98725e0_157, \19519 );
not \U$34078 ( \34421 , RI98725e0_157);
and \U$34079 ( \34422 , \34421 , \18216 );
nor \U$34080 ( \34423 , \34420 , \34422 );
not \U$34081 ( \34424 , \34423 );
or \U$34082 ( \34425 , \34424 , \4102 );
nand \U$34083 ( \34426 , \34419 , \34425 );
xnor \U$34084 ( \34427 , \34417 , \34426 );
not \U$34085 ( \34428 , \34427 );
and \U$34086 ( \34429 , \34394 , \34428 );
not \U$34087 ( \34430 , \34394 );
and \U$34088 ( \34431 , \34430 , \34427 );
nor \U$34089 ( \34432 , \34429 , \34431 );
not \U$34090 ( \34433 , \34432 );
or \U$34091 ( \34434 , \34380 , \34433 );
nand \U$34092 ( \34435 , \34394 , \34428 );
nand \U$34093 ( \34436 , \34434 , \34435 );
nand \U$34094 ( \34437 , \34370 , \34436 );
nand \U$34095 ( \34438 , \34365 , \34437 );
nand \U$34096 ( \34439 , \34296 , \34438 );
nand \U$34097 ( \34440 , \34292 , \34439 );
not \U$34098 ( \34441 , \34440 );
and \U$34099 ( \34442 , \34028 , \33948 );
not \U$34100 ( \34443 , \34028 );
not \U$34101 ( \34444 , \33948 );
and \U$34102 ( \34445 , \34443 , \34444 );
nor \U$34103 ( \34446 , \34442 , \34445 );
not \U$34104 ( \34447 , \34446 );
not \U$34105 ( \34448 , \34447 );
not \U$34106 ( \34449 , \33847 );
not \U$34107 ( \34450 , \33854 );
or \U$34108 ( \34451 , \34449 , \34450 );
nand \U$34109 ( \34452 , \33850 , \33846 );
nand \U$34110 ( \34453 , \34451 , \34452 );
not \U$34111 ( \34454 , \33888 );
and \U$34112 ( \34455 , \34453 , \34454 );
not \U$34113 ( \34456 , \34453 );
and \U$34114 ( \34457 , \34456 , \33888 );
nor \U$34115 ( \34458 , \34455 , \34457 );
not \U$34116 ( \34459 , \34458 );
not \U$34117 ( \34460 , \34459 );
or \U$34118 ( \34461 , \34448 , \34460 );
nand \U$34119 ( \34462 , \34446 , \34458 );
nand \U$34120 ( \34463 , \34461 , \34462 );
not \U$34121 ( \34464 , \34463 );
or \U$34122 ( \34465 , \34441 , \34464 );
nand \U$34123 ( \34466 , \34459 , \34446 );
nand \U$34124 ( \34467 , \34465 , \34466 );
not \U$34125 ( \34468 , \34467 );
not \U$34126 ( \34469 , \33754 );
not \U$34127 ( \34470 , \33744 );
and \U$34128 ( \34471 , \34469 , \34470 );
and \U$34129 ( \34472 , \33754 , \33744 );
nor \U$34130 ( \34473 , \34471 , \34472 );
not \U$34131 ( \34474 , \34473 );
not \U$34132 ( \34475 , \34474 );
or \U$34133 ( \34476 , \34468 , \34475 );
not \U$34134 ( \34477 , \34467 );
not \U$34135 ( \34478 , \34477 );
not \U$34136 ( \34479 , \34473 );
or \U$34137 ( \34480 , \34478 , \34479 );
not \U$34138 ( \34481 , \17263 );
not \U$34139 ( \34482 , \33819 );
or \U$34140 ( \34483 , \34481 , \34482 );
and \U$34141 ( \34484 , RI98733f0_187, \5206 );
not \U$34142 ( \34485 , RI98733f0_187);
and \U$34143 ( \34486 , \34485 , \17799 );
or \U$34144 ( \34487 , \34484 , \34486 );
nand \U$34145 ( \34488 , \34487 , \17371 );
nand \U$34146 ( \34489 , \34483 , \34488 );
not \U$34147 ( \34490 , \34489 );
not \U$34148 ( \34491 , \4922 );
not \U$34149 ( \34492 , \33976 );
or \U$34150 ( \34493 , \34491 , \34492 );
nand \U$34151 ( \34494 , \34239 , \4918 );
nand \U$34152 ( \34495 , \34493 , \34494 );
not \U$34153 ( \34496 , \34495 );
and \U$34154 ( \34497 , \27523 , \3169 );
not \U$34155 ( \34498 , \3467 );
not \U$34156 ( \34499 , \34410 );
or \U$34157 ( \34500 , \34498 , \34499 );
nand \U$34158 ( \34501 , \34215 , \3464 );
nand \U$34159 ( \34502 , \34500 , \34501 );
xor \U$34160 ( \34503 , \34497 , \34502 );
not \U$34161 ( \34504 , \4084 );
not \U$34162 ( \34505 , \34423 );
or \U$34163 ( \34506 , \34504 , \34505 );
xor \U$34164 ( \34507 , RI98725e0_157, \17702 );
nand \U$34165 ( \34508 , \34507 , \4101 );
nand \U$34166 ( \34509 , \34506 , \34508 );
and \U$34167 ( \34510 , \34503 , \34509 );
and \U$34168 ( \34511 , \34497 , \34502 );
nor \U$34169 ( \34512 , \34510 , \34511 );
not \U$34170 ( \34513 , \34512 );
and \U$34171 ( \34514 , \34496 , \34513 );
and \U$34172 ( \34515 , \34495 , \34512 );
nor \U$34173 ( \34516 , \34514 , \34515 );
not \U$34174 ( \34517 , \34516 );
not \U$34175 ( \34518 , \34517 );
not \U$34176 ( \34519 , \7338 );
not \U$34177 ( \34520 , \33783 );
or \U$34178 ( \34521 , \34519 , \34520 );
not \U$34179 ( \34522 , \7333 );
not \U$34180 ( \34523 , \12594 );
or \U$34181 ( \34524 , \34522 , \34523 );
nand \U$34182 ( \34525 , \12597 , RI98729a0_165);
nand \U$34183 ( \34526 , \34524 , \34525 );
nand \U$34184 ( \34527 , \34526 , \7325 );
nand \U$34185 ( \34528 , \34521 , \34527 );
not \U$34186 ( \34529 , \34528 );
or \U$34187 ( \34530 , \34518 , \34529 );
not \U$34188 ( \34531 , \34512 );
nand \U$34189 ( \34532 , \34531 , \34495 );
nand \U$34190 ( \34533 , \34530 , \34532 );
not \U$34191 ( \34534 , RI9873648_192);
not \U$34192 ( \34535 , \33905 );
or \U$34193 ( \34536 , \34534 , \34535 );
not \U$34194 ( \34537 , RI9873558_190);
not \U$34195 ( \34538 , \3859 );
or \U$34196 ( \34539 , \34537 , \34538 );
or \U$34197 ( \34540 , \3859 , RI9873558_190);
nand \U$34198 ( \34541 , \34539 , \34540 );
nand \U$34199 ( \34542 , \34541 , \18615 );
nand \U$34200 ( \34543 , \34536 , \34542 );
xor \U$34201 ( \34544 , \34533 , \34543 );
not \U$34202 ( \34545 , \34544 );
or \U$34203 ( \34546 , \34490 , \34545 );
nand \U$34204 ( \34547 , \34543 , \34533 );
nand \U$34205 ( \34548 , \34546 , \34547 );
not \U$34206 ( \34549 , \34548 );
not \U$34207 ( \34550 , \33866 );
xor \U$34208 ( \34551 , \34550 , \33881 );
xor \U$34209 ( \34552 , \33909 , \33941 );
xnor \U$34210 ( \34553 , \34551 , \34552 );
not \U$34211 ( \34554 , \34553 );
or \U$34212 ( \34555 , \34549 , \34554 );
nand \U$34213 ( \34556 , \33881 , \34550 );
not \U$34214 ( \34557 , \34556 );
not \U$34215 ( \34558 , \33881 );
nand \U$34216 ( \34559 , \34558 , \33866 );
not \U$34217 ( \34560 , \34559 );
or \U$34218 ( \34561 , \34557 , \34560 );
nand \U$34219 ( \34562 , \34561 , \34552 );
nand \U$34220 ( \34563 , \34555 , \34562 );
not \U$34221 ( \34564 , \34563 );
not \U$34222 ( \34565 , \22167 );
not \U$34223 ( \34566 , \33584 );
or \U$34224 ( \34567 , \34565 , \34566 );
nand \U$34225 ( \34568 , \34140 , \9249 );
nand \U$34226 ( \34569 , \34567 , \34568 );
not \U$34227 ( \34570 , \9293 );
not \U$34228 ( \34571 , \34386 );
or \U$34229 ( \34572 , \34570 , \34571 );
nand \U$34230 ( \34573 , \34060 , \9272 );
nand \U$34231 ( \34574 , \34572 , \34573 );
nor \U$34232 ( \34575 , \34569 , \34574 );
not \U$34233 ( \34576 , \8819 );
not \U$34234 ( \34577 , \34155 );
or \U$34235 ( \34578 , \34576 , \34577 );
nand \U$34236 ( \34579 , \34071 , \10624 );
nand \U$34237 ( \34580 , \34578 , \34579 );
not \U$34238 ( \34581 , \34580 );
or \U$34239 ( \34582 , \34575 , \34581 );
nand \U$34240 ( \34583 , \34569 , \34574 );
nand \U$34241 ( \34584 , \34582 , \34583 );
not \U$34242 ( \34585 , \34584 );
xor \U$34243 ( \34586 , \33588 , \34585 );
xnor \U$34244 ( \34587 , \34586 , \33604 );
and \U$34245 ( \34588 , \34077 , \34057 );
not \U$34246 ( \34589 , \34077 );
not \U$34247 ( \34590 , \34057 );
and \U$34248 ( \34591 , \34589 , \34590 );
nor \U$34249 ( \34592 , \34588 , \34591 );
nand \U$34250 ( \34593 , \34587 , \34592 );
not \U$34251 ( \34594 , \33588 );
and \U$34252 ( \34595 , \33604 , \34594 );
not \U$34253 ( \34596 , \33604 );
and \U$34254 ( \34597 , \34596 , \33588 );
or \U$34255 ( \34598 , \34595 , \34597 );
not \U$34256 ( \34599 , \34585 );
nand \U$34257 ( \34600 , \34598 , \34599 );
nand \U$34258 ( \34601 , \34593 , \34600 );
not \U$34259 ( \34602 , \19036 );
not \U$34260 ( \34603 , RI98734e0_189);
not \U$34261 ( \34604 , \11672 );
or \U$34262 ( \34605 , \34603 , \34604 );
or \U$34263 ( \34606 , \3568 , RI98734e0_189);
nand \U$34264 ( \34607 , \34605 , \34606 );
not \U$34265 ( \34608 , \34607 );
or \U$34266 ( \34609 , \34602 , \34608 );
nand \U$34267 ( \34610 , \33864 , \20147 );
nand \U$34268 ( \34611 , \34609 , \34610 );
not \U$34269 ( \34612 , \34611 );
not \U$34270 ( \34613 , \13484 );
not \U$34271 ( \34614 , \33930 );
or \U$34272 ( \34615 , \34613 , \34614 );
not \U$34273 ( \34616 , RI9873210_183);
not \U$34274 ( \34617 , \5775 );
or \U$34275 ( \34618 , \34616 , \34617 );
or \U$34276 ( \34619 , \5775 , RI9873210_183);
nand \U$34277 ( \34620 , \34618 , \34619 );
nand \U$34278 ( \34621 , \34620 , \13475 );
nand \U$34279 ( \34622 , \34615 , \34621 );
not \U$34280 ( \34623 , \34622 );
xnor \U$34281 ( \34624 , \33980 , \34004 );
not \U$34282 ( \34625 , \34624 );
and \U$34283 ( \34626 , \34623 , \34625 );
and \U$34284 ( \34627 , \34622 , \34624 );
nor \U$34285 ( \34628 , \34626 , \34627 );
not \U$34286 ( \34629 , \34628 );
not \U$34287 ( \34630 , \34629 );
or \U$34288 ( \34631 , \34612 , \34630 );
not \U$34289 ( \34632 , \34624 );
nand \U$34290 ( \34633 , \34632 , \34622 );
nand \U$34291 ( \34634 , \34631 , \34633 );
not \U$34292 ( \34635 , \34634 );
not \U$34293 ( \34636 , \18672 );
not \U$34294 ( \34637 , \14132 );
not \U$34295 ( \34638 , \18793 );
or \U$34296 ( \34639 , \34637 , \34638 );
or \U$34297 ( \34640 , \7905 , \14132 );
nand \U$34298 ( \34641 , \34639 , \34640 );
not \U$34299 ( \34642 , \34641 );
or \U$34300 ( \34643 , \34636 , \34642 );
not \U$34301 ( \34644 , \33593 );
nand \U$34302 ( \34645 , \34644 , \9937 );
nand \U$34303 ( \34646 , \34643 , \34645 );
not \U$34304 ( \34647 , \34646 );
not \U$34305 ( \34648 , \29633 );
not \U$34306 ( \34649 , \34270 );
or \U$34307 ( \34650 , \34648 , \34649 );
nand \U$34308 ( \34651 , \33918 , \22618 );
nand \U$34309 ( \34652 , \34650 , \34651 );
not \U$34310 ( \34653 , \34652 );
or \U$34311 ( \34654 , \34647 , \34653 );
or \U$34312 ( \34655 , \34652 , \34646 );
not \U$34313 ( \34656 , \19641 );
and \U$34314 ( \34657 , RI9873288_184, \4960 );
not \U$34315 ( \34658 , RI9873288_184);
and \U$34316 ( \34659 , \34658 , \23391 );
nor \U$34317 ( \34660 , \34657 , \34659 );
not \U$34318 ( \34661 , \34660 );
or \U$34319 ( \34662 , \34656 , \34661 );
nand \U$34320 ( \34663 , \33873 , \17528 );
nand \U$34321 ( \34664 , \34662 , \34663 );
nand \U$34322 ( \34665 , \34655 , \34664 );
nand \U$34323 ( \34666 , \34654 , \34665 );
not \U$34324 ( \34667 , \34666 );
xor \U$34325 ( \34668 , \34011 , \33959 );
xor \U$34326 ( \34669 , \34668 , \33970 );
not \U$34327 ( \34670 , \34669 );
or \U$34328 ( \34671 , \34667 , \34670 );
or \U$34329 ( \34672 , \34669 , \34666 );
nand \U$34330 ( \34673 , \34671 , \34672 );
not \U$34331 ( \34674 , \34673 );
or \U$34332 ( \34675 , \34635 , \34674 );
not \U$34333 ( \34676 , \34669 );
nand \U$34334 ( \34677 , \34676 , \34666 );
nand \U$34335 ( \34678 , \34675 , \34677 );
xor \U$34336 ( \34679 , \34601 , \34678 );
not \U$34337 ( \34680 , \34679 );
or \U$34338 ( \34681 , \34564 , \34680 );
not \U$34339 ( \34682 , \34600 );
not \U$34340 ( \34683 , \34593 );
or \U$34341 ( \34684 , \34682 , \34683 );
nand \U$34342 ( \34685 , \34684 , \34678 );
nand \U$34343 ( \34686 , \34681 , \34685 );
nand \U$34344 ( \34687 , \34480 , \34686 );
nand \U$34345 ( \34688 , \34476 , \34687 );
not \U$34346 ( \34689 , \34688 );
xor \U$34347 ( \34690 , \33770 , \34096 );
xor \U$34348 ( \34691 , \34690 , \33897 );
not \U$34349 ( \34692 , \34691 );
not \U$34350 ( \34693 , \34692 );
or \U$34351 ( \34694 , \34689 , \34693 );
not \U$34352 ( \34695 , \34691 );
not \U$34353 ( \34696 , \34688 );
not \U$34354 ( \34697 , \34696 );
or \U$34355 ( \34698 , \34695 , \34697 );
xnor \U$34356 ( \34699 , \33891 , \33835 );
not \U$34357 ( \34700 , \34699 );
not \U$34358 ( \34701 , \34700 );
not \U$34359 ( \34702 , \8041 );
not \U$34360 ( \34703 , \33955 );
or \U$34361 ( \34704 , \34702 , \34703 );
nand \U$34362 ( \34705 , \34204 , \8028 );
nand \U$34363 ( \34706 , \34704 , \34705 );
not \U$34364 ( \34707 , \34706 );
nand \U$34365 ( \34708 , \34417 , \34426 );
nand \U$34366 ( \34709 , \34399 , \34412 );
and \U$34367 ( \34710 , \34708 , \34709 );
not \U$34368 ( \34711 , \34710 );
not \U$34369 ( \34712 , \9196 );
not \U$34370 ( \34713 , \34172 );
or \U$34371 ( \34714 , \34712 , \34713 );
nand \U$34372 ( \34715 , \33968 , \9214 );
nand \U$34373 ( \34716 , \34714 , \34715 );
not \U$34374 ( \34717 , \34716 );
or \U$34375 ( \34718 , \34711 , \34717 );
or \U$34376 ( \34719 , \34716 , \34710 );
nand \U$34377 ( \34720 , \34718 , \34719 );
not \U$34378 ( \34721 , \34720 );
or \U$34379 ( \34722 , \34707 , \34721 );
not \U$34380 ( \34723 , \34710 );
nand \U$34381 ( \34724 , \34723 , \34716 );
nand \U$34382 ( \34725 , \34722 , \34724 );
not \U$34383 ( \34726 , \34725 );
not \U$34384 ( \34727 , \33547 );
not \U$34385 ( \34728 , \34727 );
not \U$34386 ( \34729 , \33573 );
or \U$34387 ( \34730 , \34728 , \34729 );
or \U$34388 ( \34731 , \33573 , \34727 );
nand \U$34389 ( \34732 , \34730 , \34731 );
not \U$34390 ( \34733 , \34732 );
not \U$34391 ( \34734 , \34323 );
nand \U$34392 ( \34735 , \34734 , \34314 , \34315 );
not \U$34393 ( \34736 , \34735 );
not \U$34394 ( \34737 , \34306 );
or \U$34395 ( \34738 , \34736 , \34737 );
nand \U$34396 ( \34739 , \34316 , \34323 );
nand \U$34397 ( \34740 , \34738 , \34739 );
not \U$34398 ( \34741 , \34740 );
not \U$34399 ( \34742 , \34741 );
or \U$34400 ( \34743 , \34733 , \34742 );
not \U$34401 ( \34744 , \34732 );
nand \U$34402 ( \34745 , \34744 , \34740 );
nand \U$34403 ( \34746 , \34743 , \34745 );
not \U$34404 ( \34747 , \34746 );
or \U$34405 ( \34748 , \34726 , \34747 );
nand \U$34406 ( \34749 , \34740 , \34732 );
nand \U$34407 ( \34750 , \34748 , \34749 );
xor \U$34408 ( \34751 , \34039 , \34046 );
xor \U$34409 ( \34752 , \34751 , \34082 );
xor \U$34410 ( \34753 , \34750 , \34752 );
xor \U$34411 ( \34754 , \33536 , \33577 );
xor \U$34412 ( \34755 , \34754 , \33609 );
and \U$34413 ( \34756 , \34753 , \34755 );
and \U$34414 ( \34757 , \34750 , \34752 );
or \U$34415 ( \34758 , \34756 , \34757 );
not \U$34416 ( \34759 , \34758 );
not \U$34417 ( \34760 , \34032 );
not \U$34418 ( \34761 , \34760 );
not \U$34419 ( \34762 , \34092 );
or \U$34420 ( \34763 , \34761 , \34762 );
or \U$34421 ( \34764 , \34092 , \34760 );
nand \U$34422 ( \34765 , \34763 , \34764 );
not \U$34423 ( \34766 , \34765 );
not \U$34424 ( \34767 , \34766 );
or \U$34425 ( \34768 , \34759 , \34767 );
not \U$34426 ( \34769 , \34758 );
nand \U$34427 ( \34770 , \34769 , \34765 );
nand \U$34428 ( \34771 , \34768 , \34770 );
not \U$34429 ( \34772 , \34771 );
or \U$34430 ( \34773 , \34701 , \34772 );
nand \U$34431 ( \34774 , \34765 , \34758 );
nand \U$34432 ( \34775 , \34773 , \34774 );
nand \U$34433 ( \34776 , \34698 , \34775 );
nand \U$34434 ( \34777 , \34694 , \34776 );
buf \U$34435 ( \34778 , \34777 );
not \U$34436 ( \34779 , \33465 );
and \U$34437 ( \34780 , \33644 , \34779 );
not \U$34438 ( \34781 , \33644 );
and \U$34439 ( \34782 , \34781 , \33465 );
nor \U$34440 ( \34783 , \34780 , \34782 );
not \U$34441 ( \34784 , \34783 );
nor \U$34442 ( \34785 , \34778 , \34784 );
nand \U$34443 ( \34786 , \34107 , \34103 );
and \U$34444 ( \34787 , \34786 , \33767 );
not \U$34445 ( \34788 , \34786 );
not \U$34446 ( \34789 , \33767 );
and \U$34447 ( \34790 , \34788 , \34789 );
nor \U$34448 ( \34791 , \34787 , \34790 );
or \U$34449 ( \34792 , \34785 , \34791 );
nand \U$34450 ( \34793 , \34778 , \34784 );
nand \U$34451 ( \34794 , \34792 , \34793 );
or \U$34452 ( \34795 , \34134 , \34794 );
and \U$34453 ( \34796 , \33455 , \33728 , \34128 , \34795 );
not \U$34454 ( \34797 , \32687 );
not \U$34455 ( \34798 , \32128 );
not \U$34456 ( \34799 , \32723 );
or \U$34457 ( \34800 , \34798 , \34799 );
or \U$34458 ( \34801 , \32723 , \32128 );
nand \U$34459 ( \34802 , \34800 , \34801 );
not \U$34460 ( \34803 , \34802 );
or \U$34461 ( \34804 , \34797 , \34803 );
not \U$34462 ( \34805 , \32128 );
nand \U$34463 ( \34806 , \34805 , \32724 );
nand \U$34464 ( \34807 , \34804 , \34806 );
buf \U$34465 ( \34808 , \34807 );
xor \U$34466 ( \34809 , \31366 , \31375 );
xor \U$34467 ( \34810 , \34809 , \31682 );
not \U$34468 ( \34811 , \34810 );
not \U$34469 ( \34812 , \32695 );
not \U$34470 ( \34813 , \32717 );
or \U$34471 ( \34814 , \34812 , \34813 );
not \U$34472 ( \34815 , \32712 );
nand \U$34473 ( \34816 , \34815 , \32700 );
nand \U$34474 ( \34817 , \34814 , \34816 );
not \U$34475 ( \34818 , \34817 );
not \U$34476 ( \34819 , \34818 );
or \U$34477 ( \34820 , \34811 , \34819 );
not \U$34478 ( \34821 , \34810 );
nand \U$34479 ( \34822 , \34821 , \34817 );
nand \U$34480 ( \34823 , \34820 , \34822 );
buf \U$34481 ( \34824 , \31771 );
buf \U$34482 ( \34825 , \32099 );
xor \U$34483 ( \34826 , \34824 , \34825 );
xor \U$34484 ( \34827 , \34823 , \34826 );
buf \U$34485 ( \34828 , \34827 );
nor \U$34486 ( \34829 , \34808 , \34828 );
not \U$34487 ( \34830 , \34826 );
not \U$34488 ( \34831 , \34823 );
or \U$34489 ( \34832 , \34830 , \34831 );
nand \U$34490 ( \34833 , \34817 , \34810 );
nand \U$34491 ( \34834 , \34832 , \34833 );
not \U$34492 ( \34835 , \31715 );
not \U$34493 ( \34836 , \32112 );
or \U$34494 ( \34837 , \34835 , \34836 );
or \U$34495 ( \34838 , \32112 , \31715 );
nand \U$34496 ( \34839 , \34837 , \34838 );
nor \U$34497 ( \34840 , \34834 , \34839 );
nor \U$34498 ( \34841 , \34829 , \34840 );
and \U$34499 ( \34842 , \32121 , \34796 , \34841 );
not \U$34500 ( \34843 , \7326 );
and \U$34501 ( \34844 , \17783 , \7333 );
not \U$34502 ( \34845 , \17783 );
and \U$34503 ( \34846 , \34845 , RI98729a0_165);
nor \U$34504 ( \34847 , \34844 , \34846 );
not \U$34505 ( \34848 , \34847 );
or \U$34506 ( \34849 , \34843 , \34848 );
not \U$34507 ( \34850 , RI98729a0_165);
not \U$34508 ( \34851 , \24523 );
or \U$34509 ( \34852 , \34850 , \34851 );
or \U$34510 ( \34853 , \24523 , RI98729a0_165);
nand \U$34511 ( \34854 , \34852 , \34853 );
nand \U$34512 ( \34855 , \34854 , \7338 );
nand \U$34513 ( \34856 , \34849 , \34855 );
not \U$34514 ( \34857 , \9214 );
and \U$34515 ( \34858 , RI9872b80_169, \12597 );
not \U$34516 ( \34859 , RI9872b80_169);
and \U$34517 ( \34860 , \34859 , \12594 );
or \U$34518 ( \34861 , \34858 , \34860 );
not \U$34519 ( \34862 , \34861 );
or \U$34520 ( \34863 , \34857 , \34862 );
and \U$34521 ( \34864 , RI9872b80_169, \13391 );
not \U$34522 ( \34865 , RI9872b80_169);
and \U$34523 ( \34866 , \34865 , \13876 );
or \U$34524 ( \34867 , \34864 , \34866 );
nand \U$34525 ( \34868 , \34867 , \9196 );
nand \U$34526 ( \34869 , \34863 , \34868 );
xor \U$34527 ( \34870 , \34856 , \34869 );
not \U$34528 ( \34871 , \34870 );
not \U$34529 ( \34872 , \8751 );
not \U$34530 ( \34873 , \8668 );
not \U$34531 ( \34874 , RI9872f40_177);
and \U$34532 ( \34875 , \34873 , \34874 );
and \U$34533 ( \34876 , \8668 , RI9872f40_177);
nor \U$34534 ( \34877 , \34875 , \34876 );
not \U$34535 ( \34878 , \34877 );
not \U$34536 ( \34879 , \34878 );
or \U$34537 ( \34880 , \34872 , \34879 );
xor \U$34538 ( \34881 , RI9872f40_177, \8640 );
nand \U$34539 ( \34882 , \34881 , \9526 );
nand \U$34540 ( \34883 , \34880 , \34882 );
not \U$34541 ( \34884 , \34883 );
or \U$34542 ( \34885 , \34871 , \34884 );
nand \U$34543 ( \34886 , \34869 , \34856 );
nand \U$34544 ( \34887 , \34885 , \34886 );
not \U$34545 ( \34888 , \8802 );
xor \U$34546 ( \34889 , \8722 , RI9872d60_173);
not \U$34547 ( \34890 , \34889 );
or \U$34548 ( \34891 , \34888 , \34890 );
not \U$34549 ( \34892 , \8807 );
not \U$34550 ( \34893 , \8695 );
or \U$34551 ( \34894 , \34892 , \34893 );
or \U$34552 ( \34895 , \23712 , \8811 );
nand \U$34553 ( \34896 , \34894 , \34895 );
nand \U$34554 ( \34897 , \34896 , \8819 );
nand \U$34555 ( \34898 , \34891 , \34897 );
not \U$34556 ( \34899 , \34898 );
not \U$34557 ( \34900 , \5032 );
and \U$34558 ( \34901 , RI9872478_154, \20490 );
not \U$34559 ( \34902 , RI9872478_154);
and \U$34560 ( \34903 , \34902 , \28653 );
or \U$34561 ( \34904 , \34901 , \34903 );
not \U$34562 ( \34905 , \34904 );
or \U$34563 ( \34906 , \34900 , \34905 );
not \U$34564 ( \34907 , \5025 );
not \U$34565 ( \34908 , \24854 );
or \U$34566 ( \34909 , \34907 , \34908 );
or \U$34567 ( \34910 , \24854 , \5025 );
nand \U$34568 ( \34911 , \34909 , \34910 );
nand \U$34569 ( \34912 , \34911 , \5033 );
nand \U$34570 ( \34913 , \34906 , \34912 );
not \U$34571 ( \34914 , \4922 );
not \U$34572 ( \34915 , \4902 );
not \U$34573 ( \34916 , \28671 );
or \U$34574 ( \34917 , \34915 , \34916 );
or \U$34575 ( \34918 , \23952 , \4902 );
nand \U$34576 ( \34919 , \34917 , \34918 );
not \U$34577 ( \34920 , \34919 );
or \U$34578 ( \34921 , \34914 , \34920 );
and \U$34579 ( \34922 , RI9872388_152, \19383 );
not \U$34580 ( \34923 , RI9872388_152);
and \U$34581 ( \34924 , \34923 , \24449 );
nor \U$34582 ( \34925 , \34922 , \34924 );
nand \U$34583 ( \34926 , \34925 , \4915 );
nand \U$34584 ( \34927 , \34921 , \34926 );
or \U$34585 ( \34928 , RI9872400_153, RI9872478_154);
nand \U$34586 ( \34929 , \34928 , \18704 );
nand \U$34587 ( \34930 , \34929 , \4531 );
xor \U$34588 ( \34931 , \34927 , \34930 );
not \U$34589 ( \34932 , \34931 );
xor \U$34590 ( \34933 , \34913 , \34932 );
not \U$34591 ( \34934 , \34933 );
not \U$34592 ( \34935 , \6285 );
and \U$34593 ( \34936 , RI98728b0_163, \20764 );
not \U$34594 ( \34937 , RI98728b0_163);
not \U$34595 ( \34938 , \25380 );
and \U$34596 ( \34939 , \34937 , \34938 );
or \U$34597 ( \34940 , \34936 , \34939 );
not \U$34598 ( \34941 , \34940 );
or \U$34599 ( \34942 , \34935 , \34941 );
not \U$34600 ( \34943 , RI98728b0_163);
not \U$34601 ( \34944 , \17741 );
or \U$34602 ( \34945 , \34943 , \34944 );
or \U$34603 ( \34946 , \17911 , RI98728b0_163);
nand \U$34604 ( \34947 , \34945 , \34946 );
nand \U$34605 ( \34948 , \34947 , \6282 );
nand \U$34606 ( \34949 , \34942 , \34948 );
not \U$34607 ( \34950 , \34949 );
or \U$34608 ( \34951 , \34934 , \34950 );
not \U$34609 ( \34952 , \34931 );
nand \U$34610 ( \34953 , \34952 , \34913 );
nand \U$34611 ( \34954 , \34951 , \34953 );
not \U$34612 ( \34955 , \34954 );
not \U$34613 ( \34956 , \34955 );
not \U$34614 ( \34957 , \13477 );
not \U$34615 ( \34958 , RI9873210_183);
not \U$34616 ( \34959 , \7466 );
or \U$34617 ( \34960 , \34958 , \34959 );
or \U$34618 ( \34961 , \21642 , RI9873210_183);
nand \U$34619 ( \34962 , \34960 , \34961 );
not \U$34620 ( \34963 , \34962 );
or \U$34621 ( \34964 , \34957 , \34963 );
not \U$34622 ( \34965 , RI9873210_183);
not \U$34623 ( \34966 , \8081 );
or \U$34624 ( \34967 , \34965 , \34966 );
or \U$34625 ( \34968 , \8081 , RI9873210_183);
nand \U$34626 ( \34969 , \34967 , \34968 );
nand \U$34627 ( \34970 , \34969 , \30963 );
nand \U$34628 ( \34971 , \34964 , \34970 );
not \U$34629 ( \34972 , \34971 );
or \U$34630 ( \34973 , \34956 , \34972 );
or \U$34631 ( \34974 , \34971 , \34955 );
nand \U$34632 ( \34975 , \34973 , \34974 );
not \U$34633 ( \34976 , \34975 );
or \U$34634 ( \34977 , \34899 , \34976 );
nand \U$34635 ( \34978 , \34971 , \34954 );
nand \U$34636 ( \34979 , \34977 , \34978 );
xor \U$34637 ( \34980 , \34887 , \34979 );
not \U$34638 ( \34981 , \9293 );
not \U$34639 ( \34982 , RI9872e50_175);
not \U$34640 ( \34983 , \10369 );
or \U$34641 ( \34984 , \34982 , \34983 );
or \U$34642 ( \34985 , \9761 , RI9872e50_175);
nand \U$34643 ( \34986 , \34984 , \34985 );
not \U$34644 ( \34987 , \34986 );
or \U$34645 ( \34988 , \34981 , \34987 );
not \U$34646 ( \34989 , RI9872e50_175);
not \U$34647 ( \34990 , \18312 );
not \U$34648 ( \34991 , \34990 );
or \U$34649 ( \34992 , \34989 , \34991 );
nand \U$34650 ( \34993 , \8580 , \9690 );
nand \U$34651 ( \34994 , \34992 , \34993 );
nand \U$34652 ( \34995 , \34994 , \9272 );
nand \U$34653 ( \34996 , \34988 , \34995 );
not \U$34654 ( \34997 , \17528 );
not \U$34655 ( \34998 , RI9873288_184);
not \U$34656 ( \34999 , \12805 );
or \U$34657 ( \35000 , \34998 , \34999 );
or \U$34658 ( \35001 , \8053 , RI9873288_184);
nand \U$34659 ( \35002 , \35000 , \35001 );
not \U$34660 ( \35003 , \35002 );
or \U$34661 ( \35004 , \34997 , \35003 );
not \U$34662 ( \35005 , \22715 );
not \U$34663 ( \35006 , \10412 );
or \U$34664 ( \35007 , \35005 , \35006 );
or \U$34665 ( \35008 , \10412 , \27966 );
nand \U$34666 ( \35009 , \35007 , \35008 );
nand \U$34667 ( \35010 , \35009 , \32965 );
nand \U$34668 ( \35011 , \35004 , \35010 );
xor \U$34669 ( \35012 , \34996 , \35011 );
not \U$34670 ( \35013 , \17252 );
not \U$34671 ( \35014 , RI98733f0_187);
not \U$34672 ( \35015 , \5705 );
or \U$34673 ( \35016 , \35014 , \35015 );
or \U$34674 ( \35017 , \8895 , RI98733f0_187);
nand \U$34675 ( \35018 , \35016 , \35017 );
not \U$34676 ( \35019 , \35018 );
or \U$34677 ( \35020 , \35013 , \35019 );
not \U$34678 ( \35021 , RI98733f0_187);
and \U$34679 ( \35022 , \35021 , \6480 );
not \U$34680 ( \35023 , \35021 );
and \U$34681 ( \35024 , \35023 , \5761 );
nor \U$34682 ( \35025 , \35022 , \35024 );
or \U$34683 ( \35026 , \35025 , \17620 );
nand \U$34684 ( \35027 , \35020 , \35026 );
and \U$34685 ( \35028 , \35012 , \35027 );
and \U$34686 ( \35029 , \34996 , \35011 );
or \U$34687 ( \35030 , \35028 , \35029 );
xor \U$34688 ( \35031 , \34980 , \35030 );
not \U$34689 ( \35032 , \35031 );
and \U$34690 ( \35033 , \5393 , RI98733f0_187);
not \U$34691 ( \35034 , \5393 );
and \U$34692 ( \35035 , \35034 , \35021 );
nor \U$34693 ( \35036 , \35033 , \35035 );
not \U$34694 ( \35037 , \35036 );
or \U$34695 ( \35038 , \35037 , \17620 );
or \U$34696 ( \35039 , \35025 , \18079 );
nand \U$34697 ( \35040 , \35038 , \35039 );
not \U$34698 ( \35041 , \35040 );
nand \U$34699 ( \35042 , \19383 , \4084 );
not \U$34700 ( \35043 , \35042 );
not \U$34701 ( \35044 , \4922 );
and \U$34702 ( \35045 , \17863 , RI9872388_152);
not \U$34703 ( \35046 , \17863 );
and \U$34704 ( \35047 , \35046 , \7993 );
nor \U$34705 ( \35048 , \35045 , \35047 );
not \U$34706 ( \35049 , \35048 );
or \U$34707 ( \35050 , \35044 , \35049 );
nand \U$34708 ( \35051 , \34919 , \4916 );
nand \U$34709 ( \35052 , \35050 , \35051 );
not \U$34710 ( \35053 , \35052 );
or \U$34711 ( \35054 , \35043 , \35053 );
or \U$34712 ( \35055 , \35052 , \35042 );
nand \U$34713 ( \35056 , \35054 , \35055 );
not \U$34714 ( \35057 , \34904 );
not \U$34715 ( \35058 , \35057 );
not \U$34716 ( \35059 , \7591 );
and \U$34717 ( \35060 , \35058 , \35059 );
and \U$34718 ( \35061 , RI9872478_154, \16995 );
not \U$34719 ( \35062 , RI9872478_154);
and \U$34720 ( \35063 , \35062 , \16996 );
nor \U$34721 ( \35064 , \35061 , \35063 );
and \U$34722 ( \35065 , \35064 , \5035 );
nor \U$34723 ( \35066 , \35060 , \35065 );
not \U$34724 ( \35067 , \35066 );
and \U$34725 ( \35068 , \35056 , \35067 );
not \U$34726 ( \35069 , \35056 );
and \U$34727 ( \35070 , \35069 , \35066 );
nor \U$34728 ( \35071 , \35068 , \35070 );
not \U$34729 ( \35072 , \8028 );
not \U$34730 ( \35073 , RI9872a18_166);
not \U$34731 ( \35074 , \12773 );
or \U$34732 ( \35075 , \35073 , \35074 );
or \U$34733 ( \35076 , \25847 , RI9872a18_166);
nand \U$34734 ( \35077 , \35075 , \35076 );
not \U$34735 ( \35078 , \35077 );
or \U$34736 ( \35079 , \35072 , \35078 );
not \U$34737 ( \35080 , RI9872a18_166);
not \U$34738 ( \35081 , \12784 );
or \U$34739 ( \35082 , \35080 , \35081 );
buf \U$34740 ( \35083 , \18151 );
or \U$34741 ( \35084 , \35083 , RI9872a18_166);
nand \U$34742 ( \35085 , \35082 , \35084 );
nand \U$34743 ( \35086 , \35085 , \13017 );
nand \U$34744 ( \35087 , \35079 , \35086 );
xor \U$34745 ( \35088 , \35071 , \35087 );
not \U$34746 ( \35089 , \9670 );
and \U$34747 ( \35090 , RI9872bf8_170, \9113 );
not \U$34748 ( \35091 , RI9872bf8_170);
and \U$34749 ( \35092 , \35091 , \18344 );
or \U$34750 ( \35093 , \35090 , \35092 );
not \U$34751 ( \35094 , \35093 );
or \U$34752 ( \35095 , \35089 , \35094 );
xnor \U$34753 ( \35096 , \12460 , RI9872bf8_170);
nand \U$34754 ( \35097 , \35096 , \9227 );
nand \U$34755 ( \35098 , \35095 , \35097 );
and \U$34756 ( \35099 , \35088 , \35098 );
and \U$34757 ( \35100 , \35071 , \35087 );
nor \U$34758 ( \35101 , \35099 , \35100 );
not \U$34759 ( \35102 , \35101 );
or \U$34760 ( \35103 , \35041 , \35102 );
not \U$34761 ( \35104 , \35040 );
not \U$34762 ( \35105 , \35101 );
nand \U$34763 ( \35106 , \35104 , \35105 );
nand \U$34764 ( \35107 , \35103 , \35106 );
not \U$34765 ( \35108 , \9214 );
xnor \U$34766 ( \35109 , \9114 , RI9872b80_169);
not \U$34767 ( \35110 , \35109 );
or \U$34768 ( \35111 , \35108 , \35110 );
nand \U$34769 ( \35112 , \34861 , \9196 );
nand \U$34770 ( \35113 , \35111 , \35112 );
not \U$34771 ( \35114 , \35067 );
not \U$34772 ( \35115 , \35056 );
or \U$34773 ( \35116 , \35114 , \35115 );
not \U$34774 ( \35117 , \35042 );
nand \U$34775 ( \35118 , \35117 , \35052 );
nand \U$34776 ( \35119 , \35116 , \35118 );
not \U$34777 ( \35120 , \35119 );
and \U$34778 ( \35121 , RI9872478_154, \25412 );
not \U$34779 ( \35122 , RI9872478_154);
and \U$34780 ( \35123 , \35122 , \19412 );
or \U$34781 ( \35124 , \35121 , \35123 );
not \U$34782 ( \35125 , \35124 );
not \U$34783 ( \35126 , \35125 );
not \U$34784 ( \35127 , \5795 );
and \U$34785 ( \35128 , \35126 , \35127 );
and \U$34786 ( \35129 , \35064 , \5034 );
nor \U$34787 ( \35130 , \35128 , \35129 );
not \U$34788 ( \35131 , \35130 );
and \U$34789 ( \35132 , \35120 , \35131 );
and \U$34790 ( \35133 , \35119 , \35130 );
nor \U$34791 ( \35134 , \35132 , \35133 );
xor \U$34792 ( \35135 , \35113 , \35134 );
and \U$34793 ( \35136 , \35107 , \35135 );
not \U$34794 ( \35137 , \35107 );
not \U$34795 ( \35138 , \35135 );
and \U$34796 ( \35139 , \35137 , \35138 );
nor \U$34797 ( \35140 , \35136 , \35139 );
not \U$34798 ( \35141 , \35140 );
not \U$34799 ( \35142 , \19046 );
not \U$34800 ( \35143 , RI98734e0_189);
not \U$34801 ( \35144 , \5774 );
or \U$34802 ( \35145 , \35143 , \35144 );
not \U$34803 ( \35146 , RI98734e0_189);
nand \U$34804 ( \35147 , \5392 , \35146 );
nand \U$34805 ( \35148 , \35145 , \35147 );
not \U$34806 ( \35149 , \35148 );
or \U$34807 ( \35150 , \35142 , \35149 );
not \U$34808 ( \35151 , RI98734e0_189);
not \U$34809 ( \35152 , \5761 );
or \U$34810 ( \35153 , \35151 , \35152 );
or \U$34811 ( \35154 , \6481 , RI98734e0_189);
nand \U$34812 ( \35155 , \35153 , \35154 );
nand \U$34813 ( \35156 , \35155 , \24076 );
nand \U$34814 ( \35157 , \35150 , \35156 );
not \U$34815 ( \35158 , \35157 );
not \U$34816 ( \35159 , \12507 );
not \U$34817 ( \35160 , RI9873030_179);
not \U$34818 ( \35161 , \8857 );
or \U$34819 ( \35162 , \35160 , \35161 );
or \U$34820 ( \35163 , \9882 , RI9873030_179);
nand \U$34821 ( \35164 , \35162 , \35163 );
not \U$34822 ( \35165 , \35164 );
or \U$34823 ( \35166 , \35159 , \35165 );
not \U$34824 ( \35167 , RI9873030_179);
not \U$34825 ( \35168 , \8607 );
or \U$34826 ( \35169 , \35167 , \35168 );
or \U$34827 ( \35170 , \10308 , RI9873030_179);
nand \U$34828 ( \35171 , \35169 , \35170 );
nand \U$34829 ( \35172 , \35171 , \9937 );
nand \U$34830 ( \35173 , \35166 , \35172 );
not \U$34831 ( \35174 , \35173 );
or \U$34832 ( \35175 , \35158 , \35174 );
or \U$34833 ( \35176 , \35173 , \35157 );
not \U$34834 ( \35177 , RI9873648_192);
not \U$34835 ( \35178 , RI9873558_190);
not \U$34836 ( \35179 , \7791 );
or \U$34837 ( \35180 , \35178 , \35179 );
or \U$34838 ( \35181 , \4990 , RI9873558_190);
nand \U$34839 ( \35182 , \35180 , \35181 );
not \U$34840 ( \35183 , \35182 );
or \U$34841 ( \35184 , \35177 , \35183 );
not \U$34842 ( \35185 , \18239 );
not \U$34843 ( \35186 , \9374 );
or \U$34844 ( \35187 , \35185 , \35186 );
nand \U$34845 ( \35188 , \5736 , RI9873558_190);
nand \U$34846 ( \35189 , \35187 , \35188 );
nand \U$34847 ( \35190 , \35189 , \18545 );
nand \U$34848 ( \35191 , \35184 , \35190 );
nand \U$34849 ( \35192 , \35176 , \35191 );
nand \U$34850 ( \35193 , \35175 , \35192 );
not \U$34851 ( \35194 , \35193 );
xor \U$34852 ( \35195 , \34996 , \35011 );
xor \U$34853 ( \35196 , \35195 , \35027 );
not \U$34854 ( \35197 , \35196 );
or \U$34855 ( \35198 , \35194 , \35197 );
or \U$34856 ( \35199 , \35196 , \35193 );
not \U$34857 ( \35200 , \28811 );
not \U$34858 ( \35201 , \22314 );
xor \U$34859 ( \35202 , RI98734e0_189, \35201 );
not \U$34860 ( \35203 , \35202 );
or \U$34861 ( \35204 , \35200 , \35203 );
nand \U$34862 ( \35205 , \35148 , \19243 );
nand \U$34863 ( \35206 , \35204 , \35205 );
not \U$34864 ( \35207 , \17347 );
not \U$34865 ( \35208 , \8333 );
xor \U$34866 ( \35209 , RI98730a8_180, \35208 );
not \U$34867 ( \35210 , \35209 );
or \U$34868 ( \35211 , \35207 , \35210 );
xor \U$34869 ( \35212 , RI98730a8_180, \9598 );
nand \U$34870 ( \35213 , \35212 , \13020 );
nand \U$34871 ( \35214 , \35211 , \35213 );
xor \U$34872 ( \35215 , \35206 , \35214 );
not \U$34873 ( \35216 , \18672 );
not \U$34874 ( \35217 , \35171 );
or \U$34875 ( \35218 , \35216 , \35217 );
not \U$34876 ( \35219 , RI9873030_179);
not \U$34877 ( \35220 , \12712 );
or \U$34878 ( \35221 , \35219 , \35220 );
buf \U$34879 ( \35222 , \22347 );
or \U$34880 ( \35223 , \35222 , RI9873030_179);
nand \U$34881 ( \35224 , \35221 , \35223 );
nand \U$34882 ( \35225 , \35224 , \9937 );
nand \U$34883 ( \35226 , \35218 , \35225 );
xor \U$34884 ( \35227 , \35215 , \35226 );
nand \U$34885 ( \35228 , \35199 , \35227 );
nand \U$34886 ( \35229 , \35198 , \35228 );
not \U$34887 ( \35230 , \35229 );
or \U$34888 ( \35231 , \35141 , \35230 );
or \U$34889 ( \35232 , \35229 , \35140 );
nand \U$34890 ( \35233 , \35231 , \35232 );
not \U$34891 ( \35234 , \35233 );
or \U$34892 ( \35235 , \35032 , \35234 );
not \U$34893 ( \35236 , \35140 );
nand \U$34894 ( \35237 , \35236 , \35229 );
nand \U$34895 ( \35238 , \35235 , \35237 );
not \U$34896 ( \35239 , \22664 );
and \U$34897 ( \35240 , RI9872d60_173, \13298 );
not \U$34898 ( \35241 , RI9872d60_173);
and \U$34899 ( \35242 , \35241 , \10372 );
or \U$34900 ( \35243 , \35240 , \35242 );
not \U$34901 ( \35244 , \35243 );
or \U$34902 ( \35245 , \35239 , \35244 );
and \U$34903 ( \35246 , RI9872d60_173, \19701 );
not \U$34904 ( \35247 , RI9872d60_173);
and \U$34905 ( \35248 , \35247 , \12848 );
or \U$34906 ( \35249 , \35246 , \35248 );
nand \U$34907 ( \35250 , \35249 , \10624 );
nand \U$34908 ( \35251 , \35245 , \35250 );
not \U$34909 ( \35252 , \24627 );
not \U$34910 ( \35253 , \8732 );
not \U$34911 ( \35254 , \8597 );
or \U$34912 ( \35255 , \35253 , \35254 );
nand \U$34913 ( \35256 , \10308 , RI9872f40_177);
nand \U$34914 ( \35257 , \35255 , \35256 );
not \U$34915 ( \35258 , \35257 );
or \U$34916 ( \35259 , \35252 , \35258 );
not \U$34917 ( \35260 , \8732 );
not \U$34918 ( \35261 , \10597 );
or \U$34919 ( \35262 , \35260 , \35261 );
nand \U$34920 ( \35263 , \8878 , RI9872f40_177);
nand \U$34921 ( \35264 , \35262 , \35263 );
nand \U$34922 ( \35265 , \35264 , \8751 );
nand \U$34923 ( \35266 , \35259 , \35265 );
xor \U$34924 ( \35267 , \35251 , \35266 );
not \U$34925 ( \35268 , \9686 );
not \U$34926 ( \35269 , \8650 );
not \U$34927 ( \35270 , RI9872e50_175);
and \U$34928 ( \35271 , \35269 , \35270 );
and \U$34929 ( \35272 , \8650 , RI9872e50_175);
nor \U$34930 ( \35273 , \35271 , \35272 );
not \U$34931 ( \35274 , \35273 );
not \U$34932 ( \35275 , \35274 );
or \U$34933 ( \35276 , \35268 , \35275 );
and \U$34934 ( \35277 , \9880 , \9690 );
not \U$34935 ( \35278 , \9880 );
and \U$34936 ( \35279 , \35278 , RI9872e50_175);
nor \U$34937 ( \35280 , \35277 , \35279 );
nand \U$34938 ( \35281 , \35280 , \9273 );
nand \U$34939 ( \35282 , \35276 , \35281 );
xor \U$34940 ( \35283 , \35267 , \35282 );
not \U$34941 ( \35284 , RI98728b0_163);
not \U$34942 ( \35285 , \24523 );
or \U$34943 ( \35286 , \35284 , \35285 );
nand \U$34944 ( \35287 , \13281 , \5632 );
nand \U$34945 ( \35288 , \35286 , \35287 );
not \U$34946 ( \35289 , \35288 );
or \U$34947 ( \35290 , \35289 , \6609 );
not \U$34948 ( \35291 , \6283 );
and \U$34949 ( \35292 , \20787 , \5632 );
not \U$34950 ( \35293 , \20787 );
and \U$34951 ( \35294 , \35293 , RI98728b0_163);
nor \U$34952 ( \35295 , \35292 , \35294 );
nand \U$34953 ( \35296 , \35291 , \35295 );
nand \U$34954 ( \35297 , \35290 , \35296 );
not \U$34955 ( \35298 , \7326 );
not \U$34956 ( \35299 , \7333 );
not \U$34957 ( \35300 , \12774 );
or \U$34958 ( \35301 , \35299 , \35300 );
nand \U$34959 ( \35302 , \12773 , RI98729a0_165);
nand \U$34960 ( \35303 , \35301 , \35302 );
not \U$34961 ( \35304 , \35303 );
or \U$34962 ( \35305 , \35298 , \35304 );
not \U$34963 ( \35306 , RI98729a0_165);
not \U$34964 ( \35307 , \18151 );
or \U$34965 ( \35308 , \35306 , \35307 );
or \U$34966 ( \35309 , \29808 , RI98729a0_165);
nand \U$34967 ( \35310 , \35308 , \35309 );
nand \U$34968 ( \35311 , \35310 , \7338 );
nand \U$34969 ( \35312 , \35305 , \35311 );
xor \U$34970 ( \35313 , \35297 , \35312 );
not \U$34971 ( \35314 , \13477 );
not \U$34972 ( \35315 , \28789 );
not \U$34973 ( \35316 , \7905 );
or \U$34974 ( \35317 , \35315 , \35316 );
or \U$34975 ( \35318 , \8934 , \22675 );
nand \U$34976 ( \35319 , \35317 , \35318 );
not \U$34977 ( \35320 , \35319 );
or \U$34978 ( \35321 , \35314 , \35320 );
not \U$34979 ( \35322 , RI9873210_183);
not \U$34980 ( \35323 , \8053 );
or \U$34981 ( \35324 , \35322 , \35323 );
or \U$34982 ( \35325 , \8904 , RI9873210_183);
nand \U$34983 ( \35326 , \35324 , \35325 );
nand \U$34984 ( \35327 , \35326 , \30963 );
nand \U$34985 ( \35328 , \35321 , \35327 );
xor \U$34986 ( \35329 , \35313 , \35328 );
or \U$34987 ( \35330 , \35283 , \35329 );
nand \U$34988 ( \35331 , \35283 , \35329 );
nand \U$34989 ( \35332 , \35330 , \35331 );
not \U$34990 ( \35333 , \12867 );
not \U$34991 ( \35334 , RI98730a8_180);
not \U$34992 ( \35335 , \13645 );
or \U$34993 ( \35336 , \35334 , \35335 );
or \U$34994 ( \35337 , \8081 , RI98730a8_180);
nand \U$34995 ( \35338 , \35336 , \35337 );
not \U$34996 ( \35339 , \35338 );
or \U$34997 ( \35340 , \35333 , \35339 );
and \U$34998 ( \35341 , RI98730a8_180, \7466 );
not \U$34999 ( \35342 , RI98730a8_180);
and \U$35000 ( \35343 , \35342 , \8923 );
or \U$35001 ( \35344 , \35341 , \35343 );
nand \U$35002 ( \35345 , \35344 , \24209 );
nand \U$35003 ( \35346 , \35340 , \35345 );
not \U$35004 ( \35347 , \18672 );
and \U$35005 ( \35348 , RI9873030_179, \11628 );
not \U$35006 ( \35349 , RI9873030_179);
and \U$35007 ( \35350 , \35349 , \8075 );
or \U$35008 ( \35351 , \35348 , \35350 );
not \U$35009 ( \35352 , \35351 );
or \U$35010 ( \35353 , \35347 , \35352 );
and \U$35011 ( \35354 , RI9873030_179, \8333 );
not \U$35012 ( \35355 , RI9873030_179);
and \U$35013 ( \35356 , \35355 , \8916 );
or \U$35014 ( \35357 , \35354 , \35356 );
nand \U$35015 ( \35358 , \35357 , \9937 );
nand \U$35016 ( \35359 , \35353 , \35358 );
and \U$35017 ( \35360 , \35346 , \35359 );
not \U$35018 ( \35361 , \35346 );
not \U$35019 ( \35362 , \35359 );
and \U$35020 ( \35363 , \35361 , \35362 );
nor \U$35021 ( \35364 , \35360 , \35363 );
buf \U$35022 ( \35365 , \35364 );
not \U$35023 ( \35366 , \19036 );
and \U$35024 ( \35367 , RI98734e0_189, \4960 );
not \U$35025 ( \35368 , RI98734e0_189);
and \U$35026 ( \35369 , \35368 , \4990 );
nor \U$35027 ( \35370 , \35367 , \35369 );
not \U$35028 ( \35371 , \35370 );
or \U$35029 ( \35372 , \35366 , \35371 );
and \U$35030 ( \35373 , RI98734e0_189, \4470 );
not \U$35031 ( \35374 , RI98734e0_189);
and \U$35032 ( \35375 , \35374 , \4472 );
or \U$35033 ( \35376 , \35373 , \35375 );
nand \U$35034 ( \35377 , \35376 , \20147 );
nand \U$35035 ( \35378 , \35372 , \35377 );
and \U$35036 ( \35379 , \35365 , \35378 );
not \U$35037 ( \35380 , \35365 );
not \U$35038 ( \35381 , \35378 );
and \U$35039 ( \35382 , \35380 , \35381 );
nor \U$35040 ( \35383 , \35379 , \35382 );
and \U$35041 ( \35384 , \35332 , \35383 );
not \U$35042 ( \35385 , \35332 );
not \U$35043 ( \35386 , \35383 );
and \U$35044 ( \35387 , \35385 , \35386 );
nor \U$35045 ( \35388 , \35384 , \35387 );
not \U$35046 ( \35389 , \35388 );
xor \U$35047 ( \35390 , \35206 , \35214 );
and \U$35048 ( \35391 , \35390 , \35226 );
and \U$35049 ( \35392 , \35206 , \35214 );
or \U$35050 ( \35393 , \35391 , \35392 );
not \U$35051 ( \35394 , \7338 );
not \U$35052 ( \35395 , \35303 );
or \U$35053 ( \35396 , \35394 , \35395 );
nand \U$35054 ( \35397 , \34854 , \7325 );
nand \U$35055 ( \35398 , \35396 , \35397 );
not \U$35056 ( \35399 , \35398 );
not \U$35057 ( \35400 , \35399 );
not \U$35058 ( \35401 , \9071 );
not \U$35059 ( \35402 , RI9872a18_166);
not \U$35060 ( \35403 , \10064 );
or \U$35061 ( \35404 , \35402 , \35403 );
or \U$35062 ( \35405 , \10064 , RI9872a18_166);
nand \U$35063 ( \35406 , \35404 , \35405 );
not \U$35064 ( \35407 , \35406 );
or \U$35065 ( \35408 , \35401 , \35407 );
nand \U$35066 ( \35409 , \35085 , \8027 );
nand \U$35067 ( \35410 , \35408 , \35409 );
not \U$35068 ( \35411 , \6285 );
not \U$35069 ( \35412 , \35295 );
or \U$35070 ( \35413 , \35411 , \35412 );
not \U$35071 ( \35414 , RI98728b0_163);
not \U$35072 ( \35415 , \13860 );
or \U$35073 ( \35416 , \35414 , \35415 );
or \U$35074 ( \35417 , \17015 , RI98728b0_163);
nand \U$35075 ( \35418 , \35416 , \35417 );
nand \U$35076 ( \35419 , \35418 , \6282 );
nand \U$35077 ( \35420 , \35413 , \35419 );
xor \U$35078 ( \35421 , \35410 , \35420 );
not \U$35079 ( \35422 , \35421 );
or \U$35080 ( \35423 , \35400 , \35422 );
or \U$35081 ( \35424 , \35421 , \35399 );
nand \U$35082 ( \35425 , \35423 , \35424 );
xor \U$35083 ( \35426 , \35393 , \35425 );
not \U$35084 ( \35427 , \35426 );
not \U$35085 ( \35428 , \17702 );
not \U$35086 ( \35429 , \35428 );
not \U$35087 ( \35430 , RI9872388_152);
and \U$35088 ( \35431 , \35429 , \35430 );
and \U$35089 ( \35432 , \33482 , RI9872388_152);
nor \U$35090 ( \35433 , \35431 , \35432 );
or \U$35091 ( \35434 , \35433 , \32178 );
not \U$35092 ( \35435 , \35048 );
or \U$35093 ( \35436 , \35435 , \4917 );
nand \U$35094 ( \35437 , \35434 , \35436 );
not \U$35095 ( \35438 , \35437 );
not \U$35096 ( \35439 , \4084 );
xor \U$35097 ( \35440 , \25166 , RI98725e0_157);
not \U$35098 ( \35441 , \35440 );
or \U$35099 ( \35442 , \35439 , \35441 );
xor \U$35100 ( \35443 , \18705 , RI98725e0_157);
nand \U$35101 ( \35444 , \35443 , \4101 );
nand \U$35102 ( \35445 , \35442 , \35444 );
or \U$35103 ( \35446 , RI9872388_152, RI98727c0_161);
nand \U$35104 ( \35447 , \35446 , \18705 );
nand \U$35105 ( \35448 , \35447 , \3926 );
not \U$35106 ( \35449 , \35448 );
and \U$35107 ( \35450 , \35445 , \35449 );
not \U$35108 ( \35451 , \35445 );
and \U$35109 ( \35452 , \35451 , \35448 );
or \U$35110 ( \35453 , \35450 , \35452 );
not \U$35111 ( \35454 , \35453 );
or \U$35112 ( \35455 , \35438 , \35454 );
or \U$35113 ( \35456 , \35453 , \35437 );
nand \U$35114 ( \35457 , \35455 , \35456 );
not \U$35115 ( \35458 , \5653 );
and \U$35116 ( \35459 , \25380 , \5644 );
not \U$35117 ( \35460 , \25380 );
and \U$35118 ( \35461 , \35460 , RI9872568_156);
nor \U$35119 ( \35462 , \35459 , \35461 );
not \U$35120 ( \35463 , \35462 );
or \U$35121 ( \35464 , \35458 , \35463 );
xor \U$35122 ( \35465 , \28191 , RI9872568_156);
nand \U$35123 ( \35466 , \35465 , \5641 );
nand \U$35124 ( \35467 , \35464 , \35466 );
xor \U$35125 ( \35468 , \35457 , \35467 );
not \U$35126 ( \35469 , \34877 );
not \U$35127 ( \35470 , \18284 );
and \U$35128 ( \35471 , \35469 , \35470 );
and \U$35129 ( \35472 , \35257 , \8751 );
nor \U$35130 ( \35473 , \35471 , \35472 );
xor \U$35131 ( \35474 , \35468 , \35473 );
not \U$35132 ( \35475 , \17123 );
not \U$35133 ( \35476 , \35319 );
or \U$35134 ( \35477 , \35475 , \35476 );
nand \U$35135 ( \35478 , \34969 , \13477 );
nand \U$35136 ( \35479 , \35477 , \35478 );
xnor \U$35137 ( \35480 , \35474 , \35479 );
not \U$35138 ( \35481 , \35480 );
or \U$35139 ( \35482 , \35427 , \35481 );
nand \U$35140 ( \35483 , \35393 , \35425 );
nand \U$35141 ( \35484 , \35482 , \35483 );
not \U$35142 ( \35485 , \34927 );
nor \U$35143 ( \35486 , \35485 , \34930 );
not \U$35144 ( \35487 , \6063 );
and \U$35145 ( \35488 , RI9872568_156, \27889 );
not \U$35146 ( \35489 , RI9872568_156);
and \U$35147 ( \35490 , \35489 , \19412 );
or \U$35148 ( \35491 , \35488 , \35490 );
not \U$35149 ( \35492 , \35491 );
or \U$35150 ( \35493 , \35487 , \35492 );
nand \U$35151 ( \35494 , \35465 , \5653 );
nand \U$35152 ( \35495 , \35493 , \35494 );
xor \U$35153 ( \35496 , \35486 , \35495 );
not \U$35154 ( \35497 , \6282 );
not \U$35155 ( \35498 , \34940 );
or \U$35156 ( \35499 , \35497 , \35498 );
nand \U$35157 ( \35500 , \35418 , \6285 );
nand \U$35158 ( \35501 , \35499 , \35500 );
and \U$35159 ( \35502 , \35496 , \35501 );
and \U$35160 ( \35503 , \35486 , \35495 );
nor \U$35161 ( \35504 , \35502 , \35503 );
not \U$35162 ( \35505 , \35504 );
not \U$35163 ( \35506 , \35505 );
not \U$35164 ( \35507 , \17528 );
not \U$35165 ( \35508 , \22715 );
not \U$35166 ( \35509 , \6303 );
or \U$35167 ( \35510 , \35508 , \35509 );
or \U$35168 ( \35511 , \11438 , \27966 );
nand \U$35169 ( \35512 , \35510 , \35511 );
not \U$35170 ( \35513 , \35512 );
or \U$35171 ( \35514 , \35507 , \35513 );
nand \U$35172 ( \35515 , \35002 , \18508 );
nand \U$35173 ( \35516 , \35514 , \35515 );
not \U$35174 ( \35517 , \35516 );
or \U$35175 ( \35518 , \35506 , \35517 );
not \U$35176 ( \35519 , \12867 );
not \U$35177 ( \35520 , \35344 );
or \U$35178 ( \35521 , \35519 , \35520 );
nand \U$35179 ( \35522 , \35209 , \13020 );
nand \U$35180 ( \35523 , \35521 , \35522 );
not \U$35181 ( \35524 , \35523 );
nand \U$35182 ( \35525 , \35518 , \35524 );
not \U$35183 ( \35526 , \35516 );
nand \U$35184 ( \35527 , \35526 , \35504 );
not \U$35185 ( \35528 , \4084 );
not \U$35186 ( \35529 , \4088 );
not \U$35187 ( \35530 , \34407 );
not \U$35188 ( \35531 , \35530 );
or \U$35189 ( \35532 , \35529 , \35531 );
or \U$35190 ( \35533 , \24854 , \4088 );
nand \U$35191 ( \35534 , \35532 , \35533 );
not \U$35192 ( \35535 , \35534 );
or \U$35193 ( \35536 , \35528 , \35535 );
nand \U$35194 ( \35537 , \35440 , \4101 );
nand \U$35195 ( \35538 , \35536 , \35537 );
and \U$35196 ( \35539 , \21779 , \3467 );
and \U$35197 ( \35540 , \35538 , \35539 );
not \U$35198 ( \35541 , \35538 );
not \U$35199 ( \35542 , \35539 );
and \U$35200 ( \35543 , \35541 , \35542 );
nor \U$35201 ( \35544 , \35540 , \35543 );
not \U$35202 ( \35545 , \4922 );
and \U$35203 ( \35546 , \16996 , \4902 );
not \U$35204 ( \35547 , \16996 );
and \U$35205 ( \35548 , \35547 , RI9872388_152);
nor \U$35206 ( \35549 , \35546 , \35548 );
not \U$35207 ( \35550 , \35549 );
or \U$35208 ( \35551 , \35545 , \35550 );
not \U$35209 ( \35552 , \35433 );
nand \U$35210 ( \35553 , \35552 , \4916 );
nand \U$35211 ( \35554 , \35551 , \35553 );
xor \U$35212 ( \35555 , \35544 , \35554 );
not \U$35213 ( \35556 , \8027 );
not \U$35214 ( \35557 , \35406 );
or \U$35215 ( \35558 , \35556 , \35557 );
not \U$35216 ( \35559 , \7901 );
not \U$35217 ( \35560 , \13070 );
or \U$35218 ( \35561 , \35559 , \35560 );
not \U$35219 ( \35562 , \17758 );
nand \U$35220 ( \35563 , \35562 , RI9872a18_166);
nand \U$35221 ( \35564 , \35561 , \35563 );
nand \U$35222 ( \35565 , \35564 , \8039 );
nand \U$35223 ( \35566 , \35558 , \35565 );
xor \U$35224 ( \35567 , \35555 , \35566 );
not \U$35225 ( \35568 , \9196 );
not \U$35226 ( \35569 , \35109 );
or \U$35227 ( \35570 , \35568 , \35569 );
and \U$35228 ( \35571 , RI9872b80_169, \12460 );
not \U$35229 ( \35572 , RI9872b80_169);
and \U$35230 ( \35573 , \35572 , \8708 );
or \U$35231 ( \35574 , \35571 , \35573 );
nand \U$35232 ( \35575 , \35574 , \9214 );
nand \U$35233 ( \35576 , \35570 , \35575 );
xor \U$35234 ( \35577 , \35567 , \35576 );
and \U$35235 ( \35578 , \35525 , \35527 , \35577 );
not \U$35236 ( \35579 , \35578 );
not \U$35237 ( \35580 , \35577 );
nand \U$35238 ( \35581 , \35527 , \35525 );
nand \U$35239 ( \35582 , \35580 , \35581 );
nand \U$35240 ( \35583 , \35579 , \35582 );
not \U$35241 ( \35584 , \10624 );
not \U$35242 ( \35585 , \35243 );
or \U$35243 ( \35586 , \35584 , \35585 );
nand \U$35244 ( \35587 , \34889 , \9312 );
nand \U$35245 ( \35588 , \35586 , \35587 );
not \U$35246 ( \35589 , \35588 );
not \U$35247 ( \35590 , \35273 );
not \U$35248 ( \35591 , \9272 );
not \U$35249 ( \35592 , \35591 );
and \U$35250 ( \35593 , \35590 , \35592 );
and \U$35251 ( \35594 , \34994 , \9294 );
nor \U$35252 ( \35595 , \35593 , \35594 );
not \U$35253 ( \35596 , \22167 );
not \U$35254 ( \35597 , \9185 );
not \U$35255 ( \35598 , \9750 );
or \U$35256 ( \35599 , \35597 , \35598 );
nand \U$35257 ( \35600 , \23713 , RI9872bf8_170);
nand \U$35258 ( \35601 , \35599 , \35600 );
not \U$35259 ( \35602 , \35601 );
or \U$35260 ( \35603 , \35596 , \35602 );
nand \U$35261 ( \35604 , \35096 , \9249 );
nand \U$35262 ( \35605 , \35603 , \35604 );
not \U$35263 ( \35606 , \35605 );
and \U$35264 ( \35607 , \35595 , \35606 );
not \U$35265 ( \35608 , \35595 );
and \U$35266 ( \35609 , \35608 , \35605 );
nor \U$35267 ( \35610 , \35607 , \35609 );
not \U$35268 ( \35611 , \35610 );
or \U$35269 ( \35612 , \35589 , \35611 );
not \U$35270 ( \35613 , \35595 );
nand \U$35271 ( \35614 , \35613 , \35605 );
nand \U$35272 ( \35615 , \35612 , \35614 );
and \U$35273 ( \35616 , \35583 , \35615 );
not \U$35274 ( \35617 , \35583 );
not \U$35275 ( \35618 , \35615 );
and \U$35276 ( \35619 , \35617 , \35618 );
nor \U$35277 ( \35620 , \35616 , \35619 );
not \U$35278 ( \35621 , \35620 );
and \U$35279 ( \35622 , \35484 , \35621 );
not \U$35280 ( \35623 , \35484 );
and \U$35281 ( \35624 , \35623 , \35620 );
nor \U$35282 ( \35625 , \35622 , \35624 );
not \U$35283 ( \35626 , \35625 );
or \U$35284 ( \35627 , \35389 , \35626 );
or \U$35285 ( \35628 , \35388 , \35625 );
nand \U$35286 ( \35629 , \35627 , \35628 );
or \U$35287 ( \35630 , \35238 , \35629 );
and \U$35288 ( \35631 , \35445 , \35449 );
not \U$35289 ( \35632 , \5035 );
and \U$35290 ( \35633 , RI9872478_154, \17741 );
not \U$35291 ( \35634 , RI9872478_154);
and \U$35292 ( \35635 , \35634 , \31226 );
or \U$35293 ( \35636 , \35633 , \35635 );
not \U$35294 ( \35637 , \35636 );
or \U$35295 ( \35638 , \35632 , \35637 );
nand \U$35296 ( \35639 , \35124 , \5034 );
nand \U$35297 ( \35640 , \35638 , \35639 );
xor \U$35298 ( \35641 , \35631 , \35640 );
not \U$35299 ( \35642 , \9320 );
not \U$35300 ( \35643 , \35462 );
or \U$35301 ( \35644 , \35642 , \35643 );
not \U$35302 ( \35645 , \13860 );
xor \U$35303 ( \35646 , \35645 , RI9872568_156);
nand \U$35304 ( \35647 , \35646 , \5653 );
nand \U$35305 ( \35648 , \35644 , \35647 );
xor \U$35306 ( \35649 , \35641 , \35648 );
not \U$35307 ( \35650 , \17263 );
and \U$35308 ( \35651 , RI98733f0_187, \4986 );
not \U$35309 ( \35652 , RI98733f0_187);
and \U$35310 ( \35653 , \35652 , \5739 );
or \U$35311 ( \35654 , \35651 , \35653 );
not \U$35312 ( \35655 , \35654 );
or \U$35313 ( \35656 , \35650 , \35655 );
nand \U$35314 ( \35657 , \35036 , \17251 );
nand \U$35315 ( \35658 , \35656 , \35657 );
xor \U$35316 ( \35659 , \35649 , \35658 );
not \U$35317 ( \35660 , RI9873648_192);
and \U$35318 ( \35661 , \11028 , \18239 );
not \U$35319 ( \35662 , \11028 );
and \U$35320 ( \35663 , \35662 , RI9873558_190);
nor \U$35321 ( \35664 , \35661 , \35663 );
not \U$35322 ( \35665 , \35664 );
or \U$35323 ( \35666 , \35660 , \35665 );
not \U$35324 ( \35667 , \18239 );
not \U$35325 ( \35668 , \5208 );
or \U$35326 ( \35669 , \35667 , \35668 );
nand \U$35327 ( \35670 , \5614 , RI9873558_190);
nand \U$35328 ( \35671 , \35669 , \35670 );
nand \U$35329 ( \35672 , \35671 , \20626 );
nand \U$35330 ( \35673 , \35666 , \35672 );
xor \U$35331 ( \35674 , \35659 , \35673 );
xor \U$35332 ( \35675 , \34887 , \34979 );
and \U$35333 ( \35676 , \35675 , \35030 );
and \U$35334 ( \35677 , \34887 , \34979 );
or \U$35335 ( \35678 , \35676 , \35677 );
not \U$35336 ( \35679 , \35678 );
xor \U$35337 ( \35680 , \35674 , \35679 );
nor \U$35338 ( \35681 , \35479 , \35468 );
or \U$35339 ( \35682 , \35681 , \35473 );
nand \U$35340 ( \35683 , \35479 , \35468 );
nand \U$35341 ( \35684 , \35682 , \35683 );
not \U$35342 ( \35685 , \35398 );
not \U$35343 ( \35686 , \35421 );
or \U$35344 ( \35687 , \35685 , \35686 );
nand \U$35345 ( \35688 , \35410 , \35420 );
nand \U$35346 ( \35689 , \35687 , \35688 );
not \U$35347 ( \35690 , \35134 );
not \U$35348 ( \35691 , \35690 );
not \U$35349 ( \35692 , \35113 );
or \U$35350 ( \35693 , \35691 , \35692 );
not \U$35351 ( \35694 , \35130 );
nand \U$35352 ( \35695 , \35694 , \35119 );
nand \U$35353 ( \35696 , \35693 , \35695 );
xor \U$35354 ( \35697 , \35689 , \35696 );
xnor \U$35355 ( \35698 , \35684 , \35697 );
xnor \U$35356 ( \35699 , \35680 , \35698 );
not \U$35357 ( \35700 , \35699 );
nand \U$35358 ( \35701 , \35630 , \35700 );
nand \U$35359 ( \35702 , \35238 , \35629 );
nand \U$35360 ( \35703 , \35701 , \35702 );
not \U$35361 ( \35704 , \35703 );
not \U$35362 ( \35705 , \9937 );
not \U$35363 ( \35706 , \35351 );
or \U$35364 ( \35707 , \35705 , \35706 );
nand \U$35365 ( \35708 , \35224 , \9952 );
nand \U$35366 ( \35709 , \35707 , \35708 );
not \U$35367 ( \35710 , \19046 );
not \U$35368 ( \35711 , \35370 );
or \U$35369 ( \35712 , \35710 , \35711 );
nand \U$35370 ( \35713 , \35202 , \19244 );
nand \U$35371 ( \35714 , \35712 , \35713 );
xor \U$35372 ( \35715 , \35709 , \35714 );
not \U$35373 ( \35716 , RI9873648_192);
not \U$35374 ( \35717 , \35671 );
or \U$35375 ( \35718 , \35716 , \35717 );
not \U$35376 ( \35719 , \18239 );
not \U$35377 ( \35720 , \4712 );
or \U$35378 ( \35721 , \35719 , \35720 );
nand \U$35379 ( \35722 , \4470 , RI9873558_190);
nand \U$35380 ( \35723 , \35721 , \35722 );
nand \U$35381 ( \35724 , \35723 , \18615 );
nand \U$35382 ( \35725 , \35718 , \35724 );
xor \U$35383 ( \35726 , \35715 , \35725 );
not \U$35384 ( \35727 , \35726 );
xor \U$35385 ( \35728 , \35504 , \35523 );
xnor \U$35386 ( \35729 , \35728 , \35516 );
not \U$35387 ( \35730 , \35729 );
not \U$35388 ( \35731 , \35730 );
not \U$35389 ( \35732 , \35610 );
and \U$35390 ( \35733 , \35588 , \35732 );
not \U$35391 ( \35734 , \35588 );
and \U$35392 ( \35735 , \35734 , \35610 );
nor \U$35393 ( \35736 , \35733 , \35735 );
not \U$35394 ( \35737 , \35736 );
not \U$35395 ( \35738 , \35737 );
or \U$35396 ( \35739 , \35731 , \35738 );
nand \U$35397 ( \35740 , \35736 , \35729 );
nand \U$35398 ( \35741 , \35739 , \35740 );
not \U$35399 ( \35742 , \35741 );
or \U$35400 ( \35743 , \35727 , \35742 );
not \U$35401 ( \35744 , \35736 );
nand \U$35402 ( \35745 , \35744 , \35729 );
nand \U$35403 ( \35746 , \35743 , \35745 );
not \U$35404 ( \35747 , \35457 );
not \U$35405 ( \35748 , \35467 );
or \U$35406 ( \35749 , \35747 , \35748 );
not \U$35407 ( \35750 , \35453 );
nand \U$35408 ( \35751 , \35750 , \35437 );
nand \U$35409 ( \35752 , \35749 , \35751 );
not \U$35410 ( \35753 , \9668 );
and \U$35411 ( \35754 , \22752 , \19775 );
not \U$35412 ( \35755 , \22752 );
and \U$35413 ( \35756 , \35755 , RI9872bf8_170);
nor \U$35414 ( \35757 , \35754 , \35756 );
not \U$35415 ( \35758 , \35757 );
or \U$35416 ( \35759 , \35753 , \35758 );
nand \U$35417 ( \35760 , \35601 , \9249 );
nand \U$35418 ( \35761 , \35759 , \35760 );
xor \U$35419 ( \35762 , \35752 , \35761 );
not \U$35420 ( \35763 , \18508 );
not \U$35421 ( \35764 , \35512 );
or \U$35422 ( \35765 , \35763 , \35764 );
and \U$35423 ( \35766 , \5762 , RI9873288_184);
not \U$35424 ( \35767 , \5762 );
and \U$35425 ( \35768 , \35767 , \24305 );
nor \U$35426 ( \35769 , \35766 , \35768 );
nand \U$35427 ( \35770 , \35769 , \17528 );
nand \U$35428 ( \35771 , \35765 , \35770 );
xor \U$35429 ( \35772 , \35762 , \35771 );
xor \U$35430 ( \35773 , \35709 , \35714 );
and \U$35431 ( \35774 , \35773 , \35725 );
and \U$35432 ( \35775 , \35709 , \35714 );
or \U$35433 ( \35776 , \35774 , \35775 );
xor \U$35434 ( \35777 , \35772 , \35776 );
not \U$35435 ( \35778 , \35135 );
not \U$35436 ( \35779 , \35101 );
or \U$35437 ( \35780 , \35778 , \35779 );
nand \U$35438 ( \35781 , \35780 , \35040 );
nand \U$35439 ( \35782 , \35105 , \35138 );
nand \U$35440 ( \35783 , \35781 , \35782 );
xor \U$35441 ( \35784 , \35777 , \35783 );
or \U$35442 ( \35785 , \35746 , \35784 );
not \U$35443 ( \35786 , \35785 );
not \U$35444 ( \35787 , \13475 );
and \U$35445 ( \35788 , RI9873210_183, \9898 );
not \U$35446 ( \35789 , RI9873210_183);
and \U$35447 ( \35790 , \35789 , \9895 );
nor \U$35448 ( \35791 , \35788 , \35790 );
not \U$35449 ( \35792 , \35791 );
or \U$35450 ( \35793 , \35787 , \35792 );
nand \U$35451 ( \35794 , \34962 , \30963 );
nand \U$35452 ( \35795 , \35793 , \35794 );
not \U$35453 ( \35796 , \35795 );
not \U$35454 ( \35797 , \7325 );
not \U$35455 ( \35798 , RI98729a0_165);
not \U$35456 ( \35799 , \25380 );
or \U$35457 ( \35800 , \35798 , \35799 );
or \U$35458 ( \35801 , \30320 , RI98729a0_165);
nand \U$35459 ( \35802 , \35800 , \35801 );
not \U$35460 ( \35803 , \35802 );
or \U$35461 ( \35804 , \35797 , \35803 );
xor \U$35462 ( \35805 , \35645 , RI98729a0_165);
nand \U$35463 ( \35806 , \35805 , \7338 );
nand \U$35464 ( \35807 , \35804 , \35806 );
not \U$35465 ( \35808 , \35807 );
not \U$35466 ( \35809 , \5032 );
not \U$35467 ( \35810 , RI9872478_154);
not \U$35468 ( \35811 , \21773 );
or \U$35469 ( \35812 , \35810 , \35811 );
nand \U$35470 ( \35813 , \28671 , \5025 );
nand \U$35471 ( \35814 , \35812 , \35813 );
not \U$35472 ( \35815 , \35814 );
or \U$35473 ( \35816 , \35809 , \35815 );
not \U$35474 ( \35817 , \5025 );
not \U$35475 ( \35818 , \18705 );
or \U$35476 ( \35819 , \35817 , \35818 );
or \U$35477 ( \35820 , \25394 , \5025 );
nand \U$35478 ( \35821 , \35819 , \35820 );
nand \U$35479 ( \35822 , \35821 , \5033 );
nand \U$35480 ( \35823 , \35816 , \35822 );
or \U$35481 ( \35824 , RI98724f0_155, RI9872568_156);
nand \U$35482 ( \35825 , \35824 , \18704 );
and \U$35483 ( \35826 , RI98724f0_155, RI9872568_156);
nor \U$35484 ( \35827 , \35826 , \5025 );
and \U$35485 ( \35828 , \35825 , \35827 );
nand \U$35486 ( \35829 , \35823 , \35828 );
not \U$35487 ( \35830 , \35829 );
not \U$35488 ( \35831 , \6282 );
not \U$35489 ( \35832 , RI98728b0_163);
not \U$35490 ( \35833 , \24470 );
or \U$35491 ( \35834 , \35832 , \35833 );
or \U$35492 ( \35835 , \33986 , RI98728b0_163);
nand \U$35493 ( \35836 , \35834 , \35835 );
not \U$35494 ( \35837 , \35836 );
or \U$35495 ( \35838 , \35831 , \35837 );
nand \U$35496 ( \35839 , \34947 , \6285 );
nand \U$35497 ( \35840 , \35838 , \35839 );
not \U$35498 ( \35841 , \35840 );
or \U$35499 ( \35842 , \35830 , \35841 );
or \U$35500 ( \35843 , \35840 , \35829 );
nand \U$35501 ( \35844 , \35842 , \35843 );
not \U$35502 ( \35845 , \35844 );
or \U$35503 ( \35846 , \35808 , \35845 );
not \U$35504 ( \35847 , \35829 );
nand \U$35505 ( \35848 , \35847 , \35840 );
nand \U$35506 ( \35849 , \35846 , \35848 );
not \U$35507 ( \35850 , \12867 );
not \U$35508 ( \35851 , \35212 );
or \U$35509 ( \35852 , \35850 , \35851 );
xor \U$35510 ( \35853 , RI98730a8_180, \8873 );
nand \U$35511 ( \35854 , \35853 , \24209 );
nand \U$35512 ( \35855 , \35852 , \35854 );
xor \U$35513 ( \35856 , \35849 , \35855 );
not \U$35514 ( \35857 , \35856 );
or \U$35515 ( \35858 , \35796 , \35857 );
nand \U$35516 ( \35859 , \35855 , \35849 );
nand \U$35517 ( \35860 , \35858 , \35859 );
not \U$35518 ( \35861 , \35860 );
not \U$35519 ( \35862 , \35098 );
and \U$35520 ( \35863 , \35088 , \35862 );
not \U$35521 ( \35864 , \35088 );
and \U$35522 ( \35865 , \35864 , \35098 );
nor \U$35523 ( \35866 , \35863 , \35865 );
not \U$35524 ( \35867 , \35866 );
xor \U$35525 ( \35868 , \34870 , \34883 );
not \U$35526 ( \35869 , \35868 );
or \U$35527 ( \35870 , \35867 , \35869 );
or \U$35528 ( \35871 , \35868 , \35866 );
nand \U$35529 ( \35872 , \35870 , \35871 );
not \U$35530 ( \35873 , \35872 );
or \U$35531 ( \35874 , \35861 , \35873 );
not \U$35532 ( \35875 , \35866 );
nand \U$35533 ( \35876 , \35875 , \35868 );
nand \U$35534 ( \35877 , \35874 , \35876 );
not \U$35535 ( \35878 , \35877 );
xor \U$35536 ( \35879 , \34949 , \34933 );
not \U$35537 ( \35880 , \35879 );
not \U$35538 ( \35881 , \11198 );
not \U$35539 ( \35882 , \34881 );
or \U$35540 ( \35883 , \35881 , \35882 );
not \U$35541 ( \35884 , \8732 );
not \U$35542 ( \35885 , \12848 );
or \U$35543 ( \35886 , \35884 , \35885 );
or \U$35544 ( \35887 , \8575 , \8732 );
nand \U$35545 ( \35888 , \35886 , \35887 );
nand \U$35546 ( \35889 , \35888 , \8742 );
nand \U$35547 ( \35890 , \35883 , \35889 );
not \U$35548 ( \35891 , \35890 );
nand \U$35549 ( \35892 , \35880 , \35891 );
not \U$35550 ( \35893 , \35892 );
not \U$35551 ( \35894 , \17263 );
not \U$35552 ( \35895 , \35018 );
or \U$35553 ( \35896 , \35894 , \35895 );
and \U$35554 ( \35897 , RI98733f0_187, \12805 );
not \U$35555 ( \35898 , RI98733f0_187);
and \U$35556 ( \35899 , \35898 , \6298 );
or \U$35557 ( \35900 , \35897 , \35899 );
nand \U$35558 ( \35901 , \35900 , \17251 );
nand \U$35559 ( \35902 , \35896 , \35901 );
not \U$35560 ( \35903 , \35902 );
or \U$35561 ( \35904 , \35893 , \35903 );
nand \U$35562 ( \35905 , \35890 , \35879 );
nand \U$35563 ( \35906 , \35904 , \35905 );
not \U$35564 ( \35907 , \35906 );
not \U$35565 ( \35908 , \7338 );
not \U$35566 ( \35909 , \34847 );
or \U$35567 ( \35910 , \35908 , \35909 );
nand \U$35568 ( \35911 , \35805 , \7325 );
nand \U$35569 ( \35912 , \35910 , \35911 );
not \U$35570 ( \35913 , \35912 );
not \U$35571 ( \35914 , \9214 );
not \U$35572 ( \35915 , \34867 );
or \U$35573 ( \35916 , \35914 , \35915 );
and \U$35574 ( \35917 , RI9872b80_169, \11454 );
not \U$35575 ( \35918 , RI9872b80_169);
and \U$35576 ( \35919 , \35918 , \12788 );
nor \U$35577 ( \35920 , \35917 , \35919 );
nand \U$35578 ( \35921 , \35920 , \9195 );
nand \U$35579 ( \35922 , \35916 , \35921 );
not \U$35580 ( \35923 , \35922 );
not \U$35581 ( \35924 , \8039 );
not \U$35582 ( \35925 , \35077 );
or \U$35583 ( \35926 , \35924 , \35925 );
and \U$35584 ( \35927 , RI9872a18_166, \19591 );
not \U$35585 ( \35928 , RI9872a18_166);
and \U$35586 ( \35929 , \35928 , \19594 );
or \U$35587 ( \35930 , \35927 , \35929 );
nand \U$35588 ( \35931 , \35930 , \8027 );
nand \U$35589 ( \35932 , \35926 , \35931 );
not \U$35590 ( \35933 , \35932 );
nand \U$35591 ( \35934 , \35923 , \35933 );
not \U$35592 ( \35935 , \35934 );
or \U$35593 ( \35936 , \35913 , \35935 );
nand \U$35594 ( \35937 , \35922 , \35932 );
nand \U$35595 ( \35938 , \35936 , \35937 );
not \U$35596 ( \35939 , \35938 );
not \U$35597 ( \35940 , \35939 );
not \U$35598 ( \35941 , \17528 );
not \U$35599 ( \35942 , \35009 );
or \U$35600 ( \35943 , \35941 , \35942 );
and \U$35601 ( \35944 , RI9873288_184, \8942 );
not \U$35602 ( \35945 , RI9873288_184);
and \U$35603 ( \35946 , \35945 , \20583 );
nor \U$35604 ( \35947 , \35944 , \35946 );
nand \U$35605 ( \35948 , \35947 , \19641 );
nand \U$35606 ( \35949 , \35943 , \35948 );
not \U$35607 ( \35950 , \10624 );
not \U$35608 ( \35951 , \34896 );
or \U$35609 ( \35952 , \35950 , \35951 );
and \U$35610 ( \35953 , \8811 , \9847 );
not \U$35611 ( \35954 , \8811 );
and \U$35612 ( \35955 , \35954 , \8707 );
nor \U$35613 ( \35956 , \35953 , \35955 );
nand \U$35614 ( \35957 , \35956 , \8818 );
nand \U$35615 ( \35958 , \35952 , \35957 );
nor \U$35616 ( \35959 , \35949 , \35958 );
not \U$35617 ( \35960 , \9273 );
not \U$35618 ( \35961 , \34986 );
or \U$35619 ( \35962 , \35960 , \35961 );
not \U$35620 ( \35963 , RI9872e50_175);
not \U$35621 ( \35964 , \18498 );
or \U$35622 ( \35965 , \35963 , \35964 );
or \U$35623 ( \35966 , \9924 , RI9872e50_175);
nand \U$35624 ( \35967 , \35965 , \35966 );
nand \U$35625 ( \35968 , \35967 , \18563 );
nand \U$35626 ( \35969 , \35962 , \35968 );
not \U$35627 ( \35970 , \35969 );
or \U$35628 ( \35971 , \35959 , \35970 );
nand \U$35629 ( \35972 , \35949 , \35958 );
nand \U$35630 ( \35973 , \35971 , \35972 );
not \U$35631 ( \35974 , \35973 );
or \U$35632 ( \35975 , \35940 , \35974 );
or \U$35633 ( \35976 , \35959 , \35970 );
nand \U$35634 ( \35977 , \35976 , \35938 , \35972 );
nand \U$35635 ( \35978 , \35975 , \35977 );
not \U$35636 ( \35979 , \35978 );
or \U$35637 ( \35980 , \35907 , \35979 );
not \U$35638 ( \35981 , \35939 );
nand \U$35639 ( \35982 , \35981 , \35973 );
nand \U$35640 ( \35983 , \35980 , \35982 );
not \U$35641 ( \35984 , \20626 );
not \U$35642 ( \35985 , \35182 );
or \U$35643 ( \35986 , \35984 , \35985 );
nand \U$35644 ( \35987 , \35723 , RI9873648_192);
nand \U$35645 ( \35988 , \35986 , \35987 );
not \U$35646 ( \35989 , \35988 );
xor \U$35647 ( \35990 , \35496 , \35501 );
not \U$35648 ( \35991 , \5653 );
not \U$35649 ( \35992 , \35491 );
or \U$35650 ( \35993 , \35991 , \35992 );
and \U$35651 ( \35994 , \21553 , \5644 );
not \U$35652 ( \35995 , \21553 );
and \U$35653 ( \35996 , \35995 , RI9872568_156);
nor \U$35654 ( \35997 , \35994 , \35996 );
nand \U$35655 ( \35998 , \35997 , \6063 );
nand \U$35656 ( \35999 , \35993 , \35998 );
not \U$35657 ( \36000 , \5653 );
not \U$35658 ( \36001 , \35997 );
or \U$35659 ( \36002 , \36000 , \36001 );
not \U$35660 ( \36003 , \5644 );
not \U$35661 ( \36004 , \17703 );
or \U$35662 ( \36005 , \36003 , \36004 );
not \U$35663 ( \36006 , \25179 );
nand \U$35664 ( \36007 , \36006 , RI9872568_156);
nand \U$35665 ( \36008 , \36005 , \36007 );
nand \U$35666 ( \36009 , \36008 , \5641 );
nand \U$35667 ( \36010 , \36002 , \36009 );
not \U$35668 ( \36011 , \36010 );
nand \U$35669 ( \36012 , \27523 , \4922 );
not \U$35670 ( \36013 , \36012 );
not \U$35671 ( \36014 , \5032 );
not \U$35672 ( \36015 , \34911 );
or \U$35673 ( \36016 , \36014 , \36015 );
nand \U$35674 ( \36017 , \35814 , \5033 );
nand \U$35675 ( \36018 , \36016 , \36017 );
not \U$35676 ( \36019 , \36018 );
or \U$35677 ( \36020 , \36013 , \36019 );
or \U$35678 ( \36021 , \36018 , \36012 );
nand \U$35679 ( \36022 , \36020 , \36021 );
not \U$35680 ( \36023 , \36022 );
or \U$35681 ( \36024 , \36011 , \36023 );
not \U$35682 ( \36025 , \36012 );
nand \U$35683 ( \36026 , \36025 , \36018 );
nand \U$35684 ( \36027 , \36024 , \36026 );
xor \U$35685 ( \36028 , \35999 , \36027 );
not \U$35686 ( \36029 , \32292 );
and \U$35687 ( \36030 , RI9872bf8_170, \24501 );
not \U$35688 ( \36031 , RI9872bf8_170);
and \U$35689 ( \36032 , \36031 , \13067 );
or \U$35690 ( \36033 , \36030 , \36032 );
not \U$35691 ( \36034 , \36033 );
or \U$35692 ( \36035 , \36029 , \36034 );
nand \U$35693 ( \36036 , \35093 , \9227 );
nand \U$35694 ( \36037 , \36035 , \36036 );
and \U$35695 ( \36038 , \36028 , \36037 );
and \U$35696 ( \36039 , \35999 , \36027 );
or \U$35697 ( \36040 , \36038 , \36039 );
xor \U$35698 ( \36041 , \35990 , \36040 );
not \U$35699 ( \36042 , \36041 );
or \U$35700 ( \36043 , \35989 , \36042 );
nand \U$35701 ( \36044 , \36040 , \35990 );
nand \U$35702 ( \36045 , \36043 , \36044 );
and \U$35703 ( \36046 , \35983 , \36045 );
not \U$35704 ( \36047 , \35983 );
not \U$35705 ( \36048 , \36045 );
and \U$35706 ( \36049 , \36047 , \36048 );
nor \U$35707 ( \36050 , \36046 , \36049 );
not \U$35708 ( \36051 , \36050 );
or \U$35709 ( \36052 , \35878 , \36051 );
nand \U$35710 ( \36053 , \35983 , \36045 );
nand \U$35711 ( \36054 , \36052 , \36053 );
not \U$35712 ( \36055 , \36054 );
or \U$35713 ( \36056 , \35786 , \36055 );
nand \U$35714 ( \36057 , \35746 , \35784 );
nand \U$35715 ( \36058 , \36056 , \36057 );
not \U$35716 ( \36059 , \36058 );
xor \U$35717 ( \36060 , \35772 , \35776 );
and \U$35718 ( \36061 , \36060 , \35783 );
and \U$35719 ( \36062 , \35772 , \35776 );
or \U$35720 ( \36063 , \36061 , \36062 );
not \U$35721 ( \36064 , \8802 );
not \U$35722 ( \36065 , RI9872d60_173);
not \U$35723 ( \36066 , \8650 );
or \U$35724 ( \36067 , \36065 , \36066 );
or \U$35725 ( \36068 , \8650 , RI9872d60_173);
nand \U$35726 ( \36069 , \36067 , \36068 );
not \U$35727 ( \36070 , \36069 );
or \U$35728 ( \36071 , \36064 , \36070 );
nand \U$35729 ( \36072 , \35249 , \9312 );
nand \U$35730 ( \36073 , \36071 , \36072 );
not \U$35731 ( \36074 , \36073 );
not \U$35732 ( \36075 , \36074 );
xor \U$35733 ( \36076 , \35631 , \35640 );
and \U$35734 ( \36077 , \36076 , \35648 );
and \U$35735 ( \36078 , \35631 , \35640 );
nor \U$35736 ( \36079 , \36077 , \36078 );
not \U$35737 ( \36080 , \36079 );
not \U$35738 ( \36081 , \9668 );
and \U$35739 ( \36082 , \8554 , \9185 );
not \U$35740 ( \36083 , \8554 );
and \U$35741 ( \36084 , \36083 , RI9872bf8_170);
nor \U$35742 ( \36085 , \36082 , \36084 );
not \U$35743 ( \36086 , \36085 );
or \U$35744 ( \36087 , \36081 , \36086 );
nand \U$35745 ( \36088 , \35757 , \9249 );
nand \U$35746 ( \36089 , \36087 , \36088 );
not \U$35747 ( \36090 , \36089 );
or \U$35748 ( \36091 , \36080 , \36090 );
or \U$35749 ( \36092 , \36089 , \36079 );
nand \U$35750 ( \36093 , \36091 , \36092 );
buf \U$35751 ( \36094 , \36093 );
not \U$35752 ( \36095 , \36094 );
or \U$35753 ( \36096 , \36075 , \36095 );
or \U$35754 ( \36097 , \36094 , \36074 );
nand \U$35755 ( \36098 , \36096 , \36097 );
not \U$35756 ( \36099 , \17528 );
and \U$35757 ( \36100 , \7028 , RI9873288_184);
not \U$35758 ( \36101 , \7028 );
and \U$35759 ( \36102 , \36101 , \22727 );
nor \U$35760 ( \36103 , \36100 , \36102 );
not \U$35761 ( \36104 , \36103 );
or \U$35762 ( \36105 , \36099 , \36104 );
nand \U$35763 ( \36106 , \35769 , \18508 );
nand \U$35764 ( \36107 , \36105 , \36106 );
not \U$35765 ( \36108 , \22670 );
not \U$35766 ( \36109 , RI9873210_183);
not \U$35767 ( \36110 , \28258 );
or \U$35768 ( \36111 , \36109 , \36110 );
nand \U$35769 ( \36112 , \6309 , \18012 );
nand \U$35770 ( \36113 , \36111 , \36112 );
not \U$35771 ( \36114 , \36113 );
or \U$35772 ( \36115 , \36108 , \36114 );
nand \U$35773 ( \36116 , \35326 , \18957 );
nand \U$35774 ( \36117 , \36115 , \36116 );
xor \U$35775 ( \36118 , \36107 , \36117 );
not \U$35776 ( \36119 , \20626 );
not \U$35777 ( \36120 , \35664 );
or \U$35778 ( \36121 , \36119 , \36120 );
not \U$35779 ( \36122 , \18239 );
not \U$35780 ( \36123 , \10698 );
or \U$35781 ( \36124 , \36122 , \36123 );
nand \U$35782 ( \36125 , \3568 , RI9873558_190);
nand \U$35783 ( \36126 , \36124 , \36125 );
nand \U$35784 ( \36127 , \36126 , RI9873648_192);
nand \U$35785 ( \36128 , \36121 , \36127 );
xor \U$35786 ( \36129 , \36118 , \36128 );
xor \U$35787 ( \36130 , \36098 , \36129 );
not \U$35788 ( \36131 , \13017 );
not \U$35789 ( \36132 , RI9872a18_166);
not \U$35790 ( \36133 , \31511 );
or \U$35791 ( \36134 , \36132 , \36133 );
or \U$35792 ( \36135 , \9114 , RI9872a18_166);
nand \U$35793 ( \36136 , \36134 , \36135 );
not \U$35794 ( \36137 , \36136 );
or \U$35795 ( \36138 , \36131 , \36137 );
nand \U$35796 ( \36139 , \35564 , \8027 );
nand \U$35797 ( \36140 , \36138 , \36139 );
not \U$35798 ( \36141 , \5035 );
not \U$35799 ( \36142 , \34248 );
or \U$35800 ( \36143 , \36141 , \36142 );
nand \U$35801 ( \36144 , \35636 , \5034 );
nand \U$35802 ( \36145 , \36143 , \36144 );
not \U$35803 ( \36146 , \35554 );
not \U$35804 ( \36147 , \35544 );
or \U$35805 ( \36148 , \36146 , \36147 );
nand \U$35806 ( \36149 , \35538 , \35539 );
nand \U$35807 ( \36150 , \36148 , \36149 );
xor \U$35808 ( \36151 , \36145 , \36150 );
xor \U$35809 ( \36152 , \36140 , \36151 );
not \U$35810 ( \36153 , \19282 );
xnor \U$35811 ( \36154 , \7007 , RI98733f0_187);
not \U$35812 ( \36155 , \36154 );
or \U$35813 ( \36156 , \36153 , \36155 );
nand \U$35814 ( \36157 , \35654 , \17251 );
nand \U$35815 ( \36158 , \36156 , \36157 );
xor \U$35816 ( \36159 , \36152 , \36158 );
not \U$35817 ( \36160 , \20147 );
not \U$35818 ( \36161 , \16999 );
not \U$35819 ( \36162 , \15685 );
or \U$35820 ( \36163 , \36161 , \36162 );
or \U$35821 ( \36164 , \12145 , \19361 );
nand \U$35822 ( \36165 , \36163 , \36164 );
not \U$35823 ( \36166 , \36165 );
or \U$35824 ( \36167 , \36160 , \36166 );
nand \U$35825 ( \36168 , \35376 , \19036 );
nand \U$35826 ( \36169 , \36167 , \36168 );
xor \U$35827 ( \36170 , \36159 , \36169 );
xor \U$35828 ( \36171 , \36130 , \36170 );
xor \U$35829 ( \36172 , \36063 , \36171 );
not \U$35830 ( \36173 , \35679 );
nor \U$35831 ( \36174 , \36173 , \35674 );
or \U$35832 ( \36175 , \36174 , \35698 );
nand \U$35833 ( \36176 , \36173 , \35674 );
nand \U$35834 ( \36177 , \36175 , \36176 );
xnor \U$35835 ( \36178 , \36172 , \36177 );
not \U$35836 ( \36179 , \36178 );
or \U$35837 ( \36180 , \36059 , \36179 );
or \U$35838 ( \36181 , \36178 , \36058 );
nand \U$35839 ( \36182 , \36180 , \36181 );
not \U$35840 ( \36183 , \36182 );
or \U$35841 ( \36184 , \35704 , \36183 );
or \U$35842 ( \36185 , \36182 , \35703 );
nand \U$35843 ( \36186 , \36184 , \36185 );
not \U$35844 ( \36187 , \36186 );
xnor \U$35845 ( \36188 , \36041 , \35988 );
not \U$35846 ( \36189 , \36188 );
xor \U$35847 ( \36190 , \34955 , \34898 );
xnor \U$35848 ( \36191 , \36190 , \34971 );
not \U$35849 ( \36192 , \36191 );
not \U$35850 ( \36193 , \36192 );
or \U$35851 ( \36194 , \36189 , \36193 );
xor \U$35852 ( \36195 , \35999 , \36027 );
xor \U$35853 ( \36196 , \36195 , \36037 );
not \U$35854 ( \36197 , \9071 );
not \U$35855 ( \36198 , \35930 );
or \U$35856 ( \36199 , \36197 , \36198 );
and \U$35857 ( \36200 , \8031 , \17783 );
not \U$35858 ( \36201 , \8031 );
and \U$35859 ( \36202 , \36201 , \24757 );
nor \U$35860 ( \36203 , \36200 , \36202 );
nand \U$35861 ( \36204 , \36203 , \8027 );
nand \U$35862 ( \36205 , \36199 , \36204 );
not \U$35863 ( \36206 , \36205 );
not \U$35864 ( \36207 , \36022 );
not \U$35865 ( \36208 , \36010 );
not \U$35866 ( \36209 , \36208 );
and \U$35867 ( \36210 , \36207 , \36209 );
and \U$35868 ( \36211 , \36022 , \36208 );
nor \U$35869 ( \36212 , \36210 , \36211 );
not \U$35870 ( \36213 , \36212 );
or \U$35871 ( \36214 , \36206 , \36213 );
or \U$35872 ( \36215 , \36205 , \36212 );
nand \U$35873 ( \36216 , \36214 , \36215 );
not \U$35874 ( \36217 , \36216 );
not \U$35875 ( \36218 , \22167 );
not \U$35876 ( \36219 , \36033 );
or \U$35877 ( \36220 , \36218 , \36219 );
not \U$35878 ( \36221 , \13391 );
not \U$35879 ( \36222 , RI9872bf8_170);
and \U$35880 ( \36223 , \36221 , \36222 );
and \U$35881 ( \36224 , \27588 , RI9872bf8_170);
nor \U$35882 ( \36225 , \36223 , \36224 );
not \U$35883 ( \36226 , \36225 );
nand \U$35884 ( \36227 , \36226 , \9249 );
nand \U$35885 ( \36228 , \36220 , \36227 );
not \U$35886 ( \36229 , \36228 );
or \U$35887 ( \36230 , \36217 , \36229 );
not \U$35888 ( \36231 , \36212 );
nand \U$35889 ( \36232 , \36231 , \36205 );
nand \U$35890 ( \36233 , \36230 , \36232 );
or \U$35891 ( \36234 , \36196 , \36233 );
not \U$35892 ( \36235 , \36234 );
not \U$35893 ( \36236 , \13020 );
and \U$35894 ( \36237 , \18111 , \13022 );
not \U$35895 ( \36238 , \18111 );
and \U$35896 ( \36239 , \36238 , RI98730a8_180);
nor \U$35897 ( \36240 , \36237 , \36239 );
not \U$35898 ( \36241 , \36240 );
or \U$35899 ( \36242 , \36236 , \36241 );
nand \U$35900 ( \36243 , \35853 , \12867 );
nand \U$35901 ( \36244 , \36242 , \36243 );
not \U$35902 ( \36245 , \36244 );
xor \U$35903 ( \36246 , \35823 , \35828 );
not \U$35904 ( \36247 , \36246 );
not \U$35905 ( \36248 , \5653 );
not \U$35906 ( \36249 , \36008 );
or \U$35907 ( \36250 , \36248 , \36249 );
and \U$35908 ( \36251 , \17862 , RI9872568_156);
not \U$35909 ( \36252 , \17862 );
and \U$35910 ( \36253 , \36252 , \5648 );
nor \U$35911 ( \36254 , \36251 , \36253 );
nand \U$35912 ( \36255 , \36254 , \5641 );
nand \U$35913 ( \36256 , \36250 , \36255 );
not \U$35914 ( \36257 , \36256 );
not \U$35915 ( \36258 , \36257 );
or \U$35916 ( \36259 , \36247 , \36258 );
or \U$35917 ( \36260 , \36257 , \36246 );
nand \U$35918 ( \36261 , \36259 , \36260 );
not \U$35919 ( \36262 , \36261 );
not \U$35920 ( \36263 , \7338 );
not \U$35921 ( \36264 , \35802 );
or \U$35922 ( \36265 , \36263 , \36264 );
not \U$35923 ( \36266 , \7333 );
not \U$35924 ( \36267 , \28191 );
or \U$35925 ( \36268 , \36266 , \36267 );
nand \U$35926 ( \36269 , \17911 , RI98729a0_165);
nand \U$35927 ( \36270 , \36268 , \36269 );
nand \U$35928 ( \36271 , \36270 , \7325 );
nand \U$35929 ( \36272 , \36265 , \36271 );
not \U$35930 ( \36273 , \36272 );
or \U$35931 ( \36274 , \36262 , \36273 );
nand \U$35932 ( \36275 , \36246 , \36256 );
nand \U$35933 ( \36276 , \36274 , \36275 );
not \U$35934 ( \36277 , \36276 );
not \U$35935 ( \36278 , \36277 );
not \U$35936 ( \36279 , \18508 );
not \U$35937 ( \36280 , RI9873288_184);
not \U$35938 ( \36281 , \21642 );
or \U$35939 ( \36282 , \36280 , \36281 );
or \U$35940 ( \36283 , \17440 , RI9873288_184);
nand \U$35941 ( \36284 , \36282 , \36283 );
not \U$35942 ( \36285 , \36284 );
or \U$35943 ( \36286 , \36279 , \36285 );
nand \U$35944 ( \36287 , \35947 , \17528 );
nand \U$35945 ( \36288 , \36286 , \36287 );
not \U$35946 ( \36289 , \36288 );
or \U$35947 ( \36290 , \36278 , \36289 );
or \U$35948 ( \36291 , \36288 , \36277 );
nand \U$35949 ( \36292 , \36290 , \36291 );
not \U$35950 ( \36293 , \36292 );
or \U$35951 ( \36294 , \36245 , \36293 );
not \U$35952 ( \36295 , \36277 );
nand \U$35953 ( \36296 , \36295 , \36288 );
nand \U$35954 ( \36297 , \36294 , \36296 );
not \U$35955 ( \36298 , \36297 );
or \U$35956 ( \36299 , \36235 , \36298 );
nand \U$35957 ( \36300 , \36196 , \36233 );
nand \U$35958 ( \36301 , \36299 , \36300 );
nand \U$35959 ( \36302 , \36194 , \36301 );
not \U$35960 ( \36303 , \36188 );
nand \U$35961 ( \36304 , \36303 , \36191 );
and \U$35962 ( \36305 , \36302 , \36304 );
not \U$35963 ( \36306 , \36305 );
xor \U$35964 ( \36307 , \35480 , \35426 );
not \U$35965 ( \36308 , \36307 );
not \U$35966 ( \36309 , \35726 );
not \U$35967 ( \36310 , \35741 );
not \U$35968 ( \36311 , \36310 );
or \U$35969 ( \36312 , \36309 , \36311 );
not \U$35970 ( \36313 , \35726 );
nand \U$35971 ( \36314 , \36313 , \35741 );
nand \U$35972 ( \36315 , \36312 , \36314 );
not \U$35973 ( \36316 , \36315 );
nand \U$35974 ( \36317 , \36308 , \36316 );
nand \U$35975 ( \36318 , \36306 , \36317 );
not \U$35976 ( \36319 , \36316 );
nand \U$35977 ( \36320 , \36319 , \36307 );
nand \U$35978 ( \36321 , \36318 , \36320 );
not \U$35979 ( \36322 , \36321 );
not \U$35980 ( \36323 , \35746 );
not \U$35981 ( \36324 , \35784 );
and \U$35982 ( \36325 , \36323 , \36324 );
and \U$35983 ( \36326 , \35746 , \35784 );
nor \U$35984 ( \36327 , \36325 , \36326 );
not \U$35985 ( \36328 , \36327 );
not \U$35986 ( \36329 , \36054 );
or \U$35987 ( \36330 , \36328 , \36329 );
or \U$35988 ( \36331 , \36054 , \36327 );
nand \U$35989 ( \36332 , \36330 , \36331 );
nand \U$35990 ( \36333 , \36322 , \36332 );
xor \U$35991 ( \36334 , \35872 , \35860 );
not \U$35992 ( \36335 , \36334 );
xor \U$35993 ( \36336 , \35912 , \35933 );
xnor \U$35994 ( \36337 , \36336 , \35922 );
not \U$35995 ( \36338 , \9526 );
not \U$35996 ( \36339 , RI9872f40_177);
not \U$35997 ( \36340 , \10369 );
or \U$35998 ( \36341 , \36339 , \36340 );
or \U$35999 ( \36342 , \8555 , RI9872f40_177);
nand \U$36000 ( \36343 , \36341 , \36342 );
not \U$36001 ( \36344 , \36343 );
or \U$36002 ( \36345 , \36338 , \36344 );
nand \U$36003 ( \36346 , \35888 , \11198 );
nand \U$36004 ( \36347 , \36345 , \36346 );
not \U$36005 ( \36348 , \36347 );
not \U$36006 ( \36349 , \9195 );
not \U$36007 ( \36350 , RI9872b80_169);
not \U$36008 ( \36351 , \13268 );
or \U$36009 ( \36352 , \36350 , \36351 );
or \U$36010 ( \36353 , \13268 , RI9872b80_169);
nand \U$36011 ( \36354 , \36352 , \36353 );
not \U$36012 ( \36355 , \36354 );
or \U$36013 ( \36356 , \36349 , \36355 );
nand \U$36014 ( \36357 , \35920 , \9214 );
nand \U$36015 ( \36358 , \36356 , \36357 );
not \U$36016 ( \36359 , \8817 );
and \U$36017 ( \36360 , RI9872d60_173, \17897 );
not \U$36018 ( \36361 , RI9872d60_173);
and \U$36019 ( \36362 , \36361 , \9113 );
nor \U$36020 ( \36363 , \36360 , \36362 );
not \U$36021 ( \36364 , \36363 );
or \U$36022 ( \36365 , \36359 , \36364 );
nand \U$36023 ( \36366 , \35956 , \8800 );
nand \U$36024 ( \36367 , \36365 , \36366 );
xor \U$36025 ( \36368 , \36358 , \36367 );
not \U$36026 ( \36369 , \36368 );
or \U$36027 ( \36370 , \36348 , \36369 );
nand \U$36028 ( \36371 , \36367 , \36358 );
nand \U$36029 ( \36372 , \36370 , \36371 );
not \U$36030 ( \36373 , \36372 );
and \U$36031 ( \36374 , \36337 , \36373 );
not \U$36032 ( \36375 , \36337 );
and \U$36033 ( \36376 , \36375 , \36372 );
nor \U$36034 ( \36377 , \36374 , \36376 );
not \U$36035 ( \36378 , \36377 );
not \U$36036 ( \36379 , \36378 );
not \U$36037 ( \36380 , \18562 );
not \U$36038 ( \36381 , \9690 );
not \U$36039 ( \36382 , \9750 );
or \U$36040 ( \36383 , \36381 , \36382 );
or \U$36041 ( \36384 , \9750 , \9690 );
nand \U$36042 ( \36385 , \36383 , \36384 );
not \U$36043 ( \36386 , \36385 );
or \U$36044 ( \36387 , \36380 , \36386 );
nand \U$36045 ( \36388 , \35967 , \9272 );
nand \U$36046 ( \36389 , \36387 , \36388 );
not \U$36047 ( \36390 , \13475 );
and \U$36048 ( \36391 , RI9873210_183, \13358 );
not \U$36049 ( \36392 , RI9873210_183);
and \U$36050 ( \36393 , \36392 , \11628 );
nor \U$36051 ( \36394 , \36391 , \36393 );
not \U$36052 ( \36395 , \36394 );
or \U$36053 ( \36396 , \36390 , \36395 );
nand \U$36054 ( \36397 , \35791 , \33922 );
nand \U$36055 ( \36398 , \36396 , \36397 );
xor \U$36056 ( \36399 , \36389 , \36398 );
not \U$36057 ( \36400 , RI98734e0_189);
not \U$36058 ( \36401 , \11435 );
or \U$36059 ( \36402 , \36400 , \36401 );
not \U$36060 ( \36403 , \11435 );
nand \U$36061 ( \36404 , \36403 , \16999 );
nand \U$36062 ( \36405 , \36402 , \36404 );
not \U$36063 ( \36406 , \36405 );
not \U$36064 ( \36407 , \19036 );
or \U$36065 ( \36408 , \36406 , \36407 );
nand \U$36066 ( \36409 , \35155 , \19046 );
nand \U$36067 ( \36410 , \36408 , \36409 );
and \U$36068 ( \36411 , \36399 , \36410 );
and \U$36069 ( \36412 , \36389 , \36398 );
or \U$36070 ( \36413 , \36411 , \36412 );
not \U$36071 ( \36414 , \36413 );
or \U$36072 ( \36415 , \36379 , \36414 );
not \U$36073 ( \36416 , \36373 );
nand \U$36074 ( \36417 , \36416 , \36337 );
nand \U$36075 ( \36418 , \36415 , \36417 );
not \U$36076 ( \36419 , \36418 );
not \U$36077 ( \36420 , \36419 );
not \U$36078 ( \36421 , \35795 );
not \U$36079 ( \36422 , \35856 );
not \U$36080 ( \36423 , \36422 );
or \U$36081 ( \36424 , \36421 , \36423 );
not \U$36082 ( \36425 , \35795 );
nand \U$36083 ( \36426 , \36425 , \35856 );
nand \U$36084 ( \36427 , \36424 , \36426 );
not \U$36085 ( \36428 , \36427 );
and \U$36086 ( \36429 , \35879 , \35890 );
not \U$36087 ( \36430 , \35879 );
and \U$36088 ( \36431 , \36430 , \35891 );
nor \U$36089 ( \36432 , \36429 , \36431 );
not \U$36090 ( \36433 , \36432 );
not \U$36091 ( \36434 , \36433 );
not \U$36092 ( \36435 , \35902 );
not \U$36093 ( \36436 , \36435 );
or \U$36094 ( \36437 , \36434 , \36436 );
nand \U$36095 ( \36438 , \36432 , \35902 );
nand \U$36096 ( \36439 , \36437 , \36438 );
not \U$36097 ( \36440 , \36439 );
not \U$36098 ( \36441 , \36440 );
or \U$36099 ( \36442 , \36428 , \36441 );
not \U$36100 ( \36443 , \36427 );
not \U$36101 ( \36444 , \36443 );
not \U$36102 ( \36445 , \36439 );
or \U$36103 ( \36446 , \36444 , \36445 );
xor \U$36104 ( \36447 , \35969 , \35958 );
xor \U$36105 ( \36448 , \36447 , \35949 );
nand \U$36106 ( \36449 , \36446 , \36448 );
nand \U$36107 ( \36450 , \36442 , \36449 );
not \U$36108 ( \36451 , \36450 );
or \U$36109 ( \36452 , \36420 , \36451 );
or \U$36110 ( \36453 , \36450 , \36419 );
nand \U$36111 ( \36454 , \36452 , \36453 );
not \U$36112 ( \36455 , \36454 );
or \U$36113 ( \36456 , \36335 , \36455 );
nand \U$36114 ( \36457 , \36418 , \36450 );
nand \U$36115 ( \36458 , \36456 , \36457 );
not \U$36116 ( \36459 , \36458 );
not \U$36117 ( \36460 , \36459 );
xor \U$36118 ( \36461 , \36048 , \35877 );
xor \U$36119 ( \36462 , \36461 , \35983 );
not \U$36120 ( \36463 , \36462 );
or \U$36121 ( \36464 , \36460 , \36463 );
not \U$36122 ( \36465 , \35193 );
not \U$36123 ( \36466 , \35227 );
or \U$36124 ( \36467 , \36465 , \36466 );
or \U$36125 ( \36468 , \35227 , \35193 );
nand \U$36126 ( \36469 , \36467 , \36468 );
not \U$36127 ( \36470 , \36469 );
not \U$36128 ( \36471 , \35196 );
and \U$36129 ( \36472 , \36470 , \36471 );
and \U$36130 ( \36473 , \35196 , \36469 );
nor \U$36131 ( \36474 , \36472 , \36473 );
xnor \U$36132 ( \36475 , \35978 , \35906 );
nand \U$36133 ( \36476 , \36474 , \36475 );
not \U$36134 ( \36477 , \36476 );
not \U$36135 ( \36478 , RI9873648_192);
not \U$36136 ( \36479 , \35189 );
or \U$36137 ( \36480 , \36478 , \36479 );
not \U$36138 ( \36481 , RI9873558_190);
not \U$36139 ( \36482 , \5775 );
or \U$36140 ( \36483 , \36481 , \36482 );
or \U$36141 ( \36484 , \5775 , RI9873558_190);
nand \U$36142 ( \36485 , \36483 , \36484 );
nand \U$36143 ( \36486 , \36485 , \18544 );
nand \U$36144 ( \36487 , \36480 , \36486 );
not \U$36145 ( \36488 , \36487 );
not \U$36146 ( \36489 , \17251 );
xnor \U$36147 ( \36490 , \6529 , RI98733f0_187);
not \U$36148 ( \36491 , \36490 );
or \U$36149 ( \36492 , \36489 , \36491 );
nand \U$36150 ( \36493 , \35900 , \17263 );
nand \U$36151 ( \36494 , \36492 , \36493 );
not \U$36152 ( \36495 , \13109 );
not \U$36153 ( \36496 , RI9873030_179);
not \U$36154 ( \36497 , \8650 );
or \U$36155 ( \36498 , \36496 , \36497 );
or \U$36156 ( \36499 , \8650 , RI9873030_179);
nand \U$36157 ( \36500 , \36498 , \36499 );
not \U$36158 ( \36501 , \36500 );
or \U$36159 ( \36502 , \36495 , \36501 );
nand \U$36160 ( \36503 , \35164 , \9937 );
nand \U$36161 ( \36504 , \36502 , \36503 );
or \U$36162 ( \36505 , \36494 , \36504 );
not \U$36163 ( \36506 , \36505 );
or \U$36164 ( \36507 , \36488 , \36506 );
nand \U$36165 ( \36508 , \36494 , \36504 );
nand \U$36166 ( \36509 , \36507 , \36508 );
not \U$36167 ( \36510 , \36509 );
xor \U$36168 ( \36511 , \35844 , \35807 );
not \U$36169 ( \36512 , \6285 );
and \U$36170 ( \36513 , RI98728b0_163, \23924 );
not \U$36171 ( \36514 , RI98728b0_163);
not \U$36172 ( \36515 , \21553 );
and \U$36173 ( \36516 , \36514 , \36515 );
or \U$36174 ( \36517 , \36513 , \36516 );
not \U$36175 ( \36518 , \36517 );
or \U$36176 ( \36519 , \36512 , \36518 );
not \U$36177 ( \36520 , \5632 );
not \U$36178 ( \36521 , \25179 );
or \U$36179 ( \36522 , \36520 , \36521 );
nand \U$36180 ( \36523 , \28657 , RI98728b0_163);
nand \U$36181 ( \36524 , \36522 , \36523 );
nand \U$36182 ( \36525 , \36524 , \6282 );
nand \U$36183 ( \36526 , \36519 , \36525 );
not \U$36184 ( \36527 , \36526 );
nand \U$36185 ( \36528 , \18704 , \5032 );
not \U$36186 ( \36529 , \36528 );
not \U$36187 ( \36530 , \5653 );
not \U$36188 ( \36531 , \36254 );
or \U$36189 ( \36532 , \36530 , \36531 );
xor \U$36190 ( \36533 , \23948 , RI9872568_156);
nand \U$36191 ( \36534 , \36533 , \5641 );
nand \U$36192 ( \36535 , \36532 , \36534 );
not \U$36193 ( \36536 , \36535 );
or \U$36194 ( \36537 , \36529 , \36536 );
or \U$36195 ( \36538 , \36535 , \36528 );
nand \U$36196 ( \36539 , \36537 , \36538 );
not \U$36197 ( \36540 , \36539 );
or \U$36198 ( \36541 , \36527 , \36540 );
not \U$36199 ( \36542 , \36528 );
nand \U$36200 ( \36543 , \36542 , \36535 );
nand \U$36201 ( \36544 , \36541 , \36543 );
not \U$36202 ( \36545 , \36544 );
not \U$36203 ( \36546 , \6285 );
not \U$36204 ( \36547 , \35836 );
or \U$36205 ( \36548 , \36546 , \36547 );
nand \U$36206 ( \36549 , \36517 , \6282 );
nand \U$36207 ( \36550 , \36548 , \36549 );
not \U$36208 ( \36551 , \36550 );
not \U$36209 ( \36552 , \36551 );
and \U$36210 ( \36553 , \36545 , \36552 );
and \U$36211 ( \36554 , \36544 , \36551 );
nor \U$36212 ( \36555 , \36553 , \36554 );
not \U$36213 ( \36556 , \36555 );
not \U$36214 ( \36557 , \36556 );
not \U$36215 ( \36558 , RI9872bf8_170);
not \U$36216 ( \36559 , \18151 );
or \U$36217 ( \36560 , \36558 , \36559 );
or \U$36218 ( \36561 , \18155 , RI9872bf8_170);
nand \U$36219 ( \36562 , \36560 , \36561 );
not \U$36220 ( \36563 , \36562 );
not \U$36221 ( \36564 , \9249 );
or \U$36222 ( \36565 , \36563 , \36564 );
not \U$36223 ( \36566 , \9226 );
or \U$36224 ( \36567 , \36225 , \36566 );
nand \U$36225 ( \36568 , \36565 , \36567 );
not \U$36226 ( \36569 , \36568 );
or \U$36227 ( \36570 , \36557 , \36569 );
nand \U$36228 ( \36571 , \36544 , \36550 );
nand \U$36229 ( \36572 , \36570 , \36571 );
xor \U$36230 ( \36573 , \36511 , \36572 );
not \U$36231 ( \36574 , \36203 );
not \U$36232 ( \36575 , \9071 );
or \U$36233 ( \36576 , \36574 , \36575 );
and \U$36234 ( \36577 , RI9872a18_166, \17013 );
not \U$36235 ( \36578 , RI9872a18_166);
and \U$36236 ( \36579 , \36578 , \17014 );
or \U$36237 ( \36580 , \36577 , \36579 );
not \U$36238 ( \36581 , \36580 );
not \U$36239 ( \36582 , \8027 );
or \U$36240 ( \36583 , \36581 , \36582 );
nand \U$36241 ( \36584 , \36576 , \36583 );
not \U$36242 ( \36585 , \36584 );
not \U$36243 ( \36586 , \8800 );
not \U$36244 ( \36587 , \36363 );
or \U$36245 ( \36588 , \36586 , \36587 );
xor \U$36246 ( \36589 , RI9872d60_173, \9138 );
nand \U$36247 ( \36590 , \36589 , \8818 );
nand \U$36248 ( \36591 , \36588 , \36590 );
not \U$36249 ( \36592 , \36591 );
or \U$36250 ( \36593 , \36585 , \36592 );
not \U$36251 ( \36594 , \36584 );
not \U$36252 ( \36595 , \36591 );
not \U$36253 ( \36596 , \36595 );
or \U$36254 ( \36597 , \36594 , \36596 );
or \U$36255 ( \36598 , \36595 , \36584 );
nand \U$36256 ( \36599 , \36597 , \36598 );
not \U$36257 ( \36600 , \36599 );
and \U$36258 ( \36601 , \9214 , \36354 );
not \U$36259 ( \36602 , RI9872b80_169);
not \U$36260 ( \36603 , \17090 );
or \U$36261 ( \36604 , \36602 , \36603 );
or \U$36262 ( \36605 , \24523 , RI9872b80_169);
nand \U$36263 ( \36606 , \36604 , \36605 );
and \U$36264 ( \36607 , \36606 , \9196 );
nor \U$36265 ( \36608 , \36601 , \36607 );
or \U$36266 ( \36609 , \36600 , \36608 );
nand \U$36267 ( \36610 , \36593 , \36609 );
and \U$36268 ( \36611 , \36573 , \36610 );
and \U$36269 ( \36612 , \36511 , \36572 );
or \U$36270 ( \36613 , \36611 , \36612 );
not \U$36271 ( \36614 , \36613 );
nand \U$36272 ( \36615 , \36510 , \36614 );
not \U$36273 ( \36616 , \36615 );
and \U$36274 ( \36617 , \35173 , \35157 );
not \U$36275 ( \36618 , \35173 );
not \U$36276 ( \36619 , \35157 );
and \U$36277 ( \36620 , \36618 , \36619 );
nor \U$36278 ( \36621 , \36617 , \36620 );
and \U$36279 ( \36622 , \36621 , \35191 );
not \U$36280 ( \36623 , \36621 );
not \U$36281 ( \36624 , \35191 );
and \U$36282 ( \36625 , \36623 , \36624 );
nor \U$36283 ( \36626 , \36622 , \36625 );
not \U$36284 ( \36627 , \36626 );
or \U$36285 ( \36628 , \36616 , \36627 );
nand \U$36286 ( \36629 , \36509 , \36613 );
nand \U$36287 ( \36630 , \36628 , \36629 );
not \U$36288 ( \36631 , \36630 );
or \U$36289 ( \36632 , \36477 , \36631 );
not \U$36290 ( \36633 , \36475 );
not \U$36291 ( \36634 , \36474 );
nand \U$36292 ( \36635 , \36633 , \36634 );
nand \U$36293 ( \36636 , \36632 , \36635 );
nand \U$36294 ( \36637 , \36464 , \36636 );
not \U$36295 ( \36638 , \36462 );
nand \U$36296 ( \36639 , \36638 , \36458 );
nand \U$36297 ( \36640 , \36637 , \36639 );
nand \U$36298 ( \36641 , \36333 , \36640 );
not \U$36299 ( \36642 , \36332 );
nand \U$36300 ( \36643 , \36642 , \36321 );
nand \U$36301 ( \36644 , \36641 , \36643 );
not \U$36302 ( \36645 , \36644 );
xor \U$36303 ( \36646 , \35251 , \35266 );
and \U$36304 ( \36647 , \36646 , \35282 );
and \U$36305 ( \36648 , \35251 , \35266 );
or \U$36306 ( \36649 , \36647 , \36648 );
xor \U$36307 ( \36650 , \35752 , \35761 );
and \U$36308 ( \36651 , \36650 , \35771 );
and \U$36309 ( \36652 , \35752 , \35761 );
or \U$36310 ( \36653 , \36651 , \36652 );
not \U$36311 ( \36654 , \36653 );
and \U$36312 ( \36655 , \36649 , \36654 );
not \U$36313 ( \36656 , \36649 );
and \U$36314 ( \36657 , \36656 , \36653 );
or \U$36315 ( \36658 , \36655 , \36657 );
not \U$36316 ( \36659 , \9214 );
and \U$36317 ( \36660 , RI9872b80_169, \24807 );
not \U$36318 ( \36661 , RI9872b80_169);
and \U$36319 ( \36662 , \36661 , \9750 );
or \U$36320 ( \36663 , \36660 , \36662 );
not \U$36321 ( \36664 , \36663 );
or \U$36322 ( \36665 , \36659 , \36664 );
nand \U$36323 ( \36666 , \35574 , \9195 );
nand \U$36324 ( \36667 , \36665 , \36666 );
not \U$36325 ( \36668 , \9952 );
not \U$36326 ( \36669 , \35357 );
or \U$36327 ( \36670 , \36668 , \36669 );
and \U$36328 ( \36671 , \13824 , \14132 );
not \U$36329 ( \36672 , \13824 );
and \U$36330 ( \36673 , \36672 , RI9873030_179);
nor \U$36331 ( \36674 , \36671 , \36673 );
nand \U$36332 ( \36675 , \36674 , \9937 );
nand \U$36333 ( \36676 , \36670 , \36675 );
xor \U$36334 ( \36677 , \36667 , \36676 );
not \U$36335 ( \36678 , \22618 );
not \U$36336 ( \36679 , \13022 );
not \U$36337 ( \36680 , \10412 );
or \U$36338 ( \36681 , \36679 , \36680 );
nand \U$36339 ( \36682 , \18794 , RI98730a8_180);
nand \U$36340 ( \36683 , \36681 , \36682 );
not \U$36341 ( \36684 , \36683 );
or \U$36342 ( \36685 , \36678 , \36684 );
nand \U$36343 ( \36686 , \35338 , \13020 );
nand \U$36344 ( \36687 , \36685 , \36686 );
xor \U$36345 ( \36688 , \36677 , \36687 );
not \U$36346 ( \36689 , \36688 );
and \U$36347 ( \36690 , \36658 , \36689 );
not \U$36348 ( \36691 , \36658 );
and \U$36349 ( \36692 , \36691 , \36688 );
nor \U$36350 ( \36693 , \36690 , \36692 );
not \U$36351 ( \36694 , \36693 );
xor \U$36352 ( \36695 , \35555 , \35566 );
and \U$36353 ( \36696 , \36695 , \35576 );
and \U$36354 ( \36697 , \35555 , \35566 );
nor \U$36355 ( \36698 , \36696 , \36697 );
and \U$36356 ( \36699 , \17783 , \5648 );
not \U$36357 ( \36700 , \17783 );
and \U$36358 ( \36701 , \36700 , RI9872568_156);
nor \U$36359 ( \36702 , \36699 , \36701 );
and \U$36360 ( \36703 , \5653 , \36702 );
and \U$36361 ( \36704 , \35646 , \5641 );
nor \U$36362 ( \36705 , \36703 , \36704 );
not \U$36363 ( \36706 , \36705 );
not \U$36364 ( \36707 , \7338 );
not \U$36365 ( \36708 , RI98729a0_165);
not \U$36366 ( \36709 , \27588 );
or \U$36367 ( \36710 , \36708 , \36709 );
or \U$36368 ( \36711 , \17767 , RI98729a0_165);
nand \U$36369 ( \36712 , \36710 , \36711 );
not \U$36370 ( \36713 , \36712 );
or \U$36371 ( \36714 , \36707 , \36713 );
nand \U$36372 ( \36715 , \35310 , \7325 );
nand \U$36373 ( \36716 , \36714 , \36715 );
not \U$36374 ( \36717 , \36716 );
or \U$36375 ( \36718 , \36706 , \36717 );
or \U$36376 ( \36719 , \36716 , \36705 );
nand \U$36377 ( \36720 , \36718 , \36719 );
not \U$36378 ( \36721 , \36720 );
not \U$36379 ( \36722 , \6285 );
and \U$36380 ( \36723 , RI98728b0_163, \13268 );
not \U$36381 ( \36724 , RI98728b0_163);
and \U$36382 ( \36725 , \36724 , \32173 );
or \U$36383 ( \36726 , \36723 , \36725 );
not \U$36384 ( \36727 , \36726 );
or \U$36385 ( \36728 , \36722 , \36727 );
nand \U$36386 ( \36729 , \35288 , \6282 );
nand \U$36387 ( \36730 , \36728 , \36729 );
not \U$36388 ( \36731 , \36730 );
not \U$36389 ( \36732 , \36731 );
and \U$36390 ( \36733 , \36721 , \36732 );
and \U$36391 ( \36734 , \36720 , \36731 );
nor \U$36392 ( \36735 , \36733 , \36734 );
and \U$36393 ( \36736 , \36698 , \36735 );
not \U$36394 ( \36737 , \36698 );
not \U$36395 ( \36738 , \36735 );
and \U$36396 ( \36739 , \36737 , \36738 );
nor \U$36397 ( \36740 , \36736 , \36739 );
xor \U$36398 ( \36741 , \35297 , \35312 );
and \U$36399 ( \36742 , \36741 , \35328 );
and \U$36400 ( \36743 , \35297 , \35312 );
or \U$36401 ( \36744 , \36742 , \36743 );
xnor \U$36402 ( \36745 , \36740 , \36744 );
not \U$36403 ( \36746 , \36745 );
nand \U$36404 ( \36747 , \36694 , \36746 );
nand \U$36405 ( \36748 , \36693 , \36745 );
nand \U$36406 ( \36749 , \36747 , \36748 );
xor \U$36407 ( \36750 , \35649 , \35658 );
and \U$36408 ( \36751 , \36750 , \35673 );
and \U$36409 ( \36752 , \35649 , \35658 );
or \U$36410 ( \36753 , \36751 , \36752 );
not \U$36411 ( \36754 , \36753 );
not \U$36412 ( \36755 , \36754 );
xor \U$36413 ( \36756 , \34223 , \34226 );
not \U$36414 ( \36757 , \36756 );
not \U$36415 ( \36758 , \36757 );
not \U$36416 ( \36759 , \4084 );
not \U$36417 ( \36760 , \34507 );
or \U$36418 ( \36761 , \36759 , \36760 );
nand \U$36419 ( \36762 , \35534 , \4101 );
nand \U$36420 ( \36763 , \36761 , \36762 );
not \U$36421 ( \36764 , \36763 );
not \U$36422 ( \36765 , \36764 );
or \U$36423 ( \36766 , \36758 , \36765 );
nand \U$36424 ( \36767 , \36756 , \36763 );
nand \U$36425 ( \36768 , \36766 , \36767 );
not \U$36426 ( \36769 , \36768 );
not \U$36427 ( \36770 , \4922 );
not \U$36428 ( \36771 , \34233 );
or \U$36429 ( \36772 , \36770 , \36771 );
nand \U$36430 ( \36773 , \35549 , \4918 );
nand \U$36431 ( \36774 , \36772 , \36773 );
not \U$36432 ( \36775 , \36774 );
not \U$36433 ( \36776 , \36775 );
and \U$36434 ( \36777 , \36769 , \36776 );
and \U$36435 ( \36778 , \36768 , \36775 );
nor \U$36436 ( \36779 , \36777 , \36778 );
not \U$36437 ( \36780 , \36779 );
not \U$36438 ( \36781 , \9272 );
not \U$36439 ( \36782 , RI9872e50_175);
not \U$36440 ( \36783 , \22524 );
or \U$36441 ( \36784 , \36782 , \36783 );
or \U$36442 ( \36785 , \18111 , RI9872e50_175);
nand \U$36443 ( \36786 , \36784 , \36785 );
not \U$36444 ( \36787 , \36786 );
or \U$36445 ( \36788 , \36781 , \36787 );
nand \U$36446 ( \36789 , \35280 , \18562 );
nand \U$36447 ( \36790 , \36788 , \36789 );
not \U$36448 ( \36791 , \36790 );
or \U$36449 ( \36792 , \36780 , \36791 );
or \U$36450 ( \36793 , \36790 , \36779 );
nand \U$36451 ( \36794 , \36792 , \36793 );
not \U$36452 ( \36795 , \8751 );
not \U$36453 ( \36796 , RI9872f40_177);
not \U$36454 ( \36797 , \10392 );
or \U$36455 ( \36798 , \36796 , \36797 );
or \U$36456 ( \36799 , \8074 , RI9872f40_177);
nand \U$36457 ( \36800 , \36798 , \36799 );
not \U$36458 ( \36801 , \36800 );
or \U$36459 ( \36802 , \36795 , \36801 );
nand \U$36460 ( \36803 , \35264 , \9526 );
nand \U$36461 ( \36804 , \36802 , \36803 );
xnor \U$36462 ( \36805 , \36794 , \36804 );
not \U$36463 ( \36806 , \36805 );
not \U$36464 ( \36807 , \36806 );
not \U$36465 ( \36808 , \35378 );
not \U$36466 ( \36809 , \35364 );
or \U$36467 ( \36810 , \36808 , \36809 );
nand \U$36468 ( \36811 , \35359 , \35346 );
nand \U$36469 ( \36812 , \36810 , \36811 );
not \U$36470 ( \36813 , \36812 );
not \U$36471 ( \36814 , \36813 );
or \U$36472 ( \36815 , \36807 , \36814 );
nand \U$36473 ( \36816 , \36812 , \36805 );
nand \U$36474 ( \36817 , \36815 , \36816 );
not \U$36475 ( \36818 , \36817 );
or \U$36476 ( \36819 , \36755 , \36818 );
or \U$36477 ( \36820 , \36817 , \36754 );
nand \U$36478 ( \36821 , \36819 , \36820 );
xor \U$36479 ( \36822 , \36749 , \36821 );
not \U$36480 ( \36823 , \36822 );
not \U$36481 ( \36824 , \35388 );
not \U$36482 ( \36825 , \36824 );
not \U$36483 ( \36826 , \35625 );
or \U$36484 ( \36827 , \36825 , \36826 );
nand \U$36485 ( \36828 , \35484 , \35621 );
nand \U$36486 ( \36829 , \36827 , \36828 );
not \U$36487 ( \36830 , \35578 );
nand \U$36488 ( \36831 , \35582 , \35615 );
nand \U$36489 ( \36832 , \36830 , \36831 );
or \U$36490 ( \36833 , \35283 , \35329 );
nand \U$36491 ( \36834 , \36833 , \35383 );
nand \U$36492 ( \36835 , \36834 , \35331 );
xor \U$36493 ( \36836 , \36832 , \36835 );
not \U$36494 ( \36837 , \35697 );
not \U$36495 ( \36838 , \35684 );
or \U$36496 ( \36839 , \36837 , \36838 );
nand \U$36497 ( \36840 , \35689 , \35696 );
nand \U$36498 ( \36841 , \36839 , \36840 );
xor \U$36499 ( \36842 , \36836 , \36841 );
nor \U$36500 ( \36843 , \36829 , \36842 );
not \U$36501 ( \36844 , \36843 );
nand \U$36502 ( \36845 , \36829 , \36842 );
nand \U$36503 ( \36846 , \36844 , \36845 );
not \U$36504 ( \36847 , \36846 );
or \U$36505 ( \36848 , \36823 , \36847 );
or \U$36506 ( \36849 , \36846 , \36822 );
nand \U$36507 ( \36850 , \36848 , \36849 );
not \U$36508 ( \36851 , \36850 );
and \U$36509 ( \36852 , \36645 , \36851 );
and \U$36510 ( \36853 , \36644 , \36850 );
nor \U$36511 ( \36854 , \36852 , \36853 );
not \U$36512 ( \36855 , \36854 );
or \U$36513 ( \36856 , \36187 , \36855 );
or \U$36514 ( \36857 , \36854 , \36186 );
nand \U$36515 ( \36858 , \36856 , \36857 );
not \U$36516 ( \36859 , \35700 );
not \U$36517 ( \36860 , \35238 );
not \U$36518 ( \36861 , \36860 );
or \U$36519 ( \36862 , \36859 , \36861 );
nand \U$36520 ( \36863 , \35238 , \35699 );
nand \U$36521 ( \36864 , \36862 , \36863 );
buf \U$36522 ( \36865 , \35629 );
and \U$36523 ( \36866 , \36864 , \36865 );
not \U$36524 ( \36867 , \36864 );
not \U$36525 ( \36868 , \36865 );
and \U$36526 ( \36869 , \36867 , \36868 );
nor \U$36527 ( \36870 , \36866 , \36869 );
not \U$36528 ( \36871 , \36870 );
not \U$36529 ( \36872 , \35031 );
and \U$36530 ( \36873 , \35233 , \36872 );
not \U$36531 ( \36874 , \35233 );
and \U$36532 ( \36875 , \36874 , \35031 );
nor \U$36533 ( \36876 , \36873 , \36875 );
not \U$36534 ( \36877 , \36876 );
xor \U$36535 ( \36878 , \36307 , \36315 );
xor \U$36536 ( \36879 , \36878 , \36305 );
not \U$36537 ( \36880 , \36879 );
or \U$36538 ( \36881 , \36877 , \36880 );
not \U$36539 ( \36882 , RI9873648_192);
not \U$36540 ( \36883 , \36485 );
or \U$36541 ( \36884 , \36882 , \36883 );
not \U$36542 ( \36885 , RI9873558_190);
not \U$36543 ( \36886 , \5761 );
or \U$36544 ( \36887 , \36885 , \36886 );
or \U$36545 ( \36888 , \5761 , RI9873558_190);
nand \U$36546 ( \36889 , \36887 , \36888 );
nand \U$36547 ( \36890 , \36889 , \18545 );
nand \U$36548 ( \36891 , \36884 , \36890 );
not \U$36549 ( \36892 , \9937 );
not \U$36550 ( \36893 , \36500 );
or \U$36551 ( \36894 , \36892 , \36893 );
and \U$36552 ( \36895 , RI9873030_179, \19701 );
not \U$36553 ( \36896 , RI9873030_179);
and \U$36554 ( \36897 , \36896 , \8580 );
or \U$36555 ( \36898 , \36895 , \36897 );
nand \U$36556 ( \36899 , \36898 , \18672 );
nand \U$36557 ( \36900 , \36894 , \36899 );
xor \U$36558 ( \36901 , \36891 , \36900 );
not \U$36559 ( \36902 , \32292 );
not \U$36560 ( \36903 , RI9872bf8_170);
not \U$36561 ( \36904 , \13268 );
or \U$36562 ( \36905 , \36903 , \36904 );
or \U$36563 ( \36906 , \12773 , RI9872bf8_170);
nand \U$36564 ( \36907 , \36905 , \36906 );
not \U$36565 ( \36908 , \36907 );
or \U$36566 ( \36909 , \36902 , \36908 );
nand \U$36567 ( \36910 , \36562 , \22167 );
nand \U$36568 ( \36911 , \36909 , \36910 );
not \U$36569 ( \36912 , \36911 );
xor \U$36570 ( \36913 , \36539 , \36526 );
not \U$36571 ( \36914 , \8818 );
not \U$36572 ( \36915 , \8811 );
not \U$36573 ( \36916 , \33307 );
or \U$36574 ( \36917 , \36915 , \36916 );
or \U$36575 ( \36918 , \20292 , \8807 );
nand \U$36576 ( \36919 , \36917 , \36918 );
not \U$36577 ( \36920 , \36919 );
or \U$36578 ( \36921 , \36914 , \36920 );
nand \U$36579 ( \36922 , \36589 , \8801 );
nand \U$36580 ( \36923 , \36921 , \36922 );
xor \U$36581 ( \36924 , \36913 , \36923 );
not \U$36582 ( \36925 , \36924 );
or \U$36583 ( \36926 , \36912 , \36925 );
nand \U$36584 ( \36927 , \36923 , \36913 );
nand \U$36585 ( \36928 , \36926 , \36927 );
and \U$36586 ( \36929 , \36901 , \36928 );
and \U$36587 ( \36930 , \36891 , \36900 );
or \U$36588 ( \36931 , \36929 , \36930 );
xor \U$36589 ( \36932 , \36244 , \36292 );
xor \U$36590 ( \36933 , \36931 , \36932 );
xor \U$36591 ( \36934 , \36487 , \36504 );
xor \U$36592 ( \36935 , \36934 , \36494 );
and \U$36593 ( \36936 , \36933 , \36935 );
and \U$36594 ( \36937 , \36931 , \36932 );
or \U$36595 ( \36938 , \36936 , \36937 );
not \U$36596 ( \36939 , \36938 );
not \U$36597 ( \36940 , \36448 );
not \U$36598 ( \36941 , \36940 );
not \U$36599 ( \36942 , \36427 );
not \U$36600 ( \36943 , \36439 );
or \U$36601 ( \36944 , \36942 , \36943 );
or \U$36602 ( \36945 , \36427 , \36439 );
nand \U$36603 ( \36946 , \36944 , \36945 );
not \U$36604 ( \36947 , \36946 );
or \U$36605 ( \36948 , \36941 , \36947 );
or \U$36606 ( \36949 , \36946 , \36940 );
nand \U$36607 ( \36950 , \36948 , \36949 );
not \U$36608 ( \36951 , \36950 );
xor \U$36609 ( \36952 , \36216 , \36228 );
not \U$36610 ( \36953 , \12867 );
not \U$36611 ( \36954 , \36240 );
or \U$36612 ( \36955 , \36953 , \36954 );
not \U$36613 ( \36956 , RI98730a8_180);
not \U$36614 ( \36957 , \8857 );
or \U$36615 ( \36958 , \36956 , \36957 );
or \U$36616 ( \36959 , \8857 , RI98730a8_180);
nand \U$36617 ( \36960 , \36958 , \36959 );
nand \U$36618 ( \36961 , \36960 , \24209 );
nand \U$36619 ( \36962 , \36955 , \36961 );
not \U$36620 ( \36963 , \36962 );
not \U$36621 ( \36964 , \36963 );
not \U$36622 ( \36965 , \17528 );
not \U$36623 ( \36966 , \36284 );
or \U$36624 ( \36967 , \36965 , \36966 );
not \U$36625 ( \36968 , \22727 );
not \U$36626 ( \36969 , \9898 );
or \U$36627 ( \36970 , \36968 , \36969 );
or \U$36628 ( \36971 , \12727 , \24305 );
nand \U$36629 ( \36972 , \36970 , \36971 );
nand \U$36630 ( \36973 , \36972 , \18508 );
nand \U$36631 ( \36974 , \36967 , \36973 );
not \U$36632 ( \36975 , \36974 );
not \U$36633 ( \36976 , \36975 );
or \U$36634 ( \36977 , \36964 , \36976 );
not \U$36635 ( \36978 , \17263 );
not \U$36636 ( \36979 , \36490 );
or \U$36637 ( \36980 , \36978 , \36979 );
not \U$36638 ( \36981 , \17539 );
not \U$36639 ( \36982 , \8942 );
or \U$36640 ( \36983 , \36981 , \36982 );
nand \U$36641 ( \36984 , \8081 , RI98733f0_187);
nand \U$36642 ( \36985 , \36983 , \36984 );
nand \U$36643 ( \36986 , \36985 , \17251 );
nand \U$36644 ( \36987 , \36980 , \36986 );
nand \U$36645 ( \36988 , \36977 , \36987 );
nand \U$36646 ( \36989 , \36974 , \36962 );
nand \U$36647 ( \36990 , \36988 , \36989 );
xor \U$36648 ( \36991 , \36952 , \36990 );
xor \U$36649 ( \36992 , \36389 , \36398 );
xor \U$36650 ( \36993 , \36992 , \36410 );
and \U$36651 ( \36994 , \36991 , \36993 );
and \U$36652 ( \36995 , \36952 , \36990 );
nor \U$36653 ( \36996 , \36994 , \36995 );
not \U$36654 ( \36997 , \36996 );
or \U$36655 ( \36998 , \36951 , \36997 );
or \U$36656 ( \36999 , \36996 , \36950 );
nand \U$36657 ( \37000 , \36998 , \36999 );
not \U$36658 ( \37001 , \37000 );
or \U$36659 ( \37002 , \36939 , \37001 );
not \U$36660 ( \37003 , \36996 );
nand \U$36661 ( \37004 , \37003 , \36950 );
nand \U$36662 ( \37005 , \37002 , \37004 );
not \U$36663 ( \37006 , \37005 );
and \U$36664 ( \37007 , \36413 , \36377 );
not \U$36665 ( \37008 , \36413 );
and \U$36666 ( \37009 , \37008 , \36378 );
or \U$36667 ( \37010 , \37007 , \37009 );
nand \U$36668 ( \37011 , \36300 , \36234 );
xnor \U$36669 ( \37012 , \36297 , \37011 );
xor \U$36670 ( \37013 , \37010 , \37012 );
xor \U$36671 ( \37014 , \36368 , \36347 );
not \U$36672 ( \37015 , \11198 );
not \U$36673 ( \37016 , \36343 );
or \U$36674 ( \37017 , \37015 , \37016 );
not \U$36675 ( \37018 , RI9872f40_177);
not \U$36676 ( \37019 , \20385 );
or \U$36677 ( \37020 , \37018 , \37019 );
or \U$36678 ( \37021 , \13454 , RI9872f40_177);
nand \U$36679 ( \37022 , \37020 , \37021 );
nand \U$36680 ( \37023 , \37022 , \24627 );
nand \U$36681 ( \37024 , \37017 , \37023 );
not \U$36682 ( \37025 , \37024 );
xnor \U$36683 ( \37026 , \36272 , \36261 );
not \U$36684 ( \37027 , \37026 );
not \U$36685 ( \37028 , \9272 );
not \U$36686 ( \37029 , \36385 );
or \U$36687 ( \37030 , \37028 , \37029 );
not \U$36688 ( \37031 , RI9872e50_175);
not \U$36689 ( \37032 , \9849 );
or \U$36690 ( \37033 , \37031 , \37032 );
or \U$36691 ( \37034 , \12460 , RI9872e50_175);
nand \U$36692 ( \37035 , \37033 , \37034 );
nand \U$36693 ( \37036 , \37035 , \9294 );
nand \U$36694 ( \37037 , \37030 , \37036 );
not \U$36695 ( \37038 , \37037 );
or \U$36696 ( \37039 , \37027 , \37038 );
or \U$36697 ( \37040 , \37037 , \37026 );
nand \U$36698 ( \37041 , \37039 , \37040 );
not \U$36699 ( \37042 , \37041 );
or \U$36700 ( \37043 , \37025 , \37042 );
not \U$36701 ( \37044 , \37026 );
nand \U$36702 ( \37045 , \37044 , \37037 );
nand \U$36703 ( \37046 , \37043 , \37045 );
xor \U$36704 ( \37047 , \37014 , \37046 );
not \U$36705 ( \37048 , \17234 );
not \U$36706 ( \37049 , \36394 );
or \U$36707 ( \37050 , \37048 , \37049 );
and \U$36708 ( \37051 , \9869 , RI9873210_183);
not \U$36709 ( \37052 , \9869 );
and \U$36710 ( \37053 , \37052 , \28789 );
nor \U$36711 ( \37054 , \37051 , \37053 );
nand \U$36712 ( \37055 , \37054 , \13476 );
nand \U$36713 ( \37056 , \37050 , \37055 );
not \U$36714 ( \37057 , \37056 );
not \U$36715 ( \37058 , \8027 );
not \U$36716 ( \37059 , RI9872a18_166);
not \U$36717 ( \37060 , \25380 );
or \U$36718 ( \37061 , \37059 , \37060 );
or \U$36719 ( \37062 , \18710 , RI9872a18_166);
nand \U$36720 ( \37063 , \37061 , \37062 );
not \U$36721 ( \37064 , \37063 );
or \U$36722 ( \37065 , \37058 , \37064 );
nand \U$36723 ( \37066 , \36580 , \8039 );
nand \U$36724 ( \37067 , \37065 , \37066 );
not \U$36725 ( \37068 , \37067 );
not \U$36726 ( \37069 , \7325 );
not \U$36727 ( \37070 , \7333 );
not \U$36728 ( \37071 , \22285 );
or \U$36729 ( \37072 , \37070 , \37071 );
nand \U$36730 ( \37073 , \24470 , RI98729a0_165);
nand \U$36731 ( \37074 , \37072 , \37073 );
not \U$36732 ( \37075 , \37074 );
or \U$36733 ( \37076 , \37069 , \37075 );
nand \U$36734 ( \37077 , \36270 , \7338 );
nand \U$36735 ( \37078 , \37076 , \37077 );
not \U$36736 ( \37079 , \5653 );
not \U$36737 ( \37080 , \36533 );
or \U$36738 ( \37081 , \37079 , \37080 );
and \U$36739 ( \37082 , RI9872568_156, \18704 );
not \U$36740 ( \37083 , RI9872568_156);
and \U$36741 ( \37084 , \37083 , \22278 );
nor \U$36742 ( \37085 , \37082 , \37084 );
nand \U$36743 ( \37086 , \37085 , \5641 );
nand \U$36744 ( \37087 , \37081 , \37086 );
nand \U$36745 ( \37088 , \25394 , \5633 );
nand \U$36746 ( \37089 , \37088 , \5634 , RI9872568_156);
not \U$36747 ( \37090 , \37089 );
and \U$36748 ( \37091 , \37087 , \37090 );
xnor \U$36749 ( \37092 , \37078 , \37091 );
not \U$36750 ( \37093 , \37092 );
not \U$36751 ( \37094 , \37093 );
or \U$36752 ( \37095 , \37068 , \37094 );
nand \U$36753 ( \37096 , \37078 , \37091 );
nand \U$36754 ( \37097 , \37095 , \37096 );
not \U$36755 ( \37098 , \36405 );
not \U$36756 ( \37099 , \19046 );
or \U$36757 ( \37100 , \37098 , \37099 );
not \U$36758 ( \37101 , \35146 );
not \U$36759 ( \37102 , \22516 );
or \U$36760 ( \37103 , \37101 , \37102 );
nand \U$36761 ( \37104 , \12805 , RI98734e0_189);
nand \U$36762 ( \37105 , \37103 , \37104 );
nand \U$36763 ( \37106 , \37105 , \19035 );
nand \U$36764 ( \37107 , \37100 , \37106 );
xor \U$36765 ( \37108 , \37097 , \37107 );
not \U$36766 ( \37109 , \37108 );
or \U$36767 ( \37110 , \37057 , \37109 );
nand \U$36768 ( \37111 , \37107 , \37097 );
nand \U$36769 ( \37112 , \37110 , \37111 );
and \U$36770 ( \37113 , \37047 , \37112 );
and \U$36771 ( \37114 , \37014 , \37046 );
or \U$36772 ( \37115 , \37113 , \37114 );
and \U$36773 ( \37116 , \37013 , \37115 );
and \U$36774 ( \37117 , \37010 , \37012 );
or \U$36775 ( \37118 , \37116 , \37117 );
not \U$36776 ( \37119 , \37118 );
not \U$36777 ( \37120 , \36301 );
not \U$36778 ( \37121 , \36192 );
not \U$36779 ( \37122 , \36303 );
or \U$36780 ( \37123 , \37121 , \37122 );
nand \U$36781 ( \37124 , \36188 , \36191 );
nand \U$36782 ( \37125 , \37123 , \37124 );
not \U$36783 ( \37126 , \37125 );
or \U$36784 ( \37127 , \37120 , \37126 );
or \U$36785 ( \37128 , \36301 , \37125 );
nand \U$36786 ( \37129 , \37127 , \37128 );
nand \U$36787 ( \37130 , \37119 , \37129 );
not \U$36788 ( \37131 , \37130 );
or \U$36789 ( \37132 , \37006 , \37131 );
not \U$36790 ( \37133 , \37129 );
nand \U$36791 ( \37134 , \37133 , \37118 );
nand \U$36792 ( \37135 , \37132 , \37134 );
nand \U$36793 ( \37136 , \36881 , \37135 );
not \U$36794 ( \37137 , \36879 );
not \U$36795 ( \37138 , \36876 );
nand \U$36796 ( \37139 , \37137 , \37138 );
and \U$36797 ( \37140 , \37136 , \37139 );
not \U$36798 ( \37141 , \37140 );
and \U$36799 ( \37142 , \36871 , \37141 );
and \U$36800 ( \37143 , \36870 , \37140 );
nor \U$36801 ( \37144 , \37142 , \37143 );
not \U$36802 ( \37145 , \37144 );
not \U$36803 ( \37146 , \37145 );
not \U$36804 ( \37147 , \36640 );
not \U$36805 ( \37148 , \37147 );
nand \U$36806 ( \37149 , \36643 , \36333 );
not \U$36807 ( \37150 , \37149 );
or \U$36808 ( \37151 , \37148 , \37150 );
or \U$36809 ( \37152 , \37149 , \37147 );
nand \U$36810 ( \37153 , \37151 , \37152 );
not \U$36811 ( \37154 , \37153 );
or \U$36812 ( \37155 , \37146 , \37154 );
not \U$36813 ( \37156 , \36870 );
nand \U$36814 ( \37157 , \37156 , \37140 );
nand \U$36815 ( \37158 , \37155 , \37157 );
nand \U$36816 ( \37159 , \36858 , \37158 );
not \U$36817 ( \37160 , \37153 );
not \U$36818 ( \37161 , \37144 );
or \U$36819 ( \37162 , \37160 , \37161 );
or \U$36820 ( \37163 , \37144 , \37153 );
nand \U$36821 ( \37164 , \37162 , \37163 );
and \U$36822 ( \37165 , \36879 , \36876 );
not \U$36823 ( \37166 , \36879 );
and \U$36824 ( \37167 , \37166 , \37138 );
nor \U$36825 ( \37168 , \37165 , \37167 );
not \U$36826 ( \37169 , \37168 );
not \U$36827 ( \37170 , \37135 );
or \U$36828 ( \37171 , \37169 , \37170 );
or \U$36829 ( \37172 , \37168 , \37135 );
nand \U$36830 ( \37173 , \37171 , \37172 );
not \U$36831 ( \37174 , \37173 );
nand \U$36832 ( \37175 , \36635 , \36476 );
and \U$36833 ( \37176 , \37175 , \36630 );
not \U$36834 ( \37177 , \37175 );
not \U$36835 ( \37178 , \36630 );
and \U$36836 ( \37179 , \37177 , \37178 );
nor \U$36837 ( \37180 , \37176 , \37179 );
buf \U$36838 ( \37181 , \36454 );
not \U$36839 ( \37182 , \36334 );
and \U$36840 ( \37183 , \37181 , \37182 );
not \U$36841 ( \37184 , \37181 );
and \U$36842 ( \37185 , \37184 , \36334 );
nor \U$36843 ( \37186 , \37183 , \37185 );
nand \U$36844 ( \37187 , \37180 , \37186 );
not \U$36845 ( \37188 , \37187 );
xor \U$36846 ( \37189 , \37010 , \37012 );
xor \U$36847 ( \37190 , \37189 , \37115 );
xor \U$36848 ( \37191 , \36626 , \36614 );
xnor \U$36849 ( \37192 , \37191 , \36509 );
or \U$36850 ( \37193 , \37190 , \37192 );
xor \U$36851 ( \37194 , \36991 , \36993 );
not \U$36852 ( \37195 , \37194 );
not \U$36853 ( \37196 , \37067 );
not \U$36854 ( \37197 , \37092 );
or \U$36855 ( \37198 , \37196 , \37197 );
or \U$36856 ( \37199 , \37092 , \37067 );
nand \U$36857 ( \37200 , \37198 , \37199 );
not \U$36858 ( \37201 , \12507 );
not \U$36859 ( \37202 , RI9873030_179);
not \U$36860 ( \37203 , \13298 );
or \U$36861 ( \37204 , \37202 , \37203 );
or \U$36862 ( \37205 , \8554 , RI9873030_179);
nand \U$36863 ( \37206 , \37204 , \37205 );
not \U$36864 ( \37207 , \37206 );
or \U$36865 ( \37208 , \37201 , \37207 );
nand \U$36866 ( \37209 , \36898 , \9937 );
nand \U$36867 ( \37210 , \37208 , \37209 );
xor \U$36868 ( \37211 , \37200 , \37210 );
not \U$36869 ( \37212 , \17263 );
not \U$36870 ( \37213 , \36985 );
or \U$36871 ( \37214 , \37212 , \37213 );
and \U$36872 ( \37215 , RI98733f0_187, \7466 );
not \U$36873 ( \37216 , RI98733f0_187);
and \U$36874 ( \37217 , \37216 , \19752 );
or \U$36875 ( \37218 , \37215 , \37217 );
nand \U$36876 ( \37219 , \37218 , \17251 );
nand \U$36877 ( \37220 , \37214 , \37219 );
and \U$36878 ( \37221 , \37211 , \37220 );
and \U$36879 ( \37222 , \37200 , \37210 );
or \U$36880 ( \37223 , \37221 , \37222 );
not \U$36881 ( \37224 , \36962 );
not \U$36882 ( \37225 , \36975 );
or \U$36883 ( \37226 , \37224 , \37225 );
or \U$36884 ( \37227 , \36962 , \36975 );
nand \U$36885 ( \37228 , \37226 , \37227 );
xor \U$36886 ( \37229 , \36987 , \37228 );
xor \U$36887 ( \37230 , \37223 , \37229 );
xor \U$36888 ( \37231 , \37056 , \37108 );
and \U$36889 ( \37232 , \37230 , \37231 );
and \U$36890 ( \37233 , \37223 , \37229 );
or \U$36891 ( \37234 , \37232 , \37233 );
not \U$36892 ( \37235 , \37234 );
or \U$36893 ( \37236 , \37195 , \37235 );
or \U$36894 ( \37237 , \37234 , \37194 );
not \U$36895 ( \37238 , \37041 );
not \U$36896 ( \37239 , \37024 );
not \U$36897 ( \37240 , \37239 );
and \U$36898 ( \37241 , \37238 , \37240 );
and \U$36899 ( \37242 , \37041 , \37239 );
nor \U$36900 ( \37243 , \37241 , \37242 );
not \U$36901 ( \37244 , \37243 );
not \U$36902 ( \37245 , \37244 );
not \U$36903 ( \37246 , \29633 );
not \U$36904 ( \37247 , \13022 );
not \U$36905 ( \37248 , \8642 );
or \U$36906 ( \37249 , \37247 , \37248 );
or \U$36907 ( \37250 , \8642 , \13022 );
nand \U$36908 ( \37251 , \37249 , \37250 );
not \U$36909 ( \37252 , \37251 );
or \U$36910 ( \37253 , \37246 , \37252 );
nand \U$36911 ( \37254 , \36960 , \12867 );
nand \U$36912 ( \37255 , \37253 , \37254 );
not \U$36913 ( \37256 , \37255 );
not \U$36914 ( \37257 , \18544 );
not \U$36915 ( \37258 , \18239 );
not \U$36916 ( \37259 , \36403 );
or \U$36917 ( \37260 , \37258 , \37259 );
or \U$36918 ( \37261 , \6303 , \18239 );
nand \U$36919 ( \37262 , \37260 , \37261 );
not \U$36920 ( \37263 , \37262 );
or \U$36921 ( \37264 , \37257 , \37263 );
nand \U$36922 ( \37265 , \36889 , RI9873648_192);
nand \U$36923 ( \37266 , \37264 , \37265 );
not \U$36924 ( \37267 , \37266 );
or \U$36925 ( \37268 , \37256 , \37267 );
or \U$36926 ( \37269 , \37266 , \37255 );
not \U$36927 ( \37270 , \17243 );
and \U$36928 ( \37271 , \22524 , \22675 );
not \U$36929 ( \37272 , \22524 );
and \U$36930 ( \37273 , \37272 , RI9873210_183);
nor \U$36931 ( \37274 , \37271 , \37273 );
not \U$36932 ( \37275 , \37274 );
or \U$36933 ( \37276 , \37270 , \37275 );
nand \U$36934 ( \37277 , \37054 , \30963 );
nand \U$36935 ( \37278 , \37276 , \37277 );
nand \U$36936 ( \37279 , \37269 , \37278 );
nand \U$36937 ( \37280 , \37268 , \37279 );
xnor \U$36938 ( \37281 , \36608 , \36599 );
xor \U$36939 ( \37282 , \37280 , \37281 );
not \U$36940 ( \37283 , \37282 );
or \U$36941 ( \37284 , \37245 , \37283 );
nand \U$36942 ( \37285 , \37280 , \37281 );
nand \U$36943 ( \37286 , \37284 , \37285 );
nand \U$36944 ( \37287 , \37237 , \37286 );
nand \U$36945 ( \37288 , \37236 , \37287 );
nand \U$36946 ( \37289 , \37193 , \37288 );
nand \U$36947 ( \37290 , \37190 , \37192 );
nand \U$36948 ( \37291 , \37289 , \37290 );
not \U$36949 ( \37292 , \37291 );
or \U$36950 ( \37293 , \37188 , \37292 );
not \U$36951 ( \37294 , \37180 );
not \U$36952 ( \37295 , \37186 );
nand \U$36953 ( \37296 , \37294 , \37295 );
nand \U$36954 ( \37297 , \37293 , \37296 );
not \U$36955 ( \37298 , \37297 );
xor \U$36956 ( \37299 , \36458 , \36636 );
xor \U$36957 ( \37300 , \37299 , \36462 );
not \U$36958 ( \37301 , \37300 );
or \U$36959 ( \37302 , \37298 , \37301 );
or \U$36960 ( \37303 , \37300 , \37297 );
nand \U$36961 ( \37304 , \37302 , \37303 );
not \U$36962 ( \37305 , \37304 );
or \U$36963 ( \37306 , \37174 , \37305 );
not \U$36964 ( \37307 , \37297 );
nand \U$36965 ( \37308 , \37307 , \37300 );
nand \U$36966 ( \37309 , \37306 , \37308 );
nand \U$36967 ( \37310 , \37164 , \37309 );
xor \U$36968 ( \37311 , \37173 , \37304 );
nand \U$36969 ( \37312 , \37296 , \37187 );
buf \U$36970 ( \37313 , \37291 );
not \U$36971 ( \37314 , \37313 );
and \U$36972 ( \37315 , \37312 , \37314 );
not \U$36973 ( \37316 , \37312 );
and \U$36974 ( \37317 , \37316 , \37313 );
nor \U$36975 ( \37318 , \37315 , \37317 );
not \U$36976 ( \37319 , \37318 );
not \U$36977 ( \37320 , \37319 );
not \U$36978 ( \37321 , \37129 );
not \U$36979 ( \37322 , \37119 );
or \U$36980 ( \37323 , \37321 , \37322 );
nand \U$36981 ( \37324 , \37323 , \37134 );
not \U$36982 ( \37325 , \37005 );
xor \U$36983 ( \37326 , \37324 , \37325 );
not \U$36984 ( \37327 , \37326 );
not \U$36985 ( \37328 , \37087 );
not \U$36986 ( \37329 , \37089 );
and \U$36987 ( \37330 , \37328 , \37329 );
and \U$36988 ( \37331 , \37087 , \37089 );
nor \U$36989 ( \37332 , \37330 , \37331 );
not \U$36990 ( \37333 , \6285 );
not \U$36991 ( \37334 , \36524 );
or \U$36992 ( \37335 , \37333 , \37334 );
not \U$36993 ( \37336 , \5632 );
not \U$36994 ( \37337 , \17862 );
or \U$36995 ( \37338 , \37336 , \37337 );
or \U$36996 ( \37339 , \34408 , \7049 );
nand \U$36997 ( \37340 , \37338 , \37339 );
nand \U$36998 ( \37341 , \37340 , \6282 );
nand \U$36999 ( \37342 , \37335 , \37341 );
xor \U$37000 ( \37343 , \37332 , \37342 );
not \U$37001 ( \37344 , \37343 );
not \U$37002 ( \37345 , \37344 );
not \U$37003 ( \37346 , \8039 );
not \U$37004 ( \37347 , \37063 );
or \U$37005 ( \37348 , \37346 , \37347 );
and \U$37006 ( \37349 , RI9872a18_166, \17911 );
not \U$37007 ( \37350 , RI9872a18_166);
and \U$37008 ( \37351 , \37350 , \17912 );
or \U$37009 ( \37352 , \37349 , \37351 );
nand \U$37010 ( \37353 , \37352 , \8027 );
nand \U$37011 ( \37354 , \37348 , \37353 );
not \U$37012 ( \37355 , \37354 );
or \U$37013 ( \37356 , \37345 , \37355 );
not \U$37014 ( \37357 , \37332 );
nand \U$37015 ( \37358 , \37357 , \37342 );
nand \U$37016 ( \37359 , \37356 , \37358 );
not \U$37017 ( \37360 , \17528 );
not \U$37018 ( \37361 , \36972 );
or \U$37019 ( \37362 , \37360 , \37361 );
not \U$37020 ( \37363 , \22715 );
not \U$37021 ( \37364 , \10391 );
or \U$37022 ( \37365 , \37363 , \37364 );
or \U$37023 ( \37366 , \8075 , \24305 );
nand \U$37024 ( \37367 , \37365 , \37366 );
nand \U$37025 ( \37368 , \37367 , \18508 );
nand \U$37026 ( \37369 , \37362 , \37368 );
xor \U$37027 ( \37370 , \37359 , \37369 );
not \U$37028 ( \37371 , \19036 );
not \U$37029 ( \37372 , \16999 );
not \U$37030 ( \37373 , \18793 );
or \U$37031 ( \37374 , \37372 , \37373 );
or \U$37032 ( \37375 , \7905 , \19361 );
nand \U$37033 ( \37376 , \37374 , \37375 );
not \U$37034 ( \37377 , \37376 );
or \U$37035 ( \37378 , \37371 , \37377 );
nand \U$37036 ( \37379 , \37105 , \28811 );
nand \U$37037 ( \37380 , \37378 , \37379 );
and \U$37038 ( \37381 , \37370 , \37380 );
and \U$37039 ( \37382 , \37359 , \37369 );
or \U$37040 ( \37383 , \37381 , \37382 );
not \U$37041 ( \37384 , \37383 );
not \U$37042 ( \37385 , \9294 );
not \U$37043 ( \37386 , RI9872e50_175);
not \U$37044 ( \37387 , \24729 );
or \U$37045 ( \37388 , \37386 , \37387 );
or \U$37046 ( \37389 , \9114 , RI9872e50_175);
nand \U$37047 ( \37390 , \37388 , \37389 );
not \U$37048 ( \37391 , \37390 );
or \U$37049 ( \37392 , \37385 , \37391 );
nand \U$37050 ( \37393 , \37035 , \9272 );
nand \U$37051 ( \37394 , \37392 , \37393 );
not \U$37052 ( \37395 , \9195 );
and \U$37053 ( \37396 , RI9872b80_169, \24754 );
not \U$37054 ( \37397 , RI9872b80_169);
and \U$37055 ( \37398 , \37397 , \22391 );
or \U$37056 ( \37399 , \37396 , \37398 );
not \U$37057 ( \37400 , \37399 );
or \U$37058 ( \37401 , \37395 , \37400 );
nand \U$37059 ( \37402 , \36606 , \9214 );
nand \U$37060 ( \37403 , \37401 , \37402 );
nor \U$37061 ( \37404 , \37394 , \37403 );
not \U$37062 ( \37405 , \24627 );
and \U$37063 ( \37406 , RI9872f40_177, \8695 );
not \U$37064 ( \37407 , RI9872f40_177);
and \U$37065 ( \37408 , \37407 , \24807 );
nor \U$37066 ( \37409 , \37406 , \37408 );
not \U$37067 ( \37410 , \37409 );
or \U$37068 ( \37411 , \37405 , \37410 );
nand \U$37069 ( \37412 , \37022 , \8751 );
nand \U$37070 ( \37413 , \37411 , \37412 );
not \U$37071 ( \37414 , \37413 );
or \U$37072 ( \37415 , \37404 , \37414 );
nand \U$37073 ( \37416 , \37394 , \37403 );
nand \U$37074 ( \37417 , \37415 , \37416 );
not \U$37075 ( \37418 , \36568 );
not \U$37076 ( \37419 , \36555 );
and \U$37077 ( \37420 , \37418 , \37419 );
and \U$37078 ( \37421 , \36568 , \36555 );
nor \U$37079 ( \37422 , \37420 , \37421 );
xor \U$37080 ( \37423 , \37417 , \37422 );
not \U$37081 ( \37424 , \37423 );
not \U$37082 ( \37425 , \37424 );
or \U$37083 ( \37426 , \37384 , \37425 );
not \U$37084 ( \37427 , \37422 );
nand \U$37085 ( \37428 , \37427 , \37417 );
nand \U$37086 ( \37429 , \37426 , \37428 );
xor \U$37087 ( \37430 , \36511 , \36572 );
xor \U$37088 ( \37431 , \37430 , \36610 );
nor \U$37089 ( \37432 , \37429 , \37431 );
not \U$37090 ( \37433 , \37432 );
not \U$37091 ( \37434 , \37433 );
xor \U$37092 ( \37435 , \37014 , \37046 );
xor \U$37093 ( \37436 , \37435 , \37112 );
not \U$37094 ( \37437 , \37436 );
or \U$37095 ( \37438 , \37434 , \37437 );
nand \U$37096 ( \37439 , \37429 , \37431 );
nand \U$37097 ( \37440 , \37438 , \37439 );
xor \U$37098 ( \37441 , \36891 , \36900 );
xor \U$37099 ( \37442 , \37441 , \36928 );
not \U$37100 ( \37443 , \37442 );
or \U$37101 ( \37444 , RI9872928_164, RI98729a0_165);
nand \U$37102 ( \37445 , \37444 , \18705 );
and \U$37103 ( \37446 , RI9872928_164, RI98729a0_165);
nor \U$37104 ( \37447 , \37446 , \5632 );
and \U$37105 ( \37448 , \37445 , \37447 );
not \U$37106 ( \37449 , \6285 );
and \U$37107 ( \37450 , RI98728b0_163, \23953 );
not \U$37108 ( \37451 , RI98728b0_163);
and \U$37109 ( \37452 , \37451 , \28671 );
or \U$37110 ( \37453 , \37450 , \37452 );
not \U$37111 ( \37454 , \37453 );
or \U$37112 ( \37455 , \37449 , \37454 );
xor \U$37113 ( \37456 , \18704 , RI98728b0_163);
nand \U$37114 ( \37457 , \37456 , \6282 );
nand \U$37115 ( \37458 , \37455 , \37457 );
and \U$37116 ( \37459 , \37448 , \37458 );
not \U$37117 ( \37460 , \8039 );
not \U$37118 ( \37461 , \37352 );
or \U$37119 ( \37462 , \37460 , \37461 );
not \U$37120 ( \37463 , RI9872a18_166);
not \U$37121 ( \37464 , \30350 );
or \U$37122 ( \37465 , \37463 , \37464 );
or \U$37123 ( \37466 , \25412 , RI9872a18_166);
nand \U$37124 ( \37467 , \37465 , \37466 );
nand \U$37125 ( \37468 , \37467 , \8027 );
nand \U$37126 ( \37469 , \37462 , \37468 );
xor \U$37127 ( \37470 , \37459 , \37469 );
not \U$37128 ( \37471 , \9195 );
and \U$37129 ( \37472 , RI9872b80_169, \34938 );
not \U$37130 ( \37473 , RI9872b80_169);
and \U$37131 ( \37474 , \37473 , \20765 );
nor \U$37132 ( \37475 , \37472 , \37474 );
not \U$37133 ( \37476 , \37475 );
or \U$37134 ( \37477 , \37471 , \37476 );
not \U$37135 ( \37478 , \9198 );
not \U$37136 ( \37479 , \17014 );
or \U$37137 ( \37480 , \37478 , \37479 );
or \U$37138 ( \37481 , \17014 , \11688 );
nand \U$37139 ( \37482 , \37480 , \37481 );
nand \U$37140 ( \37483 , \37482 , \9214 );
nand \U$37141 ( \37484 , \37477 , \37483 );
and \U$37142 ( \37485 , \37470 , \37484 );
and \U$37143 ( \37486 , \37459 , \37469 );
nor \U$37144 ( \37487 , \37485 , \37486 );
not \U$37145 ( \37488 , \37487 );
not \U$37146 ( \37489 , \37488 );
not \U$37147 ( \37490 , \17528 );
not \U$37148 ( \37491 , \37367 );
or \U$37149 ( \37492 , \37490 , \37491 );
and \U$37150 ( \37493 , \32967 , \8874 );
not \U$37151 ( \37494 , \32967 );
and \U$37152 ( \37495 , \37494 , \8877 );
nor \U$37153 ( \37496 , \37493 , \37495 );
nand \U$37154 ( \37497 , \37496 , \18508 );
nand \U$37155 ( \37498 , \37492 , \37497 );
buf \U$37156 ( \37499 , \37498 );
not \U$37157 ( \37500 , \37499 );
or \U$37158 ( \37501 , \37489 , \37500 );
not \U$37159 ( \37502 , \30963 );
not \U$37160 ( \37503 , \37274 );
or \U$37161 ( \37504 , \37502 , \37503 );
and \U$37162 ( \37505 , \8668 , \28789 );
not \U$37163 ( \37506 , \8668 );
and \U$37164 ( \37507 , \37506 , RI9873210_183);
nor \U$37165 ( \37508 , \37505 , \37507 );
nand \U$37166 ( \37509 , \37508 , \13477 );
nand \U$37167 ( \37510 , \37504 , \37509 );
not \U$37168 ( \37511 , \37498 );
nand \U$37169 ( \37512 , \37511 , \37487 );
nand \U$37170 ( \37513 , \37510 , \37512 );
nand \U$37171 ( \37514 , \37501 , \37513 );
not \U$37172 ( \37515 , \37514 );
xnor \U$37173 ( \37516 , \36924 , \36911 );
nand \U$37174 ( \37517 , \37515 , \37516 );
not \U$37175 ( \37518 , \37517 );
not \U$37176 ( \37519 , \12867 );
not \U$37177 ( \37520 , \37251 );
or \U$37178 ( \37521 , \37519 , \37520 );
and \U$37179 ( \37522 , \8845 , RI98730a8_180);
not \U$37180 ( \37523 , \8845 );
and \U$37181 ( \37524 , \37523 , \13022 );
nor \U$37182 ( \37525 , \37522 , \37524 );
nand \U$37183 ( \37526 , \37525 , \13020 );
nand \U$37184 ( \37527 , \37521 , \37526 );
not \U$37185 ( \37528 , \37527 );
not \U$37186 ( \37529 , \18615 );
not \U$37187 ( \37530 , RI9873558_190);
not \U$37188 ( \37531 , \8904 );
or \U$37189 ( \37532 , \37530 , \37531 );
or \U$37190 ( \37533 , \8904 , RI9873558_190);
nand \U$37191 ( \37534 , \37532 , \37533 );
not \U$37192 ( \37535 , \37534 );
or \U$37193 ( \37536 , \37529 , \37535 );
nand \U$37194 ( \37537 , \37262 , RI9873648_192);
nand \U$37195 ( \37538 , \37536 , \37537 );
not \U$37196 ( \37539 , \37538 );
or \U$37197 ( \37540 , \37528 , \37539 );
or \U$37198 ( \37541 , \37538 , \37527 );
not \U$37199 ( \37542 , \17252 );
and \U$37200 ( \37543 , RI98733f0_187, \8334 );
not \U$37201 ( \37544 , RI98733f0_187);
and \U$37202 ( \37545 , \37544 , \8916 );
or \U$37203 ( \37546 , \37543 , \37545 );
not \U$37204 ( \37547 , \37546 );
or \U$37205 ( \37548 , \37542 , \37547 );
nand \U$37206 ( \37549 , \37218 , \19282 );
nand \U$37207 ( \37550 , \37548 , \37549 );
nand \U$37208 ( \37551 , \37541 , \37550 );
nand \U$37209 ( \37552 , \37540 , \37551 );
not \U$37210 ( \37553 , \37552 );
or \U$37211 ( \37554 , \37518 , \37553 );
not \U$37212 ( \37555 , \37516 );
nand \U$37213 ( \37556 , \37555 , \37514 );
nand \U$37214 ( \37557 , \37554 , \37556 );
not \U$37215 ( \37558 , \37557 );
or \U$37216 ( \37559 , \37443 , \37558 );
or \U$37217 ( \37560 , \37557 , \37442 );
not \U$37218 ( \37561 , \9214 );
not \U$37219 ( \37562 , \37399 );
or \U$37220 ( \37563 , \37561 , \37562 );
nand \U$37221 ( \37564 , \37482 , \9195 );
nand \U$37222 ( \37565 , \37563 , \37564 );
not \U$37223 ( \37566 , \9227 );
not \U$37224 ( \37567 , \36907 );
or \U$37225 ( \37568 , \37566 , \37567 );
not \U$37226 ( \37569 , RI9872bf8_170);
not \U$37227 ( \37570 , \24523 );
or \U$37228 ( \37571 , \37569 , \37570 );
or \U$37229 ( \37572 , \24523 , RI9872bf8_170);
nand \U$37230 ( \37573 , \37571 , \37572 );
nand \U$37231 ( \37574 , \37573 , \32292 );
nand \U$37232 ( \37575 , \37568 , \37574 );
xor \U$37233 ( \37576 , \37565 , \37575 );
not \U$37234 ( \37577 , \9294 );
not \U$37235 ( \37578 , \9690 );
not \U$37236 ( \37579 , \24502 );
or \U$37237 ( \37580 , \37578 , \37579 );
or \U$37238 ( \37581 , \13070 , \9694 );
nand \U$37239 ( \37582 , \37580 , \37581 );
not \U$37240 ( \37583 , \37582 );
or \U$37241 ( \37584 , \37577 , \37583 );
nand \U$37242 ( \37585 , \37390 , \10331 );
nand \U$37243 ( \37586 , \37584 , \37585 );
and \U$37244 ( \37587 , \37576 , \37586 );
and \U$37245 ( \37588 , \37565 , \37575 );
or \U$37246 ( \37589 , \37587 , \37588 );
not \U$37247 ( \37590 , \22664 );
xor \U$37248 ( \37591 , \18152 , RI9872d60_173);
not \U$37249 ( \37592 , \37591 );
or \U$37250 ( \37593 , \37590 , \37592 );
nand \U$37251 ( \37594 , \36919 , \8800 );
nand \U$37252 ( \37595 , \37593 , \37594 );
not \U$37253 ( \37596 , \37595 );
not \U$37254 ( \37597 , \7338 );
not \U$37255 ( \37598 , \37074 );
or \U$37256 ( \37599 , \37597 , \37598 );
and \U$37257 ( \37600 , RI98729a0_165, \24867 );
not \U$37258 ( \37601 , RI98729a0_165);
and \U$37259 ( \37602 , \37601 , \24868 );
or \U$37260 ( \37603 , \37600 , \37602 );
nand \U$37261 ( \37604 , \37603 , \7325 );
nand \U$37262 ( \37605 , \37599 , \37604 );
not \U$37263 ( \37606 , \7338 );
not \U$37264 ( \37607 , \37603 );
or \U$37265 ( \37608 , \37606 , \37607 );
not \U$37266 ( \37609 , \7333 );
not \U$37267 ( \37610 , \17702 );
or \U$37268 ( \37611 , \37609 , \37610 );
nand \U$37269 ( \37612 , \18209 , RI98729a0_165);
nand \U$37270 ( \37613 , \37611 , \37612 );
nand \U$37271 ( \37614 , \37613 , \7325 );
nand \U$37272 ( \37615 , \37608 , \37614 );
not \U$37273 ( \37616 , \37615 );
and \U$37274 ( \37617 , \27523 , \5653 );
not \U$37275 ( \37618 , \6285 );
not \U$37276 ( \37619 , \37340 );
or \U$37277 ( \37620 , \37618 , \37619 );
nand \U$37278 ( \37621 , \37453 , \6282 );
nand \U$37279 ( \37622 , \37620 , \37621 );
xor \U$37280 ( \37623 , \37617 , \37622 );
not \U$37281 ( \37624 , \37623 );
or \U$37282 ( \37625 , \37616 , \37624 );
nand \U$37283 ( \37626 , \37622 , \37617 );
nand \U$37284 ( \37627 , \37625 , \37626 );
xor \U$37285 ( \37628 , \37605 , \37627 );
not \U$37286 ( \37629 , \37628 );
or \U$37287 ( \37630 , \37596 , \37629 );
nand \U$37288 ( \37631 , \37627 , \37605 );
nand \U$37289 ( \37632 , \37630 , \37631 );
nor \U$37290 ( \37633 , \37589 , \37632 );
not \U$37291 ( \37634 , \37633 );
not \U$37292 ( \37635 , \37414 );
not \U$37293 ( \37636 , \37404 );
nand \U$37294 ( \37637 , \37636 , \37416 );
not \U$37295 ( \37638 , \37637 );
or \U$37296 ( \37639 , \37635 , \37638 );
or \U$37297 ( \37640 , \37637 , \37414 );
nand \U$37298 ( \37641 , \37639 , \37640 );
nand \U$37299 ( \37642 , \37589 , \37632 );
nand \U$37300 ( \37643 , \37641 , \37642 );
nand \U$37301 ( \37644 , \37634 , \37643 );
not \U$37302 ( \37645 , \37644 );
nand \U$37303 ( \37646 , \37560 , \37645 );
nand \U$37304 ( \37647 , \37559 , \37646 );
xor \U$37305 ( \37648 , \36931 , \36932 );
xor \U$37306 ( \37649 , \37648 , \36935 );
xor \U$37307 ( \37650 , \37647 , \37649 );
not \U$37308 ( \37651 , \37423 );
not \U$37309 ( \37652 , \37383 );
or \U$37310 ( \37653 , \37651 , \37652 );
or \U$37311 ( \37654 , \37383 , \37423 );
nand \U$37312 ( \37655 , \37653 , \37654 );
xor \U$37313 ( \37656 , \37200 , \37210 );
xor \U$37314 ( \37657 , \37656 , \37220 );
not \U$37315 ( \37658 , \37657 );
xor \U$37316 ( \37659 , \37354 , \37343 );
not \U$37317 ( \37660 , \11198 );
not \U$37318 ( \37661 , \37409 );
or \U$37319 ( \37662 , \37660 , \37661 );
not \U$37320 ( \37663 , RI9872f40_177);
not \U$37321 ( \37664 , \12460 );
or \U$37322 ( \37665 , \37663 , \37664 );
or \U$37323 ( \37666 , \12460 , RI9872f40_177);
nand \U$37324 ( \37667 , \37665 , \37666 );
nand \U$37325 ( \37668 , \37667 , \8742 );
nand \U$37326 ( \37669 , \37662 , \37668 );
xnor \U$37327 ( \37670 , \37659 , \37669 );
not \U$37328 ( \37671 , \37670 );
not \U$37329 ( \37672 , \19046 );
not \U$37330 ( \37673 , \37376 );
or \U$37331 ( \37674 , \37672 , \37673 );
not \U$37332 ( \37675 , \8082 );
not \U$37333 ( \37676 , RI98734e0_189);
and \U$37334 ( \37677 , \37675 , \37676 );
and \U$37335 ( \37678 , \7003 , RI98734e0_189);
nor \U$37336 ( \37679 , \37677 , \37678 );
nand \U$37337 ( \37680 , \37679 , \24076 );
nand \U$37338 ( \37681 , \37674 , \37680 );
not \U$37339 ( \37682 , \37681 );
or \U$37340 ( \37683 , \37671 , \37682 );
not \U$37341 ( \37684 , \37659 );
nand \U$37342 ( \37685 , \37684 , \37669 );
nand \U$37343 ( \37686 , \37683 , \37685 );
not \U$37344 ( \37687 , \37686 );
or \U$37345 ( \37688 , \37658 , \37687 );
or \U$37346 ( \37689 , \37686 , \37657 );
xor \U$37347 ( \37690 , \37359 , \37369 );
xor \U$37348 ( \37691 , \37690 , \37380 );
nand \U$37349 ( \37692 , \37689 , \37691 );
nand \U$37350 ( \37693 , \37688 , \37692 );
xor \U$37351 ( \37694 , \37655 , \37693 );
not \U$37352 ( \37695 , \37243 );
not \U$37353 ( \37696 , \37282 );
or \U$37354 ( \37697 , \37695 , \37696 );
or \U$37355 ( \37698 , \37282 , \37243 );
nand \U$37356 ( \37699 , \37697 , \37698 );
and \U$37357 ( \37700 , \37694 , \37699 );
and \U$37358 ( \37701 , \37655 , \37693 );
or \U$37359 ( \37702 , \37700 , \37701 );
and \U$37360 ( \37703 , \37650 , \37702 );
and \U$37361 ( \37704 , \37647 , \37649 );
or \U$37362 ( \37705 , \37703 , \37704 );
xor \U$37363 ( \37706 , \37440 , \37705 );
xor \U$37364 ( \37707 , \37000 , \36938 );
nand \U$37365 ( \37708 , \37706 , \37707 );
not \U$37366 ( \37709 , \37708 );
and \U$37367 ( \37710 , \37440 , \37705 );
nor \U$37368 ( \37711 , \37709 , \37710 );
not \U$37369 ( \37712 , \37711 );
or \U$37370 ( \37713 , \37327 , \37712 );
not \U$37371 ( \37714 , \37710 );
not \U$37372 ( \37715 , \37714 );
not \U$37373 ( \37716 , \37708 );
or \U$37374 ( \37717 , \37715 , \37716 );
not \U$37375 ( \37718 , \37326 );
nand \U$37376 ( \37719 , \37717 , \37718 );
nand \U$37377 ( \37720 , \37713 , \37719 );
not \U$37378 ( \37721 , \37720 );
or \U$37379 ( \37722 , \37320 , \37721 );
nand \U$37380 ( \37723 , \37708 , \37718 , \37714 );
nand \U$37381 ( \37724 , \37722 , \37723 );
nand \U$37382 ( \37725 , \37311 , \37724 );
not \U$37383 ( \37726 , \37318 );
not \U$37384 ( \37727 , \37720 );
or \U$37385 ( \37728 , \37726 , \37727 );
or \U$37386 ( \37729 , \37720 , \37318 );
nand \U$37387 ( \37730 , \37728 , \37729 );
xnor \U$37388 ( \37731 , \37192 , \37190 );
xor \U$37389 ( \37732 , \37731 , \37288 );
not \U$37390 ( \37733 , \37732 );
not \U$37391 ( \37734 , \37707 );
and \U$37392 ( \37735 , \37706 , \37734 );
not \U$37393 ( \37736 , \37706 );
and \U$37394 ( \37737 , \37736 , \37707 );
nor \U$37395 ( \37738 , \37735 , \37737 );
not \U$37396 ( \37739 , \37738 );
or \U$37397 ( \37740 , \37733 , \37739 );
not \U$37398 ( \37741 , \37432 );
nand \U$37399 ( \37742 , \37741 , \37439 );
xor \U$37400 ( \37743 , \37742 , \37436 );
not \U$37401 ( \37744 , \37743 );
not \U$37402 ( \37745 , \37744 );
xor \U$37403 ( \37746 , \37286 , \37194 );
xnor \U$37404 ( \37747 , \37746 , \37234 );
not \U$37405 ( \37748 , \37747 );
not \U$37406 ( \37749 , \37748 );
or \U$37407 ( \37750 , \37745 , \37749 );
not \U$37408 ( \37751 , \37743 );
not \U$37409 ( \37752 , \37747 );
or \U$37410 ( \37753 , \37751 , \37752 );
xor \U$37411 ( \37754 , \37647 , \37649 );
xor \U$37412 ( \37755 , \37754 , \37702 );
nand \U$37413 ( \37756 , \37753 , \37755 );
nand \U$37414 ( \37757 , \37750 , \37756 );
nand \U$37415 ( \37758 , \37740 , \37757 );
not \U$37416 ( \37759 , \37732 );
not \U$37417 ( \37760 , \37738 );
nand \U$37418 ( \37761 , \37759 , \37760 );
and \U$37419 ( \37762 , \37758 , \37761 );
nand \U$37420 ( \37763 , \37730 , \37762 );
nand \U$37421 ( \37764 , \37159 , \37310 , \37725 , \37763 );
not \U$37422 ( \37765 , \37764 );
not \U$37423 ( \37766 , \22618 );
not \U$37424 ( \37767 , \8555 );
xor \U$37425 ( \37768 , RI98730a8_180, \37767 );
not \U$37426 ( \37769 , \37768 );
or \U$37427 ( \37770 , \37766 , \37769 );
and \U$37428 ( \37771 , \13022 , \22752 );
not \U$37429 ( \37772 , \13022 );
and \U$37430 ( \37773 , \37772 , \8722 );
nor \U$37431 ( \37774 , \37771 , \37773 );
nand \U$37432 ( \37775 , \37774 , \13020 );
nand \U$37433 ( \37776 , \37770 , \37775 );
not \U$37434 ( \37777 , \9937 );
and \U$37435 ( \37778 , \14132 , \9750 );
not \U$37436 ( \37779 , \14132 );
and \U$37437 ( \37780 , \37779 , \8696 );
or \U$37438 ( \37781 , \37778 , \37780 );
not \U$37439 ( \37782 , \37781 );
or \U$37440 ( \37783 , \37777 , \37782 );
and \U$37441 ( \37784 , RI9873030_179, \12460 );
not \U$37442 ( \37785 , RI9873030_179);
and \U$37443 ( \37786 , \37785 , \8708 );
or \U$37444 ( \37787 , \37784 , \37786 );
nand \U$37445 ( \37788 , \37787 , \12507 );
nand \U$37446 ( \37789 , \37783 , \37788 );
xor \U$37447 ( \37790 , \37776 , \37789 );
not \U$37448 ( \37791 , \17263 );
not \U$37449 ( \37792 , RI98733f0_187);
not \U$37450 ( \37793 , \9599 );
or \U$37451 ( \37794 , \37792 , \37793 );
or \U$37452 ( \37795 , \11628 , RI98733f0_187);
nand \U$37453 ( \37796 , \37794 , \37795 );
not \U$37454 ( \37797 , \37796 );
or \U$37455 ( \37798 , \37791 , \37797 );
and \U$37456 ( \37799 , \17539 , \35222 );
not \U$37457 ( \37800 , \17539 );
and \U$37458 ( \37801 , \37800 , \10601 );
nor \U$37459 ( \37802 , \37799 , \37801 );
nand \U$37460 ( \37803 , \37802 , \17371 );
nand \U$37461 ( \37804 , \37798 , \37803 );
and \U$37462 ( \37805 , \37790 , \37804 );
and \U$37463 ( \37806 , \37776 , \37789 );
or \U$37464 ( \37807 , \37805 , \37806 );
not \U$37465 ( \37808 , \37807 );
xor \U$37466 ( \37809 , \37623 , \37615 );
not \U$37467 ( \37810 , \9272 );
not \U$37468 ( \37811 , \37582 );
or \U$37469 ( \37812 , \37810 , \37811 );
not \U$37470 ( \37813 , \11358 );
and \U$37471 ( \37814 , RI9872e50_175, \37813 );
not \U$37472 ( \37815 , RI9872e50_175);
and \U$37473 ( \37816 , \37815 , \13876 );
or \U$37474 ( \37817 , \37814 , \37816 );
nand \U$37475 ( \37818 , \37817 , \9293 );
nand \U$37476 ( \37819 , \37812 , \37818 );
xor \U$37477 ( \37820 , \37809 , \37819 );
not \U$37478 ( \37821 , \37820 );
and \U$37479 ( \37822 , \37591 , \8801 );
and \U$37480 ( \37823 , RI9872d60_173, \12773 );
not \U$37481 ( \37824 , RI9872d60_173);
and \U$37482 ( \37825 , \37824 , \32173 );
or \U$37483 ( \37826 , \37823 , \37825 );
and \U$37484 ( \37827 , \37826 , \22664 );
nor \U$37485 ( \37828 , \37822 , \37827 );
not \U$37486 ( \37829 , \37828 );
and \U$37487 ( \37830 , \37821 , \37829 );
and \U$37488 ( \37831 , \37820 , \37828 );
nor \U$37489 ( \37832 , \37830 , \37831 );
not \U$37490 ( \37833 , \37832 );
or \U$37491 ( \37834 , \37808 , \37833 );
or \U$37492 ( \37835 , \37832 , \37807 );
nand \U$37493 ( \37836 , \37834 , \37835 );
buf \U$37494 ( \37837 , \37836 );
not \U$37495 ( \37838 , \19046 );
not \U$37496 ( \37839 , \30509 );
not \U$37497 ( \37840 , RI98734e0_189);
and \U$37498 ( \37841 , \37839 , \37840 );
and \U$37499 ( \37842 , \7467 , RI98734e0_189);
nor \U$37500 ( \37843 , \37841 , \37842 );
not \U$37501 ( \37844 , \37843 );
or \U$37502 ( \37845 , \37838 , \37844 );
and \U$37503 ( \37846 , RI98734e0_189, \9895 );
not \U$37504 ( \37847 , RI98734e0_189);
and \U$37505 ( \37848 , \37847 , \27847 );
or \U$37506 ( \37849 , \37846 , \37848 );
nand \U$37507 ( \37850 , \37849 , \24076 );
nand \U$37508 ( \37851 , \37845 , \37850 );
not \U$37509 ( \37852 , \37851 );
not \U$37510 ( \37853 , \22670 );
not \U$37511 ( \37854 , RI9873210_183);
not \U$37512 ( \37855 , \8650 );
or \U$37513 ( \37856 , \37854 , \37855 );
or \U$37514 ( \37857 , \8650 , RI9873210_183);
nand \U$37515 ( \37858 , \37856 , \37857 );
not \U$37516 ( \37859 , \37858 );
or \U$37517 ( \37860 , \37853 , \37859 );
not \U$37518 ( \37861 , RI9873210_183);
not \U$37519 ( \37862 , \8841 );
or \U$37520 ( \37863 , \37861 , \37862 );
nand \U$37521 ( \37864 , \18312 , \18012 );
nand \U$37522 ( \37865 , \37863 , \37864 );
nand \U$37523 ( \37866 , \37865 , \17243 );
nand \U$37524 ( \37867 , \37860 , \37866 );
not \U$37525 ( \37868 , \9249 );
not \U$37526 ( \37869 , \9185 );
not \U$37527 ( \37870 , \34938 );
or \U$37528 ( \37871 , \37869 , \37870 );
nand \U$37529 ( \37872 , \25380 , RI9872bf8_170);
nand \U$37530 ( \37873 , \37871 , \37872 );
not \U$37531 ( \37874 , \37873 );
or \U$37532 ( \37875 , \37868 , \37874 );
and \U$37533 ( \37876 , RI9872bf8_170, \13860 );
not \U$37534 ( \37877 , RI9872bf8_170);
and \U$37535 ( \37878 , \37877 , \13861 );
or \U$37536 ( \37879 , \37876 , \37878 );
nand \U$37537 ( \37880 , \37879 , \9226 );
nand \U$37538 ( \37881 , \37875 , \37880 );
not \U$37539 ( \37882 , \37881 );
not \U$37540 ( \37883 , \7338 );
and \U$37541 ( \37884 , RI98729a0_165, \18194 );
not \U$37542 ( \37885 , RI98729a0_165);
and \U$37543 ( \37886 , \37885 , \28671 );
or \U$37544 ( \37887 , \37884 , \37886 );
not \U$37545 ( \37888 , \37887 );
or \U$37546 ( \37889 , \37883 , \37888 );
xor \U$37547 ( \37890 , \28663 , RI98729a0_165);
nand \U$37548 ( \37891 , \37890 , \7324 );
nand \U$37549 ( \37892 , \37889 , \37891 );
or \U$37550 ( \37893 , RI9872a18_166, RI9872a90_167);
nand \U$37551 ( \37894 , \37893 , \18704 );
nand \U$37552 ( \37895 , \37894 , \7121 );
not \U$37553 ( \37896 , \37895 );
and \U$37554 ( \37897 , \37892 , \37896 );
not \U$37555 ( \37898 , \9214 );
and \U$37556 ( \37899 , RI9872b80_169, \17908 );
not \U$37557 ( \37900 , RI9872b80_169);
and \U$37558 ( \37901 , \37900 , \17744 );
or \U$37559 ( \37902 , \37899 , \37901 );
not \U$37560 ( \37903 , \37902 );
or \U$37561 ( \37904 , \37898 , \37903 );
not \U$37562 ( \37905 , \9198 );
not \U$37563 ( \37906 , \25409 );
or \U$37564 ( \37907 , \37905 , \37906 );
nand \U$37565 ( \37908 , \24470 , RI9872b80_169);
nand \U$37566 ( \37909 , \37907 , \37908 );
nand \U$37567 ( \37910 , \37909 , \9195 );
nand \U$37568 ( \37911 , \37904 , \37910 );
and \U$37569 ( \37912 , \37897 , \37911 );
not \U$37570 ( \37913 , \37897 );
not \U$37571 ( \37914 , \37911 );
and \U$37572 ( \37915 , \37913 , \37914 );
nor \U$37573 ( \37916 , \37912 , \37915 );
not \U$37574 ( \37917 , \37916 );
or \U$37575 ( \37918 , \37882 , \37917 );
not \U$37576 ( \37919 , \37914 );
nand \U$37577 ( \37920 , \37919 , \37897 );
nand \U$37578 ( \37921 , \37918 , \37920 );
xor \U$37579 ( \37922 , \37867 , \37921 );
not \U$37580 ( \37923 , \37922 );
or \U$37581 ( \37924 , \37852 , \37923 );
nand \U$37582 ( \37925 , \37867 , \37921 );
nand \U$37583 ( \37926 , \37924 , \37925 );
and \U$37584 ( \37927 , \37837 , \37926 );
not \U$37585 ( \37928 , \37837 );
not \U$37586 ( \37929 , \37926 );
and \U$37587 ( \37930 , \37928 , \37929 );
nor \U$37588 ( \37931 , \37927 , \37930 );
not \U$37589 ( \37932 , \9214 );
not \U$37590 ( \37933 , \37909 );
or \U$37591 ( \37934 , \37932 , \37933 );
and \U$37592 ( \37935 , RI9872b80_169, \21553 );
not \U$37593 ( \37936 , RI9872b80_169);
and \U$37594 ( \37937 , \37936 , \19518 );
or \U$37595 ( \37938 , \37935 , \37937 );
nand \U$37596 ( \37939 , \37938 , \9195 );
nand \U$37597 ( \37940 , \37934 , \37939 );
not \U$37598 ( \37941 , \37940 );
and \U$37599 ( \37942 , \37892 , \37895 );
not \U$37600 ( \37943 , \37892 );
and \U$37601 ( \37944 , \37943 , \37896 );
nor \U$37602 ( \37945 , \37942 , \37944 );
not \U$37603 ( \37946 , \37945 );
not \U$37604 ( \37947 , \8039 );
and \U$37605 ( \37948 , RI9872a18_166, \27541 );
not \U$37606 ( \37949 , RI9872a18_166);
and \U$37607 ( \37950 , \37949 , \17703 );
or \U$37608 ( \37951 , \37948 , \37950 );
not \U$37609 ( \37952 , \37951 );
or \U$37610 ( \37953 , \37947 , \37952 );
xor \U$37611 ( \37954 , RI9872a18_166, \17862 );
nand \U$37612 ( \37955 , \37954 , \8027 );
nand \U$37613 ( \37956 , \37953 , \37955 );
not \U$37614 ( \37957 , \37956 );
or \U$37615 ( \37958 , \37946 , \37957 );
or \U$37616 ( \37959 , \37956 , \37945 );
nand \U$37617 ( \37960 , \37958 , \37959 );
not \U$37618 ( \37961 , \37960 );
or \U$37619 ( \37962 , \37941 , \37961 );
not \U$37620 ( \37963 , \37945 );
nand \U$37621 ( \37964 , \37963 , \37956 );
nand \U$37622 ( \37965 , \37962 , \37964 );
not \U$37623 ( \37966 , \37965 );
not \U$37624 ( \37967 , \37966 );
not \U$37625 ( \37968 , \17243 );
and \U$37626 ( \37969 , RI9873210_183, \8554 );
not \U$37627 ( \37970 , RI9873210_183);
and \U$37628 ( \37971 , \37970 , \9760 );
or \U$37629 ( \37972 , \37969 , \37971 );
not \U$37630 ( \37973 , \37972 );
or \U$37631 ( \37974 , \37968 , \37973 );
nand \U$37632 ( \37975 , \37865 , \30963 );
nand \U$37633 ( \37976 , \37974 , \37975 );
not \U$37634 ( \37977 , \37976 );
not \U$37635 ( \37978 , \37977 );
or \U$37636 ( \37979 , \37967 , \37978 );
not \U$37637 ( \37980 , \19035 );
and \U$37638 ( \37981 , RI98734e0_189, \11628 );
not \U$37639 ( \37982 , RI98734e0_189);
and \U$37640 ( \37983 , \37982 , \24779 );
or \U$37641 ( \37984 , \37981 , \37983 );
not \U$37642 ( \37985 , \37984 );
or \U$37643 ( \37986 , \37980 , \37985 );
nand \U$37644 ( \37987 , \37849 , \19046 );
nand \U$37645 ( \37988 , \37986 , \37987 );
nand \U$37646 ( \37989 , \37979 , \37988 );
not \U$37647 ( \37990 , \37966 );
nand \U$37648 ( \37991 , \37990 , \37976 );
nand \U$37649 ( \37992 , \37989 , \37991 );
not \U$37650 ( \37993 , \37992 );
not \U$37651 ( \37994 , \8039 );
xnor \U$37652 ( \37995 , \21553 , RI9872a18_166);
not \U$37653 ( \37996 , \37995 );
or \U$37654 ( \37997 , \37994 , \37996 );
nand \U$37655 ( \37998 , \37951 , \8027 );
nand \U$37656 ( \37999 , \37997 , \37998 );
not \U$37657 ( \38000 , \37999 );
and \U$37658 ( \38001 , \27523 , \6285 );
not \U$37659 ( \38002 , \7338 );
not \U$37660 ( \38003 , \7333 );
not \U$37661 ( \38004 , \17863 );
or \U$37662 ( \38005 , \38003 , \38004 );
or \U$37663 ( \38006 , \17863 , \7333 );
nand \U$37664 ( \38007 , \38005 , \38006 );
not \U$37665 ( \38008 , \38007 );
or \U$37666 ( \38009 , \38002 , \38008 );
nand \U$37667 ( \38010 , \37887 , \7324 );
nand \U$37668 ( \38011 , \38009 , \38010 );
xor \U$37669 ( \38012 , \38001 , \38011 );
not \U$37670 ( \38013 , \38012 );
or \U$37671 ( \38014 , \38000 , \38013 );
nand \U$37672 ( \38015 , \38011 , \38001 );
nand \U$37673 ( \38016 , \38014 , \38015 );
not \U$37674 ( \38017 , \38016 );
not \U$37675 ( \38018 , \37467 );
nor \U$37676 ( \38019 , \38018 , \8021 );
and \U$37677 ( \38020 , \37995 , \8027 );
nor \U$37678 ( \38021 , \38019 , \38020 );
not \U$37679 ( \38022 , \38021 );
and \U$37680 ( \38023 , \38017 , \38022 );
and \U$37681 ( \38024 , \38016 , \38021 );
nor \U$37682 ( \38025 , \38023 , \38024 );
not \U$37683 ( \38026 , \38025 );
not \U$37684 ( \38027 , \9272 );
not \U$37685 ( \38028 , \37817 );
or \U$37686 ( \38029 , \38027 , \38028 );
not \U$37687 ( \38030 , \32953 );
not \U$37688 ( \38031 , \18152 );
or \U$37689 ( \38032 , \38030 , \38031 );
nand \U$37690 ( \38033 , \18151 , RI9872e50_175);
nand \U$37691 ( \38034 , \38032 , \38033 );
nand \U$37692 ( \38035 , \38034 , \18562 );
nand \U$37693 ( \38036 , \38029 , \38035 );
not \U$37694 ( \38037 , \38036 );
or \U$37695 ( \38038 , \38026 , \38037 );
or \U$37696 ( \38039 , \38036 , \38025 );
nand \U$37697 ( \38040 , \38038 , \38039 );
not \U$37698 ( \38041 , \12507 );
and \U$37699 ( \38042 , RI9873030_179, \9114 );
not \U$37700 ( \38043 , RI9873030_179);
and \U$37701 ( \38044 , \38043 , \18344 );
or \U$37702 ( \38045 , \38042 , \38044 );
not \U$37703 ( \38046 , \38045 );
or \U$37704 ( \38047 , \38041 , \38046 );
nand \U$37705 ( \38048 , \37787 , \9937 );
nand \U$37706 ( \38049 , \38047 , \38048 );
not \U$37707 ( \38050 , \38049 );
xor \U$37708 ( \38051 , \37999 , \38012 );
not \U$37709 ( \38052 , \9293 );
not \U$37710 ( \38053 , \9690 );
not \U$37711 ( \38054 , \14193 );
or \U$37712 ( \38055 , \38053 , \38054 );
nand \U$37713 ( \38056 , \13268 , RI9872e50_175);
nand \U$37714 ( \38057 , \38055 , \38056 );
not \U$37715 ( \38058 , \38057 );
or \U$37716 ( \38059 , \38052 , \38058 );
nand \U$37717 ( \38060 , \38034 , \9272 );
nand \U$37718 ( \38061 , \38059 , \38060 );
xor \U$37719 ( \38062 , \38051 , \38061 );
not \U$37720 ( \38063 , \38062 );
or \U$37721 ( \38064 , \38050 , \38063 );
nand \U$37722 ( \38065 , \38061 , \38051 );
nand \U$37723 ( \38066 , \38064 , \38065 );
xor \U$37724 ( \38067 , \38040 , \38066 );
not \U$37725 ( \38068 , \38067 );
or \U$37726 ( \38069 , \37993 , \38068 );
nand \U$37727 ( \38070 , \38066 , \38040 );
nand \U$37728 ( \38071 , \38069 , \38070 );
not \U$37729 ( \38072 , \24209 );
and \U$37730 ( \38073 , RI98730a8_180, \8696 );
not \U$37731 ( \38074 , RI98730a8_180);
and \U$37732 ( \38075 , \38074 , \8697 );
or \U$37733 ( \38076 , \38073 , \38075 );
not \U$37734 ( \38077 , \38076 );
or \U$37735 ( \38078 , \38072 , \38077 );
nand \U$37736 ( \38079 , \37774 , \12867 );
nand \U$37737 ( \38080 , \38078 , \38079 );
not \U$37738 ( \38081 , \17251 );
not \U$37739 ( \38082 , RI98733f0_187);
not \U$37740 ( \38083 , \18107 );
or \U$37741 ( \38084 , \38082 , \38083 );
or \U$37742 ( \38085 , \10308 , RI98733f0_187);
nand \U$37743 ( \38086 , \38084 , \38085 );
not \U$37744 ( \38087 , \38086 );
or \U$37745 ( \38088 , \38081 , \38087 );
nand \U$37746 ( \38089 , \37802 , \17263 );
nand \U$37747 ( \38090 , \38088 , \38089 );
xor \U$37748 ( \38091 , \38080 , \38090 );
not \U$37749 ( \38092 , \18615 );
not \U$37750 ( \38093 , \18239 );
not \U$37751 ( \38094 , \9570 );
or \U$37752 ( \38095 , \38093 , \38094 );
or \U$37753 ( \38096 , \8923 , \18239 );
nand \U$37754 ( \38097 , \38095 , \38096 );
not \U$37755 ( \38098 , \38097 );
or \U$37756 ( \38099 , \38092 , \38098 );
not \U$37757 ( \38100 , \18239 );
not \U$37758 ( \38101 , \7003 );
or \U$37759 ( \38102 , \38100 , \38101 );
nand \U$37760 ( \38103 , \27862 , RI9873558_190);
nand \U$37761 ( \38104 , \38102 , \38103 );
nand \U$37762 ( \38105 , \38104 , RI9873648_192);
nand \U$37763 ( \38106 , \38099 , \38105 );
and \U$37764 ( \38107 , \38091 , \38106 );
and \U$37765 ( \38108 , \38080 , \38090 );
or \U$37766 ( \38109 , \38107 , \38108 );
not \U$37767 ( \38110 , \38109 );
not \U$37768 ( \38111 , \17544 );
xnor \U$37769 ( \38112 , RI9873288_184, \11406 );
not \U$37770 ( \38113 , \38112 );
or \U$37771 ( \38114 , \38111 , \38113 );
not \U$37772 ( \38115 , RI9873288_184);
not \U$37773 ( \38116 , \9880 );
or \U$37774 ( \38117 , \38115 , \38116 );
or \U$37775 ( \38118 , \8857 , RI9873288_184);
nand \U$37776 ( \38119 , \38117 , \38118 );
nand \U$37777 ( \38120 , \38119 , \17528 );
nand \U$37778 ( \38121 , \38114 , \38120 );
not \U$37779 ( \38122 , \38121 );
not \U$37780 ( \38123 , \22664 );
not \U$37781 ( \38124 , \24754 );
and \U$37782 ( \38125 , RI9872d60_173, \38124 );
not \U$37783 ( \38126 , RI9872d60_173);
and \U$37784 ( \38127 , \38126 , \20787 );
nor \U$37785 ( \38128 , \38125 , \38127 );
not \U$37786 ( \38129 , \38128 );
or \U$37787 ( \38130 , \38123 , \38129 );
not \U$37788 ( \38131 , RI9872d60_173);
not \U$37789 ( \38132 , \20928 );
or \U$37790 ( \38133 , \38131 , \38132 );
or \U$37791 ( \38134 , \17090 , RI9872d60_173);
nand \U$37792 ( \38135 , \38133 , \38134 );
nand \U$37793 ( \38136 , \38135 , \8801 );
nand \U$37794 ( \38137 , \38130 , \38136 );
not \U$37795 ( \38138 , \11198 );
not \U$37796 ( \38139 , \8732 );
not \U$37797 ( \38140 , \24502 );
or \U$37798 ( \38141 , \38139 , \38140 );
nand \U$37799 ( \38142 , \17757 , RI9872f40_177);
nand \U$37800 ( \38143 , \38141 , \38142 );
not \U$37801 ( \38144 , \38143 );
or \U$37802 ( \38145 , \38138 , \38144 );
not \U$37803 ( \38146 , \11358 );
and \U$37804 ( \38147 , RI9872f40_177, \38146 );
not \U$37805 ( \38148 , RI9872f40_177);
and \U$37806 ( \38149 , \38148 , \33307 );
or \U$37807 ( \38150 , \38147 , \38149 );
nand \U$37808 ( \38151 , \38150 , \9525 );
nand \U$37809 ( \38152 , \38145 , \38151 );
and \U$37810 ( \38153 , \38137 , \38152 );
not \U$37811 ( \38154 , \38137 );
not \U$37812 ( \38155 , \38152 );
and \U$37813 ( \38156 , \38154 , \38155 );
nor \U$37814 ( \38157 , \38153 , \38156 );
not \U$37815 ( \38158 , \38157 );
or \U$37816 ( \38159 , \38122 , \38158 );
nand \U$37817 ( \38160 , \38152 , \38137 );
nand \U$37818 ( \38161 , \38159 , \38160 );
not \U$37819 ( \38162 , \38161 );
not \U$37820 ( \38163 , \8801 );
not \U$37821 ( \38164 , \37826 );
or \U$37822 ( \38165 , \38163 , \38164 );
nand \U$37823 ( \38166 , \38135 , \8818 );
nand \U$37824 ( \38167 , \38165 , \38166 );
not \U$37825 ( \38168 , \9226 );
and \U$37826 ( \38169 , \24754 , \17164 );
not \U$37827 ( \38170 , \24754 );
and \U$37828 ( \38171 , \38170 , RI9872bf8_170);
nor \U$37829 ( \38172 , \38169 , \38171 );
not \U$37830 ( \38173 , \38172 );
or \U$37831 ( \38174 , \38168 , \38173 );
nand \U$37832 ( \38175 , \37879 , \9249 );
nand \U$37833 ( \38176 , \38174 , \38175 );
not \U$37834 ( \38177 , \9525 );
not \U$37835 ( \38178 , \38143 );
or \U$37836 ( \38179 , \38177 , \38178 );
not \U$37837 ( \38180 , RI9872f40_177);
not \U$37838 ( \38181 , \31511 );
or \U$37839 ( \38182 , \38180 , \38181 );
or \U$37840 ( \38183 , \24729 , RI9872f40_177);
nand \U$37841 ( \38184 , \38182 , \38183 );
nand \U$37842 ( \38185 , \38184 , \11198 );
nand \U$37843 ( \38186 , \38179 , \38185 );
xor \U$37844 ( \38187 , \38176 , \38186 );
xor \U$37845 ( \38188 , \38167 , \38187 );
not \U$37846 ( \38189 , \38188 );
not \U$37847 ( \38190 , \38189 );
or \U$37848 ( \38191 , \38162 , \38190 );
not \U$37849 ( \38192 , \38161 );
nand \U$37850 ( \38193 , \38192 , \38188 );
nand \U$37851 ( \38194 , \38191 , \38193 );
not \U$37852 ( \38195 , \38194 );
or \U$37853 ( \38196 , \38110 , \38195 );
nand \U$37854 ( \38197 , \38188 , \38161 );
nand \U$37855 ( \38198 , \38196 , \38197 );
xor \U$37856 ( \38199 , \38071 , \38198 );
and \U$37857 ( \38200 , \37931 , \38199 );
and \U$37858 ( \38201 , \38071 , \38198 );
nor \U$37859 ( \38202 , \38200 , \38201 );
not \U$37860 ( \38203 , \18508 );
xor \U$37861 ( \38204 , \8597 , RI9873288_184);
not \U$37862 ( \38205 , \38204 );
or \U$37863 ( \38206 , \38203 , \38205 );
nand \U$37864 ( \38207 , \37496 , \17528 );
nand \U$37865 ( \38208 , \38206 , \38207 );
not \U$37866 ( \38209 , \37573 );
or \U$37867 ( \38210 , \38209 , \31277 );
not \U$37868 ( \38211 , \38172 );
not \U$37869 ( \38212 , \9249 );
or \U$37870 ( \38213 , \38211 , \38212 );
nand \U$37871 ( \38214 , \38210 , \38213 );
not \U$37872 ( \38215 , \24627 );
not \U$37873 ( \38216 , \38184 );
or \U$37874 ( \38217 , \38215 , \38216 );
nand \U$37875 ( \38218 , \37667 , \8751 );
nand \U$37876 ( \38219 , \38217 , \38218 );
xor \U$37877 ( \38220 , \38214 , \38219 );
and \U$37878 ( \38221 , \38208 , \38220 );
and \U$37879 ( \38222 , \38214 , \38219 );
nor \U$37880 ( \38223 , \38221 , \38222 );
not \U$37881 ( \38224 , \29633 );
not \U$37882 ( \38225 , \37768 );
or \U$37883 ( \38226 , \38224 , \38225 );
nand \U$37884 ( \38227 , \37525 , \17347 );
nand \U$37885 ( \38228 , \38226 , \38227 );
not \U$37886 ( \38229 , \17243 );
not \U$37887 ( \38230 , \37858 );
or \U$37888 ( \38231 , \38229 , \38230 );
nand \U$37889 ( \38232 , \37508 , \17234 );
nand \U$37890 ( \38233 , \38231 , \38232 );
xor \U$37891 ( \38234 , \38228 , \38233 );
not \U$37892 ( \38235 , \17251 );
not \U$37893 ( \38236 , \37796 );
or \U$37894 ( \38237 , \38235 , \38236 );
nand \U$37895 ( \38238 , \37546 , \17263 );
nand \U$37896 ( \38239 , \38237 , \38238 );
and \U$37897 ( \38240 , \38234 , \38239 );
and \U$37898 ( \38241 , \38228 , \38233 );
or \U$37899 ( \38242 , \38240 , \38241 );
not \U$37900 ( \38243 , \38242 );
xor \U$37901 ( \38244 , \38223 , \38243 );
not \U$37902 ( \38245 , \18615 );
not \U$37903 ( \38246 , \10412 );
not \U$37904 ( \38247 , RI9873558_190);
and \U$37905 ( \38248 , \38246 , \38247 );
and \U$37906 ( \38249 , \7905 , RI9873558_190);
nor \U$37907 ( \38250 , \38248 , \38249 );
not \U$37908 ( \38251 , \38250 );
or \U$37909 ( \38252 , \38245 , \38251 );
nand \U$37910 ( \38253 , \37534 , RI9873648_192);
nand \U$37911 ( \38254 , \38252 , \38253 );
not \U$37912 ( \38255 , \38254 );
not \U$37913 ( \38256 , \9214 );
not \U$37914 ( \38257 , \37475 );
or \U$37915 ( \38258 , \38256 , \38257 );
nand \U$37916 ( \38259 , \37902 , \9195 );
nand \U$37917 ( \38260 , \38258 , \38259 );
not \U$37918 ( \38261 , \38260 );
not \U$37919 ( \38262 , \38261 );
not \U$37920 ( \38263 , \7338 );
not \U$37921 ( \38264 , \37613 );
or \U$37922 ( \38265 , \38263 , \38264 );
nand \U$37923 ( \38266 , \38007 , \7325 );
nand \U$37924 ( \38267 , \38265 , \38266 );
xor \U$37925 ( \38268 , \37448 , \37458 );
xnor \U$37926 ( \38269 , \38267 , \38268 );
not \U$37927 ( \38270 , \38269 );
and \U$37928 ( \38271 , \38262 , \38270 );
and \U$37929 ( \38272 , \38267 , \38268 );
nor \U$37930 ( \38273 , \38271 , \38272 );
not \U$37931 ( \38274 , \38273 );
not \U$37932 ( \38275 , \38274 );
or \U$37933 ( \38276 , \38255 , \38275 );
and \U$37934 ( \38277 , \37679 , \20147 );
and \U$37935 ( \38278 , \37843 , \19243 );
nor \U$37936 ( \38279 , \38277 , \38278 );
not \U$37937 ( \38280 , \38279 );
and \U$37938 ( \38281 , \38254 , \38274 );
not \U$37939 ( \38282 , \38254 );
and \U$37940 ( \38283 , \38282 , \38273 );
nor \U$37941 ( \38284 , \38281 , \38283 );
nand \U$37942 ( \38285 , \38280 , \38284 );
nand \U$37943 ( \38286 , \38276 , \38285 );
xnor \U$37944 ( \38287 , \38244 , \38286 );
not \U$37945 ( \38288 , \38287 );
not \U$37946 ( \38289 , \38288 );
not \U$37947 ( \38290 , \9937 );
not \U$37948 ( \38291 , \37206 );
or \U$37949 ( \38292 , \38290 , \38291 );
and \U$37950 ( \38293 , RI9873030_179, \12470 );
not \U$37951 ( \38294 , RI9873030_179);
and \U$37952 ( \38295 , \38294 , \18498 );
nor \U$37953 ( \38296 , \38293 , \38295 );
nand \U$37954 ( \38297 , \38296 , \12507 );
nand \U$37955 ( \38298 , \38292 , \38297 );
not \U$37956 ( \38299 , \38298 );
not \U$37957 ( \38300 , \37595 );
not \U$37958 ( \38301 , \38300 );
not \U$37959 ( \38302 , \37628 );
and \U$37960 ( \38303 , \38301 , \38302 );
and \U$37961 ( \38304 , \38300 , \37628 );
nor \U$37962 ( \38305 , \38303 , \38304 );
not \U$37963 ( \38306 , \38305 );
or \U$37964 ( \38307 , \38299 , \38306 );
or \U$37965 ( \38308 , \38298 , \38305 );
nand \U$37966 ( \38309 , \38307 , \38308 );
not \U$37967 ( \38310 , \37828 );
not \U$37968 ( \38311 , \38310 );
not \U$37969 ( \38312 , \37820 );
or \U$37970 ( \38313 , \38311 , \38312 );
nand \U$37971 ( \38314 , \37819 , \37809 );
nand \U$37972 ( \38315 , \38313 , \38314 );
xor \U$37973 ( \38316 , \38309 , \38315 );
not \U$37974 ( \38317 , \38167 );
not \U$37975 ( \38318 , \38187 );
or \U$37976 ( \38319 , \38317 , \38318 );
nand \U$37977 ( \38320 , \38186 , \38176 );
nand \U$37978 ( \38321 , \38319 , \38320 );
not \U$37979 ( \38322 , \38269 );
not \U$37980 ( \38323 , \38260 );
or \U$37981 ( \38324 , \38322 , \38323 );
or \U$37982 ( \38325 , \38260 , \38269 );
nand \U$37983 ( \38326 , \38324 , \38325 );
not \U$37984 ( \38327 , \17528 );
not \U$37985 ( \38328 , \38204 );
or \U$37986 ( \38329 , \38327 , \38328 );
nand \U$37987 ( \38330 , \38119 , \17544 );
nand \U$37988 ( \38331 , \38329 , \38330 );
xor \U$37989 ( \38332 , \38326 , \38331 );
not \U$37990 ( \38333 , RI9873648_192);
not \U$37991 ( \38334 , \38250 );
or \U$37992 ( \38335 , \38333 , \38334 );
nand \U$37993 ( \38336 , \38104 , \18545 );
nand \U$37994 ( \38337 , \38335 , \38336 );
and \U$37995 ( \38338 , \38332 , \38337 );
and \U$37996 ( \38339 , \38326 , \38331 );
or \U$37997 ( \38340 , \38338 , \38339 );
xor \U$37998 ( \38341 , \38321 , \38340 );
xor \U$37999 ( \38342 , \38208 , \38220 );
and \U$38000 ( \38343 , \38341 , \38342 );
and \U$38001 ( \38344 , \38321 , \38340 );
nor \U$38002 ( \38345 , \38343 , \38344 );
xnor \U$38003 ( \38346 , \38316 , \38345 );
not \U$38004 ( \38347 , \38346 );
not \U$38005 ( \38348 , \38347 );
or \U$38006 ( \38349 , \38289 , \38348 );
nand \U$38007 ( \38350 , \38287 , \38346 );
nand \U$38008 ( \38351 , \38349 , \38350 );
xor \U$38009 ( \38352 , \38202 , \38351 );
not \U$38010 ( \38353 , \38025 );
not \U$38011 ( \38354 , \38353 );
not \U$38012 ( \38355 , \38036 );
or \U$38013 ( \38356 , \38354 , \38355 );
not \U$38014 ( \38357 , \38021 );
nand \U$38015 ( \38358 , \38357 , \38016 );
nand \U$38016 ( \38359 , \38356 , \38358 );
not \U$38017 ( \38360 , \38359 );
not \U$38018 ( \38361 , \38360 );
not \U$38019 ( \38362 , \9937 );
not \U$38020 ( \38363 , \38296 );
or \U$38021 ( \38364 , \38362 , \38363 );
nand \U$38022 ( \38365 , \37781 , \12507 );
nand \U$38023 ( \38366 , \38364 , \38365 );
not \U$38024 ( \38367 , \37484 );
and \U$38025 ( \38368 , \37470 , \38367 );
not \U$38026 ( \38369 , \37470 );
and \U$38027 ( \38370 , \38369 , \37484 );
nor \U$38028 ( \38371 , \38368 , \38370 );
not \U$38029 ( \38372 , \38371 );
and \U$38030 ( \38373 , \38366 , \38372 );
not \U$38031 ( \38374 , \38366 );
and \U$38032 ( \38375 , \38374 , \38371 );
nor \U$38033 ( \38376 , \38373 , \38375 );
not \U$38034 ( \38377 , \38376 );
or \U$38035 ( \38378 , \38361 , \38377 );
or \U$38036 ( \38379 , \38376 , \38360 );
nand \U$38037 ( \38380 , \38378 , \38379 );
xor \U$38038 ( \38381 , \38228 , \38233 );
xor \U$38039 ( \38382 , \38381 , \38239 );
xor \U$38040 ( \38383 , \38380 , \38382 );
xnor \U$38041 ( \38384 , \38279 , \38284 );
xor \U$38042 ( \38385 , \38383 , \38384 );
not \U$38043 ( \38386 , \38385 );
xor \U$38044 ( \38387 , \38342 , \38341 );
xor \U$38045 ( \38388 , \37776 , \37789 );
xor \U$38046 ( \38389 , \38388 , \37804 );
not \U$38047 ( \38390 , \38389 );
not \U$38048 ( \38391 , \37851 );
not \U$38049 ( \38392 , \38391 );
not \U$38050 ( \38393 , \37922 );
or \U$38051 ( \38394 , \38392 , \38393 );
or \U$38052 ( \38395 , \37922 , \38391 );
nand \U$38053 ( \38396 , \38394 , \38395 );
xor \U$38054 ( \38397 , \38326 , \38331 );
xor \U$38055 ( \38398 , \38397 , \38337 );
xor \U$38056 ( \38399 , \38396 , \38398 );
not \U$38057 ( \38400 , \38399 );
or \U$38058 ( \38401 , \38390 , \38400 );
nand \U$38059 ( \38402 , \38396 , \38398 );
nand \U$38060 ( \38403 , \38401 , \38402 );
xor \U$38061 ( \38404 , \38387 , \38403 );
not \U$38062 ( \38405 , \38404 );
or \U$38063 ( \38406 , \38386 , \38405 );
nand \U$38064 ( \38407 , \38403 , \38387 );
nand \U$38065 ( \38408 , \38406 , \38407 );
xor \U$38066 ( \38409 , \38352 , \38408 );
xor \U$38067 ( \38410 , \38380 , \38382 );
and \U$38068 ( \38411 , \38410 , \38384 );
and \U$38069 ( \38412 , \38380 , \38382 );
or \U$38070 ( \38413 , \38411 , \38412 );
and \U$38071 ( \38414 , \37499 , \37488 );
not \U$38072 ( \38415 , \37499 );
and \U$38073 ( \38416 , \38415 , \37487 );
nor \U$38074 ( \38417 , \38414 , \38416 );
xnor \U$38075 ( \38418 , \37510 , \38417 );
not \U$38076 ( \38419 , \38418 );
xor \U$38077 ( \38420 , \37565 , \37575 );
xor \U$38078 ( \38421 , \38420 , \37586 );
not \U$38079 ( \38422 , \38421 );
and \U$38080 ( \38423 , \38419 , \38422 );
and \U$38081 ( \38424 , \38418 , \38421 );
nor \U$38082 ( \38425 , \38423 , \38424 );
not \U$38083 ( \38426 , \38425 );
not \U$38084 ( \38427 , \37527 );
and \U$38085 ( \38428 , \37550 , \38427 );
not \U$38086 ( \38429 , \37550 );
and \U$38087 ( \38430 , \38429 , \37527 );
nor \U$38088 ( \38431 , \38428 , \38430 );
xnor \U$38089 ( \38432 , \37538 , \38431 );
not \U$38090 ( \38433 , \38432 );
and \U$38091 ( \38434 , \38426 , \38433 );
and \U$38092 ( \38435 , \38425 , \38432 );
nor \U$38093 ( \38436 , \38434 , \38435 );
and \U$38094 ( \38437 , \38413 , \38436 );
not \U$38095 ( \38438 , \38413 );
not \U$38096 ( \38439 , \38436 );
and \U$38097 ( \38440 , \38438 , \38439 );
nor \U$38098 ( \38441 , \38437 , \38440 );
not \U$38099 ( \38442 , \37926 );
not \U$38100 ( \38443 , \37836 );
or \U$38101 ( \38444 , \38442 , \38443 );
not \U$38102 ( \38445 , \37832 );
nand \U$38103 ( \38446 , \38445 , \37807 );
nand \U$38104 ( \38447 , \38444 , \38446 );
not \U$38105 ( \38448 , \38447 );
not \U$38106 ( \38449 , \38371 );
not \U$38107 ( \38450 , \38360 );
or \U$38108 ( \38451 , \38449 , \38450 );
not \U$38109 ( \38452 , \38366 );
not \U$38110 ( \38453 , \38371 );
nand \U$38111 ( \38454 , \38453 , \38359 );
nand \U$38112 ( \38455 , \38452 , \38454 );
nand \U$38113 ( \38456 , \38451 , \38455 );
not \U$38114 ( \38457 , \38456 );
and \U$38115 ( \38458 , \37681 , \37670 );
not \U$38116 ( \38459 , \37681 );
not \U$38117 ( \38460 , \37670 );
and \U$38118 ( \38461 , \38459 , \38460 );
nor \U$38119 ( \38462 , \38458 , \38461 );
nand \U$38120 ( \38463 , \38457 , \38462 );
not \U$38121 ( \38464 , \38462 );
nand \U$38122 ( \38465 , \38464 , \38456 );
nand \U$38123 ( \38466 , \38463 , \38465 );
not \U$38124 ( \38467 , \38466 );
and \U$38125 ( \38468 , \38448 , \38467 );
and \U$38126 ( \38469 , \38447 , \38466 );
nor \U$38127 ( \38470 , \38468 , \38469 );
and \U$38128 ( \38471 , \38441 , \38470 );
not \U$38129 ( \38472 , \38441 );
not \U$38130 ( \38473 , \38470 );
and \U$38131 ( \38474 , \38472 , \38473 );
or \U$38132 ( \38475 , \38471 , \38474 );
not \U$38133 ( \38476 , \11198 );
not \U$38134 ( \38477 , \38150 );
or \U$38135 ( \38478 , \38476 , \38477 );
not \U$38136 ( \38479 , \8732 );
not \U$38137 ( \38480 , \28628 );
or \U$38138 ( \38481 , \38479 , \38480 );
nand \U$38139 ( \38482 , \18155 , RI9872f40_177);
nand \U$38140 ( \38483 , \38481 , \38482 );
nand \U$38141 ( \38484 , \38483 , \24627 );
nand \U$38142 ( \38485 , \38478 , \38484 );
not \U$38143 ( \38486 , \38485 );
not \U$38144 ( \38487 , \8801 );
not \U$38145 ( \38488 , \38128 );
or \U$38146 ( \38489 , \38487 , \38488 );
and \U$38147 ( \38490 , RI9872d60_173, \17013 );
not \U$38148 ( \38491 , RI9872d60_173);
and \U$38149 ( \38492 , \38491 , \35645 );
or \U$38150 ( \38493 , \38490 , \38492 );
nand \U$38151 ( \38494 , \38493 , \22664 );
nand \U$38152 ( \38495 , \38489 , \38494 );
not \U$38153 ( \38496 , \38495 );
not \U$38154 ( \38497 , \9272 );
not \U$38155 ( \38498 , \38057 );
or \U$38156 ( \38499 , \38497 , \38498 );
not \U$38157 ( \38500 , \19591 );
xor \U$38158 ( \38501 , RI9872e50_175, \38500 );
nand \U$38159 ( \38502 , \38501 , \9294 );
nand \U$38160 ( \38503 , \38499 , \38502 );
not \U$38161 ( \38504 , \38503 );
not \U$38162 ( \38505 , \38504 );
or \U$38163 ( \38506 , \38496 , \38505 );
or \U$38164 ( \38507 , \38504 , \38495 );
nand \U$38165 ( \38508 , \38506 , \38507 );
not \U$38166 ( \38509 , \38508 );
or \U$38167 ( \38510 , \38486 , \38509 );
nand \U$38168 ( \38511 , \38503 , \38495 );
nand \U$38169 ( \38512 , \38510 , \38511 );
not \U$38170 ( \38513 , \38512 );
not \U$38171 ( \38514 , \37881 );
and \U$38172 ( \38515 , \37916 , \38514 );
not \U$38173 ( \38516 , \37916 );
and \U$38174 ( \38517 , \38516 , \37881 );
nor \U$38175 ( \38518 , \38515 , \38517 );
not \U$38176 ( \38519 , \38518 );
not \U$38177 ( \38520 , \38519 );
not \U$38178 ( \38521 , \9214 );
not \U$38179 ( \38522 , \37938 );
or \U$38180 ( \38523 , \38521 , \38522 );
xor \U$38181 ( \38524 , RI9872b80_169, \17702 );
nand \U$38182 ( \38525 , \38524 , \9195 );
nand \U$38183 ( \38526 , \38523 , \38525 );
not \U$38184 ( \38527 , \38526 );
and \U$38185 ( \38528 , \18704 , \7338 );
not \U$38186 ( \38529 , \8039 );
not \U$38187 ( \38530 , \37954 );
or \U$38188 ( \38531 , \38529 , \38530 );
not \U$38189 ( \38532 , \21773 );
xor \U$38190 ( \38533 , RI9872a18_166, \38532 );
nand \U$38191 ( \38534 , \38533 , \8026 );
nand \U$38192 ( \38535 , \38531 , \38534 );
xor \U$38193 ( \38536 , \38528 , \38535 );
not \U$38194 ( \38537 , \38536 );
or \U$38195 ( \38538 , \38527 , \38537 );
nand \U$38196 ( \38539 , \38535 , \38528 );
nand \U$38197 ( \38540 , \38538 , \38539 );
not \U$38198 ( \38541 , \38540 );
not \U$38199 ( \38542 , \9226 );
not \U$38200 ( \38543 , \37873 );
or \U$38201 ( \38544 , \38542 , \38543 );
and \U$38202 ( \38545 , RI9872bf8_170, \17908 );
not \U$38203 ( \38546 , RI9872bf8_170);
and \U$38204 ( \38547 , \38546 , \32208 );
or \U$38205 ( \38548 , \38545 , \38547 );
nand \U$38206 ( \38549 , \38548 , \9249 );
nand \U$38207 ( \38550 , \38544 , \38549 );
not \U$38208 ( \38551 , \38550 );
not \U$38209 ( \38552 , \38551 );
or \U$38210 ( \38553 , \38541 , \38552 );
or \U$38211 ( \38554 , \38551 , \38540 );
nand \U$38212 ( \38555 , \38553 , \38554 );
not \U$38213 ( \38556 , \38555 );
not \U$38214 ( \38557 , \12507 );
and \U$38215 ( \38558 , RI9873030_179, \35562 );
not \U$38216 ( \38559 , RI9873030_179);
and \U$38217 ( \38560 , \38559 , \13070 );
or \U$38218 ( \38561 , \38558 , \38560 );
not \U$38219 ( \38562 , \38561 );
or \U$38220 ( \38563 , \38557 , \38562 );
nand \U$38221 ( \38564 , \38045 , \9937 );
nand \U$38222 ( \38565 , \38563 , \38564 );
not \U$38223 ( \38566 , \38565 );
or \U$38224 ( \38567 , \38556 , \38566 );
nand \U$38225 ( \38568 , \38550 , \38540 );
nand \U$38226 ( \38569 , \38567 , \38568 );
not \U$38227 ( \38570 , \38569 );
not \U$38228 ( \38571 , \38570 );
or \U$38229 ( \38572 , \38520 , \38571 );
nand \U$38230 ( \38573 , \38569 , \38518 );
nand \U$38231 ( \38574 , \38572 , \38573 );
not \U$38232 ( \38575 , \38574 );
or \U$38233 ( \38576 , \38513 , \38575 );
nand \U$38234 ( \38577 , \38569 , \38519 );
nand \U$38235 ( \38578 , \38576 , \38577 );
not \U$38236 ( \38579 , \38067 );
not \U$38237 ( \38580 , \37992 );
not \U$38238 ( \38581 , \38580 );
and \U$38239 ( \38582 , \38579 , \38581 );
and \U$38240 ( \38583 , \38067 , \38580 );
nor \U$38241 ( \38584 , \38582 , \38583 );
not \U$38242 ( \38585 , \38584 );
xor \U$38243 ( \38586 , \38578 , \38585 );
not \U$38244 ( \38587 , \12867 );
not \U$38245 ( \38588 , \38076 );
or \U$38246 ( \38589 , \38587 , \38588 );
and \U$38247 ( \38590 , RI98730a8_180, \8708 );
not \U$38248 ( \38591 , RI98730a8_180);
and \U$38249 ( \38592 , \38591 , \12460 );
nor \U$38250 ( \38593 , \38590 , \38592 );
nand \U$38251 ( \38594 , \38593 , \13020 );
nand \U$38252 ( \38595 , \38589 , \38594 );
not \U$38253 ( \38596 , \30963 );
not \U$38254 ( \38597 , \37972 );
or \U$38255 ( \38598 , \38596 , \38597 );
and \U$38256 ( \38599 , RI9873210_183, \22752 );
not \U$38257 ( \38600 , RI9873210_183);
and \U$38258 ( \38601 , \38600 , \10099 );
or \U$38259 ( \38602 , \38599 , \38601 );
nand \U$38260 ( \38603 , \38602 , \13476 );
nand \U$38261 ( \38604 , \38598 , \38603 );
xor \U$38262 ( \38605 , \38595 , \38604 );
not \U$38263 ( \38606 , \18545 );
not \U$38264 ( \38607 , \18239 );
not \U$38265 ( \38608 , \12727 );
or \U$38266 ( \38609 , \38607 , \38608 );
or \U$38267 ( \38610 , \9898 , \18239 );
nand \U$38268 ( \38611 , \38609 , \38610 );
not \U$38269 ( \38612 , \38611 );
or \U$38270 ( \38613 , \38606 , \38612 );
nand \U$38271 ( \38614 , \38097 , RI9873648_192);
nand \U$38272 ( \38615 , \38613 , \38614 );
and \U$38273 ( \38616 , \38605 , \38615 );
and \U$38274 ( \38617 , \38595 , \38604 );
or \U$38275 ( \38618 , \38616 , \38617 );
xor \U$38276 ( \38619 , \38121 , \38157 );
or \U$38277 ( \38620 , \38618 , \38619 );
or \U$38278 ( \38621 , RI9872b08_168, RI9872b80_169);
nand \U$38279 ( \38622 , \38621 , \18704 );
and \U$38280 ( \38623 , \38622 , \7902 );
not \U$38281 ( \38624 , \8039 );
not \U$38282 ( \38625 , \38533 );
or \U$38283 ( \38626 , \38624 , \38625 );
xor \U$38284 ( \38627 , \18704 , RI9872a18_166);
nand \U$38285 ( \38628 , \38627 , \8026 );
nand \U$38286 ( \38629 , \38626 , \38628 );
and \U$38287 ( \38630 , \38623 , \38629 );
not \U$38288 ( \38631 , \9249 );
xnor \U$38289 ( \38632 , \17726 , RI9872bf8_170);
not \U$38290 ( \38633 , \38632 );
or \U$38291 ( \38634 , \38631 , \38633 );
nand \U$38292 ( \38635 , \38548 , \9226 );
nand \U$38293 ( \38636 , \38634 , \38635 );
xor \U$38294 ( \38637 , \38630 , \38636 );
not \U$38295 ( \38638 , \8817 );
not \U$38296 ( \38639 , RI9872d60_173);
buf \U$38297 ( \38640 , \29412 );
not \U$38298 ( \38641 , \38640 );
or \U$38299 ( \38642 , \38639 , \38641 );
or \U$38300 ( \38643 , \20450 , RI9872d60_173);
nand \U$38301 ( \38644 , \38642 , \38643 );
not \U$38302 ( \38645 , \38644 );
or \U$38303 ( \38646 , \38638 , \38645 );
nand \U$38304 ( \38647 , \38493 , \8800 );
nand \U$38305 ( \38648 , \38646 , \38647 );
and \U$38306 ( \38649 , \38637 , \38648 );
and \U$38307 ( \38650 , \38630 , \38636 );
or \U$38308 ( \38651 , \38649 , \38650 );
not \U$38309 ( \38652 , \17528 );
not \U$38310 ( \38653 , \38112 );
or \U$38311 ( \38654 , \38652 , \38653 );
not \U$38312 ( \38655 , RI9873288_184);
not \U$38313 ( \38656 , \12849 );
or \U$38314 ( \38657 , \38655 , \38656 );
not \U$38315 ( \38658 , \34990 );
nand \U$38316 ( \38659 , \38658 , \22715 );
nand \U$38317 ( \38660 , \38657 , \38659 );
nand \U$38318 ( \38661 , \38660 , \18508 );
nand \U$38319 ( \38662 , \38654 , \38661 );
xor \U$38320 ( \38663 , \38651 , \38662 );
not \U$38321 ( \38664 , \19046 );
not \U$38322 ( \38665 , \37984 );
or \U$38323 ( \38666 , \38664 , \38665 );
and \U$38324 ( \38667 , RI98734e0_189, \8874 );
not \U$38325 ( \38668 , RI98734e0_189);
and \U$38326 ( \38669 , \38668 , \8877 );
or \U$38327 ( \38670 , \38667 , \38669 );
nand \U$38328 ( \38671 , \38670 , \24076 );
nand \U$38329 ( \38672 , \38666 , \38671 );
and \U$38330 ( \38673 , \38663 , \38672 );
and \U$38331 ( \38674 , \38651 , \38662 );
or \U$38332 ( \38675 , \38673 , \38674 );
nand \U$38333 ( \38676 , \38620 , \38675 );
nand \U$38334 ( \38677 , \38618 , \38619 );
nand \U$38335 ( \38678 , \38676 , \38677 );
and \U$38336 ( \38679 , \38586 , \38678 );
and \U$38337 ( \38680 , \38578 , \38585 );
nor \U$38338 ( \38681 , \38679 , \38680 );
xnor \U$38339 ( \38682 , \38062 , \38049 );
not \U$38340 ( \38683 , \38682 );
xor \U$38341 ( \38684 , \37966 , \37976 );
xor \U$38342 ( \38685 , \38684 , \37988 );
not \U$38343 ( \38686 , \38685 );
or \U$38344 ( \38687 , \38683 , \38686 );
xor \U$38345 ( \38688 , \38080 , \38090 );
xor \U$38346 ( \38689 , \38688 , \38106 );
nand \U$38347 ( \38690 , \38687 , \38689 );
or \U$38348 ( \38691 , \38685 , \38682 );
nand \U$38349 ( \38692 , \38690 , \38691 );
not \U$38350 ( \38693 , \38692 );
not \U$38351 ( \38694 , \38109 );
and \U$38352 ( \38695 , \38194 , \38694 );
not \U$38353 ( \38696 , \38194 );
and \U$38354 ( \38697 , \38696 , \38109 );
nor \U$38355 ( \38698 , \38695 , \38697 );
not \U$38356 ( \38699 , \38698 );
not \U$38357 ( \38700 , \38699 );
or \U$38358 ( \38701 , \38693 , \38700 );
not \U$38359 ( \38702 , \38389 );
and \U$38360 ( \38703 , \38399 , \38702 );
not \U$38361 ( \38704 , \38399 );
and \U$38362 ( \38705 , \38704 , \38389 );
nor \U$38363 ( \38706 , \38703 , \38705 );
not \U$38364 ( \38707 , \38706 );
not \U$38365 ( \38708 , \38699 );
not \U$38366 ( \38709 , \38692 );
not \U$38367 ( \38710 , \38709 );
or \U$38368 ( \38711 , \38708 , \38710 );
nand \U$38369 ( \38712 , \38692 , \38698 );
nand \U$38370 ( \38713 , \38711 , \38712 );
nand \U$38371 ( \38714 , \38707 , \38713 );
nand \U$38372 ( \38715 , \38701 , \38714 );
not \U$38373 ( \38716 , \38715 );
xor \U$38374 ( \38717 , \38681 , \38716 );
not \U$38375 ( \38718 , \37931 );
not \U$38376 ( \38719 , \38718 );
not \U$38377 ( \38720 , \38199 );
and \U$38378 ( \38721 , \38719 , \38720 );
and \U$38379 ( \38722 , \38199 , \38718 );
nor \U$38380 ( \38723 , \38721 , \38722 );
and \U$38381 ( \38724 , \38717 , \38723 );
and \U$38382 ( \38725 , \38681 , \38716 );
or \U$38383 ( \38726 , \38724 , \38725 );
xor \U$38384 ( \38727 , \38475 , \38726 );
and \U$38385 ( \38728 , \38409 , \38727 );
not \U$38386 ( \38729 , \38409 );
not \U$38387 ( \38730 , \38727 );
and \U$38388 ( \38731 , \38729 , \38730 );
nor \U$38389 ( \38732 , \38728 , \38731 );
not \U$38390 ( \38733 , \38385 );
and \U$38391 ( \38734 , \38404 , \38733 );
not \U$38392 ( \38735 , \38404 );
and \U$38393 ( \38736 , \38735 , \38385 );
nor \U$38394 ( \38737 , \38734 , \38736 );
not \U$38395 ( \38738 , \38574 );
not \U$38396 ( \38739 , \38512 );
not \U$38397 ( \38740 , \38739 );
or \U$38398 ( \38741 , \38738 , \38740 );
or \U$38399 ( \38742 , \38739 , \38574 );
nand \U$38400 ( \38743 , \38741 , \38742 );
not \U$38401 ( \38744 , \24209 );
and \U$38402 ( \38745 , RI98730a8_180, \9119 );
not \U$38403 ( \38746 , RI98730a8_180);
and \U$38404 ( \38747 , \38746 , \9114 );
nor \U$38405 ( \38748 , \38745 , \38747 );
not \U$38406 ( \38749 , \38748 );
or \U$38407 ( \38750 , \38744 , \38749 );
nand \U$38408 ( \38751 , \38593 , \17347 );
nand \U$38409 ( \38752 , \38750 , \38751 );
not \U$38410 ( \38753 , \38752 );
not \U$38411 ( \38754 , \9293 );
not \U$38412 ( \38755 , RI9872e50_175);
not \U$38413 ( \38756 , \17783 );
or \U$38414 ( \38757 , \38755 , \38756 );
or \U$38415 ( \38758 , \20787 , RI9872e50_175);
nand \U$38416 ( \38759 , \38757 , \38758 );
not \U$38417 ( \38760 , \38759 );
or \U$38418 ( \38761 , \38754 , \38760 );
nand \U$38419 ( \38762 , \38501 , \9272 );
nand \U$38420 ( \38763 , \38761 , \38762 );
not \U$38421 ( \38764 , \38763 );
not \U$38422 ( \38765 , \38526 );
and \U$38423 ( \38766 , \38536 , \38765 );
not \U$38424 ( \38767 , \38536 );
and \U$38425 ( \38768 , \38767 , \38526 );
nor \U$38426 ( \38769 , \38766 , \38768 );
not \U$38427 ( \38770 , \38769 );
and \U$38428 ( \38771 , \38764 , \38770 );
and \U$38429 ( \38772 , \38763 , \38769 );
nor \U$38430 ( \38773 , \38771 , \38772 );
not \U$38431 ( \38774 , \38773 );
not \U$38432 ( \38775 , \38774 );
or \U$38433 ( \38776 , \38753 , \38775 );
not \U$38434 ( \38777 , \38769 );
nand \U$38435 ( \38778 , \38777 , \38763 );
nand \U$38436 ( \38779 , \38776 , \38778 );
not \U$38437 ( \38780 , \38779 );
xor \U$38438 ( \38781 , \37960 , \37940 );
not \U$38439 ( \38782 , \38781 );
not \U$38440 ( \38783 , \17251 );
not \U$38441 ( \38784 , RI98733f0_187);
not \U$38442 ( \38785 , \8668 );
or \U$38443 ( \38786 , \38784 , \38785 );
or \U$38444 ( \38787 , \8857 , RI98733f0_187);
nand \U$38445 ( \38788 , \38786 , \38787 );
not \U$38446 ( \38789 , \38788 );
or \U$38447 ( \38790 , \38783 , \38789 );
nand \U$38448 ( \38791 , \38086 , \17263 );
nand \U$38449 ( \38792 , \38790 , \38791 );
not \U$38450 ( \38793 , \38792 );
not \U$38451 ( \38794 , \38793 );
or \U$38452 ( \38795 , \38782 , \38794 );
or \U$38453 ( \38796 , \38793 , \38781 );
nand \U$38454 ( \38797 , \38795 , \38796 );
not \U$38455 ( \38798 , \38797 );
or \U$38456 ( \38799 , \38780 , \38798 );
not \U$38457 ( \38800 , \38793 );
nand \U$38458 ( \38801 , \38800 , \38781 );
nand \U$38459 ( \38802 , \38799 , \38801 );
xor \U$38460 ( \38803 , \38743 , \38802 );
xor \U$38461 ( \38804 , \38565 , \38555 );
xor \U$38462 ( \38805 , \38485 , \38508 );
xor \U$38463 ( \38806 , \38804 , \38805 );
not \U$38464 ( \38807 , \9226 );
not \U$38465 ( \38808 , \38632 );
or \U$38466 ( \38809 , \38807 , \38808 );
not \U$38467 ( \38810 , RI9872bf8_170);
not \U$38468 ( \38811 , \16996 );
or \U$38469 ( \38812 , \38810 , \38811 );
or \U$38470 ( \38813 , \23924 , RI9872bf8_170);
nand \U$38471 ( \38814 , \38812 , \38813 );
nand \U$38472 ( \38815 , \38814 , \9249 );
nand \U$38473 ( \38816 , \38809 , \38815 );
xor \U$38474 ( \38817 , \38623 , \38629 );
not \U$38475 ( \38818 , \38817 );
not \U$38476 ( \38819 , \9214 );
not \U$38477 ( \38820 , \38524 );
or \U$38478 ( \38821 , \38819 , \38820 );
and \U$38479 ( \38822 , RI9872b80_169, \19542 );
not \U$38480 ( \38823 , RI9872b80_169);
and \U$38481 ( \38824 , \38823 , \24854 );
or \U$38482 ( \38825 , \38822 , \38824 );
nand \U$38483 ( \38826 , \38825 , \9195 );
nand \U$38484 ( \38827 , \38821 , \38826 );
not \U$38485 ( \38828 , \38827 );
not \U$38486 ( \38829 , \38828 );
or \U$38487 ( \38830 , \38818 , \38829 );
or \U$38488 ( \38831 , \38828 , \38817 );
nand \U$38489 ( \38832 , \38830 , \38831 );
and \U$38490 ( \38833 , \38816 , \38832 );
and \U$38491 ( \38834 , \38817 , \38827 );
nor \U$38492 ( \38835 , \38833 , \38834 );
not \U$38493 ( \38836 , \38835 );
not \U$38494 ( \38837 , \17544 );
not \U$38495 ( \38838 , RI9873288_184);
not \U$38496 ( \38839 , \8555 );
or \U$38497 ( \38840 , \38838 , \38839 );
or \U$38498 ( \38841 , \13298 , RI9873288_184);
nand \U$38499 ( \38842 , \38840 , \38841 );
not \U$38500 ( \38843 , \38842 );
or \U$38501 ( \38844 , \38837 , \38843 );
nand \U$38502 ( \38845 , \38660 , \17528 );
nand \U$38503 ( \38846 , \38844 , \38845 );
not \U$38504 ( \38847 , \38846 );
not \U$38505 ( \38848 , \38847 );
or \U$38506 ( \38849 , \38836 , \38848 );
not \U$38507 ( \38850 , \24076 );
and \U$38508 ( \38851 , RI98734e0_189, \22524 );
not \U$38509 ( \38852 , RI98734e0_189);
and \U$38510 ( \38853 , \38852 , \8597 );
or \U$38511 ( \38854 , \38851 , \38853 );
not \U$38512 ( \38855 , \38854 );
or \U$38513 ( \38856 , \38850 , \38855 );
nand \U$38514 ( \38857 , \38670 , \20147 );
nand \U$38515 ( \38858 , \38856 , \38857 );
nand \U$38516 ( \38859 , \38849 , \38858 );
not \U$38517 ( \38860 , \38835 );
nand \U$38518 ( \38861 , \38860 , \38846 );
nand \U$38519 ( \38862 , \38859 , \38861 );
and \U$38520 ( \38863 , \38806 , \38862 );
and \U$38521 ( \38864 , \38804 , \38805 );
or \U$38522 ( \38865 , \38863 , \38864 );
and \U$38523 ( \38866 , \38803 , \38865 );
and \U$38524 ( \38867 , \38743 , \38802 );
or \U$38525 ( \38868 , \38866 , \38867 );
xor \U$38526 ( \38869 , \38578 , \38584 );
xnor \U$38527 ( \38870 , \38869 , \38678 );
xor \U$38528 ( \38871 , \38868 , \38870 );
not \U$38529 ( \38872 , \38706 );
not \U$38530 ( \38873 , \38713 );
or \U$38531 ( \38874 , \38872 , \38873 );
or \U$38532 ( \38875 , \38713 , \38706 );
nand \U$38533 ( \38876 , \38874 , \38875 );
and \U$38534 ( \38877 , \38871 , \38876 );
and \U$38535 ( \38878 , \38868 , \38870 );
or \U$38536 ( \38879 , \38877 , \38878 );
not \U$38537 ( \38880 , \38879 );
xor \U$38538 ( \38881 , \38737 , \38880 );
xor \U$38539 ( \38882 , \38681 , \38716 );
xor \U$38540 ( \38883 , \38882 , \38723 );
and \U$38541 ( \38884 , \38881 , \38883 );
and \U$38542 ( \38885 , \38737 , \38880 );
or \U$38543 ( \38886 , \38884 , \38885 );
nand \U$38544 ( \38887 , \38732 , \38886 );
not \U$38545 ( \38888 , \38887 );
xor \U$38546 ( \38889 , \38595 , \38604 );
xor \U$38547 ( \38890 , \38889 , \38615 );
xor \U$38548 ( \38891 , \38779 , \38797 );
xor \U$38549 ( \38892 , \38890 , \38891 );
not \U$38550 ( \38893 , \22618 );
not \U$38551 ( \38894 , \38748 );
or \U$38552 ( \38895 , \38893 , \38894 );
and \U$38553 ( \38896 , RI98730a8_180, \24502 );
not \U$38554 ( \38897 , RI98730a8_180);
and \U$38555 ( \38898 , \38897 , \12597 );
nor \U$38556 ( \38899 , \38896 , \38898 );
nand \U$38557 ( \38900 , \38899 , \13020 );
nand \U$38558 ( \38901 , \38895 , \38900 );
not \U$38559 ( \38902 , \38901 );
not \U$38560 ( \38903 , \8751 );
not \U$38561 ( \38904 , RI9872f40_177);
not \U$38562 ( \38905 , \25847 );
or \U$38563 ( \38906 , \38904 , \38905 );
or \U$38564 ( \38907 , \13268 , RI9872f40_177);
nand \U$38565 ( \38908 , \38906 , \38907 );
not \U$38566 ( \38909 , \38908 );
or \U$38567 ( \38910 , \38903 , \38909 );
xor \U$38568 ( \38911 , RI9872f40_177, \13281 );
nand \U$38569 ( \38912 , \38911 , \9525 );
nand \U$38570 ( \38913 , \38910 , \38912 );
not \U$38571 ( \38914 , \38913 );
not \U$38572 ( \38915 , \9937 );
not \U$38573 ( \38916 , RI9873030_179);
not \U$38574 ( \38917 , \17767 );
or \U$38575 ( \38918 , \38916 , \38917 );
nand \U$38576 ( \38919 , \13387 , \14132 );
nand \U$38577 ( \38920 , \38918 , \38919 );
not \U$38578 ( \38921 , \38920 );
or \U$38579 ( \38922 , \38915 , \38921 );
not \U$38580 ( \38923 , RI9873030_179);
not \U$38581 ( \38924 , \29808 );
or \U$38582 ( \38925 , \38923 , \38924 );
or \U$38583 ( \38926 , \18155 , RI9873030_179);
nand \U$38584 ( \38927 , \38925 , \38926 );
nand \U$38585 ( \38928 , \38927 , \9952 );
nand \U$38586 ( \38929 , \38922 , \38928 );
not \U$38587 ( \38930 , \38929 );
not \U$38588 ( \38931 , \38930 );
or \U$38589 ( \38932 , \38914 , \38931 );
or \U$38590 ( \38933 , \38930 , \38913 );
nand \U$38591 ( \38934 , \38932 , \38933 );
not \U$38592 ( \38935 , \38934 );
or \U$38593 ( \38936 , \38902 , \38935 );
nand \U$38594 ( \38937 , \38929 , \38913 );
nand \U$38595 ( \38938 , \38936 , \38937 );
not \U$38596 ( \38939 , \9272 );
not \U$38597 ( \38940 , \38759 );
or \U$38598 ( \38941 , \38939 , \38940 );
and \U$38599 ( \38942 , RI9872e50_175, \17013 );
not \U$38600 ( \38943 , RI9872e50_175);
and \U$38601 ( \38944 , \38943 , \13861 );
or \U$38602 ( \38945 , \38942 , \38944 );
nand \U$38603 ( \38946 , \38945 , \9293 );
nand \U$38604 ( \38947 , \38941 , \38946 );
not \U$38605 ( \38948 , \38947 );
and \U$38606 ( \38949 , \28663 , \8039 );
not \U$38607 ( \38950 , \9214 );
not \U$38608 ( \38951 , \38825 );
or \U$38609 ( \38952 , \38950 , \38951 );
and \U$38610 ( \38953 , RI9872b80_169, \25167 );
not \U$38611 ( \38954 , RI9872b80_169);
and \U$38612 ( \38955 , \38954 , \23952 );
or \U$38613 ( \38956 , \38953 , \38955 );
nand \U$38614 ( \38957 , \38956 , \9195 );
nand \U$38615 ( \38958 , \38952 , \38957 );
xor \U$38616 ( \38959 , \38949 , \38958 );
not \U$38617 ( \38960 , \9226 );
not \U$38618 ( \38961 , \38814 );
or \U$38619 ( \38962 , \38960 , \38961 );
not \U$38620 ( \38963 , \9244 );
not \U$38621 ( \38964 , \17702 );
or \U$38622 ( \38965 , \38963 , \38964 );
nand \U$38623 ( \38966 , \23934 , RI9872bf8_170);
nand \U$38624 ( \38967 , \38965 , \38966 );
nand \U$38625 ( \38968 , \38967 , \9249 );
nand \U$38626 ( \38969 , \38962 , \38968 );
and \U$38627 ( \38970 , \38959 , \38969 );
and \U$38628 ( \38971 , \38949 , \38958 );
nor \U$38629 ( \38972 , \38970 , \38971 );
not \U$38630 ( \38973 , \38972 );
not \U$38631 ( \38974 , \8800 );
not \U$38632 ( \38975 , \38644 );
or \U$38633 ( \38976 , \38974 , \38975 );
not \U$38634 ( \38977 , \8807 );
not \U$38635 ( \38978 , \17912 );
or \U$38636 ( \38979 , \38977 , \38978 );
nand \U$38637 ( \38980 , \17908 , RI9872d60_173);
nand \U$38638 ( \38981 , \38979 , \38980 );
nand \U$38639 ( \38982 , \38981 , \8817 );
nand \U$38640 ( \38983 , \38976 , \38982 );
not \U$38641 ( \38984 , \38983 );
or \U$38642 ( \38985 , \38973 , \38984 );
or \U$38643 ( \38986 , \38983 , \38972 );
nand \U$38644 ( \38987 , \38985 , \38986 );
not \U$38645 ( \38988 , \38987 );
or \U$38646 ( \38989 , \38948 , \38988 );
not \U$38647 ( \38990 , \38972 );
nand \U$38648 ( \38991 , \38990 , \38983 );
nand \U$38649 ( \38992 , \38989 , \38991 );
and \U$38650 ( \38993 , \38938 , \38992 );
not \U$38651 ( \38994 , \38938 );
not \U$38652 ( \38995 , \38992 );
and \U$38653 ( \38996 , \38994 , \38995 );
nor \U$38654 ( \38997 , \38993 , \38996 );
not \U$38655 ( \38998 , \38997 );
not \U$38656 ( \38999 , \9952 );
not \U$38657 ( \39000 , \38920 );
or \U$38658 ( \39001 , \38999 , \39000 );
nand \U$38659 ( \39002 , \38561 , \9937 );
nand \U$38660 ( \39003 , \39001 , \39002 );
not \U$38661 ( \39004 , \39003 );
not \U$38662 ( \39005 , \9525 );
not \U$38663 ( \39006 , \38908 );
or \U$38664 ( \39007 , \39005 , \39006 );
nand \U$38665 ( \39008 , \38483 , \11198 );
nand \U$38666 ( \39009 , \39007 , \39008 );
not \U$38667 ( \39010 , \39009 );
not \U$38668 ( \39011 , \39010 );
and \U$38669 ( \39012 , \39004 , \39011 );
and \U$38670 ( \39013 , \39003 , \39010 );
nor \U$38671 ( \39014 , \39012 , \39013 );
not \U$38672 ( \39015 , \39014 );
not \U$38673 ( \39016 , \19282 );
not \U$38674 ( \39017 , \38788 );
or \U$38675 ( \39018 , \39016 , \39017 );
and \U$38676 ( \39019 , RI98733f0_187, \8650 );
not \U$38677 ( \39020 , RI98733f0_187);
and \U$38678 ( \39021 , \39020 , \8642 );
or \U$38679 ( \39022 , \39019 , \39021 );
nand \U$38680 ( \39023 , \39022 , \17251 );
nand \U$38681 ( \39024 , \39018 , \39023 );
not \U$38682 ( \39025 , \39024 );
and \U$38683 ( \39026 , \39015 , \39025 );
and \U$38684 ( \39027 , \39024 , \39014 );
nor \U$38685 ( \39028 , \39026 , \39027 );
not \U$38686 ( \39029 , \39028 );
not \U$38687 ( \39030 , \39029 );
or \U$38688 ( \39031 , \38998 , \39030 );
not \U$38689 ( \39032 , \38995 );
nand \U$38690 ( \39033 , \39032 , \38938 );
nand \U$38691 ( \39034 , \39031 , \39033 );
and \U$38692 ( \39035 , \38892 , \39034 );
and \U$38693 ( \39036 , \38890 , \38891 );
or \U$38694 ( \39037 , \39035 , \39036 );
xor \U$38695 ( \39038 , \38743 , \38802 );
xor \U$38696 ( \39039 , \39038 , \38865 );
xor \U$38697 ( \39040 , \39037 , \39039 );
xor \U$38698 ( \39041 , \38804 , \38805 );
xor \U$38699 ( \39042 , \39041 , \38862 );
not \U$38700 ( \39043 , \39042 );
xor \U$38701 ( \39044 , \38630 , \38636 );
xor \U$38702 ( \39045 , \39044 , \38648 );
not \U$38703 ( \39046 , \17123 );
not \U$38704 ( \39047 , \38602 );
or \U$38705 ( \39048 , \39046 , \39047 );
not \U$38706 ( \39049 , \22675 );
not \U$38707 ( \39050 , \23711 );
or \U$38708 ( \39051 , \39049 , \39050 );
not \U$38709 ( \39052 , \8694 );
nand \U$38710 ( \39053 , \39052 , RI9873210_183);
nand \U$38711 ( \39054 , \39051 , \39053 );
nand \U$38712 ( \39055 , \39054 , \17243 );
nand \U$38713 ( \39056 , \39048 , \39055 );
xor \U$38714 ( \39057 , \39045 , \39056 );
not \U$38715 ( \39058 , RI9873648_192);
not \U$38716 ( \39059 , \38611 );
or \U$38717 ( \39060 , \39058 , \39059 );
not \U$38718 ( \39061 , \18239 );
not \U$38719 ( \39062 , \13358 );
or \U$38720 ( \39063 , \39061 , \39062 );
nand \U$38721 ( \39064 , \11628 , RI9873558_190);
nand \U$38722 ( \39065 , \39063 , \39064 );
nand \U$38723 ( \39066 , \39065 , \18544 );
nand \U$38724 ( \39067 , \39060 , \39066 );
xor \U$38725 ( \39068 , \39057 , \39067 );
not \U$38726 ( \39069 , \39068 );
xor \U$38727 ( \39070 , \38835 , \38858 );
xnor \U$38728 ( \39071 , \39070 , \38847 );
not \U$38729 ( \39072 , \39071 );
not \U$38730 ( \39073 , \39072 );
or \U$38731 ( \39074 , \39069 , \39073 );
not \U$38732 ( \39075 , \39068 );
nand \U$38733 ( \39076 , \39075 , \39071 );
not \U$38734 ( \39077 , \13476 );
and \U$38735 ( \39078 , \31511 , \28789 );
not \U$38736 ( \39079 , \31511 );
and \U$38737 ( \39080 , \39079 , RI9873210_183);
nor \U$38738 ( \39081 , \39078 , \39080 );
not \U$38739 ( \39082 , \39081 );
or \U$38740 ( \39083 , \39077 , \39082 );
and \U$38741 ( \39084 , RI9873210_183, \9849 );
not \U$38742 ( \39085 , RI9873210_183);
and \U$38743 ( \39086 , \39085 , \8707 );
or \U$38744 ( \39087 , \39084 , \39086 );
nand \U$38745 ( \39088 , \39087 , \33922 );
nand \U$38746 ( \39089 , \39083 , \39088 );
not \U$38747 ( \39090 , \39089 );
xor \U$38748 ( \39091 , \38969 , \38959 );
not \U$38749 ( \39092 , \8742 );
and \U$38750 ( \39093 , \18350 , \9529 );
not \U$38751 ( \39094 , \18350 );
and \U$38752 ( \39095 , \39094 , RI9872f40_177);
nor \U$38753 ( \39096 , \39093 , \39095 );
not \U$38754 ( \39097 , \39096 );
or \U$38755 ( \39098 , \39092 , \39097 );
nand \U$38756 ( \39099 , \38911 , \11198 );
nand \U$38757 ( \39100 , \39098 , \39099 );
xor \U$38758 ( \39101 , \39091 , \39100 );
not \U$38759 ( \39102 , \39101 );
or \U$38760 ( \39103 , \39090 , \39102 );
nand \U$38761 ( \39104 , \39100 , \39091 );
nand \U$38762 ( \39105 , \39103 , \39104 );
not \U$38763 ( \39106 , \39105 );
not \U$38764 ( \39107 , RI9873648_192);
not \U$38765 ( \39108 , \39065 );
or \U$38766 ( \39109 , \39107 , \39108 );
and \U$38767 ( \39110 , RI9873558_190, \9869 );
not \U$38768 ( \39111 , RI9873558_190);
and \U$38769 ( \39112 , \39111 , \12712 );
nor \U$38770 ( \39113 , \39110 , \39112 );
nand \U$38771 ( \39114 , \39113 , \18545 );
nand \U$38772 ( \39115 , \39109 , \39114 );
not \U$38773 ( \39116 , \39115 );
not \U$38774 ( \39117 , \39116 );
not \U$38775 ( \39118 , \38987 );
not \U$38776 ( \39119 , \38947 );
not \U$38777 ( \39120 , \39119 );
and \U$38778 ( \39121 , \39118 , \39120 );
and \U$38779 ( \39122 , \38987 , \39119 );
nor \U$38780 ( \39123 , \39121 , \39122 );
not \U$38781 ( \39124 , \39123 );
not \U$38782 ( \39125 , \39124 );
or \U$38783 ( \39126 , \39117 , \39125 );
nand \U$38784 ( \39127 , \39115 , \39123 );
nand \U$38785 ( \39128 , \39126 , \39127 );
not \U$38786 ( \39129 , \39128 );
or \U$38787 ( \39130 , \39106 , \39129 );
nand \U$38788 ( \39131 , \39115 , \39124 );
nand \U$38789 ( \39132 , \39130 , \39131 );
nand \U$38790 ( \39133 , \39076 , \39132 );
nand \U$38791 ( \39134 , \39074 , \39133 );
not \U$38792 ( \39135 , \39134 );
or \U$38793 ( \39136 , \39043 , \39135 );
or \U$38794 ( \39137 , \39134 , \39042 );
not \U$38795 ( \39138 , \9293 );
and \U$38796 ( \39139 , \17004 , \18862 );
not \U$38797 ( \39140 , \17004 );
and \U$38798 ( \39141 , \39140 , RI9872e50_175);
nor \U$38799 ( \39142 , \39139 , \39141 );
not \U$38800 ( \39143 , \39142 );
or \U$38801 ( \39144 , \39138 , \39143 );
nand \U$38802 ( \39145 , \38945 , \9272 );
nand \U$38803 ( \39146 , \39144 , \39145 );
not \U$38804 ( \39147 , \39146 );
and \U$38805 ( \39148 , \24450 , \9187 );
nor \U$38806 ( \39149 , \39148 , \16014 );
not \U$38807 ( \39150 , \9214 );
not \U$38808 ( \39151 , \38956 );
or \U$38809 ( \39152 , \39150 , \39151 );
xnor \U$38810 ( \39153 , \21778 , RI9872b80_169);
nand \U$38811 ( \39154 , \39153 , \9194 );
nand \U$38812 ( \39155 , \39152 , \39154 );
and \U$38813 ( \39156 , \39149 , \39155 );
not \U$38814 ( \39157 , \8800 );
not \U$38815 ( \39158 , \38981 );
or \U$38816 ( \39159 , \39157 , \39158 );
not \U$38817 ( \39160 , \8807 );
not \U$38818 ( \39161 , \25409 );
or \U$38819 ( \39162 , \39160 , \39161 );
nand \U$38820 ( \39163 , \24470 , RI9872d60_173);
nand \U$38821 ( \39164 , \39162 , \39163 );
nand \U$38822 ( \39165 , \39164 , \8817 );
nand \U$38823 ( \39166 , \39159 , \39165 );
xor \U$38824 ( \39167 , \39156 , \39166 );
not \U$38825 ( \39168 , \39167 );
or \U$38826 ( \39169 , \39147 , \39168 );
nand \U$38827 ( \39170 , \39166 , \39156 );
nand \U$38828 ( \39171 , \39169 , \39170 );
not \U$38829 ( \39172 , \17528 );
not \U$38830 ( \39173 , \38842 );
or \U$38831 ( \39174 , \39172 , \39173 );
xnor \U$38832 ( \39175 , \8723 , RI9873288_184);
nand \U$38833 ( \39176 , \39175 , \17544 );
nand \U$38834 ( \39177 , \39174 , \39176 );
xor \U$38835 ( \39178 , \39171 , \39177 );
not \U$38836 ( \39179 , \19036 );
and \U$38837 ( \39180 , \8857 , \16999 );
not \U$38838 ( \39181 , \8857 );
and \U$38839 ( \39182 , \39181 , RI98734e0_189);
nor \U$38840 ( \39183 , \39180 , \39182 );
not \U$38841 ( \39184 , \39183 );
or \U$38842 ( \39185 , \39179 , \39184 );
nand \U$38843 ( \39186 , \38854 , \19046 );
nand \U$38844 ( \39187 , \39185 , \39186 );
and \U$38845 ( \39188 , \39178 , \39187 );
and \U$38846 ( \39189 , \39171 , \39177 );
or \U$38847 ( \39190 , \39188 , \39189 );
not \U$38848 ( \39191 , \39190 );
and \U$38849 ( \39192 , \38752 , \38773 );
not \U$38850 ( \39193 , \38752 );
and \U$38851 ( \39194 , \39193 , \38774 );
or \U$38852 ( \39195 , \39192 , \39194 );
not \U$38853 ( \39196 , \39195 );
not \U$38854 ( \39197 , \17263 );
not \U$38855 ( \39198 , \39022 );
or \U$38856 ( \39199 , \39197 , \39198 );
and \U$38857 ( \39200 , RI98733f0_187, \34990 );
not \U$38858 ( \39201 , RI98733f0_187);
and \U$38859 ( \39202 , \39201 , \18308 );
or \U$38860 ( \39203 , \39200 , \39202 );
nand \U$38861 ( \39204 , \39203 , \17251 );
nand \U$38862 ( \39205 , \39199 , \39204 );
not \U$38863 ( \39206 , \39205 );
xor \U$38864 ( \39207 , \38832 , \38816 );
not \U$38865 ( \39208 , \39207 );
not \U$38866 ( \39209 , \17123 );
not \U$38867 ( \39210 , \39054 );
or \U$38868 ( \39211 , \39209 , \39210 );
nand \U$38869 ( \39212 , \39087 , \17243 );
nand \U$38870 ( \39213 , \39211 , \39212 );
not \U$38871 ( \39214 , \39213 );
not \U$38872 ( \39215 , \39214 );
or \U$38873 ( \39216 , \39208 , \39215 );
or \U$38874 ( \39217 , \39214 , \39207 );
nand \U$38875 ( \39218 , \39216 , \39217 );
not \U$38876 ( \39219 , \39218 );
or \U$38877 ( \39220 , \39206 , \39219 );
nand \U$38878 ( \39221 , \39213 , \39207 );
nand \U$38879 ( \39222 , \39220 , \39221 );
not \U$38880 ( \39223 , \39222 );
not \U$38881 ( \39224 , \39223 );
or \U$38882 ( \39225 , \39196 , \39224 );
not \U$38883 ( \39226 , \39195 );
nand \U$38884 ( \39227 , \39226 , \39222 );
nand \U$38885 ( \39228 , \39225 , \39227 );
not \U$38886 ( \39229 , \39228 );
or \U$38887 ( \39230 , \39191 , \39229 );
nand \U$38888 ( \39231 , \39222 , \39195 );
nand \U$38889 ( \39232 , \39230 , \39231 );
nand \U$38890 ( \39233 , \39137 , \39232 );
nand \U$38891 ( \39234 , \39136 , \39233 );
xor \U$38892 ( \39235 , \39040 , \39234 );
not \U$38893 ( \39236 , \39235 );
xor \U$38894 ( \39237 , \39045 , \39056 );
and \U$38895 ( \39238 , \39237 , \39067 );
and \U$38896 ( \39239 , \39045 , \39056 );
or \U$38897 ( \39240 , \39238 , \39239 );
not \U$38898 ( \39241 , \39014 );
not \U$38899 ( \39242 , \39241 );
not \U$38900 ( \39243 , \39024 );
or \U$38901 ( \39244 , \39242 , \39243 );
nand \U$38902 ( \39245 , \39003 , \39009 );
nand \U$38903 ( \39246 , \39244 , \39245 );
or \U$38904 ( \39247 , \39240 , \39246 );
xor \U$38905 ( \39248 , \38651 , \38662 );
xor \U$38906 ( \39249 , \39248 , \38672 );
and \U$38907 ( \39250 , \39247 , \39249 );
and \U$38908 ( \39251 , \39240 , \39246 );
nor \U$38909 ( \39252 , \39250 , \39251 );
xor \U$38910 ( \39253 , \38682 , \38685 );
xnor \U$38911 ( \39254 , \39253 , \38689 );
xor \U$38912 ( \39255 , \39252 , \39254 );
xor \U$38913 ( \39256 , \38619 , \38618 );
xnor \U$38914 ( \39257 , \39256 , \38675 );
xor \U$38915 ( \39258 , \39255 , \39257 );
not \U$38916 ( \39259 , \39258 );
xor \U$38917 ( \39260 , \39240 , \39246 );
xor \U$38918 ( \39261 , \39260 , \39249 );
not \U$38919 ( \39262 , \38997 );
not \U$38920 ( \39263 , \39028 );
and \U$38921 ( \39264 , \39262 , \39263 );
and \U$38922 ( \39265 , \38997 , \39028 );
nor \U$38923 ( \39266 , \39264 , \39265 );
not \U$38924 ( \39267 , \39266 );
not \U$38925 ( \39268 , \39267 );
not \U$38926 ( \39269 , \39228 );
not \U$38927 ( \39270 , \39190 );
not \U$38928 ( \39271 , \39270 );
and \U$38929 ( \39272 , \39269 , \39271 );
and \U$38930 ( \39273 , \39228 , \39270 );
nor \U$38931 ( \39274 , \39272 , \39273 );
not \U$38932 ( \39275 , \39274 );
not \U$38933 ( \39276 , \39275 );
or \U$38934 ( \39277 , \39268 , \39276 );
not \U$38935 ( \39278 , \39274 );
not \U$38936 ( \39279 , \39266 );
or \U$38937 ( \39280 , \39278 , \39279 );
not \U$38938 ( \39281 , \18615 );
not \U$38939 ( \39282 , RI9873558_190);
not \U$38940 ( \39283 , \10308 );
or \U$38941 ( \39284 , \39282 , \39283 );
or \U$38942 ( \39285 , \24842 , RI9873558_190);
nand \U$38943 ( \39286 , \39284 , \39285 );
not \U$38944 ( \39287 , \39286 );
or \U$38945 ( \39288 , \39281 , \39287 );
nand \U$38946 ( \39289 , \39113 , RI9873648_192);
nand \U$38947 ( \39290 , \39288 , \39289 );
not \U$38948 ( \39291 , \39290 );
not \U$38949 ( \39292 , \17251 );
and \U$38950 ( \39293 , \10369 , \17539 );
not \U$38951 ( \39294 , \10369 );
and \U$38952 ( \39295 , \39294 , RI98733f0_187);
nor \U$38953 ( \39296 , \39293 , \39295 );
not \U$38954 ( \39297 , \39296 );
or \U$38955 ( \39298 , \39292 , \39297 );
nand \U$38956 ( \39299 , \39203 , \17263 );
nand \U$38957 ( \39300 , \39298 , \39299 );
not \U$38958 ( \39301 , \19036 );
xnor \U$38959 ( \39302 , \8650 , RI98734e0_189);
not \U$38960 ( \39303 , \39302 );
or \U$38961 ( \39304 , \39301 , \39303 );
nand \U$38962 ( \39305 , \39183 , \19046 );
nand \U$38963 ( \39306 , \39304 , \39305 );
xor \U$38964 ( \39307 , \39300 , \39306 );
not \U$38965 ( \39308 , \39307 );
or \U$38966 ( \39309 , \39291 , \39308 );
nand \U$38967 ( \39310 , \39306 , \39300 );
nand \U$38968 ( \39311 , \39309 , \39310 );
not \U$38969 ( \39312 , \39311 );
not \U$38970 ( \39313 , \17528 );
not \U$38971 ( \39314 , \39175 );
or \U$38972 ( \39315 , \39313 , \39314 );
xor \U$38973 ( \39316 , RI9873288_184, \9750 );
nand \U$38974 ( \39317 , \39316 , \19641 );
nand \U$38975 ( \39318 , \39315 , \39317 );
buf \U$38976 ( \39319 , \39318 );
not \U$38977 ( \39320 , \39319 );
not \U$38978 ( \39321 , \12507 );
not \U$38979 ( \39322 , RI9873030_179);
not \U$38980 ( \39323 , \12773 );
or \U$38981 ( \39324 , \39322 , \39323 );
or \U$38982 ( \39325 , \12773 , RI9873030_179);
nand \U$38983 ( \39326 , \39324 , \39325 );
not \U$38984 ( \39327 , \39326 );
or \U$38985 ( \39328 , \39321 , \39327 );
nand \U$38986 ( \39329 , \38927 , \9937 );
nand \U$38987 ( \39330 , \39328 , \39329 );
not \U$38988 ( \39331 , \13020 );
and \U$38989 ( \39332 , \10064 , \13022 );
not \U$38990 ( \39333 , \10064 );
and \U$38991 ( \39334 , \39333 , RI98730a8_180);
nor \U$38992 ( \39335 , \39332 , \39334 );
not \U$38993 ( \39336 , \39335 );
or \U$38994 ( \39337 , \39331 , \39336 );
nand \U$38995 ( \39338 , \38899 , \17347 );
nand \U$38996 ( \39339 , \39337 , \39338 );
xor \U$38997 ( \39340 , \39330 , \39339 );
not \U$38998 ( \39341 , \39340 );
or \U$38999 ( \39342 , \39320 , \39341 );
nand \U$39000 ( \39343 , \39339 , \39330 );
nand \U$39001 ( \39344 , \39342 , \39343 );
xor \U$39002 ( \39345 , \38901 , \38934 );
nand \U$39003 ( \39346 , \39344 , \39345 );
not \U$39004 ( \39347 , \39346 );
not \U$39005 ( \39348 , \39347 );
and \U$39006 ( \39349 , \39312 , \39348 );
nor \U$39007 ( \39350 , \39344 , \39345 );
nor \U$39008 ( \39351 , \39349 , \39350 );
nand \U$39009 ( \39352 , \39280 , \39351 );
nand \U$39010 ( \39353 , \39277 , \39352 );
xor \U$39011 ( \39354 , \39261 , \39353 );
xor \U$39012 ( \39355 , \38890 , \38891 );
xor \U$39013 ( \39356 , \39355 , \39034 );
and \U$39014 ( \39357 , \39354 , \39356 );
and \U$39015 ( \39358 , \39261 , \39353 );
or \U$39016 ( \39359 , \39357 , \39358 );
not \U$39017 ( \39360 , \39359 );
or \U$39018 ( \39361 , \39259 , \39360 );
or \U$39019 ( \39362 , \39258 , \39359 );
nand \U$39020 ( \39363 , \39361 , \39362 );
not \U$39021 ( \39364 , \39363 );
or \U$39022 ( \39365 , \39236 , \39364 );
or \U$39023 ( \39366 , \39363 , \39235 );
nand \U$39024 ( \39367 , \39365 , \39366 );
xor \U$39025 ( \39368 , \39068 , \39072 );
xor \U$39026 ( \39369 , \39368 , \39132 );
xor \U$39027 ( \39370 , \39205 , \39218 );
xor \U$39028 ( \39371 , \39146 , \39167 );
xor \U$39029 ( \39372 , \39149 , \39155 );
not \U$39030 ( \39373 , \39372 );
not \U$39031 ( \39374 , \9226 );
not \U$39032 ( \39375 , \38967 );
or \U$39033 ( \39376 , \39374 , \39375 );
not \U$39034 ( \39377 , RI9872bf8_170);
not \U$39035 ( \39378 , \19542 );
or \U$39036 ( \39379 , \39377 , \39378 );
nand \U$39037 ( \39380 , \24854 , \9185 );
nand \U$39038 ( \39381 , \39379 , \39380 );
nand \U$39039 ( \39382 , \39381 , \9249 );
nand \U$39040 ( \39383 , \39376 , \39382 );
not \U$39041 ( \39384 , \39383 );
not \U$39042 ( \39385 , \39384 );
or \U$39043 ( \39386 , \39373 , \39385 );
or \U$39044 ( \39387 , \39384 , \39372 );
nand \U$39045 ( \39388 , \39386 , \39387 );
not \U$39046 ( \39389 , \39388 );
not \U$39047 ( \39390 , \9272 );
not \U$39048 ( \39391 , \39142 );
or \U$39049 ( \39392 , \39390 , \39391 );
not \U$39050 ( \39393 , \19394 );
xor \U$39051 ( \39394 , RI9872e50_175, \39393 );
nand \U$39052 ( \39395 , \39394 , \9293 );
nand \U$39053 ( \39396 , \39392 , \39395 );
not \U$39054 ( \39397 , \39396 );
or \U$39055 ( \39398 , \39389 , \39397 );
nand \U$39056 ( \39399 , \39372 , \39383 );
nand \U$39057 ( \39400 , \39398 , \39399 );
xor \U$39058 ( \39401 , \39371 , \39400 );
not \U$39059 ( \39402 , \39401 );
not \U$39060 ( \39403 , \30963 );
not \U$39061 ( \39404 , \39081 );
or \U$39062 ( \39405 , \39403 , \39404 );
not \U$39063 ( \39406 , \28789 );
not \U$39064 ( \39407 , \33539 );
or \U$39065 ( \39408 , \39406 , \39407 );
nand \U$39066 ( \39409 , \13066 , RI9873210_183);
nand \U$39067 ( \39410 , \39408 , \39409 );
nand \U$39068 ( \39411 , \39410 , \18957 );
nand \U$39069 ( \39412 , \39405 , \39411 );
not \U$39070 ( \39413 , \39412 );
not \U$39071 ( \39414 , \9937 );
not \U$39072 ( \39415 , \39326 );
or \U$39073 ( \39416 , \39414 , \39415 );
not \U$39074 ( \39417 , RI9873030_179);
not \U$39075 ( \39418 , \17090 );
or \U$39076 ( \39419 , \39417 , \39418 );
or \U$39077 ( \39420 , \24523 , RI9873030_179);
nand \U$39078 ( \39421 , \39419 , \39420 );
nand \U$39079 ( \39422 , \39421 , \9952 );
nand \U$39080 ( \39423 , \39416 , \39422 );
not \U$39081 ( \39424 , \39423 );
not \U$39082 ( \39425 , \39424 );
not \U$39083 ( \39426 , \22618 );
not \U$39084 ( \39427 , \39335 );
or \U$39085 ( \39428 , \39426 , \39427 );
not \U$39086 ( \39429 , RI98730a8_180);
not \U$39087 ( \39430 , \11455 );
or \U$39088 ( \39431 , \39429 , \39430 );
or \U$39089 ( \39432 , \35083 , RI98730a8_180);
nand \U$39090 ( \39433 , \39431 , \39432 );
nand \U$39091 ( \39434 , \39433 , \11350 );
nand \U$39092 ( \39435 , \39428 , \39434 );
not \U$39093 ( \39436 , \39435 );
or \U$39094 ( \39437 , \39425 , \39436 );
or \U$39095 ( \39438 , \39435 , \39424 );
nand \U$39096 ( \39439 , \39437 , \39438 );
not \U$39097 ( \39440 , \39439 );
or \U$39098 ( \39441 , \39413 , \39440 );
nand \U$39099 ( \39442 , \39435 , \39423 );
nand \U$39100 ( \39443 , \39441 , \39442 );
not \U$39101 ( \39444 , \39443 );
or \U$39102 ( \39445 , \39402 , \39444 );
nand \U$39103 ( \39446 , \39371 , \39400 );
nand \U$39104 ( \39447 , \39445 , \39446 );
xor \U$39105 ( \39448 , \39370 , \39447 );
xor \U$39106 ( \39449 , \39171 , \39177 );
xor \U$39107 ( \39450 , \39449 , \39187 );
and \U$39108 ( \39451 , \39448 , \39450 );
and \U$39109 ( \39452 , \39370 , \39447 );
or \U$39110 ( \39453 , \39451 , \39452 );
or \U$39111 ( \39454 , \39369 , \39453 );
not \U$39112 ( \39455 , \39454 );
xor \U$39113 ( \39456 , \39290 , \39307 );
not \U$39114 ( \39457 , \39456 );
not \U$39115 ( \39458 , \18615 );
and \U$39116 ( \39459 , RI9873558_190, \9881 );
not \U$39117 ( \39460 , RI9873558_190);
and \U$39118 ( \39461 , \39460 , \9882 );
nor \U$39119 ( \39462 , \39459 , \39461 );
not \U$39120 ( \39463 , \39462 );
or \U$39121 ( \39464 , \39458 , \39463 );
nand \U$39122 ( \39465 , \39286 , RI9873648_192);
nand \U$39123 ( \39466 , \39464 , \39465 );
not \U$39124 ( \39467 , \17528 );
not \U$39125 ( \39468 , \39316 );
or \U$39126 ( \39469 , \39467 , \39468 );
and \U$39127 ( \39470 , RI9873288_184, \9850 );
not \U$39128 ( \39471 , RI9873288_184);
and \U$39129 ( \39472 , \39471 , \8708 );
or \U$39130 ( \39473 , \39470 , \39472 );
nand \U$39131 ( \39474 , \39473 , \17544 );
nand \U$39132 ( \39475 , \39469 , \39474 );
nor \U$39133 ( \39476 , \39466 , \39475 );
not \U$39134 ( \39477 , \19046 );
not \U$39135 ( \39478 , \39302 );
or \U$39136 ( \39479 , \39477 , \39478 );
not \U$39137 ( \39480 , \19701 );
not \U$39138 ( \39481 , RI98734e0_189);
and \U$39139 ( \39482 , \39480 , \39481 );
and \U$39140 ( \39483 , \8842 , RI98734e0_189);
nor \U$39141 ( \39484 , \39482 , \39483 );
not \U$39142 ( \39485 , \39484 );
nand \U$39143 ( \39486 , \39485 , \19036 );
nand \U$39144 ( \39487 , \39479 , \39486 );
not \U$39145 ( \39488 , \39487 );
or \U$39146 ( \39489 , \39476 , \39488 );
nand \U$39147 ( \39490 , \39466 , \39475 );
nand \U$39148 ( \39491 , \39489 , \39490 );
xnor \U$39149 ( \39492 , \39101 , \39089 );
or \U$39150 ( \39493 , \39491 , \39492 );
nand \U$39151 ( \39494 , \39491 , \39492 );
nand \U$39152 ( \39495 , \39493 , \39494 );
not \U$39153 ( \39496 , \39495 );
or \U$39154 ( \39497 , \39457 , \39496 );
not \U$39155 ( \39498 , \39492 );
nand \U$39156 ( \39499 , \39498 , \39491 );
nand \U$39157 ( \39500 , \39497 , \39499 );
not \U$39158 ( \39501 , \39500 );
xor \U$39159 ( \39502 , \39105 , \39128 );
not \U$39160 ( \39503 , \39502 );
not \U$39161 ( \39504 , \17263 );
not \U$39162 ( \39505 , \39296 );
or \U$39163 ( \39506 , \39504 , \39505 );
and \U$39164 ( \39507 , RI98733f0_187, \20385 );
not \U$39165 ( \39508 , RI98733f0_187);
and \U$39166 ( \39509 , \39508 , \10099 );
or \U$39167 ( \39510 , \39507 , \39509 );
nand \U$39168 ( \39511 , \39510 , \17251 );
nand \U$39169 ( \39512 , \39506 , \39511 );
not \U$39170 ( \39513 , \39512 );
xor \U$39171 ( \39514 , \39396 , \39388 );
not \U$39172 ( \39515 , \39514 );
not \U$39173 ( \39516 , \8741 );
not \U$39174 ( \39517 , RI9872f40_177);
not \U$39175 ( \39518 , \38640 );
or \U$39176 ( \39519 , \39517 , \39518 );
not \U$39177 ( \39520 , \18709 );
or \U$39178 ( \39521 , \39520 , RI9872f40_177);
nand \U$39179 ( \39522 , \39519 , \39521 );
not \U$39180 ( \39523 , \39522 );
or \U$39181 ( \39524 , \39516 , \39523 );
not \U$39182 ( \39525 , \9529 );
not \U$39183 ( \39526 , \24439 );
or \U$39184 ( \39527 , \39525 , \39526 );
or \U$39185 ( \39528 , \13861 , \8732 );
nand \U$39186 ( \39529 , \39527 , \39528 );
nand \U$39187 ( \39530 , \39529 , \8751 );
nand \U$39188 ( \39531 , \39524 , \39530 );
not \U$39189 ( \39532 , \39531 );
not \U$39190 ( \39533 , \15428 );
not \U$39191 ( \39534 , \9243 );
not \U$39192 ( \39535 , \8811 );
or \U$39193 ( \39536 , \39534 , \39535 );
nand \U$39194 ( \39537 , \39536 , \24450 );
nand \U$39195 ( \39538 , \39533 , \39537 );
not \U$39196 ( \39539 , \39538 );
not \U$39197 ( \39540 , \9226 );
and \U$39198 ( \39541 , RI9872bf8_170, \21773 );
not \U$39199 ( \39542 , RI9872bf8_170);
and \U$39200 ( \39543 , \39542 , \25166 );
or \U$39201 ( \39544 , \39541 , \39543 );
not \U$39202 ( \39545 , \39544 );
or \U$39203 ( \39546 , \39540 , \39545 );
not \U$39204 ( \39547 , RI9872bf8_170);
not \U$39205 ( \39548 , \22278 );
or \U$39206 ( \39549 , \39547 , \39548 );
or \U$39207 ( \39550 , \22278 , RI9872bf8_170);
nand \U$39208 ( \39551 , \39549 , \39550 );
nand \U$39209 ( \39552 , \39551 , \9248 );
nand \U$39210 ( \39553 , \39546 , \39552 );
nand \U$39211 ( \39554 , \39539 , \39553 );
not \U$39212 ( \39555 , \39554 );
not \U$39213 ( \39556 , \9293 );
not \U$39214 ( \39557 , RI9872e50_175);
not \U$39215 ( \39558 , \31875 );
or \U$39216 ( \39559 , \39557 , \39558 );
or \U$39217 ( \39560 , \17868 , RI9872e50_175);
nand \U$39218 ( \39561 , \39559 , \39560 );
not \U$39219 ( \39562 , \39561 );
or \U$39220 ( \39563 , \39556 , \39562 );
nand \U$39221 ( \39564 , \9272 , \39394 );
nand \U$39222 ( \39565 , \39563 , \39564 );
not \U$39223 ( \39566 , \39565 );
or \U$39224 ( \39567 , \39555 , \39566 );
or \U$39225 ( \39568 , \39565 , \39554 );
nand \U$39226 ( \39569 , \39567 , \39568 );
not \U$39227 ( \39570 , \39569 );
or \U$39228 ( \39571 , \39532 , \39570 );
not \U$39229 ( \39572 , \39554 );
nand \U$39230 ( \39573 , \39572 , \39565 );
nand \U$39231 ( \39574 , \39571 , \39573 );
not \U$39232 ( \39575 , \39574 );
not \U$39233 ( \39576 , \39575 );
or \U$39234 ( \39577 , \39515 , \39576 );
not \U$39235 ( \39578 , \39514 );
nand \U$39236 ( \39579 , \39578 , \39574 );
nand \U$39237 ( \39580 , \39577 , \39579 );
not \U$39238 ( \39581 , \39580 );
or \U$39239 ( \39582 , \39513 , \39581 );
nand \U$39240 ( \39583 , \39574 , \39514 );
nand \U$39241 ( \39584 , \39582 , \39583 );
not \U$39242 ( \39585 , \39584 );
not \U$39243 ( \39586 , \11198 );
not \U$39244 ( \39587 , \39096 );
or \U$39245 ( \39588 , \39586 , \39587 );
nand \U$39246 ( \39589 , \39529 , \9525 );
nand \U$39247 ( \39590 , \39588 , \39589 );
not \U$39248 ( \39591 , \39590 );
not \U$39249 ( \39592 , \8800 );
not \U$39250 ( \39593 , \39164 );
or \U$39251 ( \39594 , \39592 , \39593 );
not \U$39252 ( \39595 , \18216 );
not \U$39253 ( \39596 , RI9872d60_173);
and \U$39254 ( \39597 , \39595 , \39596 );
and \U$39255 ( \39598 , \23924 , RI9872d60_173);
nor \U$39256 ( \39599 , \39597 , \39598 );
not \U$39257 ( \39600 , \39599 );
nand \U$39258 ( \39601 , \39600 , \8817 );
nand \U$39259 ( \39602 , \39594 , \39601 );
not \U$39260 ( \39603 , \39602 );
and \U$39261 ( \39604 , \28663 , \9214 );
not \U$39262 ( \39605 , \9226 );
not \U$39263 ( \39606 , \39381 );
or \U$39264 ( \39607 , \39605 , \39606 );
nand \U$39265 ( \39608 , \39544 , \9249 );
nand \U$39266 ( \39609 , \39607 , \39608 );
xor \U$39267 ( \39610 , \39604 , \39609 );
not \U$39268 ( \39611 , \8817 );
not \U$39269 ( \39612 , RI9872d60_173);
not \U$39270 ( \39613 , \23933 );
not \U$39271 ( \39614 , \39613 );
or \U$39272 ( \39615 , \39612 , \39614 );
or \U$39273 ( \39616 , \20490 , RI9872d60_173);
nand \U$39274 ( \39617 , \39615 , \39616 );
not \U$39275 ( \39618 , \39617 );
or \U$39276 ( \39619 , \39611 , \39618 );
not \U$39277 ( \39620 , \8800 );
or \U$39278 ( \39621 , \39599 , \39620 );
nand \U$39279 ( \39622 , \39619 , \39621 );
and \U$39280 ( \39623 , \39610 , \39622 );
and \U$39281 ( \39624 , \39604 , \39609 );
nor \U$39282 ( \39625 , \39623 , \39624 );
not \U$39283 ( \39626 , \39625 );
or \U$39284 ( \39627 , \39603 , \39626 );
or \U$39285 ( \39628 , \39625 , \39602 );
nand \U$39286 ( \39629 , \39627 , \39628 );
not \U$39287 ( \39630 , \39629 );
or \U$39288 ( \39631 , \39591 , \39630 );
not \U$39289 ( \39632 , \39625 );
nand \U$39290 ( \39633 , \39632 , \39602 );
nand \U$39291 ( \39634 , \39631 , \39633 );
xor \U$39292 ( \39635 , \39318 , \39634 );
xor \U$39293 ( \39636 , \39635 , \39340 );
not \U$39294 ( \39637 , \39636 );
or \U$39295 ( \39638 , \39585 , \39637 );
xor \U$39296 ( \39639 , \39319 , \39340 );
nand \U$39297 ( \39640 , \39639 , \39634 );
nand \U$39298 ( \39641 , \39638 , \39640 );
not \U$39299 ( \39642 , \39641 );
not \U$39300 ( \39643 , \39642 );
or \U$39301 ( \39644 , \39503 , \39643 );
not \U$39302 ( \39645 , \39502 );
nand \U$39303 ( \39646 , \39645 , \39641 );
nand \U$39304 ( \39647 , \39644 , \39646 );
not \U$39305 ( \39648 , \39647 );
or \U$39306 ( \39649 , \39501 , \39648 );
not \U$39307 ( \39650 , \39642 );
nand \U$39308 ( \39651 , \39650 , \39502 );
nand \U$39309 ( \39652 , \39649 , \39651 );
not \U$39310 ( \39653 , \39652 );
or \U$39311 ( \39654 , \39455 , \39653 );
nand \U$39312 ( \39655 , \39369 , \39453 );
nand \U$39313 ( \39656 , \39654 , \39655 );
not \U$39314 ( \39657 , \39232 );
not \U$39315 ( \39658 , \39657 );
xor \U$39316 ( \39659 , \39134 , \39042 );
not \U$39317 ( \39660 , \39659 );
or \U$39318 ( \39661 , \39658 , \39660 );
not \U$39319 ( \39662 , \39659 );
nand \U$39320 ( \39663 , \39662 , \39232 );
nand \U$39321 ( \39664 , \39661 , \39663 );
or \U$39322 ( \39665 , \39656 , \39664 );
xor \U$39323 ( \39666 , \39261 , \39353 );
xor \U$39324 ( \39667 , \39666 , \39356 );
nand \U$39325 ( \39668 , \39665 , \39667 );
nand \U$39326 ( \39669 , \39656 , \39664 );
and \U$39327 ( \39670 , \39668 , \39669 );
nor \U$39328 ( \39671 , \39367 , \39670 );
not \U$39329 ( \39672 , \39671 );
xor \U$39330 ( \39673 , \39252 , \39254 );
and \U$39331 ( \39674 , \39673 , \39257 );
and \U$39332 ( \39675 , \39252 , \39254 );
or \U$39333 ( \39676 , \39674 , \39675 );
not \U$39334 ( \39677 , \39676 );
not \U$39335 ( \39678 , \39677 );
not \U$39336 ( \39679 , \39234 );
not \U$39337 ( \39680 , \39039 );
or \U$39338 ( \39681 , \39679 , \39680 );
or \U$39339 ( \39682 , \39234 , \39039 );
nand \U$39340 ( \39683 , \39682 , \39037 );
nand \U$39341 ( \39684 , \39681 , \39683 );
not \U$39342 ( \39685 , \39684 );
not \U$39343 ( \39686 , \39685 );
or \U$39344 ( \39687 , \39678 , \39686 );
or \U$39345 ( \39688 , \39685 , \39677 );
nand \U$39346 ( \39689 , \39687 , \39688 );
not \U$39347 ( \39690 , \39689 );
xor \U$39348 ( \39691 , \38868 , \38870 );
xor \U$39349 ( \39692 , \39691 , \38876 );
not \U$39350 ( \39693 , \39692 );
or \U$39351 ( \39694 , \39690 , \39693 );
or \U$39352 ( \39695 , \39692 , \39689 );
nand \U$39353 ( \39696 , \39694 , \39695 );
not \U$39354 ( \39697 , \39235 );
not \U$39355 ( \39698 , \39697 );
not \U$39356 ( \39699 , \39363 );
or \U$39357 ( \39700 , \39698 , \39699 );
not \U$39358 ( \39701 , \39359 );
nand \U$39359 ( \39702 , \39701 , \39258 );
nand \U$39360 ( \39703 , \39700 , \39702 );
nand \U$39361 ( \39704 , \39696 , \39703 );
not \U$39362 ( \39705 , \39704 );
or \U$39363 ( \39706 , \39672 , \39705 );
not \U$39364 ( \39707 , \39696 );
not \U$39365 ( \39708 , \39703 );
nand \U$39366 ( \39709 , \39707 , \39708 );
nand \U$39367 ( \39710 , \39706 , \39709 );
not \U$39368 ( \39711 , \39710 );
xor \U$39369 ( \39712 , \38737 , \38880 );
xor \U$39370 ( \39713 , \39712 , \38883 );
not \U$39371 ( \39714 , \39689 );
not \U$39372 ( \39715 , \39692 );
not \U$39373 ( \39716 , \39715 );
or \U$39374 ( \39717 , \39714 , \39716 );
nand \U$39375 ( \39718 , \39685 , \39676 );
nand \U$39376 ( \39719 , \39717 , \39718 );
nand \U$39377 ( \39720 , \39713 , \39719 );
not \U$39378 ( \39721 , \39720 );
or \U$39379 ( \39722 , \39711 , \39721 );
or \U$39380 ( \39723 , \39713 , \39719 );
nand \U$39381 ( \39724 , \39722 , \39723 );
not \U$39382 ( \39725 , \39724 );
or \U$39383 ( \39726 , \38888 , \39725 );
or \U$39384 ( \39727 , \38732 , \38886 );
nand \U$39385 ( \39728 , \39726 , \39727 );
not \U$39386 ( \39729 , \39728 );
xor \U$39387 ( \39730 , \39370 , \39447 );
xor \U$39388 ( \39731 , \39730 , \39450 );
not \U$39389 ( \39732 , \39731 );
not \U$39390 ( \39733 , \39311 );
not \U$39391 ( \39734 , \39350 );
nand \U$39392 ( \39735 , \39734 , \39346 );
not \U$39393 ( \39736 , \39735 );
and \U$39394 ( \39737 , \39733 , \39736 );
and \U$39395 ( \39738 , \39311 , \39735 );
nor \U$39396 ( \39739 , \39737 , \39738 );
nand \U$39397 ( \39740 , \39732 , \39739 );
not \U$39398 ( \39741 , \39740 );
not \U$39399 ( \39742 , \39647 );
not \U$39400 ( \39743 , \39500 );
not \U$39401 ( \39744 , \39743 );
and \U$39402 ( \39745 , \39742 , \39744 );
and \U$39403 ( \39746 , \39647 , \39743 );
nor \U$39404 ( \39747 , \39745 , \39746 );
not \U$39405 ( \39748 , \39747 );
not \U$39406 ( \39749 , \39748 );
or \U$39407 ( \39750 , \39741 , \39749 );
not \U$39408 ( \39751 , \39739 );
nand \U$39409 ( \39752 , \39731 , \39751 );
nand \U$39410 ( \39753 , \39750 , \39752 );
not \U$39411 ( \39754 , \39753 );
not \U$39412 ( \39755 , \39754 );
and \U$39413 ( \39756 , \39351 , \39266 );
not \U$39414 ( \39757 , \39351 );
and \U$39415 ( \39758 , \39757 , \39267 );
or \U$39416 ( \39759 , \39756 , \39758 );
xnor \U$39417 ( \39760 , \39275 , \39759 );
not \U$39418 ( \39761 , \39760 );
xor \U$39419 ( \39762 , \39369 , \39453 );
not \U$39420 ( \39763 , \39762 );
not \U$39421 ( \39764 , \39652 );
and \U$39422 ( \39765 , \39763 , \39764 );
and \U$39423 ( \39766 , \39652 , \39762 );
nor \U$39424 ( \39767 , \39765 , \39766 );
not \U$39425 ( \39768 , \39767 );
or \U$39426 ( \39769 , \39761 , \39768 );
or \U$39427 ( \39770 , \39767 , \39760 );
nand \U$39428 ( \39771 , \39769 , \39770 );
not \U$39429 ( \39772 , \39771 );
not \U$39430 ( \39773 , \39772 );
or \U$39431 ( \39774 , \39755 , \39773 );
nand \U$39432 ( \39775 , \39771 , \39753 );
nand \U$39433 ( \39776 , \39774 , \39775 );
nand \U$39434 ( \39777 , \39752 , \39740 );
and \U$39435 ( \39778 , \39777 , \39748 );
not \U$39436 ( \39779 , \39777 );
and \U$39437 ( \39780 , \39779 , \39747 );
nor \U$39438 ( \39781 , \39778 , \39780 );
xor \U$39439 ( \39782 , \39495 , \39456 );
not \U$39440 ( \39783 , \39782 );
xnor \U$39441 ( \39784 , \39401 , \39443 );
and \U$39442 ( \39785 , \39439 , \39412 );
not \U$39443 ( \39786 , \39439 );
not \U$39444 ( \39787 , \39412 );
and \U$39445 ( \39788 , \39786 , \39787 );
nor \U$39446 ( \39789 , \39785 , \39788 );
not \U$39447 ( \39790 , \39789 );
xor \U$39448 ( \39791 , \39590 , \39629 );
not \U$39449 ( \39792 , \18508 );
xnor \U$39450 ( \39793 , RI9873288_184, \11371 );
not \U$39451 ( \39794 , \39793 );
or \U$39452 ( \39795 , \39792 , \39794 );
nand \U$39453 ( \39796 , \39473 , \17528 );
nand \U$39454 ( \39797 , \39795 , \39796 );
not \U$39455 ( \39798 , \39797 );
xor \U$39456 ( \39799 , \39604 , \39609 );
xor \U$39457 ( \39800 , \39799 , \39622 );
not \U$39458 ( \39801 , \39800 );
not \U$39459 ( \39802 , \17243 );
and \U$39460 ( \39803 , RI9873210_183, \38146 );
not \U$39461 ( \39804 , RI9873210_183);
and \U$39462 ( \39805 , \39804 , \33307 );
or \U$39463 ( \39806 , \39803 , \39805 );
not \U$39464 ( \39807 , \39806 );
or \U$39465 ( \39808 , \39802 , \39807 );
nand \U$39466 ( \39809 , \39410 , \17123 );
nand \U$39467 ( \39810 , \39808 , \39809 );
not \U$39468 ( \39811 , \39810 );
not \U$39469 ( \39812 , \39811 );
or \U$39470 ( \39813 , \39801 , \39812 );
or \U$39471 ( \39814 , \39811 , \39800 );
nand \U$39472 ( \39815 , \39813 , \39814 );
not \U$39473 ( \39816 , \39815 );
or \U$39474 ( \39817 , \39798 , \39816 );
nand \U$39475 ( \39818 , \39810 , \39800 );
nand \U$39476 ( \39819 , \39817 , \39818 );
xor \U$39477 ( \39820 , \39791 , \39819 );
not \U$39478 ( \39821 , \39820 );
or \U$39479 ( \39822 , \39790 , \39821 );
nand \U$39480 ( \39823 , \39819 , \39791 );
nand \U$39481 ( \39824 , \39822 , \39823 );
xnor \U$39482 ( \39825 , \39784 , \39824 );
not \U$39483 ( \39826 , \39825 );
or \U$39484 ( \39827 , \39783 , \39826 );
not \U$39485 ( \39828 , \39784 );
nand \U$39486 ( \39829 , \39828 , \39824 );
nand \U$39487 ( \39830 , \39827 , \39829 );
not \U$39488 ( \39831 , \8800 );
not \U$39489 ( \39832 , \39617 );
or \U$39490 ( \39833 , \39831 , \39832 );
not \U$39491 ( \39834 , RI9872d60_173);
not \U$39492 ( \39835 , \19542 );
or \U$39493 ( \39836 , \39834 , \39835 );
nand \U$39494 ( \39837 , \17863 , \8811 );
nand \U$39495 ( \39838 , \39836 , \39837 );
nand \U$39496 ( \39839 , \39838 , \8817 );
nand \U$39497 ( \39840 , \39833 , \39839 );
not \U$39498 ( \39841 , \39840 );
not \U$39499 ( \39842 , \39553 );
not \U$39500 ( \39843 , \39538 );
and \U$39501 ( \39844 , \39842 , \39843 );
and \U$39502 ( \39845 , \39553 , \39538 );
nor \U$39503 ( \39846 , \39844 , \39845 );
not \U$39504 ( \39847 , \39846 );
or \U$39505 ( \39848 , \39841 , \39847 );
or \U$39506 ( \39849 , \39840 , \39846 );
nand \U$39507 ( \39850 , \39848 , \39849 );
not \U$39508 ( \39851 , \39850 );
not \U$39509 ( \39852 , \8751 );
not \U$39510 ( \39853 , \39522 );
or \U$39511 ( \39854 , \39852 , \39853 );
not \U$39512 ( \39855 , RI9872f40_177);
not \U$39513 ( \39856 , \17741 );
or \U$39514 ( \39857 , \39855 , \39856 );
or \U$39515 ( \39858 , \17908 , RI9872f40_177);
nand \U$39516 ( \39859 , \39857 , \39858 );
nand \U$39517 ( \39860 , \39859 , \8741 );
nand \U$39518 ( \39861 , \39854 , \39860 );
not \U$39519 ( \39862 , \39861 );
or \U$39520 ( \39863 , \39851 , \39862 );
not \U$39521 ( \39864 , \39846 );
nand \U$39522 ( \39865 , \39864 , \39840 );
nand \U$39523 ( \39866 , \39863 , \39865 );
not \U$39524 ( \39867 , \17251 );
and \U$39525 ( \39868 , \8695 , RI98733f0_187);
not \U$39526 ( \39869 , \8695 );
and \U$39527 ( \39870 , \39869 , \17522 );
nor \U$39528 ( \39871 , \39868 , \39870 );
not \U$39529 ( \39872 , \39871 );
or \U$39530 ( \39873 , \39867 , \39872 );
nand \U$39531 ( \39874 , \39510 , \17263 );
nand \U$39532 ( \39875 , \39873 , \39874 );
xor \U$39533 ( \39876 , \39866 , \39875 );
not \U$39534 ( \39877 , RI9873648_192);
not \U$39535 ( \39878 , \39462 );
or \U$39536 ( \39879 , \39877 , \39878 );
and \U$39537 ( \39880 , RI9873558_190, \8650 );
not \U$39538 ( \39881 , RI9873558_190);
and \U$39539 ( \39882 , \39881 , \8642 );
or \U$39540 ( \39883 , \39880 , \39882 );
nand \U$39541 ( \39884 , \39883 , \18615 );
nand \U$39542 ( \39885 , \39879 , \39884 );
and \U$39543 ( \39886 , \39876 , \39885 );
and \U$39544 ( \39887 , \39866 , \39875 );
or \U$39545 ( \39888 , \39886 , \39887 );
not \U$39546 ( \39889 , \39888 );
not \U$39547 ( \39890 , RI98734e0_189);
not \U$39548 ( \39891 , \8554 );
or \U$39549 ( \39892 , \39890 , \39891 );
or \U$39550 ( \39893 , \8554 , RI98734e0_189);
nand \U$39551 ( \39894 , \39892 , \39893 );
not \U$39552 ( \39895 , \39894 );
not \U$39553 ( \39896 , \19036 );
or \U$39554 ( \39897 , \39895 , \39896 );
not \U$39555 ( \39898 , \28811 );
or \U$39556 ( \39899 , \39484 , \39898 );
nand \U$39557 ( \39900 , \39897 , \39899 );
not \U$39558 ( \39901 , \39900 );
not \U$39559 ( \39902 , \24209 );
and \U$39560 ( \39903 , \27572 , RI98730a8_180);
not \U$39561 ( \39904 , \27572 );
and \U$39562 ( \39905 , \39904 , \13022 );
nor \U$39563 ( \39906 , \39903 , \39905 );
not \U$39564 ( \39907 , \39906 );
or \U$39565 ( \39908 , \39902 , \39907 );
nand \U$39566 ( \39909 , \39433 , \12867 );
nand \U$39567 ( \39910 , \39908 , \39909 );
not \U$39568 ( \39911 , \39910 );
not \U$39569 ( \39912 , \9937 );
not \U$39570 ( \39913 , \39421 );
or \U$39571 ( \39914 , \39912 , \39913 );
not \U$39572 ( \39915 , RI9873030_179);
not \U$39573 ( \39916 , \17783 );
or \U$39574 ( \39917 , \39915 , \39916 );
or \U$39575 ( \39918 , \17783 , RI9873030_179);
nand \U$39576 ( \39919 , \39917 , \39918 );
nand \U$39577 ( \39920 , \39919 , \12507 );
nand \U$39578 ( \39921 , \39914 , \39920 );
not \U$39579 ( \39922 , \39921 );
nand \U$39580 ( \39923 , \39911 , \39922 );
not \U$39581 ( \39924 , \39923 );
or \U$39582 ( \39925 , \39901 , \39924 );
nand \U$39583 ( \39926 , \39910 , \39921 );
nand \U$39584 ( \39927 , \39925 , \39926 );
not \U$39585 ( \39928 , \39927 );
and \U$39586 ( \39929 , \39580 , \39512 );
not \U$39587 ( \39930 , \39580 );
not \U$39588 ( \39931 , \39512 );
and \U$39589 ( \39932 , \39930 , \39931 );
nor \U$39590 ( \39933 , \39929 , \39932 );
not \U$39591 ( \39934 , \39933 );
not \U$39592 ( \39935 , \39934 );
or \U$39593 ( \39936 , \39928 , \39935 );
not \U$39594 ( \39937 , \39927 );
nand \U$39595 ( \39938 , \39937 , \39933 );
nand \U$39596 ( \39939 , \39936 , \39938 );
not \U$39597 ( \39940 , \39939 );
or \U$39598 ( \39941 , \39889 , \39940 );
not \U$39599 ( \39942 , \39934 );
nand \U$39600 ( \39943 , \39942 , \39927 );
nand \U$39601 ( \39944 , \39941 , \39943 );
not \U$39602 ( \39945 , \39944 );
not \U$39603 ( \39946 , \39584 );
and \U$39604 ( \39947 , \39636 , \39946 );
not \U$39605 ( \39948 , \39636 );
and \U$39606 ( \39949 , \39948 , \39584 );
nor \U$39607 ( \39950 , \39947 , \39949 );
nand \U$39608 ( \39951 , \39945 , \39950 );
not \U$39609 ( \39952 , \39951 );
not \U$39610 ( \39953 , \9272 );
not \U$39611 ( \39954 , \39561 );
or \U$39612 ( \39955 , \39953 , \39954 );
and \U$39613 ( \39956 , \18216 , \32953 );
not \U$39614 ( \39957 , \18216 );
and \U$39615 ( \39958 , \39957 , RI9872e50_175);
nor \U$39616 ( \39959 , \39956 , \39958 );
nand \U$39617 ( \39960 , \39959 , \9293 );
nand \U$39618 ( \39961 , \39955 , \39960 );
not \U$39619 ( \39962 , \9272 );
not \U$39620 ( \39963 , \39959 );
or \U$39621 ( \39964 , \39962 , \39963 );
not \U$39622 ( \39965 , RI9872e50_175);
not \U$39623 ( \39966 , \20490 );
or \U$39624 ( \39967 , \39965 , \39966 );
or \U$39625 ( \39968 , \28657 , RI9872e50_175);
nand \U$39626 ( \39969 , \39967 , \39968 );
nand \U$39627 ( \39970 , \39969 , \9293 );
nand \U$39628 ( \39971 , \39964 , \39970 );
not \U$39629 ( \39972 , \39971 );
and \U$39630 ( \39973 , \21779 , \9226 );
not \U$39631 ( \39974 , \8800 );
not \U$39632 ( \39975 , \39838 );
or \U$39633 ( \39976 , \39974 , \39975 );
and \U$39634 ( \39977 , RI9872d60_173, \18193 );
not \U$39635 ( \39978 , RI9872d60_173);
and \U$39636 ( \39979 , \39978 , \23952 );
or \U$39637 ( \39980 , \39977 , \39979 );
nand \U$39638 ( \39981 , \39980 , \8817 );
nand \U$39639 ( \39982 , \39976 , \39981 );
xor \U$39640 ( \39983 , \39973 , \39982 );
not \U$39641 ( \39984 , \39983 );
or \U$39642 ( \39985 , \39972 , \39984 );
nand \U$39643 ( \39986 , \39982 , \39973 );
nand \U$39644 ( \39987 , \39985 , \39986 );
xor \U$39645 ( \39988 , \39961 , \39987 );
not \U$39646 ( \39989 , \39988 );
not \U$39647 ( \39990 , \17528 );
not \U$39648 ( \39991 , \39793 );
or \U$39649 ( \39992 , \39990 , \39991 );
not \U$39650 ( \39993 , \32967 );
not \U$39651 ( \39994 , \13070 );
or \U$39652 ( \39995 , \39993 , \39994 );
nand \U$39653 ( \39996 , \12597 , RI9873288_184);
nand \U$39654 ( \39997 , \39995 , \39996 );
nand \U$39655 ( \39998 , \39997 , \17544 );
nand \U$39656 ( \39999 , \39992 , \39998 );
not \U$39657 ( \40000 , \39999 );
or \U$39658 ( \40001 , \39989 , \40000 );
nand \U$39659 ( \40002 , \39987 , \39961 );
nand \U$39660 ( \40003 , \40001 , \40002 );
not \U$39661 ( \40004 , \40003 );
buf \U$39662 ( \40005 , \39569 );
buf \U$39663 ( \40006 , \39531 );
xnor \U$39664 ( \40007 , \40005 , \40006 );
not \U$39665 ( \40008 , \40007 );
not \U$39666 ( \40009 , \9937 );
not \U$39667 ( \40010 , \39919 );
or \U$39668 ( \40011 , \40009 , \40010 );
not \U$39669 ( \40012 , RI9873030_179);
not \U$39670 ( \40013 , \13860 );
or \U$39671 ( \40014 , \40012 , \40013 );
nand \U$39672 ( \40015 , \13861 , \17560 );
nand \U$39673 ( \40016 , \40014 , \40015 );
nand \U$39674 ( \40017 , \40016 , \12507 );
nand \U$39675 ( \40018 , \40011 , \40017 );
not \U$39676 ( \40019 , \40018 );
not \U$39677 ( \40020 , \11342 );
not \U$39678 ( \40021 , \39906 );
or \U$39679 ( \40022 , \40020 , \40021 );
and \U$39680 ( \40023 , RI98730a8_180, \13281 );
not \U$39681 ( \40024 , RI98730a8_180);
and \U$39682 ( \40025 , \40024 , \19595 );
nor \U$39683 ( \40026 , \40023 , \40025 );
nand \U$39684 ( \40027 , \40026 , \11350 );
nand \U$39685 ( \40028 , \40022 , \40027 );
not \U$39686 ( \40029 , \40028 );
or \U$39687 ( \40030 , \40019 , \40029 );
or \U$39688 ( \40031 , \40028 , \40018 );
not \U$39689 ( \40032 , \13483 );
not \U$39690 ( \40033 , \39806 );
or \U$39691 ( \40034 , \40032 , \40033 );
not \U$39692 ( \40035 , \28789 );
not \U$39693 ( \40036 , \12783 );
or \U$39694 ( \40037 , \40035 , \40036 );
nand \U$39695 ( \40038 , \12788 , RI9873210_183);
nand \U$39696 ( \40039 , \40037 , \40038 );
nand \U$39697 ( \40040 , \40039 , \13475 );
nand \U$39698 ( \40041 , \40034 , \40040 );
nand \U$39699 ( \40042 , \40031 , \40041 );
nand \U$39700 ( \40043 , \40030 , \40042 );
not \U$39701 ( \40044 , \40043 );
or \U$39702 ( \40045 , \40008 , \40044 );
or \U$39703 ( \40046 , \40043 , \40007 );
nand \U$39704 ( \40047 , \40045 , \40046 );
not \U$39705 ( \40048 , \40047 );
or \U$39706 ( \40049 , \40004 , \40048 );
not \U$39707 ( \40050 , \40007 );
nand \U$39708 ( \40051 , \40050 , \40043 );
nand \U$39709 ( \40052 , \40049 , \40051 );
xor \U$39710 ( \40053 , \39475 , \39487 );
xor \U$39711 ( \40054 , \40053 , \39466 );
nor \U$39712 ( \40055 , \40052 , \40054 );
not \U$39713 ( \40056 , \40055 );
not \U$39714 ( \40057 , \40056 );
and \U$39715 ( \40058 , \39926 , \39923 );
xor \U$39716 ( \40059 , \40058 , \39900 );
not \U$39717 ( \40060 , \40059 );
not \U$39718 ( \40061 , RI9873648_192);
not \U$39719 ( \40062 , \39883 );
or \U$39720 ( \40063 , \40061 , \40062 );
not \U$39721 ( \40064 , RI9873558_190);
not \U$39722 ( \40065 , \8842 );
or \U$39723 ( \40066 , \40064 , \40065 );
nand \U$39724 ( \40067 , \12848 , \18239 );
nand \U$39725 ( \40068 , \40066 , \40067 );
nand \U$39726 ( \40069 , \40068 , \18545 );
nand \U$39727 ( \40070 , \40063 , \40069 );
not \U$39728 ( \40071 , \40070 );
xor \U$39729 ( \40072 , \39850 , \39861 );
not \U$39730 ( \40073 , \40072 );
not \U$39731 ( \40074 , \28811 );
not \U$39732 ( \40075 , \39894 );
or \U$39733 ( \40076 , \40074 , \40075 );
and \U$39734 ( \40077 , RI98734e0_189, \13454 );
not \U$39735 ( \40078 , RI98734e0_189);
and \U$39736 ( \40079 , \40078 , \8722 );
or \U$39737 ( \40080 , \40077 , \40079 );
nand \U$39738 ( \40081 , \40080 , \24076 );
nand \U$39739 ( \40082 , \40076 , \40081 );
not \U$39740 ( \40083 , \40082 );
not \U$39741 ( \40084 , \40083 );
or \U$39742 ( \40085 , \40073 , \40084 );
or \U$39743 ( \40086 , \40083 , \40072 );
nand \U$39744 ( \40087 , \40085 , \40086 );
not \U$39745 ( \40088 , \40087 );
or \U$39746 ( \40089 , \40071 , \40088 );
not \U$39747 ( \40090 , \40083 );
nand \U$39748 ( \40091 , \40090 , \40072 );
nand \U$39749 ( \40092 , \40089 , \40091 );
xor \U$39750 ( \40093 , \39797 , \39815 );
xor \U$39751 ( \40094 , \40092 , \40093 );
not \U$39752 ( \40095 , \40094 );
or \U$39753 ( \40096 , \40060 , \40095 );
nand \U$39754 ( \40097 , \40093 , \40092 );
nand \U$39755 ( \40098 , \40096 , \40097 );
not \U$39756 ( \40099 , \40098 );
or \U$39757 ( \40100 , \40057 , \40099 );
nand \U$39758 ( \40101 , \40052 , \40054 );
nand \U$39759 ( \40102 , \40100 , \40101 );
not \U$39760 ( \40103 , \40102 );
or \U$39761 ( \40104 , \39952 , \40103 );
not \U$39762 ( \40105 , \39950 );
nand \U$39763 ( \40106 , \39944 , \40105 );
nand \U$39764 ( \40107 , \40104 , \40106 );
nor \U$39765 ( \40108 , \39830 , \40107 );
or \U$39766 ( \40109 , \39781 , \40108 );
nand \U$39767 ( \40110 , \39830 , \40107 );
and \U$39768 ( \40111 , \40109 , \40110 );
nand \U$39769 ( \40112 , \39776 , \40111 );
not \U$39770 ( \40113 , \39781 );
not \U$39771 ( \40114 , \40108 );
nand \U$39772 ( \40115 , \40114 , \40110 );
not \U$39773 ( \40116 , \40115 );
or \U$39774 ( \40117 , \40113 , \40116 );
or \U$39775 ( \40118 , \40115 , \39781 );
nand \U$39776 ( \40119 , \40117 , \40118 );
not \U$39777 ( \40120 , \39988 );
not \U$39778 ( \40121 , \39999 );
not \U$39779 ( \40122 , \40121 );
or \U$39780 ( \40123 , \40120 , \40122 );
or \U$39781 ( \40124 , \40121 , \39988 );
nand \U$39782 ( \40125 , \40123 , \40124 );
not \U$39783 ( \40126 , \40125 );
not \U$39784 ( \40127 , \17263 );
not \U$39785 ( \40128 , \39871 );
or \U$39786 ( \40129 , \40127 , \40128 );
and \U$39787 ( \40130 , RI98733f0_187, \12460 );
not \U$39788 ( \40131 , RI98733f0_187);
and \U$39789 ( \40132 , \40131 , \8708 );
or \U$39790 ( \40133 , \40130 , \40132 );
nand \U$39791 ( \40134 , \40133 , \17251 );
nand \U$39792 ( \40135 , \40129 , \40134 );
not \U$39793 ( \40136 , \12507 );
not \U$39794 ( \40137 , RI9873030_179);
not \U$39795 ( \40138 , \25380 );
or \U$39796 ( \40139 , \40137 , \40138 );
or \U$39797 ( \40140 , \25380 , RI9873030_179);
nand \U$39798 ( \40141 , \40139 , \40140 );
not \U$39799 ( \40142 , \40141 );
or \U$39800 ( \40143 , \40136 , \40142 );
nand \U$39801 ( \40144 , \40016 , \9937 );
nand \U$39802 ( \40145 , \40143 , \40144 );
not \U$39803 ( \40146 , \40145 );
not \U$39804 ( \40147 , \8751 );
not \U$39805 ( \40148 , \39859 );
or \U$39806 ( \40149 , \40147 , \40148 );
not \U$39807 ( \40150 , RI9872f40_177);
not \U$39808 ( \40151 , \33986 );
or \U$39809 ( \40152 , \40150 , \40151 );
or \U$39810 ( \40153 , \24470 , RI9872f40_177);
nand \U$39811 ( \40154 , \40152 , \40153 );
nand \U$39812 ( \40155 , \40154 , \8741 );
nand \U$39813 ( \40156 , \40149 , \40155 );
not \U$39814 ( \40157 , \40156 );
or \U$39815 ( \40158 , RI9872dd8_174, RI9872e50_175);
nand \U$39816 ( \40159 , \40158 , \24450 );
nand \U$39817 ( \40160 , \40159 , \14398 );
not \U$39818 ( \40161 , \40160 );
not \U$39819 ( \40162 , \8800 );
not \U$39820 ( \40163 , \39980 );
or \U$39821 ( \40164 , \40162 , \40163 );
not \U$39822 ( \40165 , \8811 );
not \U$39823 ( \40166 , \24450 );
or \U$39824 ( \40167 , \40165 , \40166 );
or \U$39825 ( \40168 , \21779 , \8807 );
nand \U$39826 ( \40169 , \40167 , \40168 );
nand \U$39827 ( \40170 , \40169 , \8816 );
nand \U$39828 ( \40171 , \40164 , \40170 );
nand \U$39829 ( \40172 , \40161 , \40171 );
not \U$39830 ( \40173 , \40172 );
and \U$39831 ( \40174 , \40157 , \40173 );
and \U$39832 ( \40175 , \40156 , \40172 );
nor \U$39833 ( \40176 , \40174 , \40175 );
not \U$39834 ( \40177 , \40176 );
not \U$39835 ( \40178 , \40177 );
or \U$39836 ( \40179 , \40146 , \40178 );
not \U$39837 ( \40180 , \40172 );
nand \U$39838 ( \40181 , \40180 , \40156 );
nand \U$39839 ( \40182 , \40179 , \40181 );
and \U$39840 ( \40183 , \40135 , \40182 );
not \U$39841 ( \40184 , \40135 );
not \U$39842 ( \40185 , \40182 );
and \U$39843 ( \40186 , \40184 , \40185 );
nor \U$39844 ( \40187 , \40183 , \40186 );
not \U$39845 ( \40188 , \40187 );
or \U$39846 ( \40189 , \40126 , \40188 );
not \U$39847 ( \40190 , \40185 );
nand \U$39848 ( \40191 , \40190 , \40135 );
nand \U$39849 ( \40192 , \40189 , \40191 );
xor \U$39850 ( \40193 , \39866 , \39875 );
xor \U$39851 ( \40194 , \40193 , \39885 );
nor \U$39852 ( \40195 , \40192 , \40194 );
not \U$39853 ( \40196 , \40195 );
not \U$39854 ( \40197 , \40196 );
not \U$39855 ( \40198 , \24209 );
not \U$39856 ( \40199 , RI98730a8_180);
not \U$39857 ( \40200 , \17783 );
or \U$39858 ( \40201 , \40199 , \40200 );
or \U$39859 ( \40202 , \24754 , RI98730a8_180);
nand \U$39860 ( \40203 , \40201 , \40202 );
not \U$39861 ( \40204 , \40203 );
or \U$39862 ( \40205 , \40198 , \40204 );
nand \U$39863 ( \40206 , \40026 , \22618 );
nand \U$39864 ( \40207 , \40205 , \40206 );
not \U$39865 ( \40208 , \17251 );
and \U$39866 ( \40209 , \9113 , \17539 );
not \U$39867 ( \40210 , \9113 );
and \U$39868 ( \40211 , \40210 , RI98733f0_187);
nor \U$39869 ( \40212 , \40209 , \40211 );
not \U$39870 ( \40213 , \40212 );
or \U$39871 ( \40214 , \40208 , \40213 );
nand \U$39872 ( \40215 , \40133 , \17263 );
nand \U$39873 ( \40216 , \40214 , \40215 );
xor \U$39874 ( \40217 , \40207 , \40216 );
not \U$39875 ( \40218 , \19035 );
and \U$39876 ( \40219 , \8697 , RI98734e0_189);
not \U$39877 ( \40220 , \8697 );
and \U$39878 ( \40221 , \40220 , \16999 );
nor \U$39879 ( \40222 , \40219 , \40221 );
not \U$39880 ( \40223 , \40222 );
or \U$39881 ( \40224 , \40218 , \40223 );
nand \U$39882 ( \40225 , \40080 , \20147 );
nand \U$39883 ( \40226 , \40224 , \40225 );
and \U$39884 ( \40227 , \40217 , \40226 );
and \U$39885 ( \40228 , \40207 , \40216 );
or \U$39886 ( \40229 , \40227 , \40228 );
not \U$39887 ( \40230 , \40229 );
xor \U$39888 ( \40231 , \39971 , \39983 );
not \U$39889 ( \40232 , \17243 );
and \U$39890 ( \40233 , RI9873210_183, \13268 );
not \U$39891 ( \40234 , RI9873210_183);
and \U$39892 ( \40235 , \40234 , \12774 );
or \U$39893 ( \40236 , \40233 , \40235 );
not \U$39894 ( \40237 , \40236 );
or \U$39895 ( \40238 , \40232 , \40237 );
nand \U$39896 ( \40239 , \40039 , \17123 );
nand \U$39897 ( \40240 , \40238 , \40239 );
xor \U$39898 ( \40241 , \40231 , \40240 );
not \U$39899 ( \40242 , \17528 );
not \U$39900 ( \40243 , \39997 );
or \U$39901 ( \40244 , \40242 , \40243 );
and \U$39902 ( \40245 , RI9873288_184, \17767 );
not \U$39903 ( \40246 , RI9873288_184);
and \U$39904 ( \40247 , \40246 , \20292 );
or \U$39905 ( \40248 , \40245 , \40247 );
nand \U$39906 ( \40249 , \40248 , \18508 );
nand \U$39907 ( \40250 , \40244 , \40249 );
and \U$39908 ( \40251 , \40241 , \40250 );
and \U$39909 ( \40252 , \40231 , \40240 );
or \U$39910 ( \40253 , \40251 , \40252 );
not \U$39911 ( \40254 , \40253 );
xor \U$39912 ( \40255 , \40018 , \40028 );
xnor \U$39913 ( \40256 , \40255 , \40041 );
not \U$39914 ( \40257 , \40256 );
or \U$39915 ( \40258 , \40254 , \40257 );
or \U$39916 ( \40259 , \40256 , \40253 );
nand \U$39917 ( \40260 , \40258 , \40259 );
not \U$39918 ( \40261 , \40260 );
or \U$39919 ( \40262 , \40230 , \40261 );
not \U$39920 ( \40263 , \40256 );
nand \U$39921 ( \40264 , \40263 , \40253 );
nand \U$39922 ( \40265 , \40262 , \40264 );
not \U$39923 ( \40266 , \40265 );
or \U$39924 ( \40267 , \40197 , \40266 );
nand \U$39925 ( \40268 , \40192 , \40194 );
nand \U$39926 ( \40269 , \40267 , \40268 );
not \U$39927 ( \40270 , \40269 );
not \U$39928 ( \40271 , \39789 );
and \U$39929 ( \40272 , \39820 , \40271 );
not \U$39930 ( \40273 , \39820 );
and \U$39931 ( \40274 , \40273 , \39789 );
nor \U$39932 ( \40275 , \40272 , \40274 );
and \U$39933 ( \40276 , \39939 , \39888 );
not \U$39934 ( \40277 , \39939 );
not \U$39935 ( \40278 , \39888 );
and \U$39936 ( \40279 , \40277 , \40278 );
nor \U$39937 ( \40280 , \40276 , \40279 );
xnor \U$39938 ( \40281 , \40275 , \40280 );
not \U$39939 ( \40282 , \40281 );
or \U$39940 ( \40283 , \40270 , \40282 );
not \U$39941 ( \40284 , \40275 );
nand \U$39942 ( \40285 , \40284 , \40280 );
nand \U$39943 ( \40286 , \40283 , \40285 );
not \U$39944 ( \40287 , \40286 );
not \U$39945 ( \40288 , \40102 );
and \U$39946 ( \40289 , \39945 , \39950 );
not \U$39947 ( \40290 , \39945 );
and \U$39948 ( \40291 , \40290 , \40105 );
nor \U$39949 ( \40292 , \40289 , \40291 );
not \U$39950 ( \40293 , \40292 );
or \U$39951 ( \40294 , \40288 , \40293 );
or \U$39952 ( \40295 , \40102 , \40292 );
nand \U$39953 ( \40296 , \40294 , \40295 );
xor \U$39954 ( \40297 , \40287 , \40296 );
xnor \U$39955 ( \40298 , \39825 , \39782 );
and \U$39956 ( \40299 , \40297 , \40298 );
and \U$39957 ( \40300 , \40287 , \40296 );
or \U$39958 ( \40301 , \40299 , \40300 );
nand \U$39959 ( \40302 , \40119 , \40301 );
not \U$39960 ( \40303 , \40302 );
xor \U$39961 ( \40304 , \40287 , \40296 );
xor \U$39962 ( \40305 , \40304 , \40298 );
not \U$39963 ( \40306 , \40055 );
nand \U$39964 ( \40307 , \40306 , \40101 );
xor \U$39965 ( \40308 , \40307 , \40098 );
not \U$39966 ( \40309 , \18615 );
and \U$39967 ( \40310 , \8555 , \18239 );
not \U$39968 ( \40311 , \8555 );
and \U$39969 ( \40312 , \40311 , RI9873558_190);
nor \U$39970 ( \40313 , \40310 , \40312 );
not \U$39971 ( \40314 , \40313 );
or \U$39972 ( \40315 , \40309 , \40314 );
nand \U$39973 ( \40316 , \40068 , RI9873648_192);
nand \U$39974 ( \40317 , \40315 , \40316 );
not \U$39975 ( \40318 , \40317 );
and \U$39976 ( \40319 , \40145 , \40176 );
not \U$39977 ( \40320 , \40145 );
and \U$39978 ( \40321 , \40320 , \40177 );
or \U$39979 ( \40322 , \40319 , \40321 );
not \U$39980 ( \40323 , \8751 );
not \U$39981 ( \40324 , \40154 );
or \U$39982 ( \40325 , \40323 , \40324 );
xor \U$39983 ( \40326 , RI9872f40_177, \19518 );
nand \U$39984 ( \40327 , \40326 , \8741 );
nand \U$39985 ( \40328 , \40325 , \40327 );
not \U$39986 ( \40329 , \40328 );
not \U$39987 ( \40330 , \9272 );
not \U$39988 ( \40331 , \39969 );
or \U$39989 ( \40332 , \40330 , \40331 );
and \U$39990 ( \40333 , RI9872e50_175, \19542 );
not \U$39991 ( \40334 , RI9872e50_175);
and \U$39992 ( \40335 , \40334 , \17862 );
or \U$39993 ( \40336 , \40333 , \40335 );
nand \U$39994 ( \40337 , \40336 , \9293 );
nand \U$39995 ( \40338 , \40332 , \40337 );
not \U$39996 ( \40339 , \40338 );
not \U$39997 ( \40340 , \40171 );
not \U$39998 ( \40341 , \40160 );
and \U$39999 ( \40342 , \40340 , \40341 );
and \U$40000 ( \40343 , \40171 , \40160 );
nor \U$40001 ( \40344 , \40342 , \40343 );
not \U$40002 ( \40345 , \40344 );
or \U$40003 ( \40346 , \40339 , \40345 );
or \U$40004 ( \40347 , \40338 , \40344 );
nand \U$40005 ( \40348 , \40346 , \40347 );
not \U$40006 ( \40349 , \40348 );
or \U$40007 ( \40350 , \40329 , \40349 );
not \U$40008 ( \40351 , \40344 );
nand \U$40009 ( \40352 , \40351 , \40338 );
nand \U$40010 ( \40353 , \40350 , \40352 );
and \U$40011 ( \40354 , \40322 , \40353 );
not \U$40012 ( \40355 , \40322 );
not \U$40013 ( \40356 , \40353 );
and \U$40014 ( \40357 , \40355 , \40356 );
nor \U$40015 ( \40358 , \40354 , \40357 );
not \U$40016 ( \40359 , \40358 );
or \U$40017 ( \40360 , \40318 , \40359 );
nand \U$40018 ( \40361 , \40322 , \40353 );
nand \U$40019 ( \40362 , \40360 , \40361 );
not \U$40020 ( \40363 , \40362 );
xor \U$40021 ( \40364 , \40125 , \40187 );
not \U$40022 ( \40365 , \40364 );
or \U$40023 ( \40366 , \40363 , \40365 );
or \U$40024 ( \40367 , \40364 , \40362 );
xor \U$40025 ( \40368 , \40087 , \40070 );
nand \U$40026 ( \40369 , \40367 , \40368 );
nand \U$40027 ( \40370 , \40366 , \40369 );
and \U$40028 ( \40371 , \40047 , \40003 );
not \U$40029 ( \40372 , \40047 );
not \U$40030 ( \40373 , \40003 );
and \U$40031 ( \40374 , \40372 , \40373 );
nor \U$40032 ( \40375 , \40371 , \40374 );
or \U$40033 ( \40376 , \40370 , \40375 );
and \U$40034 ( \40377 , \40094 , \40059 );
not \U$40035 ( \40378 , \40094 );
not \U$40036 ( \40379 , \40059 );
and \U$40037 ( \40380 , \40378 , \40379 );
nor \U$40038 ( \40381 , \40377 , \40380 );
nand \U$40039 ( \40382 , \40376 , \40381 );
nand \U$40040 ( \40383 , \40370 , \40375 );
and \U$40041 ( \40384 , \40382 , \40383 );
xor \U$40042 ( \40385 , \40308 , \40384 );
not \U$40043 ( \40386 , \40269 );
and \U$40044 ( \40387 , \40281 , \40386 );
not \U$40045 ( \40388 , \40281 );
and \U$40046 ( \40389 , \40388 , \40269 );
nor \U$40047 ( \40390 , \40387 , \40389 );
and \U$40048 ( \40391 , \40385 , \40390 );
and \U$40049 ( \40392 , \40308 , \40384 );
or \U$40050 ( \40393 , \40391 , \40392 );
nor \U$40051 ( \40394 , \40305 , \40393 );
not \U$40052 ( \40395 , \40394 );
or \U$40053 ( \40396 , \40303 , \40395 );
or \U$40054 ( \40397 , \40119 , \40301 );
nand \U$40055 ( \40398 , \40396 , \40397 );
nand \U$40056 ( \40399 , \40112 , \40398 );
not \U$40057 ( \40400 , \40399 );
or \U$40058 ( \40401 , \39776 , \40111 );
not \U$40059 ( \40402 , \40401 );
or \U$40060 ( \40403 , \40400 , \40402 );
not \U$40061 ( \40404 , \39754 );
not \U$40062 ( \40405 , \39771 );
or \U$40063 ( \40406 , \40404 , \40405 );
not \U$40064 ( \40407 , \39767 );
nand \U$40065 ( \40408 , \40407 , \39760 );
nand \U$40066 ( \40409 , \40406 , \40408 );
xor \U$40067 ( \40410 , \39664 , \39656 );
xnor \U$40068 ( \40411 , \40410 , \39667 );
nand \U$40069 ( \40412 , \40409 , \40411 );
nand \U$40070 ( \40413 , \40403 , \40412 );
not \U$40071 ( \40414 , RI9873648_192);
not \U$40072 ( \40415 , \40313 );
or \U$40073 ( \40416 , \40414 , \40415 );
not \U$40074 ( \40417 , \18239 );
not \U$40075 ( \40418 , \10099 );
or \U$40076 ( \40419 , \40417 , \40418 );
nand \U$40077 ( \40420 , \12471 , RI9873558_190);
nand \U$40078 ( \40421 , \40419 , \40420 );
nand \U$40079 ( \40422 , \40421 , \18615 );
nand \U$40080 ( \40423 , \40416 , \40422 );
not \U$40081 ( \40424 , \40423 );
and \U$40082 ( \40425 , \19383 , \8800 );
not \U$40083 ( \40426 , \40425 );
not \U$40084 ( \40427 , \9271 );
not \U$40085 ( \40428 , \40336 );
or \U$40086 ( \40429 , \40427 , \40428 );
not \U$40087 ( \40430 , \9690 );
not \U$40088 ( \40431 , \23948 );
or \U$40089 ( \40432 , \40430 , \40431 );
nand \U$40090 ( \40433 , \21773 , RI9872e50_175);
nand \U$40091 ( \40434 , \40432 , \40433 );
nand \U$40092 ( \40435 , \40434 , \9293 );
nand \U$40093 ( \40436 , \40429 , \40435 );
not \U$40094 ( \40437 , \40436 );
not \U$40095 ( \40438 , \40437 );
or \U$40096 ( \40439 , \40426 , \40438 );
not \U$40097 ( \40440 , \40436 );
or \U$40098 ( \40441 , \40440 , \40425 );
nand \U$40099 ( \40442 , \40439 , \40441 );
not \U$40100 ( \40443 , \8751 );
not \U$40101 ( \40444 , \40326 );
or \U$40102 ( \40445 , \40443 , \40444 );
and \U$40103 ( \40446 , RI9872f40_177, \20490 );
not \U$40104 ( \40447 , RI9872f40_177);
and \U$40105 ( \40448 , \40447 , \17702 );
or \U$40106 ( \40449 , \40446 , \40448 );
nand \U$40107 ( \40450 , \40449 , \8741 );
nand \U$40108 ( \40451 , \40445 , \40450 );
xor \U$40109 ( \40452 , \40442 , \40451 );
not \U$40110 ( \40453 , \13475 );
not \U$40111 ( \40454 , RI9873210_183);
not \U$40112 ( \40455 , \13624 );
or \U$40113 ( \40456 , \40454 , \40455 );
or \U$40114 ( \40457 , \29137 , RI9873210_183);
nand \U$40115 ( \40458 , \40456 , \40457 );
not \U$40116 ( \40459 , \40458 );
or \U$40117 ( \40460 , \40453 , \40459 );
xnor \U$40118 ( \40461 , RI9873210_183, \19591 );
nand \U$40119 ( \40462 , \40461 , \13483 );
nand \U$40120 ( \40463 , \40460 , \40462 );
xor \U$40121 ( \40464 , \40452 , \40463 );
not \U$40122 ( \40465 , \19641 );
not \U$40123 ( \40466 , RI9873288_184);
not \U$40124 ( \40467 , \25847 );
or \U$40125 ( \40468 , \40466 , \40467 );
or \U$40126 ( \40469 , \13268 , RI9873288_184);
nand \U$40127 ( \40470 , \40468 , \40469 );
not \U$40128 ( \40471 , \40470 );
or \U$40129 ( \40472 , \40465 , \40471 );
not \U$40130 ( \40473 , RI9873288_184);
not \U$40131 ( \40474 , \11455 );
or \U$40132 ( \40475 , \40473 , \40474 );
nand \U$40133 ( \40476 , \12787 , \22727 );
nand \U$40134 ( \40477 , \40475 , \40476 );
nand \U$40135 ( \40478 , \40477 , \17528 );
nand \U$40136 ( \40479 , \40472 , \40478 );
and \U$40137 ( \40480 , \40464 , \40479 );
and \U$40138 ( \40481 , \40452 , \40463 );
or \U$40139 ( \40482 , \40480 , \40481 );
not \U$40140 ( \40483 , \40482 );
not \U$40141 ( \40484 , \40483 );
not \U$40142 ( \40485 , \17528 );
not \U$40143 ( \40486 , \40248 );
or \U$40144 ( \40487 , \40485 , \40486 );
nand \U$40145 ( \40488 , \40477 , \19641 );
nand \U$40146 ( \40489 , \40487 , \40488 );
not \U$40147 ( \40490 , \9936 );
not \U$40148 ( \40491 , \40141 );
or \U$40149 ( \40492 , \40490 , \40491 );
not \U$40150 ( \40493 , \14132 );
not \U$40151 ( \40494 , \32208 );
or \U$40152 ( \40495 , \40493 , \40494 );
nand \U$40153 ( \40496 , \17911 , RI9873030_179);
nand \U$40154 ( \40497 , \40495 , \40496 );
nand \U$40155 ( \40498 , \40497 , \9951 );
nand \U$40156 ( \40499 , \40492 , \40498 );
not \U$40157 ( \40500 , \40499 );
not \U$40158 ( \40501 , \40451 );
not \U$40159 ( \40502 , \40442 );
or \U$40160 ( \40503 , \40501 , \40502 );
not \U$40161 ( \40504 , \40440 );
nand \U$40162 ( \40505 , \40504 , \40425 );
nand \U$40163 ( \40506 , \40503 , \40505 );
not \U$40164 ( \40507 , \40506 );
not \U$40165 ( \40508 , \40507 );
and \U$40166 ( \40509 , \40500 , \40508 );
not \U$40167 ( \40510 , \40506 );
and \U$40168 ( \40511 , \40499 , \40510 );
nor \U$40169 ( \40512 , \40509 , \40511 );
nor \U$40170 ( \40513 , \40489 , \40512 );
not \U$40171 ( \40514 , \40513 );
nand \U$40172 ( \40515 , \40512 , \40489 );
nand \U$40173 ( \40516 , \40514 , \40515 );
not \U$40174 ( \40517 , \40516 );
or \U$40175 ( \40518 , \40484 , \40517 );
not \U$40176 ( \40519 , \40482 );
or \U$40177 ( \40520 , \40516 , \40519 );
nand \U$40178 ( \40521 , \40518 , \40520 );
not \U$40179 ( \40522 , \40521 );
or \U$40180 ( \40523 , \40424 , \40522 );
nand \U$40181 ( \40524 , \40516 , \40482 );
nand \U$40182 ( \40525 , \40523 , \40524 );
not \U$40183 ( \40526 , \40512 );
not \U$40184 ( \40527 , \40526 );
not \U$40185 ( \40528 , \40489 );
or \U$40186 ( \40529 , \40527 , \40528 );
not \U$40187 ( \40530 , \40510 );
nand \U$40188 ( \40531 , \40530 , \40499 );
nand \U$40189 ( \40532 , \40529 , \40531 );
not \U$40190 ( \40533 , \17252 );
not \U$40191 ( \40534 , \17539 );
not \U$40192 ( \40535 , \13067 );
or \U$40193 ( \40536 , \40534 , \40535 );
nand \U$40194 ( \40537 , \12597 , RI98733f0_187);
nand \U$40195 ( \40538 , \40536 , \40537 );
not \U$40196 ( \40539 , \40538 );
or \U$40197 ( \40540 , \40533 , \40539 );
nand \U$40198 ( \40541 , \40212 , \17263 );
nand \U$40199 ( \40542 , \40540 , \40541 );
xor \U$40200 ( \40543 , RI98730a8_180, \13860 );
not \U$40201 ( \40544 , \40543 );
not \U$40202 ( \40545 , \11351 );
and \U$40203 ( \40546 , \40544 , \40545 );
and \U$40204 ( \40547 , \40203 , \11342 );
nor \U$40205 ( \40548 , \40546 , \40547 );
not \U$40206 ( \40549 , \40548 );
or \U$40207 ( \40550 , \40542 , \40549 );
not \U$40208 ( \40551 , \17123 );
not \U$40209 ( \40552 , \40236 );
or \U$40210 ( \40553 , \40551 , \40552 );
nand \U$40211 ( \40554 , \40461 , \17243 );
nand \U$40212 ( \40555 , \40553 , \40554 );
nand \U$40213 ( \40556 , \40550 , \40555 );
nand \U$40214 ( \40557 , \40542 , \40549 );
nand \U$40215 ( \40558 , \40556 , \40557 );
xor \U$40216 ( \40559 , \40532 , \40558 );
xor \U$40217 ( \40560 , \40231 , \40240 );
xor \U$40218 ( \40561 , \40560 , \40250 );
xor \U$40219 ( \40562 , \40559 , \40561 );
nor \U$40220 ( \40563 , \40525 , \40562 );
xor \U$40221 ( \40564 , \40548 , \40555 );
xnor \U$40222 ( \40565 , \40564 , \40542 );
not \U$40223 ( \40566 , \19046 );
not \U$40224 ( \40567 , \40222 );
or \U$40225 ( \40568 , \40566 , \40567 );
not \U$40226 ( \40569 , RI98734e0_189);
not \U$40227 ( \40570 , \12460 );
or \U$40228 ( \40571 , \40569 , \40570 );
or \U$40229 ( \40572 , \9850 , RI98734e0_189);
nand \U$40230 ( \40573 , \40571 , \40572 );
nand \U$40231 ( \40574 , \40573 , \19035 );
nand \U$40232 ( \40575 , \40568 , \40574 );
not \U$40233 ( \40576 , \40575 );
not \U$40234 ( \40577 , \40576 );
not \U$40235 ( \40578 , \40328 );
not \U$40236 ( \40579 , \40578 );
not \U$40237 ( \40580 , \40348 );
or \U$40238 ( \40581 , \40579 , \40580 );
or \U$40239 ( \40582 , \40348 , \40578 );
nand \U$40240 ( \40583 , \40581 , \40582 );
not \U$40241 ( \40584 , \40583 );
not \U$40242 ( \40585 , \11350 );
not \U$40243 ( \40586 , RI98730a8_180);
not \U$40244 ( \40587 , \20764 );
or \U$40245 ( \40588 , \40586 , \40587 );
or \U$40246 ( \40589 , \39520 , RI98730a8_180);
nand \U$40247 ( \40590 , \40588 , \40589 );
not \U$40248 ( \40591 , \40590 );
or \U$40249 ( \40592 , \40585 , \40591 );
not \U$40250 ( \40593 , \40543 );
nand \U$40251 ( \40594 , \40593 , \11342 );
nand \U$40252 ( \40595 , \40592 , \40594 );
not \U$40253 ( \40596 , \40595 );
not \U$40254 ( \40597 , \9271 );
not \U$40255 ( \40598 , \40434 );
or \U$40256 ( \40599 , \40597 , \40598 );
not \U$40257 ( \40600 , \9690 );
not \U$40258 ( \40601 , \24450 );
or \U$40259 ( \40602 , \40600 , \40601 );
or \U$40260 ( \40603 , \21779 , \32953 );
nand \U$40261 ( \40604 , \40602 , \40603 );
nand \U$40262 ( \40605 , \40604 , \9293 );
nand \U$40263 ( \40606 , \40599 , \40605 );
or \U$40264 ( \40607 , RI9872ec8_176, RI9872f40_177);
nand \U$40265 ( \40608 , \40607 , \18704 );
nand \U$40266 ( \40609 , \40608 , \10814 );
not \U$40267 ( \40610 , \40609 );
nand \U$40268 ( \40611 , \40606 , \40610 );
not \U$40269 ( \40612 , \40611 );
not \U$40270 ( \40613 , \9951 );
and \U$40271 ( \40614 , \25412 , \14132 );
not \U$40272 ( \40615 , \25412 );
and \U$40273 ( \40616 , \40615 , RI9873030_179);
nor \U$40274 ( \40617 , \40614 , \40616 );
not \U$40275 ( \40618 , \40617 );
or \U$40276 ( \40619 , \40613 , \40618 );
nand \U$40277 ( \40620 , \40497 , \9936 );
nand \U$40278 ( \40621 , \40619 , \40620 );
not \U$40279 ( \40622 , \40621 );
or \U$40280 ( \40623 , \40612 , \40622 );
or \U$40281 ( \40624 , \40621 , \40611 );
nand \U$40282 ( \40625 , \40623 , \40624 );
not \U$40283 ( \40626 , \40625 );
or \U$40284 ( \40627 , \40596 , \40626 );
not \U$40285 ( \40628 , \40611 );
nand \U$40286 ( \40629 , \40628 , \40621 );
nand \U$40287 ( \40630 , \40627 , \40629 );
not \U$40288 ( \40631 , \40630 );
not \U$40289 ( \40632 , \40631 );
or \U$40290 ( \40633 , \40584 , \40632 );
not \U$40291 ( \40634 , \40583 );
nand \U$40292 ( \40635 , \40634 , \40630 );
nand \U$40293 ( \40636 , \40633 , \40635 );
not \U$40294 ( \40637 , \40636 );
or \U$40295 ( \40638 , \40577 , \40637 );
or \U$40296 ( \40639 , \40636 , \40576 );
nand \U$40297 ( \40640 , \40638 , \40639 );
xor \U$40298 ( \40641 , \40565 , \40640 );
not \U$40299 ( \40642 , \18615 );
and \U$40300 ( \40643 , \8695 , RI9873558_190);
not \U$40301 ( \40644 , \8695 );
and \U$40302 ( \40645 , \40644 , \18239 );
nor \U$40303 ( \40646 , \40643 , \40645 );
not \U$40304 ( \40647 , \40646 );
or \U$40305 ( \40648 , \40642 , \40647 );
nand \U$40306 ( \40649 , \40421 , RI9873648_192);
nand \U$40307 ( \40650 , \40648 , \40649 );
not \U$40308 ( \40651 , \40650 );
not \U$40309 ( \40652 , \19036 );
and \U$40310 ( \40653 , RI98734e0_189, \9722 );
not \U$40311 ( \40654 , RI98734e0_189);
and \U$40312 ( \40655 , \40654 , \18344 );
or \U$40313 ( \40656 , \40653 , \40655 );
not \U$40314 ( \40657 , \40656 );
or \U$40315 ( \40658 , \40652 , \40657 );
nand \U$40316 ( \40659 , \40573 , \28811 );
nand \U$40317 ( \40660 , \40658 , \40659 );
not \U$40318 ( \40661 , \40660 );
not \U$40319 ( \40662 , \17251 );
not \U$40320 ( \40663 , RI98733f0_187);
not \U$40321 ( \40664 , \13391 );
or \U$40322 ( \40665 , \40663 , \40664 );
nand \U$40323 ( \40666 , \33307 , \17539 );
nand \U$40324 ( \40667 , \40665 , \40666 );
not \U$40325 ( \40668 , \40667 );
or \U$40326 ( \40669 , \40662 , \40668 );
nand \U$40327 ( \40670 , \40538 , \17263 );
nand \U$40328 ( \40671 , \40669 , \40670 );
not \U$40329 ( \40672 , \40671 );
not \U$40330 ( \40673 , \40672 );
or \U$40331 ( \40674 , \40661 , \40673 );
or \U$40332 ( \40675 , \40672 , \40660 );
nand \U$40333 ( \40676 , \40674 , \40675 );
not \U$40334 ( \40677 , \40676 );
or \U$40335 ( \40678 , \40651 , \40677 );
nand \U$40336 ( \40679 , \40671 , \40660 );
nand \U$40337 ( \40680 , \40678 , \40679 );
and \U$40338 ( \40681 , \40641 , \40680 );
and \U$40339 ( \40682 , \40565 , \40640 );
or \U$40340 ( \40683 , \40681 , \40682 );
not \U$40341 ( \40684 , \40683 );
or \U$40342 ( \40685 , \40563 , \40684 );
nand \U$40343 ( \40686 , \40525 , \40562 );
nand \U$40344 ( \40687 , \40685 , \40686 );
not \U$40345 ( \40688 , \40687 );
not \U$40346 ( \40689 , \40364 );
xor \U$40347 ( \40690 , \40368 , \40362 );
not \U$40348 ( \40691 , \40690 );
or \U$40349 ( \40692 , \40689 , \40691 );
or \U$40350 ( \40693 , \40364 , \40690 );
nand \U$40351 ( \40694 , \40692 , \40693 );
not \U$40352 ( \40695 , \40694 );
and \U$40353 ( \40696 , \40688 , \40695 );
and \U$40354 ( \40697 , \40687 , \40694 );
nor \U$40355 ( \40698 , \40696 , \40697 );
not \U$40356 ( \40699 , \40698 );
not \U$40357 ( \40700 , \40699 );
xor \U$40358 ( \40701 , \40532 , \40558 );
and \U$40359 ( \40702 , \40701 , \40561 );
and \U$40360 ( \40703 , \40532 , \40558 );
or \U$40361 ( \40704 , \40702 , \40703 );
xor \U$40362 ( \40705 , \40229 , \40260 );
xor \U$40363 ( \40706 , \40704 , \40705 );
not \U$40364 ( \40707 , \40706 );
not \U$40365 ( \40708 , \40575 );
not \U$40366 ( \40709 , \40636 );
or \U$40367 ( \40710 , \40708 , \40709 );
nand \U$40368 ( \40711 , \40630 , \40583 );
nand \U$40369 ( \40712 , \40710 , \40711 );
xor \U$40370 ( \40713 , \40207 , \40216 );
xor \U$40371 ( \40714 , \40713 , \40226 );
nor \U$40372 ( \40715 , \40712 , \40714 );
not \U$40373 ( \40716 , \40317 );
and \U$40374 ( \40717 , \40358 , \40716 );
not \U$40375 ( \40718 , \40358 );
and \U$40376 ( \40719 , \40718 , \40317 );
nor \U$40377 ( \40720 , \40717 , \40719 );
or \U$40378 ( \40721 , \40715 , \40720 );
nand \U$40379 ( \40722 , \40712 , \40714 );
nand \U$40380 ( \40723 , \40721 , \40722 );
not \U$40381 ( \40724 , \40723 );
not \U$40382 ( \40725 , \40724 );
and \U$40383 ( \40726 , \40707 , \40725 );
and \U$40384 ( \40727 , \40706 , \40724 );
nor \U$40385 ( \40728 , \40726 , \40727 );
not \U$40386 ( \40729 , \40728 );
not \U$40387 ( \40730 , \40729 );
or \U$40388 ( \40731 , \40700 , \40730 );
nand \U$40389 ( \40732 , \40728 , \40698 );
nand \U$40390 ( \40733 , \40731 , \40732 );
not \U$40391 ( \40734 , \40715 );
nand \U$40392 ( \40735 , \40734 , \40722 );
not \U$40393 ( \40736 , \40720 );
and \U$40394 ( \40737 , \40735 , \40736 );
not \U$40395 ( \40738 , \40735 );
and \U$40396 ( \40739 , \40738 , \40720 );
nor \U$40397 ( \40740 , \40737 , \40739 );
not \U$40398 ( \40741 , \9937 );
not \U$40399 ( \40742 , \40617 );
or \U$40400 ( \40743 , \40741 , \40742 );
and \U$40401 ( \40744 , RI9873030_179, \24867 );
not \U$40402 ( \40745 , RI9873030_179);
and \U$40403 ( \40746 , \40745 , \16995 );
or \U$40404 ( \40747 , \40744 , \40746 );
nand \U$40405 ( \40748 , \40747 , \9951 );
nand \U$40406 ( \40749 , \40743 , \40748 );
and \U$40407 ( \40750 , \18705 , \9272 );
not \U$40408 ( \40751 , \8751 );
not \U$40409 ( \40752 , \17863 );
not \U$40410 ( \40753 , RI9872f40_177);
and \U$40411 ( \40754 , \40752 , \40753 );
and \U$40412 ( \40755 , \24854 , RI9872f40_177);
nor \U$40413 ( \40756 , \40754 , \40755 );
not \U$40414 ( \40757 , \40756 );
or \U$40415 ( \40758 , \40751 , \40757 );
and \U$40416 ( \40759 , RI9872f40_177, \21773 );
not \U$40417 ( \40760 , RI9872f40_177);
and \U$40418 ( \40761 , \40760 , \23952 );
or \U$40419 ( \40762 , \40759 , \40761 );
nand \U$40420 ( \40763 , \40762 , \8741 );
nand \U$40421 ( \40764 , \40758 , \40763 );
xor \U$40422 ( \40765 , \40750 , \40764 );
not \U$40423 ( \40766 , \9936 );
not \U$40424 ( \40767 , \40747 );
or \U$40425 ( \40768 , \40766 , \40767 );
and \U$40426 ( \40769 , RI9873030_179, \27541 );
not \U$40427 ( \40770 , RI9873030_179);
and \U$40428 ( \40771 , \40770 , \17703 );
or \U$40429 ( \40772 , \40769 , \40771 );
nand \U$40430 ( \40773 , \40772 , \9951 );
nand \U$40431 ( \40774 , \40768 , \40773 );
and \U$40432 ( \40775 , \40765 , \40774 );
and \U$40433 ( \40776 , \40750 , \40764 );
nor \U$40434 ( \40777 , \40775 , \40776 );
xnor \U$40435 ( \40778 , \40749 , \40777 );
not \U$40436 ( \40779 , \40778 );
not \U$40437 ( \40780 , \17528 );
not \U$40438 ( \40781 , \40470 );
or \U$40439 ( \40782 , \40780 , \40781 );
not \U$40440 ( \40783 , RI9873288_184);
not \U$40441 ( \40784 , \24523 );
or \U$40442 ( \40785 , \40783 , \40784 );
or \U$40443 ( \40786 , \20928 , RI9873288_184);
nand \U$40444 ( \40787 , \40785 , \40786 );
nand \U$40445 ( \40788 , \40787 , \17544 );
nand \U$40446 ( \40789 , \40782 , \40788 );
not \U$40447 ( \40790 , \40789 );
or \U$40448 ( \40791 , \40779 , \40790 );
not \U$40449 ( \40792 , \40777 );
nand \U$40450 ( \40793 , \40792 , \40749 );
nand \U$40451 ( \40794 , \40791 , \40793 );
not \U$40452 ( \40795 , \40794 );
not \U$40453 ( \40796 , \40595 );
and \U$40454 ( \40797 , \40625 , \40796 );
not \U$40455 ( \40798 , \40625 );
and \U$40456 ( \40799 , \40798 , \40595 );
nor \U$40457 ( \40800 , \40797 , \40799 );
not \U$40458 ( \40801 , \40800 );
not \U$40459 ( \40802 , \40801 );
and \U$40460 ( \40803 , \40606 , \40609 );
not \U$40461 ( \40804 , \40606 );
and \U$40462 ( \40805 , \40804 , \40610 );
or \U$40463 ( \40806 , \40803 , \40805 );
not \U$40464 ( \40807 , \8751 );
not \U$40465 ( \40808 , \40449 );
or \U$40466 ( \40809 , \40807 , \40808 );
nand \U$40467 ( \40810 , \40756 , \8741 );
nand \U$40468 ( \40811 , \40809 , \40810 );
xor \U$40469 ( \40812 , \40806 , \40811 );
not \U$40470 ( \40813 , \40812 );
not \U$40471 ( \40814 , \11342 );
not \U$40472 ( \40815 , \40590 );
or \U$40473 ( \40816 , \40814 , \40815 );
and \U$40474 ( \40817 , \32208 , \13022 );
not \U$40475 ( \40818 , \32208 );
and \U$40476 ( \40819 , \40818 , RI98730a8_180);
or \U$40477 ( \40820 , \40817 , \40819 );
nand \U$40478 ( \40821 , \40820 , \11350 );
nand \U$40479 ( \40822 , \40816 , \40821 );
not \U$40480 ( \40823 , \40822 );
or \U$40481 ( \40824 , \40813 , \40823 );
nand \U$40482 ( \40825 , \40806 , \40811 );
nand \U$40483 ( \40826 , \40824 , \40825 );
not \U$40484 ( \40827 , \40826 );
not \U$40485 ( \40828 , \40827 );
or \U$40486 ( \40829 , \40802 , \40828 );
nand \U$40487 ( \40830 , \40800 , \40826 );
nand \U$40488 ( \40831 , \40829 , \40830 );
not \U$40489 ( \40832 , \40831 );
or \U$40490 ( \40833 , \40795 , \40832 );
nand \U$40491 ( \40834 , \40801 , \40826 );
nand \U$40492 ( \40835 , \40833 , \40834 );
not \U$40493 ( \40836 , \40423 );
not \U$40494 ( \40837 , \40836 );
not \U$40495 ( \40838 , \40521 );
or \U$40496 ( \40839 , \40837 , \40838 );
or \U$40497 ( \40840 , \40521 , \40836 );
nand \U$40498 ( \40841 , \40839 , \40840 );
xor \U$40499 ( \40842 , \40835 , \40841 );
not \U$40500 ( \40843 , \40458 );
not \U$40501 ( \40844 , \17123 );
or \U$40502 ( \40845 , \40843 , \40844 );
and \U$40503 ( \40846 , RI9873210_183, \13860 );
not \U$40504 ( \40847 , RI9873210_183);
and \U$40505 ( \40848 , \40847 , \17014 );
or \U$40506 ( \40849 , \40846 , \40848 );
not \U$40507 ( \40850 , \40849 );
or \U$40508 ( \40851 , \40850 , \13474 );
nand \U$40509 ( \40852 , \40845 , \40851 );
not \U$40510 ( \40853 , \17263 );
not \U$40511 ( \40854 , \40667 );
or \U$40512 ( \40855 , \40853 , \40854 );
and \U$40513 ( \40856 , \18155 , \17539 );
not \U$40514 ( \40857 , \18155 );
and \U$40515 ( \40858 , \40857 , RI98733f0_187);
nor \U$40516 ( \40859 , \40856 , \40858 );
nand \U$40517 ( \40860 , \40859 , \17251 );
nand \U$40518 ( \40861 , \40855 , \40860 );
xor \U$40519 ( \40862 , \40852 , \40861 );
not \U$40520 ( \40863 , \19035 );
not \U$40521 ( \40864 , \16999 );
not \U$40522 ( \40865 , \13067 );
or \U$40523 ( \40866 , \40864 , \40865 );
or \U$40524 ( \40867 , \13071 , \19361 );
nand \U$40525 ( \40868 , \40866 , \40867 );
not \U$40526 ( \40869 , \40868 );
or \U$40527 ( \40870 , \40863 , \40869 );
nand \U$40528 ( \40871 , \40656 , \19046 );
nand \U$40529 ( \40872 , \40870 , \40871 );
and \U$40530 ( \40873 , \40862 , \40872 );
and \U$40531 ( \40874 , \40852 , \40861 );
or \U$40532 ( \40875 , \40873 , \40874 );
not \U$40533 ( \40876 , \40875 );
xor \U$40534 ( \40877 , \40676 , \40650 );
not \U$40535 ( \40878 , \40877 );
or \U$40536 ( \40879 , \40876 , \40878 );
or \U$40537 ( \40880 , \40877 , \40875 );
not \U$40538 ( \40881 , RI9873648_192);
not \U$40539 ( \40882 , \40646 );
or \U$40540 ( \40883 , \40881 , \40882 );
and \U$40541 ( \40884 , \9849 , \18239 );
not \U$40542 ( \40885 , \9849 );
and \U$40543 ( \40886 , \40885 , RI9873558_190);
nor \U$40544 ( \40887 , \40884 , \40886 );
nand \U$40545 ( \40888 , \40887 , \18545 );
nand \U$40546 ( \40889 , \40883 , \40888 );
not \U$40547 ( \40890 , \40889 );
not \U$40548 ( \40891 , \40812 );
not \U$40549 ( \40892 , \40891 );
not \U$40550 ( \40893 , \40822 );
or \U$40551 ( \40894 , \40892 , \40893 );
or \U$40552 ( \40895 , \40822 , \40891 );
nand \U$40553 ( \40896 , \40894 , \40895 );
not \U$40554 ( \40897 , \40896 );
not \U$40555 ( \40898 , \8751 );
not \U$40556 ( \40899 , \40762 );
or \U$40557 ( \40900 , \40898 , \40899 );
and \U$40558 ( \40901 , RI9872f40_177, \18704 );
not \U$40559 ( \40902 , RI9872f40_177);
and \U$40560 ( \40903 , \40902 , \24449 );
nor \U$40561 ( \40904 , \40901 , \40903 );
nand \U$40562 ( \40905 , \40904 , \8740 );
nand \U$40563 ( \40906 , \40900 , \40905 );
not \U$40564 ( \40907 , \40906 );
or \U$40565 ( \40908 , RI9872fb8_178, RI9873030_179);
nand \U$40566 ( \40909 , \40908 , \25394 );
nand \U$40567 ( \40910 , \40909 , \8956 );
nor \U$40568 ( \40911 , \40907 , \40910 );
not \U$40569 ( \40912 , \11350 );
xnor \U$40570 ( \40913 , \24470 , RI98730a8_180);
not \U$40571 ( \40914 , \40913 );
or \U$40572 ( \40915 , \40912 , \40914 );
nand \U$40573 ( \40916 , \40820 , \11342 );
nand \U$40574 ( \40917 , \40915 , \40916 );
xor \U$40575 ( \40918 , \40911 , \40917 );
not \U$40576 ( \40919 , \20765 );
not \U$40577 ( \40920 , RI9873210_183);
and \U$40578 ( \40921 , \40919 , \40920 );
and \U$40579 ( \40922 , \13934 , RI9873210_183);
nor \U$40580 ( \40923 , \40921 , \40922 );
or \U$40581 ( \40924 , \40923 , \13474 );
nand \U$40582 ( \40925 , \40849 , \13483 );
nand \U$40583 ( \40926 , \40924 , \40925 );
and \U$40584 ( \40927 , \40918 , \40926 );
and \U$40585 ( \40928 , \40911 , \40917 );
nor \U$40586 ( \40929 , \40927 , \40928 );
not \U$40587 ( \40930 , \40929 );
or \U$40588 ( \40931 , \40897 , \40930 );
or \U$40589 ( \40932 , \40929 , \40896 );
nand \U$40590 ( \40933 , \40931 , \40932 );
not \U$40591 ( \40934 , \40933 );
or \U$40592 ( \40935 , \40890 , \40934 );
not \U$40593 ( \40936 , \40929 );
nand \U$40594 ( \40937 , \40936 , \40896 );
nand \U$40595 ( \40938 , \40935 , \40937 );
nand \U$40596 ( \40939 , \40880 , \40938 );
nand \U$40597 ( \40940 , \40879 , \40939 );
and \U$40598 ( \40941 , \40842 , \40940 );
and \U$40599 ( \40942 , \40835 , \40841 );
or \U$40600 ( \40943 , \40941 , \40942 );
not \U$40601 ( \40944 , \40943 );
xor \U$40602 ( \40945 , \40740 , \40944 );
not \U$40603 ( \40946 , \40563 );
nand \U$40604 ( \40947 , \40946 , \40686 );
and \U$40605 ( \40948 , \40947 , \40683 );
not \U$40606 ( \40949 , \40947 );
and \U$40607 ( \40950 , \40949 , \40684 );
nor \U$40608 ( \40951 , \40948 , \40950 );
and \U$40609 ( \40952 , \40945 , \40951 );
and \U$40610 ( \40953 , \40740 , \40944 );
or \U$40611 ( \40954 , \40952 , \40953 );
nand \U$40612 ( \40955 , \40733 , \40954 );
xor \U$40613 ( \40956 , \40740 , \40944 );
xor \U$40614 ( \40957 , \40956 , \40951 );
not \U$40615 ( \40958 , \18508 );
and \U$40616 ( \40959 , RI9873288_184, \22392 );
not \U$40617 ( \40960 , RI9873288_184);
and \U$40618 ( \40961 , \40960 , \38124 );
or \U$40619 ( \40962 , \40959 , \40961 );
not \U$40620 ( \40963 , \40962 );
or \U$40621 ( \40964 , \40958 , \40963 );
nand \U$40622 ( \40965 , \40787 , \17528 );
nand \U$40623 ( \40966 , \40964 , \40965 );
not \U$40624 ( \40967 , \40966 );
not \U$40625 ( \40968 , \40774 );
xor \U$40626 ( \40969 , \40765 , \40968 );
not \U$40627 ( \40970 , \40969 );
and \U$40628 ( \40971 , \40967 , \40970 );
and \U$40629 ( \40972 , \40966 , \40969 );
nor \U$40630 ( \40973 , \40971 , \40972 );
not \U$40631 ( \40974 , \40973 );
not \U$40632 ( \40975 , \18615 );
not \U$40633 ( \40976 , RI9873558_190);
not \U$40634 ( \40977 , \9114 );
or \U$40635 ( \40978 , \40976 , \40977 );
or \U$40636 ( \40979 , \11371 , RI9873558_190);
nand \U$40637 ( \40980 , \40978 , \40979 );
not \U$40638 ( \40981 , \40980 );
or \U$40639 ( \40982 , \40975 , \40981 );
nand \U$40640 ( \40983 , \40887 , RI9873648_192);
nand \U$40641 ( \40984 , \40982 , \40983 );
nand \U$40642 ( \40985 , \40974 , \40984 );
not \U$40643 ( \40986 , \40969 );
nand \U$40644 ( \40987 , \40986 , \40966 );
and \U$40645 ( \40988 , \40985 , \40987 );
not \U$40646 ( \40989 , \40988 );
not \U$40647 ( \40990 , \40989 );
xor \U$40648 ( \40991 , \40778 , \40789 );
not \U$40649 ( \40992 , \40991 );
not \U$40650 ( \40993 , \11342 );
not \U$40651 ( \40994 , \40913 );
or \U$40652 ( \40995 , \40993 , \40994 );
and \U$40653 ( \40996 , RI98730a8_180, \21553 );
not \U$40654 ( \40997 , RI98730a8_180);
and \U$40655 ( \40998 , \40997 , \19519 );
nor \U$40656 ( \40999 , \40996 , \40998 );
not \U$40657 ( \41000 , \40999 );
nand \U$40658 ( \41001 , \41000 , \11350 );
nand \U$40659 ( \41002 , \40995 , \41001 );
not \U$40660 ( \41003 , \41002 );
not \U$40661 ( \41004 , \9936 );
not \U$40662 ( \41005 , \40772 );
or \U$40663 ( \41006 , \41004 , \41005 );
not \U$40664 ( \41007 , \17560 );
not \U$40665 ( \41008 , \17863 );
or \U$40666 ( \41009 , \41007 , \41008 );
or \U$40667 ( \41010 , \24854 , \14132 );
nand \U$40668 ( \41011 , \41009 , \41010 );
nand \U$40669 ( \41012 , \41011 , \9951 );
nand \U$40670 ( \41013 , \41006 , \41012 );
not \U$40671 ( \41014 , \41013 );
not \U$40672 ( \41015 , \40906 );
not \U$40673 ( \41016 , \40910 );
and \U$40674 ( \41017 , \41015 , \41016 );
and \U$40675 ( \41018 , \40906 , \40910 );
nor \U$40676 ( \41019 , \41017 , \41018 );
not \U$40677 ( \41020 , \41019 );
or \U$40678 ( \41021 , \41014 , \41020 );
or \U$40679 ( \41022 , \41013 , \41019 );
nand \U$40680 ( \41023 , \41021 , \41022 );
not \U$40681 ( \41024 , \41023 );
or \U$40682 ( \41025 , \41003 , \41024 );
not \U$40683 ( \41026 , \41019 );
nand \U$40684 ( \41027 , \41026 , \41013 );
nand \U$40685 ( \41028 , \41025 , \41027 );
not \U$40686 ( \41029 , \17251 );
xnor \U$40687 ( \41030 , \13268 , RI98733f0_187);
not \U$40688 ( \41031 , \41030 );
or \U$40689 ( \41032 , \41029 , \41031 );
nand \U$40690 ( \41033 , \40859 , \17263 );
nand \U$40691 ( \41034 , \41032 , \41033 );
xor \U$40692 ( \41035 , \41028 , \41034 );
not \U$40693 ( \41036 , \24076 );
and \U$40694 ( \41037 , RI98734e0_189, \20292 );
not \U$40695 ( \41038 , RI98734e0_189);
and \U$40696 ( \41039 , \41038 , \17767 );
nor \U$40697 ( \41040 , \41037 , \41039 );
not \U$40698 ( \41041 , \41040 );
or \U$40699 ( \41042 , \41036 , \41041 );
nand \U$40700 ( \41043 , \40868 , \19046 );
nand \U$40701 ( \41044 , \41042 , \41043 );
and \U$40702 ( \41045 , \41035 , \41044 );
and \U$40703 ( \41046 , \41028 , \41034 );
nor \U$40704 ( \41047 , \41045 , \41046 );
not \U$40705 ( \41048 , \41047 );
or \U$40706 ( \41049 , \40992 , \41048 );
or \U$40707 ( \41050 , \41047 , \40991 );
nand \U$40708 ( \41051 , \41049 , \41050 );
not \U$40709 ( \41052 , \41051 );
or \U$40710 ( \41053 , \40990 , \41052 );
not \U$40711 ( \41054 , \41047 );
nand \U$40712 ( \41055 , \41054 , \40991 );
nand \U$40713 ( \41056 , \41053 , \41055 );
and \U$40714 ( \41057 , \40831 , \40794 );
not \U$40715 ( \41058 , \40831 );
not \U$40716 ( \41059 , \40794 );
and \U$40717 ( \41060 , \41058 , \41059 );
nor \U$40718 ( \41061 , \41057 , \41060 );
xor \U$40719 ( \41062 , \40452 , \40463 );
xor \U$40720 ( \41063 , \41062 , \40479 );
and \U$40721 ( \41064 , \41061 , \41063 );
or \U$40722 ( \41065 , \41056 , \41064 );
not \U$40723 ( \41066 , \41063 );
not \U$40724 ( \41067 , \41061 );
nand \U$40725 ( \41068 , \41066 , \41067 );
nand \U$40726 ( \41069 , \41065 , \41068 );
not \U$40727 ( \41070 , \41069 );
xor \U$40728 ( \41071 , \40565 , \40640 );
xor \U$40729 ( \41072 , \41071 , \40680 );
not \U$40730 ( \41073 , \41072 );
and \U$40731 ( \41074 , \41070 , \41073 );
not \U$40732 ( \41075 , \41070 );
and \U$40733 ( \41076 , \41075 , \41072 );
nor \U$40734 ( \41077 , \41074 , \41076 );
xor \U$40735 ( \41078 , \40835 , \40841 );
xor \U$40736 ( \41079 , \41078 , \40940 );
or \U$40737 ( \41080 , \41077 , \41079 );
or \U$40738 ( \41081 , \41070 , \41072 );
nand \U$40739 ( \41082 , \41080 , \41081 );
nand \U$40740 ( \41083 , \40957 , \41082 );
and \U$40741 ( \41084 , \40955 , \41083 );
not \U$40742 ( \41085 , \40268 );
nor \U$40743 ( \41086 , \41085 , \40195 );
not \U$40744 ( \41087 , \41086 );
not \U$40745 ( \41088 , \40265 );
or \U$40746 ( \41089 , \41087 , \41088 );
or \U$40747 ( \41090 , \40265 , \41086 );
nand \U$40748 ( \41091 , \41089 , \41090 );
not \U$40749 ( \41092 , \40723 );
not \U$40750 ( \41093 , \40706 );
or \U$40751 ( \41094 , \41092 , \41093 );
nand \U$40752 ( \41095 , \40705 , \40704 );
nand \U$40753 ( \41096 , \41094 , \41095 );
not \U$40754 ( \41097 , \41096 );
xor \U$40755 ( \41098 , \41091 , \41097 );
xor \U$40756 ( \41099 , \40375 , \40370 );
xnor \U$40757 ( \41100 , \41099 , \40381 );
xor \U$40758 ( \41101 , \41098 , \41100 );
not \U$40759 ( \41102 , \40687 );
nand \U$40760 ( \41103 , \41102 , \40694 );
not \U$40761 ( \41104 , \41103 );
not \U$40762 ( \41105 , \40729 );
or \U$40763 ( \41106 , \41104 , \41105 );
not \U$40764 ( \41107 , \40694 );
nand \U$40765 ( \41108 , \41107 , \40687 );
nand \U$40766 ( \41109 , \41106 , \41108 );
not \U$40767 ( \41110 , \41109 );
nand \U$40768 ( \41111 , \41101 , \41110 );
xor \U$40769 ( \41112 , \41091 , \41097 );
and \U$40770 ( \41113 , \41112 , \41100 );
and \U$40771 ( \41114 , \41091 , \41097 );
or \U$40772 ( \41115 , \41113 , \41114 );
xor \U$40773 ( \41116 , \40308 , \40384 );
xor \U$40774 ( \41117 , \41116 , \40390 );
nand \U$40775 ( \41118 , \41115 , \41117 );
and \U$40776 ( \41119 , \41084 , \41111 , \41118 );
not \U$40777 ( \41120 , \41056 );
not \U$40778 ( \41121 , \41068 );
nor \U$40779 ( \41122 , \41121 , \41064 );
not \U$40780 ( \41123 , \41122 );
and \U$40781 ( \41124 , \41120 , \41123 );
and \U$40782 ( \41125 , \41056 , \41122 );
nor \U$40783 ( \41126 , \41124 , \41125 );
not \U$40784 ( \41127 , \41126 );
xor \U$40785 ( \41128 , \40875 , \40938 );
xnor \U$40786 ( \41129 , \41128 , \40877 );
xor \U$40787 ( \41130 , \40926 , \40918 );
or \U$40788 ( \41131 , \40999 , \11343 );
not \U$40789 ( \41132 , \13022 );
not \U$40790 ( \41133 , \28653 );
or \U$40791 ( \41134 , \41132 , \41133 );
not \U$40792 ( \41135 , \13022 );
nand \U$40793 ( \41136 , \41135 , \27541 );
nand \U$40794 ( \41137 , \41134 , \41136 );
not \U$40795 ( \41138 , \41137 );
or \U$40796 ( \41139 , \41138 , \11351 );
nand \U$40797 ( \41140 , \41131 , \41139 );
not \U$40798 ( \41141 , \41140 );
nand \U$40799 ( \41142 , \27523 , \8751 );
not \U$40800 ( \41143 , \41142 );
not \U$40801 ( \41144 , \9936 );
not \U$40802 ( \41145 , \41011 );
or \U$40803 ( \41146 , \41144 , \41145 );
and \U$40804 ( \41147 , RI9873030_179, \18194 );
not \U$40805 ( \41148 , RI9873030_179);
and \U$40806 ( \41149 , \41148 , \28671 );
or \U$40807 ( \41150 , \41147 , \41149 );
nand \U$40808 ( \41151 , \41150 , \9951 );
nand \U$40809 ( \41152 , \41146 , \41151 );
not \U$40810 ( \41153 , \41152 );
or \U$40811 ( \41154 , \41143 , \41153 );
or \U$40812 ( \41155 , \41152 , \41142 );
nand \U$40813 ( \41156 , \41154 , \41155 );
not \U$40814 ( \41157 , \41156 );
or \U$40815 ( \41158 , \41141 , \41157 );
not \U$40816 ( \41159 , \41142 );
nand \U$40817 ( \41160 , \41159 , \41152 );
nand \U$40818 ( \41161 , \41158 , \41160 );
not \U$40819 ( \41162 , \17243 );
and \U$40820 ( \41163 , RI9873210_183, \28191 );
not \U$40821 ( \41164 , RI9873210_183);
and \U$40822 ( \41165 , \41164 , \17908 );
nor \U$40823 ( \41166 , \41163 , \41165 );
not \U$40824 ( \41167 , \41166 );
or \U$40825 ( \41168 , \41162 , \41167 );
not \U$40826 ( \41169 , \40923 );
nand \U$40827 ( \41170 , \41169 , \17123 );
nand \U$40828 ( \41171 , \41168 , \41170 );
xor \U$40829 ( \41172 , \41161 , \41171 );
not \U$40830 ( \41173 , \17528 );
not \U$40831 ( \41174 , \40962 );
or \U$40832 ( \41175 , \41173 , \41174 );
and \U$40833 ( \41176 , RI9873288_184, \17015 );
not \U$40834 ( \41177 , RI9873288_184);
and \U$40835 ( \41178 , \41177 , \17883 );
or \U$40836 ( \41179 , \41176 , \41178 );
not \U$40837 ( \41180 , \41179 );
not \U$40838 ( \41181 , \19641 );
or \U$40839 ( \41182 , \41180 , \41181 );
nand \U$40840 ( \41183 , \41175 , \41182 );
and \U$40841 ( \41184 , \41172 , \41183 );
and \U$40842 ( \41185 , \41161 , \41171 );
or \U$40843 ( \41186 , \41184 , \41185 );
xor \U$40844 ( \41187 , \41130 , \41186 );
not \U$40845 ( \41188 , \17263 );
not \U$40846 ( \41189 , \41030 );
or \U$40847 ( \41190 , \41188 , \41189 );
and \U$40848 ( \41191 , RI98733f0_187, \20928 );
not \U$40849 ( \41192 , RI98733f0_187);
and \U$40850 ( \41193 , \41192 , \13281 );
nor \U$40851 ( \41194 , \41191 , \41193 );
not \U$40852 ( \41195 , \41194 );
nand \U$40853 ( \41196 , \41195 , \17252 );
nand \U$40854 ( \41197 , \41190 , \41196 );
not \U$40855 ( \41198 , \41197 );
not \U$40856 ( \41199 , RI9873648_192);
not \U$40857 ( \41200 , \40980 );
or \U$40858 ( \41201 , \41199 , \41200 );
xor \U$40859 ( \41202 , RI9873558_190, \9138 );
nand \U$40860 ( \41203 , \41202 , \18545 );
nand \U$40861 ( \41204 , \41201 , \41203 );
not \U$40862 ( \41205 , \41204 );
or \U$40863 ( \41206 , \41198 , \41205 );
or \U$40864 ( \41207 , \41204 , \41197 );
not \U$40865 ( \41208 , \20147 );
not \U$40866 ( \41209 , \41040 );
or \U$40867 ( \41210 , \41208 , \41209 );
not \U$40868 ( \41211 , RI98734e0_189);
not \U$40869 ( \41212 , \11455 );
or \U$40870 ( \41213 , \41211 , \41212 );
or \U$40871 ( \41214 , \12784 , RI98734e0_189);
nand \U$40872 ( \41215 , \41213 , \41214 );
nand \U$40873 ( \41216 , \41215 , \19035 );
nand \U$40874 ( \41217 , \41210 , \41216 );
nand \U$40875 ( \41218 , \41207 , \41217 );
nand \U$40876 ( \41219 , \41206 , \41218 );
and \U$40877 ( \41220 , \41187 , \41219 );
and \U$40878 ( \41221 , \41130 , \41186 );
or \U$40879 ( \41222 , \41220 , \41221 );
not \U$40880 ( \41223 , \41222 );
xor \U$40881 ( \41224 , \40852 , \40861 );
xor \U$40882 ( \41225 , \41224 , \40872 );
not \U$40883 ( \41226 , \41225 );
not \U$40884 ( \41227 , \41226 );
not \U$40885 ( \41228 , \40933 );
not \U$40886 ( \41229 , \40889 );
not \U$40887 ( \41230 , \41229 );
and \U$40888 ( \41231 , \41228 , \41230 );
and \U$40889 ( \41232 , \40933 , \41229 );
nor \U$40890 ( \41233 , \41231 , \41232 );
not \U$40891 ( \41234 , \41233 );
not \U$40892 ( \41235 , \41234 );
or \U$40893 ( \41236 , \41227 , \41235 );
nand \U$40894 ( \41237 , \41233 , \41225 );
nand \U$40895 ( \41238 , \41236 , \41237 );
not \U$40896 ( \41239 , \41238 );
or \U$40897 ( \41240 , \41223 , \41239 );
nand \U$40898 ( \41241 , \41234 , \41225 );
nand \U$40899 ( \41242 , \41240 , \41241 );
and \U$40900 ( \41243 , \41129 , \41242 );
not \U$40901 ( \41244 , \41129 );
not \U$40902 ( \41245 , \41242 );
and \U$40903 ( \41246 , \41244 , \41245 );
or \U$40904 ( \41247 , \41243 , \41246 );
not \U$40905 ( \41248 , \41247 );
or \U$40906 ( \41249 , \41127 , \41248 );
or \U$40907 ( \41250 , \41247 , \41126 );
nand \U$40908 ( \41251 , \41249 , \41250 );
xor \U$40909 ( \41252 , \41023 , \41002 );
not \U$40910 ( \41253 , \19641 );
and \U$40911 ( \41254 , \18710 , \22719 );
not \U$40912 ( \41255 , \18710 );
and \U$40913 ( \41256 , \41255 , RI9873288_184);
nor \U$40914 ( \41257 , \41254 , \41256 );
not \U$40915 ( \41258 , \41257 );
or \U$40916 ( \41259 , \41253 , \41258 );
nand \U$40917 ( \41260 , \41179 , \17528 );
nand \U$40918 ( \41261 , \41259 , \41260 );
not \U$40919 ( \41262 , \41261 );
not \U$40920 ( \41263 , \13483 );
not \U$40921 ( \41264 , \41166 );
or \U$40922 ( \41265 , \41263 , \41264 );
not \U$40923 ( \41266 , RI9873210_183);
not \U$40924 ( \41267 , \17868 );
or \U$40925 ( \41268 , \41266 , \41267 );
or \U$40926 ( \41269 , \17868 , RI9873210_183);
nand \U$40927 ( \41270 , \41268 , \41269 );
nand \U$40928 ( \41271 , \41270 , \17243 );
nand \U$40929 ( \41272 , \41265 , \41271 );
not \U$40930 ( \41273 , \41272 );
nor \U$40931 ( \41274 , \18706 , \9935 );
or \U$40932 ( \41275 , \41274 , \9423 );
not \U$40933 ( \41276 , \41275 );
not \U$40934 ( \41277 , \9936 );
not \U$40935 ( \41278 , \41150 );
or \U$40936 ( \41279 , \41277 , \41278 );
or \U$40937 ( \41280 , \28663 , \9946 );
or \U$40938 ( \41281 , \24449 , RI9873030_179);
nand \U$40939 ( \41282 , \41280 , \41281 );
nand \U$40940 ( \41283 , \41282 , \9950 );
nand \U$40941 ( \41284 , \41279 , \41283 );
nand \U$40942 ( \41285 , \41276 , \41284 );
not \U$40943 ( \41286 , \41285 );
and \U$40944 ( \41287 , \41273 , \41286 );
and \U$40945 ( \41288 , \41272 , \41285 );
nor \U$40946 ( \41289 , \41287 , \41288 );
not \U$40947 ( \41290 , \41289 );
not \U$40948 ( \41291 , \41290 );
or \U$40949 ( \41292 , \41262 , \41291 );
not \U$40950 ( \41293 , \41285 );
nand \U$40951 ( \41294 , \41293 , \41272 );
nand \U$40952 ( \41295 , \41292 , \41294 );
or \U$40953 ( \41296 , \41252 , \41295 );
not \U$40954 ( \41297 , \41296 );
not \U$40955 ( \41298 , \24076 );
not \U$40956 ( \41299 , RI98734e0_189);
not \U$40957 ( \41300 , \13268 );
or \U$40958 ( \41301 , \41299 , \41300 );
or \U$40959 ( \41302 , \12773 , RI98734e0_189);
nand \U$40960 ( \41303 , \41301 , \41302 );
not \U$40961 ( \41304 , \41303 );
or \U$40962 ( \41305 , \41298 , \41304 );
nand \U$40963 ( \41306 , \41215 , \28811 );
nand \U$40964 ( \41307 , \41305 , \41306 );
not \U$40965 ( \41308 , \41307 );
not \U$40966 ( \41309 , \41140 );
and \U$40967 ( \41310 , \41156 , \41309 );
not \U$40968 ( \41311 , \41156 );
and \U$40969 ( \41312 , \41311 , \41140 );
nor \U$40970 ( \41313 , \41310 , \41312 );
not \U$40971 ( \41314 , \41313 );
and \U$40972 ( \41315 , \41308 , \41314 );
and \U$40973 ( \41316 , \41307 , \41313 );
nor \U$40974 ( \41317 , \41315 , \41316 );
or \U$40975 ( \41318 , \41194 , \17620 );
xor \U$40976 ( \41319 , \18350 , RI98733f0_187);
or \U$40977 ( \41320 , \41319 , \30886 );
nand \U$40978 ( \41321 , \41318 , \41320 );
not \U$40979 ( \41322 , \41321 );
or \U$40980 ( \41323 , \41317 , \41322 );
not \U$40981 ( \41324 , \41313 );
nand \U$40982 ( \41325 , \41324 , \41307 );
nand \U$40983 ( \41326 , \41323 , \41325 );
not \U$40984 ( \41327 , \41326 );
or \U$40985 ( \41328 , \41297 , \41327 );
nand \U$40986 ( \41329 , \41295 , \41252 );
nand \U$40987 ( \41330 , \41328 , \41329 );
not \U$40988 ( \41331 , \41044 );
and \U$40989 ( \41332 , \41035 , \41331 );
not \U$40990 ( \41333 , \41035 );
and \U$40991 ( \41334 , \41333 , \41044 );
nor \U$40992 ( \41335 , \41332 , \41334 );
not \U$40993 ( \41336 , \40973 );
not \U$40994 ( \41337 , \40984 );
and \U$40995 ( \41338 , \41336 , \41337 );
and \U$40996 ( \41339 , \40973 , \40984 );
nor \U$40997 ( \41340 , \41338 , \41339 );
nand \U$40998 ( \41341 , \41335 , \41340 );
and \U$40999 ( \41342 , \41330 , \41341 );
nor \U$41000 ( \41343 , \41335 , \41340 );
nor \U$41001 ( \41344 , \41342 , \41343 );
not \U$41002 ( \41345 , \41051 );
not \U$41003 ( \41346 , \40988 );
and \U$41004 ( \41347 , \41345 , \41346 );
and \U$41005 ( \41348 , \41051 , \40988 );
nor \U$41006 ( \41349 , \41347 , \41348 );
xor \U$41007 ( \41350 , \41344 , \41349 );
not \U$41008 ( \41351 , \41222 );
and \U$41009 ( \41352 , \41238 , \41351 );
not \U$41010 ( \41353 , \41238 );
and \U$41011 ( \41354 , \41353 , \41222 );
nor \U$41012 ( \41355 , \41352 , \41354 );
and \U$41013 ( \41356 , \41350 , \41355 );
and \U$41014 ( \41357 , \41344 , \41349 );
or \U$41015 ( \41358 , \41356 , \41357 );
or \U$41016 ( \41359 , \41251 , \41358 );
not \U$41017 ( \41360 , \41359 );
xor \U$41018 ( \41361 , \41340 , \41335 );
not \U$41019 ( \41362 , \41361 );
not \U$41020 ( \41363 , \41330 );
and \U$41021 ( \41364 , \41362 , \41363 );
and \U$41022 ( \41365 , \41361 , \41330 );
nor \U$41023 ( \41366 , \41364 , \41365 );
not \U$41024 ( \41367 , \41366 );
xor \U$41025 ( \41368 , \41130 , \41186 );
xor \U$41026 ( \41369 , \41368 , \41219 );
not \U$41027 ( \41370 , \41369 );
not \U$41028 ( \41371 , \41370 );
xor \U$41029 ( \41372 , \41197 , \41204 );
xnor \U$41030 ( \41373 , \41372 , \41217 );
not \U$41031 ( \41374 , \41373 );
xor \U$41032 ( \41375 , \41161 , \41171 );
xor \U$41033 ( \41376 , \41375 , \41183 );
not \U$41034 ( \41377 , \41376 );
not \U$41035 ( \41378 , \41261 );
not \U$41036 ( \41379 , \41289 );
or \U$41037 ( \41380 , \41378 , \41379 );
or \U$41038 ( \41381 , \41289 , \41261 );
nand \U$41039 ( \41382 , \41380 , \41381 );
not \U$41040 ( \41383 , \41382 );
not \U$41041 ( \41384 , RI9873648_192);
not \U$41042 ( \41385 , \41202 );
or \U$41043 ( \41386 , \41384 , \41385 );
and \U$41044 ( \41387 , RI9873558_190, \37813 );
not \U$41045 ( \41388 , RI9873558_190);
not \U$41046 ( \41389 , \10064 );
and \U$41047 ( \41390 , \41388 , \41389 );
or \U$41048 ( \41391 , \41387 , \41390 );
nand \U$41049 ( \41392 , \41391 , \18544 );
nand \U$41050 ( \41393 , \41386 , \41392 );
not \U$41051 ( \41394 , \13483 );
not \U$41052 ( \41395 , \41270 );
or \U$41053 ( \41396 , \41394 , \41395 );
and \U$41054 ( \41397 , RI9873210_183, \16996 );
not \U$41055 ( \41398 , RI9873210_183);
and \U$41056 ( \41399 , \41398 , \36515 );
or \U$41057 ( \41400 , \41397 , \41399 );
nand \U$41058 ( \41401 , \41400 , \17243 );
nand \U$41059 ( \41402 , \41396 , \41401 );
not \U$41060 ( \41403 , \41402 );
not \U$41061 ( \41404 , \11342 );
not \U$41062 ( \41405 , \41137 );
or \U$41063 ( \41406 , \41404 , \41405 );
not \U$41064 ( \41407 , \13022 );
not \U$41065 ( \41408 , \35530 );
or \U$41066 ( \41409 , \41407 , \41408 );
or \U$41067 ( \41410 , \24854 , \13022 );
nand \U$41068 ( \41411 , \41409 , \41410 );
nand \U$41069 ( \41412 , \41411 , \11350 );
nand \U$41070 ( \41413 , \41406 , \41412 );
not \U$41071 ( \41414 , \41413 );
not \U$41072 ( \41415 , \41284 );
not \U$41073 ( \41416 , \41275 );
and \U$41074 ( \41417 , \41415 , \41416 );
and \U$41075 ( \41418 , \41284 , \41275 );
nor \U$41076 ( \41419 , \41417 , \41418 );
not \U$41077 ( \41420 , \41419 );
or \U$41078 ( \41421 , \41414 , \41420 );
or \U$41079 ( \41422 , \41413 , \41419 );
nand \U$41080 ( \41423 , \41421 , \41422 );
not \U$41081 ( \41424 , \41423 );
or \U$41082 ( \41425 , \41403 , \41424 );
not \U$41083 ( \41426 , \41419 );
nand \U$41084 ( \41427 , \41426 , \41413 );
nand \U$41085 ( \41428 , \41425 , \41427 );
xor \U$41086 ( \41429 , \41393 , \41428 );
not \U$41087 ( \41430 , \41429 );
or \U$41088 ( \41431 , \41383 , \41430 );
nand \U$41089 ( \41432 , \41393 , \41428 );
nand \U$41090 ( \41433 , \41431 , \41432 );
not \U$41091 ( \41434 , \41433 );
not \U$41092 ( \41435 , \41434 );
or \U$41093 ( \41436 , \41377 , \41435 );
or \U$41094 ( \41437 , \41434 , \41376 );
nand \U$41095 ( \41438 , \41436 , \41437 );
not \U$41096 ( \41439 , \41438 );
or \U$41097 ( \41440 , \41374 , \41439 );
not \U$41098 ( \41441 , \41376 );
nand \U$41099 ( \41442 , \41441 , \41434 );
nand \U$41100 ( \41443 , \41440 , \41442 );
not \U$41101 ( \41444 , \41443 );
not \U$41102 ( \41445 , \41444 );
or \U$41103 ( \41446 , \41371 , \41445 );
nand \U$41104 ( \41447 , \41443 , \41369 );
nand \U$41105 ( \41448 , \41446 , \41447 );
not \U$41106 ( \41449 , \41448 );
or \U$41107 ( \41450 , \41367 , \41449 );
or \U$41108 ( \41451 , \41448 , \41366 );
nand \U$41109 ( \41452 , \41450 , \41451 );
nand \U$41110 ( \41453 , \41296 , \41329 );
xor \U$41111 ( \41454 , \41326 , \41453 );
and \U$41112 ( \41455 , \41303 , \28811 );
not \U$41113 ( \41456 , \19035 );
and \U$41114 ( \41457 , RI98734e0_189, \24523 );
not \U$41115 ( \41458 , RI98734e0_189);
and \U$41116 ( \41459 , \41458 , \13281 );
nor \U$41117 ( \41460 , \41457 , \41459 );
nor \U$41118 ( \41461 , \41456 , \41460 );
nor \U$41119 ( \41462 , \41455 , \41461 );
not \U$41120 ( \41463 , \41462 );
not \U$41121 ( \41464 , \41463 );
not \U$41122 ( \41465 , \17243 );
not \U$41123 ( \41466 , \22675 );
not \U$41124 ( \41467 , \28653 );
or \U$41125 ( \41468 , \41466 , \41467 );
nand \U$41126 ( \41469 , \39613 , RI9873210_183);
nand \U$41127 ( \41470 , \41468 , \41469 );
not \U$41128 ( \41471 , \41470 );
or \U$41129 ( \41472 , \41465 , \41471 );
nand \U$41130 ( \41473 , \41400 , \13483 );
nand \U$41131 ( \41474 , \41472 , \41473 );
not \U$41132 ( \41475 , \41474 );
nand \U$41133 ( \41476 , \28663 , \9936 );
not \U$41134 ( \41477 , \41476 );
not \U$41135 ( \41478 , \11342 );
not \U$41136 ( \41479 , \41411 );
or \U$41137 ( \41480 , \41478 , \41479 );
and \U$41138 ( \41481 , RI98730a8_180, \23953 );
not \U$41139 ( \41482 , RI98730a8_180);
and \U$41140 ( \41483 , \41482 , \23948 );
or \U$41141 ( \41484 , \41481 , \41483 );
nand \U$41142 ( \41485 , \41484 , \11350 );
nand \U$41143 ( \41486 , \41480 , \41485 );
not \U$41144 ( \41487 , \41486 );
or \U$41145 ( \41488 , \41477 , \41487 );
or \U$41146 ( \41489 , \41486 , \41476 );
nand \U$41147 ( \41490 , \41488 , \41489 );
not \U$41148 ( \41491 , \41490 );
or \U$41149 ( \41492 , \41475 , \41491 );
not \U$41150 ( \41493 , \41476 );
nand \U$41151 ( \41494 , \41493 , \41486 );
nand \U$41152 ( \41495 , \41492 , \41494 );
not \U$41153 ( \41496 , \41495 );
not \U$41154 ( \41497 , \17528 );
not \U$41155 ( \41498 , \41257 );
or \U$41156 ( \41499 , \41497 , \41498 );
and \U$41157 ( \41500 , \17741 , \17538 );
not \U$41158 ( \41501 , \17741 );
and \U$41159 ( \41502 , \41501 , RI9873288_184);
nor \U$41160 ( \41503 , \41500 , \41502 );
nand \U$41161 ( \41504 , \41503 , \17543 );
nand \U$41162 ( \41505 , \41499 , \41504 );
not \U$41163 ( \41506 , \41505 );
not \U$41164 ( \41507 , \41506 );
or \U$41165 ( \41508 , \41496 , \41507 );
not \U$41166 ( \41509 , \41495 );
nand \U$41167 ( \41510 , \41509 , \41505 );
nand \U$41168 ( \41511 , \41508 , \41510 );
not \U$41169 ( \41512 , \41511 );
or \U$41170 ( \41513 , \41464 , \41512 );
nand \U$41171 ( \41514 , \41495 , \41505 );
nand \U$41172 ( \41515 , \41513 , \41514 );
and \U$41173 ( \41516 , \41317 , \41322 );
not \U$41174 ( \41517 , \41317 );
and \U$41175 ( \41518 , \41517 , \41321 );
nor \U$41176 ( \41519 , \41516 , \41518 );
xor \U$41177 ( \41520 , \41515 , \41519 );
or \U$41178 ( \41521 , \41319 , \17620 );
xor \U$41179 ( \41522 , \35645 , RI98733f0_187);
not \U$41180 ( \41523 , \41522 );
or \U$41181 ( \41524 , \41523 , \30886 );
nand \U$41182 ( \41525 , \41521 , \41524 );
not \U$41183 ( \41526 , \41525 );
xor \U$41184 ( \41527 , \41423 , \41402 );
not \U$41185 ( \41528 , RI9873648_192);
not \U$41186 ( \41529 , \41391 );
or \U$41187 ( \41530 , \41528 , \41529 );
and \U$41188 ( \41531 , RI9873558_190, \13601 );
not \U$41189 ( \41532 , RI9873558_190);
and \U$41190 ( \41533 , \41532 , \12788 );
nor \U$41191 ( \41534 , \41531 , \41533 );
nand \U$41192 ( \41535 , \41534 , \18544 );
nand \U$41193 ( \41536 , \41530 , \41535 );
not \U$41194 ( \41537 , \41536 );
and \U$41195 ( \41538 , \41527 , \41537 );
not \U$41196 ( \41539 , \41527 );
and \U$41197 ( \41540 , \41539 , \41536 );
or \U$41198 ( \41541 , \41538 , \41540 );
not \U$41199 ( \41542 , \41541 );
or \U$41200 ( \41543 , \41526 , \41542 );
nand \U$41201 ( \41544 , \41536 , \41527 );
nand \U$41202 ( \41545 , \41543 , \41544 );
and \U$41203 ( \41546 , \41520 , \41545 );
and \U$41204 ( \41547 , \41515 , \41519 );
nor \U$41205 ( \41548 , \41546 , \41547 );
xor \U$41206 ( \41549 , \41454 , \41548 );
not \U$41207 ( \41550 , \41373 );
and \U$41208 ( \41551 , \41438 , \41550 );
not \U$41209 ( \41552 , \41438 );
and \U$41210 ( \41553 , \41552 , \41373 );
or \U$41211 ( \41554 , \41551 , \41553 );
and \U$41212 ( \41555 , \41549 , \41554 );
and \U$41213 ( \41556 , \41454 , \41548 );
or \U$41214 ( \41557 , \41555 , \41556 );
nor \U$41215 ( \41558 , \41452 , \41557 );
not \U$41216 ( \41559 , \41558 );
xor \U$41217 ( \41560 , \41344 , \41349 );
xor \U$41218 ( \41561 , \41560 , \41355 );
not \U$41219 ( \41562 , \41366 );
not \U$41220 ( \41563 , \41562 );
not \U$41221 ( \41564 , \41448 );
or \U$41222 ( \41565 , \41563 , \41564 );
nand \U$41223 ( \41566 , \41443 , \41370 );
nand \U$41224 ( \41567 , \41565 , \41566 );
nand \U$41225 ( \41568 , \41561 , \41567 );
not \U$41226 ( \41569 , \41568 );
or \U$41227 ( \41570 , \41559 , \41569 );
or \U$41228 ( \41571 , \41567 , \41561 );
nand \U$41229 ( \41572 , \41570 , \41571 );
nand \U$41230 ( \41573 , \41251 , \41358 );
nand \U$41231 ( \41574 , \41572 , \41573 );
not \U$41232 ( \41575 , \41574 );
or \U$41233 ( \41576 , \41360 , \41575 );
and \U$41234 ( \41577 , \41077 , \41079 );
not \U$41235 ( \41578 , \41077 );
not \U$41236 ( \41579 , \41079 );
and \U$41237 ( \41580 , \41578 , \41579 );
nor \U$41238 ( \41581 , \41577 , \41580 );
not \U$41239 ( \41582 , \41126 );
not \U$41240 ( \41583 , \41582 );
not \U$41241 ( \41584 , \41247 );
or \U$41242 ( \41585 , \41583 , \41584 );
nand \U$41243 ( \41586 , \41245 , \41129 );
nand \U$41244 ( \41587 , \41585 , \41586 );
nand \U$41245 ( \41588 , \41581 , \41587 );
nand \U$41246 ( \41589 , \41576 , \41588 );
xor \U$41247 ( \41590 , \41454 , \41548 );
xor \U$41248 ( \41591 , \41590 , \41554 );
xnor \U$41249 ( \41592 , \41429 , \41382 );
or \U$41250 ( \41593 , RI9873198_182, RI9873210_183);
nand \U$41251 ( \41594 , \41593 , \21779 );
and \U$41252 ( \41595 , RI9873198_182, RI9873210_183);
nor \U$41253 ( \41596 , \41595 , \13022 );
and \U$41254 ( \41597 , \41594 , \41596 );
not \U$41255 ( \41598 , \11342 );
not \U$41256 ( \41599 , \41484 );
or \U$41257 ( \41600 , \41598 , \41599 );
xor \U$41258 ( \41601 , \18704 , RI98730a8_180);
nand \U$41259 ( \41602 , \41601 , \11350 );
nand \U$41260 ( \41603 , \41600 , \41602 );
and \U$41261 ( \41604 , \41597 , \41603 );
not \U$41262 ( \41605 , \17528 );
not \U$41263 ( \41606 , \41503 );
or \U$41264 ( \41607 , \41605 , \41606 );
not \U$41265 ( \41608 , \22715 );
not \U$41266 ( \41609 , \19412 );
or \U$41267 ( \41610 , \41608 , \41609 );
nand \U$41268 ( \41611 , \17726 , RI9873288_184);
nand \U$41269 ( \41612 , \41610 , \41611 );
nand \U$41270 ( \41613 , \41612 , \17543 );
nand \U$41271 ( \41614 , \41607 , \41613 );
xor \U$41272 ( \41615 , \41604 , \41614 );
not \U$41273 ( \41616 , \17251 );
not \U$41274 ( \41617 , RI98733f0_187);
not \U$41275 ( \41618 , \13934 );
or \U$41276 ( \41619 , \41617 , \41618 );
or \U$41277 ( \41620 , \18710 , RI98733f0_187);
nand \U$41278 ( \41621 , \41619 , \41620 );
not \U$41279 ( \41622 , \41621 );
or \U$41280 ( \41623 , \41616 , \41622 );
nand \U$41281 ( \41624 , \41522 , \17263 );
nand \U$41282 ( \41625 , \41623 , \41624 );
and \U$41283 ( \41626 , \41615 , \41625 );
and \U$41284 ( \41627 , \41604 , \41614 );
or \U$41285 ( \41628 , \41626 , \41627 );
not \U$41286 ( \41629 , \41628 );
not \U$41287 ( \41630 , \41629 );
not \U$41288 ( \41631 , \41462 );
not \U$41289 ( \41632 , \41511 );
or \U$41290 ( \41633 , \41631 , \41632 );
or \U$41291 ( \41634 , \41462 , \41511 );
nand \U$41292 ( \41635 , \41633 , \41634 );
not \U$41293 ( \41636 , \41635 );
or \U$41294 ( \41637 , \41630 , \41636 );
or \U$41295 ( \41638 , \41635 , \41629 );
nand \U$41296 ( \41639 , \41637 , \41638 );
not \U$41297 ( \41640 , \41639 );
xor \U$41298 ( \41641 , \41474 , \41490 );
not \U$41299 ( \41642 , \18544 );
xor \U$41300 ( \41643 , \32173 , RI9873558_190);
not \U$41301 ( \41644 , \41643 );
or \U$41302 ( \41645 , \41642 , \41644 );
nand \U$41303 ( \41646 , \41534 , RI9873648_192);
nand \U$41304 ( \41647 , \41645 , \41646 );
xor \U$41305 ( \41648 , \41641 , \41647 );
not \U$41306 ( \41649 , \41460 );
not \U$41307 ( \41650 , \39898 );
and \U$41308 ( \41651 , \41649 , \41650 );
not \U$41309 ( \41652 , \18350 );
not \U$41310 ( \41653 , RI98734e0_189);
or \U$41311 ( \41654 , \41652 , \41653 );
or \U$41312 ( \41655 , \29137 , RI98734e0_189);
nand \U$41313 ( \41656 , \41654 , \41655 );
and \U$41314 ( \41657 , \41656 , \19243 );
nor \U$41315 ( \41658 , \41651 , \41657 );
not \U$41316 ( \41659 , \41658 );
and \U$41317 ( \41660 , \41648 , \41659 );
and \U$41318 ( \41661 , \41641 , \41647 );
nor \U$41319 ( \41662 , \41660 , \41661 );
not \U$41320 ( \41663 , \41662 );
not \U$41321 ( \41664 , \41663 );
or \U$41322 ( \41665 , \41640 , \41664 );
nand \U$41323 ( \41666 , \41628 , \41635 );
nand \U$41324 ( \41667 , \41665 , \41666 );
not \U$41325 ( \41668 , \41667 );
xor \U$41326 ( \41669 , \41592 , \41668 );
not \U$41327 ( \41670 , \41545 );
and \U$41328 ( \41671 , \41520 , \41670 );
not \U$41329 ( \41672 , \41520 );
and \U$41330 ( \41673 , \41672 , \41545 );
nor \U$41331 ( \41674 , \41671 , \41673 );
and \U$41332 ( \41675 , \41669 , \41674 );
and \U$41333 ( \41676 , \41592 , \41668 );
or \U$41334 ( \41677 , \41675 , \41676 );
nand \U$41335 ( \41678 , \41591 , \41677 );
not \U$41336 ( \41679 , \41678 );
xor \U$41337 ( \41680 , \41592 , \41668 );
xor \U$41338 ( \41681 , \41680 , \41674 );
xor \U$41339 ( \41682 , \41604 , \41614 );
xor \U$41340 ( \41683 , \41682 , \41625 );
not \U$41341 ( \41684 , \41683 );
not \U$41342 ( \41685 , \41684 );
and \U$41343 ( \41686 , \41612 , \17528 );
not \U$41344 ( \41687 , \32967 );
not \U$41345 ( \41688 , \16995 );
or \U$41346 ( \41689 , \41687 , \41688 );
or \U$41347 ( \41690 , \16995 , \32967 );
nand \U$41348 ( \41691 , \41689 , \41690 );
and \U$41349 ( \41692 , \41691 , \17543 );
nor \U$41350 ( \41693 , \41686 , \41692 );
not \U$41351 ( \41694 , \41693 );
xor \U$41352 ( \41695 , \41597 , \41603 );
not \U$41353 ( \41696 , \41695 );
not \U$41354 ( \41697 , \13483 );
not \U$41355 ( \41698 , \41470 );
or \U$41356 ( \41699 , \41697 , \41698 );
and \U$41357 ( \41700 , RI9873210_183, \17862 );
not \U$41358 ( \41701 , RI9873210_183);
and \U$41359 ( \41702 , \41701 , \19542 );
nor \U$41360 ( \41703 , \41700 , \41702 );
nand \U$41361 ( \41704 , \41703 , \17243 );
nand \U$41362 ( \41705 , \41699 , \41704 );
not \U$41363 ( \41706 , \41705 );
not \U$41364 ( \41707 , \41706 );
or \U$41365 ( \41708 , \41696 , \41707 );
or \U$41366 ( \41709 , \41706 , \41695 );
nand \U$41367 ( \41710 , \41708 , \41709 );
nand \U$41368 ( \41711 , \41694 , \41710 );
nand \U$41369 ( \41712 , \41695 , \41705 );
and \U$41370 ( \41713 , \41711 , \41712 );
not \U$41371 ( \41714 , \41713 );
or \U$41372 ( \41715 , \41685 , \41714 );
not \U$41373 ( \41716 , \17543 );
not \U$41374 ( \41717 , RI9873288_184);
not \U$41375 ( \41718 , \23934 );
or \U$41376 ( \41719 , \41717 , \41718 );
or \U$41377 ( \41720 , \35428 , RI9873288_184);
nand \U$41378 ( \41721 , \41719 , \41720 );
not \U$41379 ( \41722 , \41721 );
or \U$41380 ( \41723 , \41716 , \41722 );
nand \U$41381 ( \41724 , \41691 , \17528 );
nand \U$41382 ( \41725 , \41723 , \41724 );
not \U$41383 ( \41726 , \41725 );
and \U$41384 ( \41727 , \21779 , \11342 );
not \U$41385 ( \41728 , \13482 );
not \U$41386 ( \41729 , \41703 );
or \U$41387 ( \41730 , \41728 , \41729 );
not \U$41388 ( \41731 , \22675 );
not \U$41389 ( \41732 , \23947 );
not \U$41390 ( \41733 , \41732 );
or \U$41391 ( \41734 , \41731 , \41733 );
or \U$41392 ( \41735 , \25166 , \22675 );
nand \U$41393 ( \41736 , \41734 , \41735 );
nand \U$41394 ( \41737 , \41736 , \17243 );
nand \U$41395 ( \41738 , \41730 , \41737 );
xor \U$41396 ( \41739 , \41727 , \41738 );
not \U$41397 ( \41740 , \41739 );
or \U$41398 ( \41741 , \41726 , \41740 );
nand \U$41399 ( \41742 , \41738 , \41727 );
nand \U$41400 ( \41743 , \41741 , \41742 );
not \U$41401 ( \41744 , \17263 );
not \U$41402 ( \41745 , \41621 );
or \U$41403 ( \41746 , \41744 , \41745 );
and \U$41404 ( \41747 , RI98733f0_187, \17741 );
not \U$41405 ( \41748 , RI98733f0_187);
and \U$41406 ( \41749 , \41748 , \32208 );
or \U$41407 ( \41750 , \41747 , \41749 );
nand \U$41408 ( \41751 , \41750 , \17251 );
nand \U$41409 ( \41752 , \41746 , \41751 );
xor \U$41410 ( \41753 , \41743 , \41752 );
not \U$41411 ( \41754 , \19045 );
not \U$41412 ( \41755 , \41656 );
or \U$41413 ( \41756 , \41754 , \41755 );
xnor \U$41414 ( \41757 , RI98734e0_189, \13860 );
nand \U$41415 ( \41758 , \41757 , \24076 );
nand \U$41416 ( \41759 , \41756 , \41758 );
and \U$41417 ( \41760 , \41753 , \41759 );
and \U$41418 ( \41761 , \41743 , \41752 );
or \U$41419 ( \41762 , \41760 , \41761 );
nand \U$41420 ( \41763 , \41715 , \41762 );
not \U$41421 ( \41764 , \41713 );
nand \U$41422 ( \41765 , \41764 , \41683 );
and \U$41423 ( \41766 , \41763 , \41765 );
not \U$41424 ( \41767 , \41541 );
not \U$41425 ( \41768 , \41525 );
not \U$41426 ( \41769 , \41768 );
and \U$41427 ( \41770 , \41767 , \41769 );
and \U$41428 ( \41771 , \41541 , \41768 );
nor \U$41429 ( \41772 , \41770 , \41771 );
xor \U$41430 ( \41773 , \41766 , \41772 );
not \U$41431 ( \41774 , \41639 );
not \U$41432 ( \41775 , \41662 );
and \U$41433 ( \41776 , \41774 , \41775 );
and \U$41434 ( \41777 , \41639 , \41662 );
nor \U$41435 ( \41778 , \41776 , \41777 );
and \U$41436 ( \41779 , \41773 , \41778 );
and \U$41437 ( \41780 , \41766 , \41772 );
or \U$41438 ( \41781 , \41779 , \41780 );
nand \U$41439 ( \41782 , \41681 , \41781 );
not \U$41440 ( \41783 , \41782 );
not \U$41441 ( \41784 , \41713 );
not \U$41442 ( \41785 , \41683 );
or \U$41443 ( \41786 , \41784 , \41785 );
or \U$41444 ( \41787 , \41683 , \41713 );
nand \U$41445 ( \41788 , \41786 , \41787 );
xor \U$41446 ( \41789 , \41788 , \41762 );
not \U$41447 ( \41790 , \41789 );
not \U$41448 ( \41791 , \41648 );
not \U$41449 ( \41792 , \41658 );
and \U$41450 ( \41793 , \41791 , \41792 );
and \U$41451 ( \41794 , \41648 , \41658 );
nor \U$41452 ( \41795 , \41793 , \41794 );
not \U$41453 ( \41796 , \41795 );
not \U$41454 ( \41797 , \41796 );
or \U$41455 ( \41798 , \41790 , \41797 );
or \U$41456 ( \41799 , \41796 , \41789 );
not \U$41457 ( \41800 , \41693 );
not \U$41458 ( \41801 , \41710 );
or \U$41459 ( \41802 , \41800 , \41801 );
or \U$41460 ( \41803 , \41710 , \41693 );
nand \U$41461 ( \41804 , \41802 , \41803 );
not \U$41462 ( \41805 , \13482 );
not \U$41463 ( \41806 , \41736 );
or \U$41464 ( \41807 , \41805 , \41806 );
xor \U$41465 ( \41808 , RI9873210_183, \18704 );
nand \U$41466 ( \41809 , \41808 , \13475 );
nand \U$41467 ( \41810 , \41807 , \41809 );
not \U$41468 ( \41811 , \13471 );
and \U$41469 ( \41812 , \18704 , \41811 );
nor \U$41470 ( \41813 , \41812 , \13381 );
nand \U$41471 ( \41814 , \41810 , \41813 );
not \U$41472 ( \41815 , \41814 );
not \U$41473 ( \41816 , \41815 );
not \U$41474 ( \41817 , \17251 );
not \U$41475 ( \41818 , \17539 );
not \U$41476 ( \41819 , \19412 );
or \U$41477 ( \41820 , \41818 , \41819 );
or \U$41478 ( \41821 , \27888 , \17539 );
nand \U$41479 ( \41822 , \41820 , \41821 );
not \U$41480 ( \41823 , \41822 );
or \U$41481 ( \41824 , \41817 , \41823 );
nand \U$41482 ( \41825 , \41750 , \17263 );
nand \U$41483 ( \41826 , \41824 , \41825 );
not \U$41484 ( \41827 , \41826 );
or \U$41485 ( \41828 , \41816 , \41827 );
or \U$41486 ( \41829 , \41826 , \41815 );
not \U$41487 ( \41830 , \24076 );
and \U$41488 ( \41831 , RI98734e0_189, \25380 );
not \U$41489 ( \41832 , RI98734e0_189);
and \U$41490 ( \41833 , \41832 , \13933 );
or \U$41491 ( \41834 , \41831 , \41833 );
not \U$41492 ( \41835 , \41834 );
or \U$41493 ( \41836 , \41830 , \41835 );
nand \U$41494 ( \41837 , \41757 , \19045 );
nand \U$41495 ( \41838 , \41836 , \41837 );
nand \U$41496 ( \41839 , \41829 , \41838 );
nand \U$41497 ( \41840 , \41828 , \41839 );
xor \U$41498 ( \41841 , \41804 , \41840 );
not \U$41499 ( \41842 , RI9873648_192);
not \U$41500 ( \41843 , \41643 );
or \U$41501 ( \41844 , \41842 , \41843 );
and \U$41502 ( \41845 , \19594 , RI9873558_190);
not \U$41503 ( \41846 , \19594 );
and \U$41504 ( \41847 , \41846 , \18239 );
nor \U$41505 ( \41848 , \41845 , \41847 );
nand \U$41506 ( \41849 , \18544 , \41848 );
nand \U$41507 ( \41850 , \41844 , \41849 );
and \U$41508 ( \41851 , \41841 , \41850 );
and \U$41509 ( \41852 , \41804 , \41840 );
or \U$41510 ( \41853 , \41851 , \41852 );
nand \U$41511 ( \41854 , \41799 , \41853 );
nand \U$41512 ( \41855 , \41798 , \41854 );
not \U$41513 ( \41856 , \41855 );
xor \U$41514 ( \41857 , \41766 , \41772 );
xor \U$41515 ( \41858 , \41857 , \41778 );
nand \U$41516 ( \41859 , \41856 , \41858 );
not \U$41517 ( \41860 , \41859 );
not \U$41518 ( \41861 , \17263 );
not \U$41519 ( \41862 , \41822 );
or \U$41520 ( \41863 , \41861 , \41862 );
xor \U$41521 ( \41864 , RI98733f0_187, \19518 );
nand \U$41522 ( \41865 , \41864 , \17251 );
nand \U$41523 ( \41866 , \41863 , \41865 );
not \U$41524 ( \41867 , \17263 );
not \U$41525 ( \41868 , \41864 );
or \U$41526 ( \41869 , \41867 , \41868 );
not \U$41527 ( \41870 , RI98733f0_187);
not \U$41528 ( \41871 , \20489 );
or \U$41529 ( \41872 , \41870 , \41871 );
or \U$41530 ( \41873 , \20489 , RI98733f0_187);
nand \U$41531 ( \41874 , \41872 , \41873 );
nand \U$41532 ( \41875 , \41874 , \17251 );
nand \U$41533 ( \41876 , \41869 , \41875 );
not \U$41534 ( \41877 , \41876 );
not \U$41535 ( \41878 , \17527 );
not \U$41536 ( \41879 , RI9873288_184);
not \U$41537 ( \41880 , \19542 );
or \U$41538 ( \41881 , \41879 , \41880 );
or \U$41539 ( \41882 , \19542 , RI9873288_184);
nand \U$41540 ( \41883 , \41881 , \41882 );
not \U$41541 ( \41884 , \41883 );
or \U$41542 ( \41885 , \41878 , \41884 );
not \U$41543 ( \41886 , RI9873288_184);
not \U$41544 ( \41887 , \21772 );
or \U$41545 ( \41888 , \41886 , \41887 );
or \U$41546 ( \41889 , \18193 , RI9873288_184);
nand \U$41547 ( \41890 , \41888 , \41889 );
nand \U$41548 ( \41891 , \41890 , \17542 );
nand \U$41549 ( \41892 , \41885 , \41891 );
not \U$41550 ( \41893 , \41892 );
nand \U$41551 ( \41894 , \18705 , \13482 );
not \U$41552 ( \41895 , \41894 );
and \U$41553 ( \41896 , \41893 , \41895 );
and \U$41554 ( \41897 , \41892 , \41894 );
nor \U$41555 ( \41898 , \41896 , \41897 );
not \U$41556 ( \41899 , \41898 );
not \U$41557 ( \41900 , \41899 );
or \U$41558 ( \41901 , \41877 , \41900 );
not \U$41559 ( \41902 , \41894 );
nand \U$41560 ( \41903 , \41902 , \41892 );
nand \U$41561 ( \41904 , \41901 , \41903 );
xor \U$41562 ( \41905 , \41866 , \41904 );
not \U$41563 ( \41906 , RI9873648_192);
not \U$41564 ( \41907 , RI9873558_190);
not \U$41565 ( \41908 , \18350 );
or \U$41566 ( \41909 , \41907 , \41908 );
or \U$41567 ( \41910 , \17783 , RI9873558_190);
nand \U$41568 ( \41911 , \41909 , \41910 );
not \U$41569 ( \41912 , \41911 );
or \U$41570 ( \41913 , \41906 , \41912 );
not \U$41571 ( \41914 , RI9873558_190);
not \U$41572 ( \41915 , \17013 );
or \U$41573 ( \41916 , \41914 , \41915 );
or \U$41574 ( \41917 , \17013 , RI9873558_190);
nand \U$41575 ( \41918 , \41916 , \41917 );
nand \U$41576 ( \41919 , \41918 , \18543 );
nand \U$41577 ( \41920 , \41913 , \41919 );
and \U$41578 ( \41921 , \41905 , \41920 );
and \U$41579 ( \41922 , \41866 , \41904 );
or \U$41580 ( \41923 , \41921 , \41922 );
not \U$41581 ( \41924 , \41923 );
not \U$41582 ( \41925 , \41826 );
not \U$41583 ( \41926 , \41814 );
and \U$41584 ( \41927 , \41925 , \41926 );
and \U$41585 ( \41928 , \41826 , \41814 );
nor \U$41586 ( \41929 , \41927 , \41928 );
and \U$41587 ( \41930 , \41929 , \41838 );
not \U$41588 ( \41931 , \41929 );
not \U$41589 ( \41932 , \41838 );
and \U$41590 ( \41933 , \41931 , \41932 );
nor \U$41591 ( \41934 , \41930 , \41933 );
not \U$41592 ( \41935 , \41934 );
not \U$41593 ( \41936 , \41935 );
or \U$41594 ( \41937 , \41924 , \41936 );
or \U$41595 ( \41938 , \41935 , \41923 );
or \U$41596 ( \41939 , \41810 , \41813 );
nand \U$41597 ( \41940 , \41939 , \41814 );
not \U$41598 ( \41941 , \41940 );
not \U$41599 ( \41942 , \17528 );
not \U$41600 ( \41943 , \41721 );
or \U$41601 ( \41944 , \41942 , \41943 );
nand \U$41602 ( \41945 , \41883 , \17543 );
nand \U$41603 ( \41946 , \41944 , \41945 );
nor \U$41604 ( \41947 , \41941 , \41946 );
not \U$41605 ( \41948 , \41947 );
not \U$41606 ( \41949 , \41948 );
not \U$41607 ( \41950 , \19045 );
not \U$41608 ( \41951 , \41834 );
or \U$41609 ( \41952 , \41950 , \41951 );
xnor \U$41610 ( \41953 , RI98734e0_189, \19394 );
nand \U$41611 ( \41954 , \41953 , \19034 );
nand \U$41612 ( \41955 , \41952 , \41954 );
not \U$41613 ( \41956 , \41955 );
or \U$41614 ( \41957 , \41949 , \41956 );
not \U$41615 ( \41958 , \41940 );
nand \U$41616 ( \41959 , \41958 , \41946 );
nand \U$41617 ( \41960 , \41957 , \41959 );
not \U$41618 ( \41961 , \41960 );
not \U$41619 ( \41962 , \41961 );
xor \U$41620 ( \41963 , \41725 , \41739 );
not \U$41621 ( \41964 , \18543 );
not \U$41622 ( \41965 , \41911 );
or \U$41623 ( \41966 , \41964 , \41965 );
nand \U$41624 ( \41967 , \41848 , RI9873648_192);
nand \U$41625 ( \41968 , \41966 , \41967 );
xor \U$41626 ( \41969 , \41963 , \41968 );
not \U$41627 ( \41970 , \41969 );
or \U$41628 ( \41971 , \41962 , \41970 );
or \U$41629 ( \41972 , \41969 , \41961 );
nand \U$41630 ( \41973 , \41971 , \41972 );
nand \U$41631 ( \41974 , \41938 , \41973 );
nand \U$41632 ( \41975 , \41937 , \41974 );
not \U$41633 ( \41976 , \41975 );
and \U$41634 ( \41977 , \41963 , \41968 );
or \U$41635 ( \41978 , \41977 , \41960 );
or \U$41636 ( \41979 , \41963 , \41968 );
nand \U$41637 ( \41980 , \41978 , \41979 );
not \U$41638 ( \41981 , \41980 );
xor \U$41639 ( \41982 , \41743 , \41752 );
xor \U$41640 ( \41983 , \41982 , \41759 );
not \U$41641 ( \41984 , \41983 );
or \U$41642 ( \41985 , \41981 , \41984 );
or \U$41643 ( \41986 , \41980 , \41983 );
nand \U$41644 ( \41987 , \41985 , \41986 );
not \U$41645 ( \41988 , \41987 );
xor \U$41646 ( \41989 , \41804 , \41840 );
xor \U$41647 ( \41990 , \41989 , \41850 );
not \U$41648 ( \41991 , \41990 );
or \U$41649 ( \41992 , \41988 , \41991 );
or \U$41650 ( \41993 , \41990 , \41987 );
nand \U$41651 ( \41994 , \41992 , \41993 );
nand \U$41652 ( \41995 , \41976 , \41994 );
not \U$41653 ( \41996 , \41995 );
not \U$41654 ( \41997 , \41973 );
not \U$41655 ( \41998 , \41923 );
not \U$41656 ( \41999 , \41934 );
or \U$41657 ( \42000 , \41998 , \41999 );
or \U$41658 ( \42001 , \41923 , \41934 );
nand \U$41659 ( \42002 , \42000 , \42001 );
not \U$41660 ( \42003 , \42002 );
or \U$41661 ( \42004 , \41997 , \42003 );
or \U$41662 ( \42005 , \42002 , \41973 );
nand \U$41663 ( \42006 , \42004 , \42005 );
xor \U$41664 ( \42007 , \41866 , \41904 );
xor \U$41665 ( \42008 , \42007 , \41920 );
not \U$41666 ( \42009 , \42008 );
not \U$41667 ( \42010 , \42009 );
not \U$41668 ( \42011 , \18543 );
not \U$41669 ( \42012 , RI9873558_190);
not \U$41670 ( \42013 , \20449 );
or \U$41671 ( \42014 , \42012 , \42013 );
or \U$41672 ( \42015 , \25380 , RI9873558_190);
nand \U$41673 ( \42016 , \42014 , \42015 );
not \U$41674 ( \42017 , \42016 );
or \U$41675 ( \42018 , \42011 , \42017 );
nand \U$41676 ( \42019 , \41918 , RI9873648_192);
nand \U$41677 ( \42020 , \42018 , \42019 );
not \U$41678 ( \42021 , \42020 );
not \U$41679 ( \42022 , \19044 );
not \U$41680 ( \42023 , \41953 );
or \U$41681 ( \42024 , \42022 , \42023 );
and \U$41682 ( \42025 , RI98734e0_189, \19411 );
not \U$41683 ( \42026 , RI98734e0_189);
and \U$41684 ( \42027 , \42026 , \17725 );
or \U$41685 ( \42028 , \42025 , \42027 );
nand \U$41686 ( \42029 , \42028 , \19034 );
nand \U$41687 ( \42030 , \42024 , \42029 );
not \U$41688 ( \42031 , \17527 );
not \U$41689 ( \42032 , \41890 );
or \U$41690 ( \42033 , \42031 , \42032 );
xor \U$41691 ( \42034 , \18704 , RI9873288_184);
nand \U$41692 ( \42035 , \42034 , \17542 );
nand \U$41693 ( \42036 , \42033 , \42035 );
not \U$41694 ( \42037 , \42036 );
or \U$41695 ( \42038 , RI9873378_186, RI98733f0_187);
nand \U$41696 ( \42039 , \42038 , \18704 );
nand \U$41697 ( \42040 , \42039 , \13865 );
nor \U$41698 ( \42041 , \42037 , \42040 );
nand \U$41699 ( \42042 , \42030 , \42041 );
buf \U$41700 ( \42043 , \42042 );
and \U$41701 ( \42044 , \42021 , \42043 );
nor \U$41702 ( \42045 , \42030 , \42041 );
nor \U$41703 ( \42046 , \42044 , \42045 );
not \U$41704 ( \42047 , \42046 );
not \U$41705 ( \42048 , \41947 );
nand \U$41706 ( \42049 , \42048 , \41959 );
xor \U$41707 ( \42050 , \42049 , \41955 );
not \U$41708 ( \42051 , \42050 );
or \U$41709 ( \42052 , \42047 , \42051 );
or \U$41710 ( \42053 , \42046 , \42050 );
nand \U$41711 ( \42054 , \42052 , \42053 );
not \U$41712 ( \42055 , \42054 );
or \U$41713 ( \42056 , \42010 , \42055 );
not \U$41714 ( \42057 , \42046 );
nand \U$41715 ( \42058 , \42057 , \42050 );
nand \U$41716 ( \42059 , \42056 , \42058 );
nand \U$41717 ( \42060 , \42006 , \42059 );
not \U$41718 ( \42061 , \42060 );
and \U$41719 ( \42062 , \17539 , \23947 );
not \U$41720 ( \42063 , \17539 );
and \U$41721 ( \42064 , \42063 , \25166 );
nor \U$41722 ( \42065 , \42062 , \42064 );
not \U$41723 ( \42066 , \42065 );
or \U$41724 ( \42067 , \42066 , \17262 );
and \U$41725 ( \42068 , \24449 , RI98733f0_187);
and \U$41726 ( \42069 , \18704 , \17539 );
nor \U$41727 ( \42070 , \42068 , \42069 );
or \U$41728 ( \42071 , \42070 , \17250 );
nand \U$41729 ( \42072 , \42067 , \42071 );
not \U$41730 ( \42073 , \42072 );
or \U$41731 ( \42074 , RI9873468_188, RI98734e0_189);
nand \U$41732 ( \42075 , \42074 , \18704 );
nand \U$41733 ( \42076 , \42075 , \21054 );
nor \U$41734 ( \42077 , \42073 , \42076 );
not \U$41735 ( \42078 , \19044 );
not \U$41736 ( \42079 , \16999 );
not \U$41737 ( \42080 , \19518 );
or \U$41738 ( \42081 , \42079 , \42080 );
or \U$41739 ( \42082 , \16995 , \22709 );
nand \U$41740 ( \42083 , \42081 , \42082 );
not \U$41741 ( \42084 , \42083 );
or \U$41742 ( \42085 , \42078 , \42084 );
not \U$41743 ( \42086 , RI98734e0_189);
not \U$41744 ( \42087 , \20489 );
or \U$41745 ( \42088 , \42086 , \42087 );
or \U$41746 ( \42089 , \23934 , RI98734e0_189);
nand \U$41747 ( \42090 , \42088 , \42089 );
nand \U$41748 ( \42091 , \42090 , \19034 );
nand \U$41749 ( \42092 , \42085 , \42091 );
not \U$41750 ( \42093 , \42092 );
not \U$41751 ( \42094 , \42093 );
and \U$41752 ( \42095 , \18704 , \17527 );
not \U$41753 ( \42096 , \17263 );
not \U$41754 ( \42097 , RI98733f0_187);
not \U$41755 ( \42098 , \19542 );
or \U$41756 ( \42099 , \42097 , \42098 );
or \U$41757 ( \42100 , \19542 , RI98733f0_187);
nand \U$41758 ( \42101 , \42099 , \42100 );
not \U$41759 ( \42102 , \42101 );
or \U$41760 ( \42103 , \42096 , \42102 );
nand \U$41761 ( \42104 , \42065 , \17251 );
nand \U$41762 ( \42105 , \42103 , \42104 );
xor \U$41763 ( \42106 , \42095 , \42105 );
not \U$41764 ( \42107 , \42106 );
or \U$41765 ( \42108 , \42094 , \42107 );
not \U$41766 ( \42109 , \42106 );
nand \U$41767 ( \42110 , \42109 , \42092 );
nand \U$41768 ( \42111 , \42108 , \42110 );
xor \U$41769 ( \42112 , \42077 , \42111 );
not \U$41770 ( \42113 , \18543 );
not \U$41771 ( \42114 , RI9873558_190);
not \U$41772 ( \42115 , \31875 );
or \U$41773 ( \42116 , \42114 , \42115 );
or \U$41774 ( \42117 , \17868 , RI9873558_190);
nand \U$41775 ( \42118 , \42116 , \42117 );
not \U$41776 ( \42119 , \42118 );
or \U$41777 ( \42120 , \42113 , \42119 );
not \U$41778 ( \42121 , RI9873558_190);
not \U$41779 ( \42122 , \17911 );
or \U$41780 ( \42123 , \42121 , \42122 );
or \U$41781 ( \42124 , \17908 , RI9873558_190);
nand \U$41782 ( \42125 , \42123 , \42124 );
nand \U$41783 ( \42126 , \42125 , RI9873648_192);
nand \U$41784 ( \42127 , \42120 , \42126 );
and \U$41785 ( \42128 , \42112 , \42127 );
and \U$41786 ( \42129 , \42077 , \42111 );
or \U$41787 ( \42130 , \42128 , \42129 );
not \U$41788 ( \42131 , \42130 );
and \U$41789 ( \42132 , \42106 , \42092 );
and \U$41790 ( \42133 , \42095 , \42105 );
nor \U$41791 ( \42134 , \42132 , \42133 );
not \U$41792 ( \42135 , \42016 );
not \U$41793 ( \42136 , \42135 );
not \U$41794 ( \42137 , \18542 );
and \U$41795 ( \42138 , \42136 , \42137 );
not \U$41796 ( \42139 , \42125 );
not \U$41797 ( \42140 , \18543 );
nor \U$41798 ( \42141 , \42139 , \42140 );
nor \U$41799 ( \42142 , \42138 , \42141 );
xor \U$41800 ( \42143 , \42134 , \42142 );
not \U$41801 ( \42144 , \17263 );
not \U$41802 ( \42145 , \41874 );
or \U$41803 ( \42146 , \42144 , \42145 );
nand \U$41804 ( \42147 , \42101 , \17251 );
nand \U$41805 ( \42148 , \42146 , \42147 );
not \U$41806 ( \42149 , \42148 );
not \U$41807 ( \42150 , \42036 );
not \U$41808 ( \42151 , \42040 );
and \U$41809 ( \42152 , \42150 , \42151 );
and \U$41810 ( \42153 , \42036 , \42040 );
nor \U$41811 ( \42154 , \42152 , \42153 );
not \U$41812 ( \42155 , \42154 );
or \U$41813 ( \42156 , \42149 , \42155 );
or \U$41814 ( \42157 , \42148 , \42154 );
nand \U$41815 ( \42158 , \42156 , \42157 );
not \U$41816 ( \42159 , \19044 );
not \U$41817 ( \42160 , \42028 );
or \U$41818 ( \42161 , \42159 , \42160 );
nand \U$41819 ( \42162 , \42083 , \19034 );
nand \U$41820 ( \42163 , \42161 , \42162 );
not \U$41821 ( \42164 , \42163 );
and \U$41822 ( \42165 , \42158 , \42164 );
not \U$41823 ( \42166 , \42158 );
and \U$41824 ( \42167 , \42166 , \42163 );
nor \U$41825 ( \42168 , \42165 , \42167 );
xor \U$41826 ( \42169 , \42143 , \42168 );
not \U$41827 ( \42170 , \42169 );
not \U$41828 ( \42171 , \42170 );
or \U$41829 ( \42172 , \42131 , \42171 );
xor \U$41830 ( \42173 , \42134 , \42142 );
and \U$41831 ( \42174 , \42173 , \42168 );
and \U$41832 ( \42175 , \42134 , \42142 );
or \U$41833 ( \42176 , \42174 , \42175 );
not \U$41834 ( \42177 , \42176 );
xor \U$41835 ( \42178 , \41898 , \41876 );
not \U$41836 ( \42179 , \42178 );
not \U$41837 ( \42180 , \42163 );
not \U$41838 ( \42181 , \42158 );
or \U$41839 ( \42182 , \42180 , \42181 );
not \U$41840 ( \42183 , \42154 );
nand \U$41841 ( \42184 , \42183 , \42148 );
nand \U$41842 ( \42185 , \42182 , \42184 );
not \U$41843 ( \42186 , \42185 );
or \U$41844 ( \42187 , \42179 , \42186 );
or \U$41845 ( \42188 , \42185 , \42178 );
nand \U$41846 ( \42189 , \42187 , \42188 );
not \U$41847 ( \42190 , \42189 );
not \U$41848 ( \42191 , \42045 );
nand \U$41849 ( \42192 , \42191 , \42042 );
not \U$41850 ( \42193 , \42192 );
not \U$41851 ( \42194 , \42020 );
and \U$41852 ( \42195 , \42193 , \42194 );
and \U$41853 ( \42196 , \42192 , \42020 );
nor \U$41854 ( \42197 , \42195 , \42196 );
not \U$41855 ( \42198 , \42197 );
or \U$41856 ( \42199 , \42190 , \42198 );
or \U$41857 ( \42200 , \42189 , \42197 );
nand \U$41858 ( \42201 , \42199 , \42200 );
nand \U$41859 ( \42202 , \42177 , \42201 );
nand \U$41860 ( \42203 , \42172 , \42202 );
not \U$41861 ( \42204 , \42203 );
not \U$41862 ( \42205 , \42130 );
nand \U$41863 ( \42206 , \42205 , \42169 );
xor \U$41864 ( \42207 , \42077 , \42111 );
xor \U$41865 ( \42208 , \42207 , \42127 );
not \U$41866 ( \42209 , RI9873648_192);
not \U$41867 ( \42210 , \42118 );
or \U$41868 ( \42211 , \42209 , \42210 );
and \U$41869 ( \42212 , RI9873558_190, \19519 );
not \U$41870 ( \42213 , RI9873558_190);
and \U$41871 ( \42214 , \42213 , \24867 );
nor \U$41872 ( \42215 , \42212 , \42214 );
nand \U$41873 ( \42216 , \42215 , \18543 );
nand \U$41874 ( \42217 , \42211 , \42216 );
not \U$41875 ( \42218 , \42217 );
not \U$41876 ( \42219 , RI98734e0_189);
not \U$41877 ( \42220 , \19542 );
or \U$41878 ( \42221 , \42219 , \42220 );
or \U$41879 ( \42222 , \19542 , RI98734e0_189);
nand \U$41880 ( \42223 , \42221 , \42222 );
not \U$41881 ( \42224 , \42223 );
not \U$41882 ( \42225 , \19034 );
or \U$41883 ( \42226 , \42224 , \42225 );
not \U$41884 ( \42227 , \19032 );
nand \U$41885 ( \42228 , \42227 , \42090 );
nand \U$41886 ( \42229 , \42226 , \42228 );
not \U$41887 ( \42230 , \42229 );
not \U$41888 ( \42231 , \42072 );
not \U$41889 ( \42232 , \42076 );
and \U$41890 ( \42233 , \42231 , \42232 );
and \U$41891 ( \42234 , \42072 , \42076 );
nor \U$41892 ( \42235 , \42233 , \42234 );
not \U$41893 ( \42236 , \42235 );
or \U$41894 ( \42237 , \42230 , \42236 );
or \U$41895 ( \42238 , \42235 , \42229 );
nand \U$41896 ( \42239 , \42237 , \42238 );
not \U$41897 ( \42240 , \42239 );
or \U$41898 ( \42241 , \42218 , \42240 );
not \U$41899 ( \42242 , \42235 );
nand \U$41900 ( \42243 , \42242 , \42229 );
nand \U$41901 ( \42244 , \42241 , \42243 );
nand \U$41902 ( \42245 , \42208 , \42244 );
not \U$41903 ( \42246 , RI9873648_192);
not \U$41904 ( \42247 , \42215 );
or \U$41905 ( \42248 , \42246 , \42247 );
and \U$41906 ( \42249 , RI9873558_190, \39613 );
not \U$41907 ( \42250 , RI9873558_190);
and \U$41908 ( \42251 , \42250 , \17702 );
or \U$41909 ( \42252 , \42249 , \42251 );
nand \U$41910 ( \42253 , \42252 , \18543 );
nand \U$41911 ( \42254 , \42248 , \42253 );
not \U$41912 ( \42255 , \42254 );
not \U$41913 ( \42256 , \19044 );
not \U$41914 ( \42257 , \42223 );
or \U$41915 ( \42258 , \42256 , \42257 );
and \U$41916 ( \42259 , RI98734e0_189, \28671 );
not \U$41917 ( \42260 , RI98734e0_189);
and \U$41918 ( \42261 , \42260 , \23949 );
nor \U$41919 ( \42262 , \42259 , \42261 );
nand \U$41920 ( \42263 , \42262 , \19034 );
nand \U$41921 ( \42264 , \42258 , \42263 );
and \U$41922 ( \42265 , \21779 , \17263 );
or \U$41923 ( \42266 , \42264 , \42265 );
not \U$41924 ( \42267 , \42266 );
or \U$41925 ( \42268 , \42255 , \42267 );
nand \U$41926 ( \42269 , \42264 , \42265 );
nand \U$41927 ( \42270 , \42268 , \42269 );
not \U$41928 ( \42271 , \42270 );
not \U$41929 ( \42272 , \42239 );
not \U$41930 ( \42273 , \42217 );
not \U$41931 ( \42274 , \42273 );
and \U$41932 ( \42275 , \42272 , \42274 );
and \U$41933 ( \42276 , \42239 , \42273 );
nor \U$41934 ( \42277 , \42275 , \42276 );
nand \U$41935 ( \42278 , \42271 , \42277 );
not \U$41936 ( \42279 , \19044 );
not \U$41937 ( \42280 , \42262 );
or \U$41938 ( \42281 , \42279 , \42280 );
not \U$41939 ( \42282 , \35146 );
not \U$41940 ( \42283 , \21779 );
or \U$41941 ( \42284 , \42282 , \42283 );
or \U$41942 ( \42285 , \18705 , \16999 );
nand \U$41943 ( \42286 , \42284 , \42285 );
nand \U$41944 ( \42287 , \42286 , \19034 );
nand \U$41945 ( \42288 , \42281 , \42287 );
or \U$41946 ( \42289 , RI9873558_190, RI98735d0_191);
nand \U$41947 ( \42290 , \42289 , \18704 );
nand \U$41948 ( \42291 , \42290 , \17000 );
not \U$41949 ( \42292 , \42291 );
nand \U$41950 ( \42293 , \42288 , \42292 );
not \U$41951 ( \42294 , \42293 );
not \U$41952 ( \42295 , \42294 );
not \U$41953 ( \42296 , \18543 );
and \U$41954 ( \42297 , \19542 , \18239 );
not \U$41955 ( \42298 , \19542 );
and \U$41956 ( \42299 , \42298 , RI9873558_190);
nor \U$41957 ( \42300 , \42297 , \42299 );
not \U$41958 ( \42301 , \42300 );
or \U$41959 ( \42302 , \42296 , \42301 );
nand \U$41960 ( \42303 , \42252 , RI9873648_192);
nand \U$41961 ( \42304 , \42302 , \42303 );
not \U$41962 ( \42305 , \42304 );
and \U$41963 ( \42306 , \42288 , \42291 );
not \U$41964 ( \42307 , \42288 );
and \U$41965 ( \42308 , \42307 , \42292 );
or \U$41966 ( \42309 , \42306 , \42308 );
not \U$41967 ( \42310 , \42309 );
or \U$41968 ( \42311 , \42305 , \42310 );
or \U$41969 ( \42312 , \42309 , \42304 );
not \U$41970 ( \42313 , RI9873648_192);
not \U$41971 ( \42314 , \42300 );
or \U$41972 ( \42315 , \42313 , \42314 );
nand \U$41973 ( \42316 , \42315 , \42140 );
nand \U$41974 ( \42317 , \18705 , RI9873648_192);
and \U$41975 ( \42318 , \18195 , \42317 );
and \U$41976 ( \42319 , \21778 , \18239 );
and \U$41977 ( \42320 , \28663 , \19032 );
nor \U$41978 ( \42321 , \42318 , \42319 , \42320 );
and \U$41979 ( \42322 , \42316 , \42321 );
nand \U$41980 ( \42323 , \42312 , \42322 );
nand \U$41981 ( \42324 , \42311 , \42323 );
not \U$41982 ( \42325 , \42324 );
or \U$41983 ( \42326 , \42295 , \42325 );
nand \U$41984 ( \42327 , \42266 , \42269 );
and \U$41985 ( \42328 , \42327 , \42254 );
not \U$41986 ( \42329 , \42327 );
not \U$41987 ( \42330 , \42254 );
and \U$41988 ( \42331 , \42329 , \42330 );
nor \U$41989 ( \42332 , \42328 , \42331 );
nand \U$41990 ( \42333 , \42326 , \42332 );
not \U$41991 ( \42334 , \42324 );
nand \U$41992 ( \42335 , \42334 , \42293 );
nand \U$41993 ( \42336 , \42278 , \42333 , \42335 );
not \U$41994 ( \42337 , \42277 );
nand \U$41995 ( \42338 , \42337 , \42270 );
nand \U$41996 ( \42339 , \42245 , \42336 , \42338 );
not \U$41997 ( \42340 , \42208 );
not \U$41998 ( \42341 , \42244 );
nand \U$41999 ( \42342 , \42340 , \42341 );
and \U$42000 ( \42343 , \42206 , \42339 , \42342 );
not \U$42001 ( \42344 , \42343 );
and \U$42002 ( \42345 , \42204 , \42344 );
not \U$42003 ( \42346 , \42201 );
and \U$42004 ( \42347 , \42346 , \42176 );
nor \U$42005 ( \42348 , \42345 , \42347 );
not \U$42006 ( \42349 , \42008 );
not \U$42007 ( \42350 , \42054 );
or \U$42008 ( \42351 , \42349 , \42350 );
or \U$42009 ( \42352 , \42054 , \42008 );
nand \U$42010 ( \42353 , \42351 , \42352 );
not \U$42011 ( \42354 , \42185 );
not \U$42012 ( \42355 , \42354 );
not \U$42013 ( \42356 , \42178 );
and \U$42014 ( \42357 , \42355 , \42356 );
not \U$42015 ( \42358 , \42197 );
and \U$42016 ( \42359 , \42189 , \42358 );
nor \U$42017 ( \42360 , \42357 , \42359 );
nand \U$42018 ( \42361 , \42353 , \42360 );
nand \U$42019 ( \42362 , \42348 , \42361 );
or \U$42020 ( \42363 , \42360 , \42353 );
nand \U$42021 ( \42364 , \42362 , \42363 );
not \U$42022 ( \42365 , \42364 );
or \U$42023 ( \42366 , \42061 , \42365 );
or \U$42024 ( \42367 , \42059 , \42006 );
nand \U$42025 ( \42368 , \42366 , \42367 );
not \U$42026 ( \42369 , \42368 );
or \U$42027 ( \42370 , \41996 , \42369 );
not \U$42028 ( \42371 , \41994 );
nand \U$42029 ( \42372 , \41975 , \42371 );
nand \U$42030 ( \42373 , \42370 , \42372 );
not \U$42031 ( \42374 , \42373 );
not \U$42032 ( \42375 , \41789 );
not \U$42033 ( \42376 , \41796 );
not \U$42034 ( \42377 , \41853 );
not \U$42035 ( \42378 , \42377 );
or \U$42036 ( \42379 , \42376 , \42378 );
nand \U$42037 ( \42380 , \41795 , \41853 );
nand \U$42038 ( \42381 , \42379 , \42380 );
not \U$42039 ( \42382 , \42381 );
or \U$42040 ( \42383 , \42375 , \42382 );
or \U$42041 ( \42384 , \42381 , \41789 );
nand \U$42042 ( \42385 , \42383 , \42384 );
not \U$42043 ( \42386 , \41980 );
not \U$42044 ( \42387 , \41983 );
not \U$42045 ( \42388 , \42387 );
or \U$42046 ( \42389 , \42386 , \42388 );
not \U$42047 ( \42390 , \41990 );
nand \U$42048 ( \42391 , \42390 , \41987 );
nand \U$42049 ( \42392 , \42389 , \42391 );
nand \U$42050 ( \42393 , \42385 , \42392 );
not \U$42051 ( \42394 , \42393 );
or \U$42052 ( \42395 , \42374 , \42394 );
not \U$42053 ( \42396 , \42385 );
not \U$42054 ( \42397 , \42392 );
nand \U$42055 ( \42398 , \42396 , \42397 );
nand \U$42056 ( \42399 , \42395 , \42398 );
not \U$42057 ( \42400 , \42399 );
or \U$42058 ( \42401 , \41860 , \42400 );
not \U$42059 ( \42402 , \41858 );
nand \U$42060 ( \42403 , \42402 , \41855 );
nand \U$42061 ( \42404 , \42401 , \42403 );
not \U$42062 ( \42405 , \42404 );
or \U$42063 ( \42406 , \41783 , \42405 );
not \U$42064 ( \42407 , \41681 );
not \U$42065 ( \42408 , \41781 );
nand \U$42066 ( \42409 , \42407 , \42408 );
nand \U$42067 ( \42410 , \42406 , \42409 );
not \U$42068 ( \42411 , \42410 );
or \U$42069 ( \42412 , \41679 , \42411 );
nor \U$42070 ( \42413 , \41591 , \41677 );
not \U$42071 ( \42414 , \42413 );
nand \U$42072 ( \42415 , \42412 , \42414 );
not \U$42073 ( \42416 , \41573 );
nand \U$42074 ( \42417 , \41452 , \41557 );
nand \U$42075 ( \42418 , \42417 , \41568 );
nor \U$42076 ( \42419 , \42416 , \42418 );
nand \U$42077 ( \42420 , \42415 , \42419 , \41588 );
or \U$42078 ( \42421 , \41581 , \41587 );
nand \U$42079 ( \42422 , \41589 , \42420 , \42421 );
nand \U$42080 ( \42423 , \41119 , \42422 );
nor \U$42081 ( \42424 , \40957 , \41082 );
nand \U$42082 ( \42425 , \40955 , \42424 );
not \U$42083 ( \42426 , \40733 );
not \U$42084 ( \42427 , \40954 );
nand \U$42085 ( \42428 , \42426 , \42427 );
nand \U$42086 ( \42429 , \42425 , \42428 );
nand \U$42087 ( \42430 , \42429 , \41111 );
not \U$42088 ( \42431 , \42430 );
not \U$42089 ( \42432 , \41101 );
nand \U$42090 ( \42433 , \42432 , \41109 );
not \U$42091 ( \42434 , \42433 );
or \U$42092 ( \42435 , \42431 , \42434 );
nand \U$42093 ( \42436 , \42435 , \41118 );
or \U$42094 ( \42437 , \41117 , \41115 );
nand \U$42095 ( \42438 , \42423 , \42436 , \42437 );
nand \U$42096 ( \42439 , \40305 , \40393 );
and \U$42097 ( \42440 , \40302 , \42439 );
nand \U$42098 ( \42441 , \42438 , \40112 , \40412 , \42440 );
or \U$42099 ( \42442 , \40409 , \40411 );
nand \U$42100 ( \42443 , \40413 , \42441 , \42442 );
nand \U$42101 ( \42444 , \39367 , \39670 );
and \U$42102 ( \42445 , \39704 , \42444 );
and \U$42103 ( \42446 , \39720 , \42445 , \38887 );
nand \U$42104 ( \42447 , \42443 , \42446 );
nand \U$42105 ( \42448 , \39729 , \42447 );
and \U$42106 ( \42449 , \37442 , \37644 );
not \U$42107 ( \42450 , \37442 );
and \U$42108 ( \42451 , \42450 , \37645 );
nor \U$42109 ( \42452 , \42449 , \42451 );
not \U$42110 ( \42453 , \37557 );
and \U$42111 ( \42454 , \42452 , \42453 );
not \U$42112 ( \42455 , \42452 );
and \U$42113 ( \42456 , \42455 , \37557 );
nor \U$42114 ( \42457 , \42454 , \42456 );
xor \U$42115 ( \42458 , \37655 , \37693 );
xor \U$42116 ( \42459 , \42458 , \37699 );
xor \U$42117 ( \42460 , \42457 , \42459 );
xor \U$42118 ( \42461 , \37657 , \37686 );
xor \U$42119 ( \42462 , \42461 , \37691 );
not \U$42120 ( \42463 , \38465 );
not \U$42121 ( \42464 , \38447 );
or \U$42122 ( \42465 , \42463 , \42464 );
nand \U$42123 ( \42466 , \42465 , \38463 );
xor \U$42124 ( \42467 , \42462 , \42466 );
not \U$42125 ( \42468 , \37633 );
nand \U$42126 ( \42469 , \42468 , \37642 );
xnor \U$42127 ( \42470 , \42469 , \37641 );
not \U$42128 ( \42471 , \42470 );
xor \U$42129 ( \42472 , \37255 , \37278 );
xnor \U$42130 ( \42473 , \42472 , \37266 );
not \U$42131 ( \42474 , \42473 );
not \U$42132 ( \42475 , \38309 );
not \U$42133 ( \42476 , \38315 );
or \U$42134 ( \42477 , \42475 , \42476 );
not \U$42135 ( \42478 , \38305 );
nand \U$42136 ( \42479 , \42478 , \38298 );
nand \U$42137 ( \42480 , \42477 , \42479 );
not \U$42138 ( \42481 , \42480 );
or \U$42139 ( \42482 , \42474 , \42481 );
or \U$42140 ( \42483 , \42480 , \42473 );
nand \U$42141 ( \42484 , \42482 , \42483 );
not \U$42142 ( \42485 , \42484 );
or \U$42143 ( \42486 , \42471 , \42485 );
or \U$42144 ( \42487 , \42484 , \42470 );
nand \U$42145 ( \42488 , \42486 , \42487 );
and \U$42146 ( \42489 , \42467 , \42488 );
and \U$42147 ( \42490 , \42462 , \42466 );
or \U$42148 ( \42491 , \42489 , \42490 );
and \U$42149 ( \42492 , \42460 , \42491 );
not \U$42150 ( \42493 , \42460 );
not \U$42151 ( \42494 , \42491 );
and \U$42152 ( \42495 , \42493 , \42494 );
nor \U$42153 ( \42496 , \42492 , \42495 );
not \U$42154 ( \42497 , \42496 );
not \U$42155 ( \42498 , \38288 );
not \U$42156 ( \42499 , \38346 );
or \U$42157 ( \42500 , \42498 , \42499 );
not \U$42158 ( \42501 , \38345 );
nand \U$42159 ( \42502 , \42501 , \38316 );
nand \U$42160 ( \42503 , \42500 , \42502 );
not \U$42161 ( \42504 , \38439 );
not \U$42162 ( \42505 , \38473 );
or \U$42163 ( \42506 , \42504 , \42505 );
not \U$42164 ( \42507 , \38436 );
not \U$42165 ( \42508 , \38470 );
or \U$42166 ( \42509 , \42507 , \42508 );
nand \U$42167 ( \42510 , \42509 , \38413 );
nand \U$42168 ( \42511 , \42506 , \42510 );
or \U$42169 ( \42512 , \42503 , \42511 );
xor \U$42170 ( \42513 , \37514 , \37516 );
xnor \U$42171 ( \42514 , \42513 , \37552 );
not \U$42172 ( \42515 , \38432 );
not \U$42173 ( \42516 , \38425 );
not \U$42174 ( \42517 , \42516 );
or \U$42175 ( \42518 , \42515 , \42517 );
not \U$42176 ( \42519 , \38418 );
nand \U$42177 ( \42520 , \42519 , \38421 );
nand \U$42178 ( \42521 , \42518 , \42520 );
xor \U$42179 ( \42522 , \42514 , \42521 );
not \U$42180 ( \42523 , \38242 );
not \U$42181 ( \42524 , \38223 );
not \U$42182 ( \42525 , \38286 );
or \U$42183 ( \42526 , \42524 , \42525 );
or \U$42184 ( \42527 , \38286 , \38223 );
nand \U$42185 ( \42528 , \42526 , \42527 );
not \U$42186 ( \42529 , \42528 );
or \U$42187 ( \42530 , \42523 , \42529 );
not \U$42188 ( \42531 , \38223 );
nand \U$42189 ( \42532 , \42531 , \38286 );
nand \U$42190 ( \42533 , \42530 , \42532 );
xor \U$42191 ( \42534 , \42522 , \42533 );
nand \U$42192 ( \42535 , \42512 , \42534 );
nand \U$42193 ( \42536 , \42503 , \42511 );
nand \U$42194 ( \42537 , \42535 , \42536 );
not \U$42195 ( \42538 , \42537 );
xor \U$42196 ( \42539 , \42514 , \42521 );
and \U$42197 ( \42540 , \42539 , \42533 );
and \U$42198 ( \42541 , \42514 , \42521 );
or \U$42199 ( \42542 , \42540 , \42541 );
xor \U$42200 ( \42543 , \37223 , \37229 );
xor \U$42201 ( \42544 , \42543 , \37231 );
not \U$42202 ( \42545 , \42470 );
not \U$42203 ( \42546 , \42545 );
not \U$42204 ( \42547 , \42484 );
or \U$42205 ( \42548 , \42546 , \42547 );
not \U$42206 ( \42549 , \42473 );
nand \U$42207 ( \42550 , \42549 , \42480 );
nand \U$42208 ( \42551 , \42548 , \42550 );
and \U$42209 ( \42552 , \42544 , \42551 );
not \U$42210 ( \42553 , \42544 );
not \U$42211 ( \42554 , \42551 );
and \U$42212 ( \42555 , \42553 , \42554 );
nor \U$42213 ( \42556 , \42552 , \42555 );
xnor \U$42214 ( \42557 , \42542 , \42556 );
nand \U$42215 ( \42558 , \42538 , \42557 );
not \U$42216 ( \42559 , \42558 );
or \U$42217 ( \42560 , \42497 , \42559 );
not \U$42218 ( \42561 , \42557 );
nand \U$42219 ( \42562 , \42561 , \42537 );
nand \U$42220 ( \42563 , \42560 , \42562 );
not \U$42221 ( \42564 , \42563 );
buf \U$42222 ( \42565 , \42460 );
not \U$42223 ( \42566 , \42494 );
and \U$42224 ( \42567 , \42565 , \42566 );
and \U$42225 ( \42568 , \42457 , \42459 );
nor \U$42226 ( \42569 , \42567 , \42568 );
not \U$42227 ( \42570 , \42544 );
nand \U$42228 ( \42571 , \42570 , \42554 );
not \U$42229 ( \42572 , \42571 );
not \U$42230 ( \42573 , \42542 );
or \U$42231 ( \42574 , \42572 , \42573 );
nand \U$42232 ( \42575 , \42544 , \42551 );
nand \U$42233 ( \42576 , \42574 , \42575 );
not \U$42234 ( \42577 , \42576 );
xor \U$42235 ( \42578 , \42569 , \42577 );
and \U$42236 ( \42579 , \37743 , \37747 );
not \U$42237 ( \42580 , \37743 );
and \U$42238 ( \42581 , \42580 , \37748 );
or \U$42239 ( \42582 , \42579 , \42581 );
xor \U$42240 ( \42583 , \42582 , \37755 );
xor \U$42241 ( \42584 , \42578 , \42583 );
nand \U$42242 ( \42585 , \42564 , \42584 );
xor \U$42243 ( \42586 , \42496 , \42557 );
xnor \U$42244 ( \42587 , \42586 , \42537 );
not \U$42245 ( \42588 , \42587 );
not \U$42246 ( \42589 , \42511 );
not \U$42247 ( \42590 , \42503 );
or \U$42248 ( \42591 , \42589 , \42590 );
or \U$42249 ( \42592 , \42503 , \42511 );
nand \U$42250 ( \42593 , \42591 , \42592 );
not \U$42251 ( \42594 , \42593 );
not \U$42252 ( \42595 , \42534 );
and \U$42253 ( \42596 , \42594 , \42595 );
and \U$42254 ( \42597 , \42593 , \42534 );
nor \U$42255 ( \42598 , \42596 , \42597 );
not \U$42256 ( \42599 , \42598 );
not \U$42257 ( \42600 , \42599 );
xor \U$42258 ( \42601 , \42462 , \42466 );
xor \U$42259 ( \42602 , \42601 , \42488 );
not \U$42260 ( \42603 , \42602 );
not \U$42261 ( \42604 , \38202 );
or \U$42262 ( \42605 , \38351 , \42604 );
nand \U$42263 ( \42606 , \42605 , \38408 );
nand \U$42264 ( \42607 , \38351 , \42604 );
nand \U$42265 ( \42608 , \42606 , \42607 );
not \U$42266 ( \42609 , \42608 );
not \U$42267 ( \42610 , \42609 );
or \U$42268 ( \42611 , \42603 , \42610 );
not \U$42269 ( \42612 , \42602 );
nand \U$42270 ( \42613 , \42612 , \42608 );
nand \U$42271 ( \42614 , \42611 , \42613 );
not \U$42272 ( \42615 , \42614 );
or \U$42273 ( \42616 , \42600 , \42615 );
nand \U$42274 ( \42617 , \42608 , \42602 );
nand \U$42275 ( \42618 , \42616 , \42617 );
not \U$42276 ( \42619 , \42618 );
nand \U$42277 ( \42620 , \42588 , \42619 );
not \U$42278 ( \42621 , \42598 );
not \U$42279 ( \42622 , \42614 );
or \U$42280 ( \42623 , \42621 , \42622 );
or \U$42281 ( \42624 , \42614 , \42598 );
nand \U$42282 ( \42625 , \42623 , \42624 );
and \U$42283 ( \42626 , \38475 , \38726 );
or \U$42284 ( \42627 , \38409 , \42626 );
or \U$42285 ( \42628 , \38726 , \38475 );
nand \U$42286 ( \42629 , \42627 , \42628 );
or \U$42287 ( \42630 , \42625 , \42629 );
not \U$42288 ( \42631 , \37760 );
not \U$42289 ( \42632 , \37757 );
not \U$42290 ( \42633 , \37732 );
or \U$42291 ( \42634 , \42632 , \42633 );
or \U$42292 ( \42635 , \37757 , \37732 );
nand \U$42293 ( \42636 , \42634 , \42635 );
not \U$42294 ( \42637 , \42636 );
or \U$42295 ( \42638 , \42631 , \42637 );
or \U$42296 ( \42639 , \42636 , \37760 );
nand \U$42297 ( \42640 , \42638 , \42639 );
xor \U$42298 ( \42641 , \42569 , \42577 );
and \U$42299 ( \42642 , \42641 , \42583 );
and \U$42300 ( \42643 , \42569 , \42577 );
or \U$42301 ( \42644 , \42642 , \42643 );
nand \U$42302 ( \42645 , \42640 , \42644 );
and \U$42303 ( \42646 , \42585 , \42620 , \42630 , \42645 );
nand \U$42304 ( \42647 , \37765 , \42448 , \42646 );
not \U$42305 ( \42648 , \42647 );
not \U$42306 ( \42649 , \8028 );
not \U$42307 ( \42650 , \36136 );
or \U$42308 ( \42651 , \42649 , \42650 );
nand \U$42309 ( \42652 , \34207 , \9071 );
nand \U$42310 ( \42653 , \42651 , \42652 );
not \U$42311 ( \42654 , \42653 );
not \U$42312 ( \42655 , \34509 );
xor \U$42313 ( \42656 , \34503 , \42655 );
not \U$42314 ( \42657 , \42656 );
not \U$42315 ( \42658 , \5641 );
not \U$42316 ( \42659 , \36702 );
or \U$42317 ( \42660 , \42658 , \42659 );
nand \U$42318 ( \42661 , \34336 , \5653 );
nand \U$42319 ( \42662 , \42660 , \42661 );
not \U$42320 ( \42663 , \42662 );
or \U$42321 ( \42664 , \42657 , \42663 );
or \U$42322 ( \42665 , \42662 , \42656 );
nand \U$42323 ( \42666 , \42664 , \42665 );
not \U$42324 ( \42667 , \42666 );
or \U$42325 ( \42668 , \42654 , \42667 );
not \U$42326 ( \42669 , \42656 );
nand \U$42327 ( \42670 , \42669 , \42662 );
nand \U$42328 ( \42671 , \42668 , \42670 );
not \U$42329 ( \42672 , \42671 );
xor \U$42330 ( \42673 , \34528 , \34516 );
not \U$42331 ( \42674 , \42673 );
not \U$42332 ( \42675 , \34355 );
not \U$42333 ( \42676 , \34361 );
or \U$42334 ( \42677 , \42675 , \42676 );
or \U$42335 ( \42678 , \34361 , \34355 );
nand \U$42336 ( \42679 , \42677 , \42678 );
not \U$42337 ( \42680 , \42679 );
or \U$42338 ( \42681 , \42674 , \42680 );
or \U$42339 ( \42682 , \42679 , \42673 );
nand \U$42340 ( \42683 , \42681 , \42682 );
not \U$42341 ( \42684 , \42683 );
or \U$42342 ( \42685 , \42672 , \42684 );
not \U$42343 ( \42686 , \42673 );
nand \U$42344 ( \42687 , \42679 , \42686 );
nand \U$42345 ( \42688 , \42685 , \42687 );
xnor \U$42346 ( \42689 , \34611 , \34628 );
or \U$42347 ( \42690 , \42688 , \42689 );
not \U$42348 ( \42691 , \42690 );
not \U$42349 ( \42692 , \9670 );
not \U$42350 ( \42693 , \36085 );
or \U$42351 ( \42694 , \42692 , \42693 );
not \U$42352 ( \42695 , \34146 );
or \U$42353 ( \42696 , \42695 , \10486 );
nand \U$42354 ( \42697 , \42694 , \42696 );
not \U$42355 ( \42698 , \42697 );
not \U$42356 ( \42699 , \9294 );
not \U$42357 ( \42700 , \36786 );
or \U$42358 ( \42701 , \42699 , \42700 );
nand \U$42359 ( \42702 , \34392 , \9273 );
nand \U$42360 ( \42703 , \42701 , \42702 );
not \U$42361 ( \42704 , \42703 );
not \U$42362 ( \42705 , \8819 );
not \U$42363 ( \42706 , \36069 );
or \U$42364 ( \42707 , \42705 , \42706 );
nand \U$42365 ( \42708 , \34162 , \8802 );
nand \U$42366 ( \42709 , \42707 , \42708 );
not \U$42367 ( \42710 , \42709 );
not \U$42368 ( \42711 , \42710 );
or \U$42369 ( \42712 , \42704 , \42711 );
or \U$42370 ( \42713 , \42710 , \42703 );
nand \U$42371 ( \42714 , \42712 , \42713 );
not \U$42372 ( \42715 , \42714 );
or \U$42373 ( \42716 , \42698 , \42715 );
nand \U$42374 ( \42717 , \42709 , \42703 );
nand \U$42375 ( \42718 , \42716 , \42717 );
not \U$42376 ( \42719 , \42718 );
not \U$42377 ( \42720 , \6282 );
not \U$42378 ( \42721 , \36726 );
or \U$42379 ( \42722 , \42720 , \42721 );
nand \U$42380 ( \42723 , \34353 , \6285 );
nand \U$42381 ( \42724 , \42722 , \42723 );
not \U$42382 ( \42725 , \42724 );
not \U$42383 ( \42726 , \7338 );
not \U$42384 ( \42727 , \34526 );
or \U$42385 ( \42728 , \42726 , \42727 );
nand \U$42386 ( \42729 , \36712 , \7325 );
nand \U$42387 ( \42730 , \42728 , \42729 );
not \U$42388 ( \42731 , \42730 );
not \U$42389 ( \42732 , \42731 );
or \U$42390 ( \42733 , \42725 , \42732 );
not \U$42391 ( \42734 , \42724 );
nand \U$42392 ( \42735 , \42734 , \42730 );
nand \U$42393 ( \42736 , \42733 , \42735 );
not \U$42394 ( \42737 , \42736 );
not \U$42395 ( \42738 , \24627 );
not \U$42396 ( \42739 , \36800 );
or \U$42397 ( \42740 , \42738 , \42739 );
nand \U$42398 ( \42741 , \34375 , \8752 );
nand \U$42399 ( \42742 , \42740 , \42741 );
not \U$42400 ( \42743 , \42742 );
or \U$42401 ( \42744 , \42737 , \42743 );
nand \U$42402 ( \42745 , \42730 , \42724 );
nand \U$42403 ( \42746 , \42744 , \42745 );
not \U$42404 ( \42747 , \42746 );
not \U$42405 ( \42748 , \13020 );
not \U$42406 ( \42749 , \36683 );
or \U$42407 ( \42750 , \42748 , \42749 );
nand \U$42408 ( \42751 , \34277 , \22618 );
nand \U$42409 ( \42752 , \42750 , \42751 );
not \U$42410 ( \42753 , \36774 );
not \U$42411 ( \42754 , \36768 );
or \U$42412 ( \42755 , \42753 , \42754 );
nand \U$42413 ( \42756 , \36757 , \36763 );
nand \U$42414 ( \42757 , \42755 , \42756 );
not \U$42415 ( \42758 , \42757 );
not \U$42416 ( \42759 , \42758 );
not \U$42417 ( \42760 , \9196 );
not \U$42418 ( \42761 , \36663 );
or \U$42419 ( \42762 , \42760 , \42761 );
nand \U$42420 ( \42763 , \34179 , \9214 );
nand \U$42421 ( \42764 , \42762 , \42763 );
not \U$42422 ( \42765 , \42764 );
or \U$42423 ( \42766 , \42759 , \42765 );
or \U$42424 ( \42767 , \42764 , \42758 );
nand \U$42425 ( \42768 , \42766 , \42767 );
nand \U$42426 ( \42769 , \42752 , \42768 );
nand \U$42427 ( \42770 , \42764 , \42757 );
and \U$42428 ( \42771 , \42769 , \42770 );
not \U$42429 ( \42772 , \42771 );
or \U$42430 ( \42773 , \42747 , \42772 );
not \U$42431 ( \42774 , \42770 );
not \U$42432 ( \42775 , \42769 );
or \U$42433 ( \42776 , \42774 , \42775 );
not \U$42434 ( \42777 , \42746 );
nand \U$42435 ( \42778 , \42776 , \42777 );
nand \U$42436 ( \42779 , \42773 , \42778 );
not \U$42437 ( \42780 , \42779 );
or \U$42438 ( \42781 , \42719 , \42780 );
not \U$42439 ( \42782 , \42770 );
not \U$42440 ( \42783 , \42769 );
or \U$42441 ( \42784 , \42782 , \42783 );
nand \U$42442 ( \42785 , \42784 , \42746 );
nand \U$42443 ( \42786 , \42781 , \42785 );
not \U$42444 ( \42787 , \42786 );
or \U$42445 ( \42788 , \42691 , \42787 );
nand \U$42446 ( \42789 , \42688 , \42689 );
nand \U$42447 ( \42790 , \42788 , \42789 );
not \U$42448 ( \42791 , \42790 );
and \U$42449 ( \42792 , \34438 , \34293 );
not \U$42450 ( \42793 , \34438 );
and \U$42451 ( \42794 , \42793 , \34286 );
or \U$42452 ( \42795 , \42792 , \42794 );
and \U$42453 ( \42796 , \42795 , \34289 );
not \U$42454 ( \42797 , \42795 );
and \U$42455 ( \42798 , \42797 , \34290 );
nor \U$42456 ( \42799 , \42796 , \42798 );
not \U$42457 ( \42800 , \42799 );
not \U$42458 ( \42801 , \42800 );
or \U$42459 ( \42802 , \42791 , \42801 );
or \U$42460 ( \42803 , \42800 , \42790 );
not \U$42461 ( \42804 , \34363 );
not \U$42462 ( \42805 , \34368 );
or \U$42463 ( \42806 , \42804 , \42805 );
not \U$42464 ( \42807 , \34363 );
nand \U$42465 ( \42808 , \42807 , \34328 );
nand \U$42466 ( \42809 , \42806 , \42808 );
xnor \U$42467 ( \42810 , \42809 , \34436 );
xor \U$42468 ( \42811 , \34191 , \34196 );
xor \U$42469 ( \42812 , \42811 , \34284 );
nand \U$42470 ( \42813 , \42810 , \42812 );
not \U$42471 ( \42814 , \42813 );
not \U$42472 ( \42815 , \34263 );
not \U$42473 ( \42816 , \34279 );
not \U$42474 ( \42817 , \42816 );
or \U$42475 ( \42818 , \42815 , \42817 );
not \U$42476 ( \42819 , \34263 );
nand \U$42477 ( \42820 , \42819 , \34279 );
nand \U$42478 ( \42821 , \42818 , \42820 );
not \U$42479 ( \42822 , \42821 );
xnor \U$42480 ( \42823 , \34432 , \34379 );
nand \U$42481 ( \42824 , \42822 , \42823 );
not \U$42482 ( \42825 , \42824 );
not \U$42483 ( \42826 , \18508 );
not \U$42484 ( \42827 , \36103 );
or \U$42485 ( \42828 , \42826 , \42827 );
and \U$42486 ( \42829 , RI9873288_184, \33926 );
not \U$42487 ( \42830 , RI9873288_184);
and \U$42488 ( \42831 , \42830 , \24185 );
or \U$42489 ( \42832 , \42829 , \42831 );
nand \U$42490 ( \42833 , \42832 , \17528 );
nand \U$42491 ( \42834 , \42828 , \42833 );
not \U$42492 ( \42835 , \42834 );
not \U$42493 ( \42836 , \9937 );
not \U$42494 ( \42837 , \14132 );
not \U$42495 ( \42838 , \8082 );
or \U$42496 ( \42839 , \42837 , \42838 );
nand \U$42497 ( \42840 , \8948 , RI9873030_179);
nand \U$42498 ( \42841 , \42839 , \42840 );
not \U$42499 ( \42842 , \42841 );
or \U$42500 ( \42843 , \42836 , \42842 );
nand \U$42501 ( \42844 , \36674 , \18672 );
nand \U$42502 ( \42845 , \42843 , \42844 );
not \U$42503 ( \42846 , \13477 );
not \U$42504 ( \42847 , \36113 );
or \U$42505 ( \42848 , \42846 , \42847 );
and \U$42506 ( \42849 , \6481 , \28789 );
not \U$42507 ( \42850 , \6481 );
and \U$42508 ( \42851 , \42850 , RI9873210_183);
nor \U$42509 ( \42852 , \42849 , \42851 );
nand \U$42510 ( \42853 , \42852 , \22670 );
nand \U$42511 ( \42854 , \42848 , \42853 );
xor \U$42512 ( \42855 , \42845 , \42854 );
not \U$42513 ( \42856 , \42855 );
or \U$42514 ( \42857 , \42835 , \42856 );
nand \U$42515 ( \42858 , \42854 , \42845 );
nand \U$42516 ( \42859 , \42857 , \42858 );
not \U$42517 ( \42860 , \42859 );
or \U$42518 ( \42861 , \42825 , \42860 );
not \U$42519 ( \42862 , \42823 );
nand \U$42520 ( \42863 , \42862 , \42821 );
nand \U$42521 ( \42864 , \42861 , \42863 );
not \U$42522 ( \42865 , \42864 );
or \U$42523 ( \42866 , \42814 , \42865 );
nor \U$42524 ( \42867 , \42812 , \42810 );
not \U$42525 ( \42868 , \42867 );
nand \U$42526 ( \42869 , \42866 , \42868 );
nand \U$42527 ( \42870 , \42803 , \42869 );
nand \U$42528 ( \42871 , \42802 , \42870 );
not \U$42529 ( \42872 , \42871 );
xor \U$42530 ( \42873 , \33775 , \33777 );
xor \U$42531 ( \42874 , \42873 , \33832 );
xor \U$42532 ( \42875 , \34725 , \34746 );
not \U$42533 ( \42876 , \17528 );
not \U$42534 ( \42877 , \34660 );
or \U$42535 ( \42878 , \42876 , \42877 );
nand \U$42536 ( \42879 , \42832 , \17544 );
nand \U$42537 ( \42880 , \42878 , \42879 );
not \U$42538 ( \42881 , \9937 );
not \U$42539 ( \42882 , \34641 );
or \U$42540 ( \42883 , \42881 , \42882 );
nand \U$42541 ( \42884 , \42841 , \9952 );
nand \U$42542 ( \42885 , \42883 , \42884 );
xor \U$42543 ( \42886 , \42880 , \42885 );
not \U$42544 ( \42887 , \19036 );
not \U$42545 ( \42888 , RI98734e0_189);
not \U$42546 ( \42889 , \5595 );
or \U$42547 ( \42890 , \42888 , \42889 );
or \U$42548 ( \42891 , \5595 , RI98734e0_189);
nand \U$42549 ( \42892 , \42890 , \42891 );
not \U$42550 ( \42893 , \42892 );
or \U$42551 ( \42894 , \42887 , \42893 );
nand \U$42552 ( \42895 , \34607 , \19046 );
nand \U$42553 ( \42896 , \42894 , \42895 );
and \U$42554 ( \42897 , \42886 , \42896 );
and \U$42555 ( \42898 , \42880 , \42885 );
or \U$42556 ( \42899 , \42897 , \42898 );
not \U$42557 ( \42900 , \34574 );
not \U$42558 ( \42901 , \34569 );
or \U$42559 ( \42902 , \42900 , \42901 );
or \U$42560 ( \42903 , \34569 , \34574 );
nand \U$42561 ( \42904 , \42902 , \42903 );
xor \U$42562 ( \42905 , \42904 , \34581 );
nor \U$42563 ( \42906 , \42899 , \42905 );
buf \U$42564 ( \42907 , \34664 );
not \U$42565 ( \42908 , \42907 );
xor \U$42566 ( \42909 , \34652 , \34646 );
not \U$42567 ( \42910 , \42909 );
or \U$42568 ( \42911 , \42908 , \42910 );
or \U$42569 ( \42912 , \42909 , \42907 );
nand \U$42570 ( \42913 , \42911 , \42912 );
or \U$42571 ( \42914 , \42906 , \42913 );
nand \U$42572 ( \42915 , \42899 , \42905 );
nand \U$42573 ( \42916 , \42914 , \42915 );
xor \U$42574 ( \42917 , \42875 , \42916 );
xor \U$42575 ( \42918 , \34634 , \34673 );
and \U$42576 ( \42919 , \42917 , \42918 );
and \U$42577 ( \42920 , \42875 , \42916 );
or \U$42578 ( \42921 , \42919 , \42920 );
xor \U$42579 ( \42922 , \42874 , \42921 );
xor \U$42580 ( \42923 , \34750 , \34752 );
xor \U$42581 ( \42924 , \42923 , \34755 );
xor \U$42582 ( \42925 , \42922 , \42924 );
not \U$42583 ( \42926 , \42925 );
or \U$42584 ( \42927 , \42872 , \42926 );
not \U$42585 ( \42928 , \36730 );
not \U$42586 ( \42929 , \36720 );
or \U$42587 ( \42930 , \42928 , \42929 );
not \U$42588 ( \42931 , \36705 );
nand \U$42589 ( \42932 , \42931 , \36716 );
nand \U$42590 ( \42933 , \42930 , \42932 );
not \U$42591 ( \42934 , \42933 );
not \U$42592 ( \42935 , \36151 );
not \U$42593 ( \42936 , \36140 );
or \U$42594 ( \42937 , \42935 , \42936 );
nand \U$42595 ( \42938 , \36145 , \36150 );
nand \U$42596 ( \42939 , \42937 , \42938 );
not \U$42597 ( \42940 , \42939 );
nand \U$42598 ( \42941 , \42934 , \42940 );
not \U$42599 ( \42942 , \42941 );
not \U$42600 ( \42943 , \42939 );
not \U$42601 ( \42944 , \42933 );
or \U$42602 ( \42945 , \42943 , \42944 );
not \U$42603 ( \42946 , \17371 );
not \U$42604 ( \42947 , \36154 );
or \U$42605 ( \42948 , \42946 , \42947 );
and \U$42606 ( \42949 , \4711 , \17539 );
not \U$42607 ( \42950 , \4711 );
and \U$42608 ( \42951 , \42950 , RI98733f0_187);
nor \U$42609 ( \42952 , \42949 , \42951 );
nand \U$42610 ( \42953 , \42952 , \19282 );
nand \U$42611 ( \42954 , \42948 , \42953 );
not \U$42612 ( \42955 , \42954 );
nand \U$42613 ( \42956 , \42945 , \42955 );
not \U$42614 ( \42957 , \42956 );
or \U$42615 ( \42958 , \42942 , \42957 );
xor \U$42616 ( \42959 , \34164 , \34148 );
and \U$42617 ( \42960 , \42959 , \34181 );
not \U$42618 ( \42961 , \42959 );
not \U$42619 ( \42962 , \34181 );
and \U$42620 ( \42963 , \42961 , \42962 );
nor \U$42621 ( \42964 , \42960 , \42963 );
not \U$42622 ( \42965 , \42964 );
nand \U$42623 ( \42966 , \42958 , \42965 );
not \U$42624 ( \42967 , \42966 );
xor \U$42625 ( \42968 , \34227 , \34241 );
xor \U$42626 ( \42969 , \42968 , \34256 );
not \U$42627 ( \42970 , \18615 );
not \U$42628 ( \42971 , \36126 );
or \U$42629 ( \42972 , \42970 , \42971 );
not \U$42630 ( \42973 , \18239 );
not \U$42631 ( \42974 , \3537 );
or \U$42632 ( \42975 , \42973 , \42974 );
or \U$42633 ( \42976 , \3537 , \18239 );
nand \U$42634 ( \42977 , \42975 , \42976 );
nand \U$42635 ( \42978 , \42977 , RI9873648_192);
nand \U$42636 ( \42979 , \42972 , \42978 );
xor \U$42637 ( \42980 , \42969 , \42979 );
not \U$42638 ( \42981 , \20147 );
not \U$42639 ( \42982 , \42892 );
or \U$42640 ( \42983 , \42981 , \42982 );
nand \U$42641 ( \42984 , \36165 , \19243 );
nand \U$42642 ( \42985 , \42983 , \42984 );
and \U$42643 ( \42986 , \42980 , \42985 );
and \U$42644 ( \42987 , \42969 , \42979 );
nor \U$42645 ( \42988 , \42986 , \42987 );
or \U$42646 ( \42989 , \42967 , \42988 );
and \U$42647 ( \42990 , \42956 , \42941 , \42964 );
not \U$42648 ( \42991 , \42990 );
nand \U$42649 ( \42992 , \42989 , \42991 );
not \U$42650 ( \42993 , \42906 );
nand \U$42651 ( \42994 , \42993 , \42915 );
not \U$42652 ( \42995 , \42994 );
not \U$42653 ( \42996 , \42913 );
and \U$42654 ( \42997 , \42995 , \42996 );
and \U$42655 ( \42998 , \42994 , \42913 );
nor \U$42656 ( \42999 , \42997 , \42998 );
xor \U$42657 ( \43000 , \42992 , \42999 );
xor \U$42658 ( \43001 , \34710 , \34706 );
xor \U$42659 ( \43002 , \43001 , \34716 );
not \U$42660 ( \43003 , \13484 );
not \U$42661 ( \43004 , \34620 );
or \U$42662 ( \43005 , \43003 , \43004 );
nand \U$42663 ( \43006 , \42852 , \13476 );
nand \U$42664 ( \43007 , \43005 , \43006 );
not \U$42665 ( \43008 , \43007 );
not \U$42666 ( \43009 , RI9873648_192);
not \U$42667 ( \43010 , \34541 );
or \U$42668 ( \43011 , \43009 , \43010 );
nand \U$42669 ( \43012 , \42977 , \18545 );
nand \U$42670 ( \43013 , \43011 , \43012 );
not \U$42671 ( \43014 , \43013 );
or \U$42672 ( \43015 , \43008 , \43014 );
xor \U$42673 ( \43016 , \43013 , \43007 );
not \U$42674 ( \43017 , \17263 );
not \U$42675 ( \43018 , \34487 );
or \U$42676 ( \43019 , \43017 , \43018 );
nand \U$42677 ( \43020 , \42952 , \17252 );
nand \U$42678 ( \43021 , \43019 , \43020 );
nand \U$42679 ( \43022 , \43016 , \43021 );
nand \U$42680 ( \43023 , \43015 , \43022 );
xor \U$42681 ( \43024 , \43002 , \43023 );
xor \U$42682 ( \43025 , \34544 , \34489 );
xnor \U$42683 ( \43026 , \43024 , \43025 );
and \U$42684 ( \43027 , \43000 , \43026 );
and \U$42685 ( \43028 , \42992 , \42999 );
or \U$42686 ( \43029 , \43027 , \43028 );
xor \U$42687 ( \43030 , \42875 , \42916 );
xor \U$42688 ( \43031 , \43030 , \42918 );
or \U$42689 ( \43032 , \43029 , \43031 );
xor \U$42690 ( \43033 , \34599 , \34592 );
xor \U$42691 ( \43034 , \33599 , \34594 );
xnor \U$42692 ( \43035 , \43034 , \33607 );
xnor \U$42693 ( \43036 , \43033 , \43035 );
not \U$42694 ( \43037 , \34548 );
and \U$42695 ( \43038 , \34553 , \43037 );
not \U$42696 ( \43039 , \34553 );
and \U$42697 ( \43040 , \43039 , \34548 );
or \U$42698 ( \43041 , \43038 , \43040 );
xor \U$42699 ( \43042 , \43036 , \43041 );
not \U$42700 ( \43043 , \43025 );
not \U$42701 ( \43044 , \43002 );
not \U$42702 ( \43045 , \43023 );
or \U$42703 ( \43046 , \43044 , \43045 );
or \U$42704 ( \43047 , \43023 , \43002 );
nand \U$42705 ( \43048 , \43046 , \43047 );
not \U$42706 ( \43049 , \43048 );
or \U$42707 ( \43050 , \43043 , \43049 );
not \U$42708 ( \43051 , \43002 );
nand \U$42709 ( \43052 , \43051 , \43023 );
nand \U$42710 ( \43053 , \43050 , \43052 );
xnor \U$42711 ( \43054 , \43042 , \43053 );
and \U$42712 ( \43055 , \43032 , \43054 );
and \U$42713 ( \43056 , \43031 , \43029 );
nor \U$42714 ( \43057 , \43055 , \43056 );
nand \U$42715 ( \43058 , \42927 , \43057 );
not \U$42716 ( \43059 , \42871 );
not \U$42717 ( \43060 , \42925 );
nand \U$42718 ( \43061 , \43059 , \43060 );
and \U$42719 ( \43062 , \43058 , \43061 );
xor \U$42720 ( \43063 , \34686 , \34467 );
xor \U$42721 ( \43064 , \43063 , \34474 );
and \U$42722 ( \43065 , \43062 , \43064 );
not \U$42723 ( \43066 , \43062 );
not \U$42724 ( \43067 , \43064 );
and \U$42725 ( \43068 , \43066 , \43067 );
nor \U$42726 ( \43069 , \43065 , \43068 );
not \U$42727 ( \43070 , \43069 );
not \U$42728 ( \43071 , \43070 );
xor \U$42729 ( \43072 , \42874 , \42921 );
and \U$42730 ( \43073 , \43072 , \42924 );
and \U$42731 ( \43074 , \42874 , \42921 );
or \U$42732 ( \43075 , \43073 , \43074 );
and \U$42733 ( \43076 , \34463 , \34440 );
not \U$42734 ( \43077 , \34463 );
not \U$42735 ( \43078 , \34440 );
and \U$42736 ( \43079 , \43077 , \43078 );
nor \U$42737 ( \43080 , \43076 , \43079 );
not \U$42738 ( \43081 , \43036 );
not \U$42739 ( \43082 , \43081 );
not \U$42740 ( \43083 , \43041 );
or \U$42741 ( \43084 , \43082 , \43083 );
or \U$42742 ( \43085 , \43041 , \43081 );
nand \U$42743 ( \43086 , \43085 , \43053 );
nand \U$42744 ( \43087 , \43084 , \43086 );
xor \U$42745 ( \43088 , \43080 , \43087 );
not \U$42746 ( \43089 , \34563 );
not \U$42747 ( \43090 , \43089 );
not \U$42748 ( \43091 , \34679 );
or \U$42749 ( \43092 , \43090 , \43091 );
or \U$42750 ( \43093 , \34679 , \43089 );
nand \U$42751 ( \43094 , \43092 , \43093 );
and \U$42752 ( \43095 , \43088 , \43094 );
and \U$42753 ( \43096 , \43080 , \43087 );
or \U$42754 ( \43097 , \43095 , \43096 );
xor \U$42755 ( \43098 , \43075 , \43097 );
xnor \U$42756 ( \43099 , \34699 , \34771 );
xor \U$42757 ( \43100 , \43098 , \43099 );
not \U$42758 ( \43101 , \43100 );
not \U$42759 ( \43102 , \43101 );
or \U$42760 ( \43103 , \43071 , \43102 );
nand \U$42761 ( \43104 , \43100 , \43069 );
nand \U$42762 ( \43105 , \43103 , \43104 );
xor \U$42763 ( \43106 , \42871 , \43060 );
xor \U$42764 ( \43107 , \43106 , \43057 );
not \U$42765 ( \43108 , \43107 );
not \U$42766 ( \43109 , \43108 );
xor \U$42767 ( \43110 , \43080 , \43087 );
xor \U$42768 ( \43111 , \43110 , \43094 );
not \U$42769 ( \43112 , \43111 );
xor \U$42770 ( \43113 , \42790 , \42799 );
xor \U$42771 ( \43114 , \43113 , \42869 );
not \U$42772 ( \43115 , \43114 );
xor \U$42773 ( \43116 , \42688 , \42689 );
xnor \U$42774 ( \43117 , \43116 , \42786 );
xor \U$42775 ( \43118 , \42880 , \42885 );
xor \U$42776 ( \43119 , \43118 , \42896 );
xor \U$42777 ( \43120 , \43016 , \43021 );
xor \U$42778 ( \43121 , \43119 , \43120 );
not \U$42779 ( \43122 , \36073 );
not \U$42780 ( \43123 , \36093 );
or \U$42781 ( \43124 , \43122 , \43123 );
not \U$42782 ( \43125 , \36079 );
nand \U$42783 ( \43126 , \43125 , \36089 );
nand \U$42784 ( \43127 , \43124 , \43126 );
not \U$42785 ( \43128 , \43127 );
xor \U$42786 ( \43129 , \42666 , \42653 );
and \U$42787 ( \43130 , \42736 , \42742 );
not \U$42788 ( \43131 , \42736 );
not \U$42789 ( \43132 , \42742 );
and \U$42790 ( \43133 , \43131 , \43132 );
nor \U$42791 ( \43134 , \43130 , \43133 );
xor \U$42792 ( \43135 , \43129 , \43134 );
not \U$42793 ( \43136 , \43135 );
or \U$42794 ( \43137 , \43128 , \43136 );
nand \U$42795 ( \43138 , \43134 , \43129 );
nand \U$42796 ( \43139 , \43137 , \43138 );
and \U$42797 ( \43140 , \43121 , \43139 );
and \U$42798 ( \43141 , \43119 , \43120 );
or \U$42799 ( \43142 , \43140 , \43141 );
not \U$42800 ( \43143 , \43142 );
xor \U$42801 ( \43144 , \43117 , \43143 );
xor \U$42802 ( \43145 , \42671 , \42686 );
xnor \U$42803 ( \43146 , \43145 , \42679 );
not \U$42804 ( \43147 , \42779 );
not \U$42805 ( \43148 , \42718 );
not \U$42806 ( \43149 , \43148 );
and \U$42807 ( \43150 , \43147 , \43149 );
and \U$42808 ( \43151 , \42779 , \43148 );
nor \U$42809 ( \43152 , \43150 , \43151 );
xor \U$42810 ( \43153 , \43146 , \43152 );
xor \U$42811 ( \43154 , \36107 , \36117 );
and \U$42812 ( \43155 , \43154 , \36128 );
and \U$42813 ( \43156 , \36107 , \36117 );
or \U$42814 ( \43157 , \43155 , \43156 );
xor \U$42815 ( \43158 , \42752 , \42768 );
xor \U$42816 ( \43159 , \42697 , \42714 );
xor \U$42817 ( \43160 , \43158 , \43159 );
and \U$42818 ( \43161 , \43157 , \43160 );
and \U$42819 ( \43162 , \43158 , \43159 );
nor \U$42820 ( \43163 , \43161 , \43162 );
and \U$42821 ( \43164 , \43153 , \43163 );
and \U$42822 ( \43165 , \43146 , \43152 );
or \U$42823 ( \43166 , \43164 , \43165 );
and \U$42824 ( \43167 , \43144 , \43166 );
and \U$42825 ( \43168 , \43117 , \43143 );
or \U$42826 ( \43169 , \43167 , \43168 );
not \U$42827 ( \43170 , \43169 );
or \U$42828 ( \43171 , \43115 , \43170 );
not \U$42829 ( \43172 , \42867 );
nand \U$42830 ( \43173 , \43172 , \42813 );
not \U$42831 ( \43174 , \43173 );
xor \U$42832 ( \43175 , \42864 , \43174 );
not \U$42833 ( \43176 , \42821 );
not \U$42834 ( \43177 , \42823 );
or \U$42835 ( \43178 , \43176 , \43177 );
or \U$42836 ( \43179 , \42823 , \42821 );
nand \U$42837 ( \43180 , \43178 , \43179 );
not \U$42838 ( \43181 , \43180 );
not \U$42839 ( \43182 , \43181 );
not \U$42840 ( \43183 , \42859 );
not \U$42841 ( \43184 , \43183 );
or \U$42842 ( \43185 , \43182 , \43184 );
nand \U$42843 ( \43186 , \43180 , \42859 );
nand \U$42844 ( \43187 , \43185 , \43186 );
not \U$42845 ( \43188 , \43187 );
xor \U$42846 ( \43189 , \42834 , \42845 );
xor \U$42847 ( \43190 , \43189 , \42854 );
not \U$42848 ( \43191 , \43190 );
not \U$42849 ( \43192 , \36804 );
not \U$42850 ( \43193 , \36794 );
or \U$42851 ( \43194 , \43192 , \43193 );
not \U$42852 ( \43195 , \36779 );
nand \U$42853 ( \43196 , \43195 , \36790 );
nand \U$42854 ( \43197 , \43194 , \43196 );
not \U$42855 ( \43198 , \36687 );
not \U$42856 ( \43199 , \36677 );
or \U$42857 ( \43200 , \43198 , \43199 );
nand \U$42858 ( \43201 , \36676 , \36667 );
nand \U$42859 ( \43202 , \43200 , \43201 );
and \U$42860 ( \43203 , \43197 , \43202 );
not \U$42861 ( \43204 , \43197 );
not \U$42862 ( \43205 , \43202 );
and \U$42863 ( \43206 , \43204 , \43205 );
nor \U$42864 ( \43207 , \43203 , \43206 );
not \U$42865 ( \43208 , \43207 );
or \U$42866 ( \43209 , \43191 , \43208 );
nand \U$42867 ( \43210 , \43202 , \43197 );
nand \U$42868 ( \43211 , \43209 , \43210 );
not \U$42869 ( \43212 , \43211 );
not \U$42870 ( \43213 , \43212 );
or \U$42871 ( \43214 , \43188 , \43213 );
not \U$42872 ( \43215 , \42990 );
nand \U$42873 ( \43216 , \43215 , \42966 );
xor \U$42874 ( \43217 , \43216 , \42988 );
nand \U$42875 ( \43218 , \43214 , \43217 );
not \U$42876 ( \43219 , \43187 );
nand \U$42877 ( \43220 , \43219 , \43211 );
nand \U$42878 ( \43221 , \43218 , \43220 );
xor \U$42879 ( \43222 , \43175 , \43221 );
xor \U$42880 ( \43223 , \42992 , \42999 );
xor \U$42881 ( \43224 , \43223 , \43026 );
and \U$42882 ( \43225 , \43222 , \43224 );
and \U$42883 ( \43226 , \43175 , \43221 );
or \U$42884 ( \43227 , \43225 , \43226 );
nand \U$42885 ( \43228 , \43171 , \43227 );
or \U$42886 ( \43229 , \43169 , \43114 );
nand \U$42887 ( \43230 , \43228 , \43229 );
not \U$42888 ( \43231 , \43230 );
not \U$42889 ( \43232 , \43231 );
or \U$42890 ( \43233 , \43112 , \43232 );
or \U$42891 ( \43234 , \43231 , \43111 );
nand \U$42892 ( \43235 , \43233 , \43234 );
not \U$42893 ( \43236 , \43235 );
or \U$42894 ( \43237 , \43109 , \43236 );
not \U$42895 ( \43238 , \43111 );
nand \U$42896 ( \43239 , \43238 , \43231 );
nand \U$42897 ( \43240 , \43237 , \43239 );
nand \U$42898 ( \43241 , \43105 , \43240 );
not \U$42899 ( \43242 , \33738 );
not \U$42900 ( \43243 , \33759 );
or \U$42901 ( \43244 , \43242 , \43243 );
nand \U$42902 ( \43245 , \43244 , \33766 );
and \U$42903 ( \43246 , \43245 , \33763 );
not \U$42904 ( \43247 , \43245 );
not \U$42905 ( \43248 , \33763 );
and \U$42906 ( \43249 , \43247 , \43248 );
nor \U$42907 ( \43250 , \43246 , \43249 );
not \U$42908 ( \43251 , \43250 );
xor \U$42909 ( \43252 , \34688 , \34691 );
xor \U$42910 ( \43253 , \43252 , \34775 );
not \U$42911 ( \43254 , \43253 );
or \U$42912 ( \43255 , \43251 , \43254 );
not \U$42913 ( \43256 , \43075 );
not \U$42914 ( \43257 , \43099 );
or \U$42915 ( \43258 , \43256 , \43257 );
or \U$42916 ( \43259 , \43099 , \43075 );
nand \U$42917 ( \43260 , \43259 , \43097 );
nand \U$42918 ( \43261 , \43258 , \43260 );
nand \U$42919 ( \43262 , \43255 , \43261 );
not \U$42920 ( \43263 , \43253 );
not \U$42921 ( \43264 , \43250 );
nand \U$42922 ( \43265 , \43263 , \43264 );
nand \U$42923 ( \43266 , \43262 , \43265 );
not \U$42924 ( \43267 , \43266 );
xor \U$42925 ( \43268 , \34783 , \34777 );
xnor \U$42926 ( \43269 , \43268 , \34791 );
nand \U$42927 ( \43270 , \43267 , \43269 );
not \U$42928 ( \43271 , \43261 );
not \U$42929 ( \43272 , \43250 );
or \U$42930 ( \43273 , \43271 , \43272 );
or \U$42931 ( \43274 , \43261 , \43250 );
nand \U$42932 ( \43275 , \43273 , \43274 );
and \U$42933 ( \43276 , \43275 , \43253 );
not \U$42934 ( \43277 , \43275 );
and \U$42935 ( \43278 , \43277 , \43263 );
nor \U$42936 ( \43279 , \43276 , \43278 );
not \U$42937 ( \43280 , \43069 );
not \U$42938 ( \43281 , \43101 );
or \U$42939 ( \43282 , \43280 , \43281 );
not \U$42940 ( \43283 , \43061 );
not \U$42941 ( \43284 , \43058 );
or \U$42942 ( \43285 , \43283 , \43284 );
nand \U$42943 ( \43286 , \43285 , \43067 );
nand \U$42944 ( \43287 , \43282 , \43286 );
nand \U$42945 ( \43288 , \43279 , \43287 );
and \U$42946 ( \43289 , \43235 , \43107 );
not \U$42947 ( \43290 , \43235 );
and \U$42948 ( \43291 , \43290 , \43108 );
or \U$42949 ( \43292 , \43289 , \43291 );
xor \U$42950 ( \43293 , \43169 , \43114 );
xnor \U$42951 ( \43294 , \43293 , \43227 );
not \U$42952 ( \43295 , \43294 );
xor \U$42953 ( \43296 , \43119 , \43120 );
xor \U$42954 ( \43297 , \43296 , \43139 );
not \U$42955 ( \43298 , \36753 );
not \U$42956 ( \43299 , \36817 );
or \U$42957 ( \43300 , \43298 , \43299 );
nand \U$42958 ( \43301 , \36812 , \36806 );
nand \U$42959 ( \43302 , \43300 , \43301 );
not \U$42960 ( \43303 , \43302 );
not \U$42961 ( \43304 , \36649 );
not \U$42962 ( \43305 , \43304 );
not \U$42963 ( \43306 , \36654 );
or \U$42964 ( \43307 , \43305 , \43306 );
nand \U$42965 ( \43308 , \43307 , \36688 );
xor \U$42966 ( \43309 , \42940 , \42954 );
xnor \U$42967 ( \43310 , \43309 , \42934 );
nand \U$42968 ( \43311 , \36653 , \36649 );
nand \U$42969 ( \43312 , \43308 , \43310 , \43311 );
not \U$42970 ( \43313 , \43312 );
or \U$42971 ( \43314 , \43303 , \43313 );
not \U$42972 ( \43315 , \43310 );
nand \U$42973 ( \43316 , \43308 , \43311 );
nand \U$42974 ( \43317 , \43315 , \43316 );
nand \U$42975 ( \43318 , \43314 , \43317 );
xor \U$42976 ( \43319 , \43297 , \43318 );
not \U$42977 ( \43320 , \42985 );
and \U$42978 ( \43321 , \42980 , \43320 );
not \U$42979 ( \43322 , \42980 );
and \U$42980 ( \43323 , \43322 , \42985 );
or \U$42981 ( \43324 , \43321 , \43323 );
not \U$42982 ( \43325 , \43324 );
not \U$42983 ( \43326 , \36735 );
not \U$42984 ( \43327 , \36698 );
or \U$42985 ( \43328 , \43326 , \43327 );
nand \U$42986 ( \43329 , \43328 , \36744 );
not \U$42987 ( \43330 , \36698 );
nand \U$42988 ( \43331 , \43330 , \36738 );
nand \U$42989 ( \43332 , \43329 , \43331 );
buf \U$42990 ( \43333 , \43332 );
not \U$42991 ( \43334 , \43333 );
buf \U$42992 ( \43335 , \36152 );
xor \U$42993 ( \43336 , \43335 , \36169 );
and \U$42994 ( \43337 , \43336 , \36158 );
and \U$42995 ( \43338 , \43335 , \36169 );
nor \U$42996 ( \43339 , \43337 , \43338 );
not \U$42997 ( \43340 , \43339 );
or \U$42998 ( \43341 , \43334 , \43340 );
or \U$42999 ( \43342 , \43339 , \43333 );
nand \U$43000 ( \43343 , \43341 , \43342 );
not \U$43001 ( \43344 , \43343 );
or \U$43002 ( \43345 , \43325 , \43344 );
not \U$43003 ( \43346 , \43339 );
nand \U$43004 ( \43347 , \43346 , \43333 );
nand \U$43005 ( \43348 , \43345 , \43347 );
and \U$43006 ( \43349 , \43319 , \43348 );
and \U$43007 ( \43350 , \43297 , \43318 );
or \U$43008 ( \43351 , \43349 , \43350 );
not \U$43009 ( \43352 , \43351 );
not \U$43010 ( \43353 , \43352 );
xor \U$43011 ( \43354 , \43117 , \43143 );
xor \U$43012 ( \43355 , \43354 , \43166 );
not \U$43013 ( \43356 , \43355 );
or \U$43014 ( \43357 , \43353 , \43356 );
xor \U$43015 ( \43358 , \43211 , \43187 );
xor \U$43016 ( \43359 , \43358 , \43217 );
not \U$43017 ( \43360 , \43359 );
not \U$43018 ( \43361 , \43360 );
xor \U$43019 ( \43362 , \43146 , \43152 );
xor \U$43020 ( \43363 , \43362 , \43163 );
not \U$43021 ( \43364 , \43363 );
not \U$43022 ( \43365 , \43364 );
or \U$43023 ( \43366 , \43361 , \43365 );
not \U$43024 ( \43367 , \43363 );
not \U$43025 ( \43368 , \43359 );
or \U$43026 ( \43369 , \43367 , \43368 );
xor \U$43027 ( \43370 , \36098 , \36129 );
and \U$43028 ( \43371 , \43370 , \36170 );
and \U$43029 ( \43372 , \36098 , \36129 );
or \U$43030 ( \43373 , \43371 , \43372 );
not \U$43031 ( \43374 , \43373 );
not \U$43032 ( \43375 , \43135 );
not \U$43033 ( \43376 , \43127 );
not \U$43034 ( \43377 , \43376 );
and \U$43035 ( \43378 , \43375 , \43377 );
and \U$43036 ( \43379 , \43135 , \43376 );
nor \U$43037 ( \43380 , \43378 , \43379 );
not \U$43038 ( \43381 , \43380 );
xor \U$43039 ( \43382 , \43207 , \43190 );
not \U$43040 ( \43383 , \43382 );
or \U$43041 ( \43384 , \43381 , \43383 );
or \U$43042 ( \43385 , \43382 , \43380 );
nand \U$43043 ( \43386 , \43384 , \43385 );
not \U$43044 ( \43387 , \43386 );
or \U$43045 ( \43388 , \43374 , \43387 );
not \U$43046 ( \43389 , \43380 );
nand \U$43047 ( \43390 , \43389 , \43382 );
nand \U$43048 ( \43391 , \43388 , \43390 );
nand \U$43049 ( \43392 , \43369 , \43391 );
nand \U$43050 ( \43393 , \43366 , \43392 );
nand \U$43051 ( \43394 , \43357 , \43393 );
not \U$43052 ( \43395 , \43355 );
buf \U$43053 ( \43396 , \43351 );
nand \U$43054 ( \43397 , \43395 , \43396 );
and \U$43055 ( \43398 , \43394 , \43397 );
not \U$43056 ( \43399 , \43054 );
xor \U$43057 ( \43400 , \43031 , \43029 );
not \U$43058 ( \43401 , \43400 );
and \U$43059 ( \43402 , \43399 , \43401 );
and \U$43060 ( \43403 , \43054 , \43400 );
nor \U$43061 ( \43404 , \43402 , \43403 );
not \U$43062 ( \43405 , \43404 );
and \U$43063 ( \43406 , \43398 , \43405 );
not \U$43064 ( \43407 , \43398 );
and \U$43065 ( \43408 , \43407 , \43404 );
nor \U$43066 ( \43409 , \43406 , \43408 );
not \U$43067 ( \43410 , \43409 );
or \U$43068 ( \43411 , \43295 , \43410 );
nand \U$43069 ( \43412 , \43405 , \43394 , \43397 );
nand \U$43070 ( \43413 , \43411 , \43412 );
nand \U$43071 ( \43414 , \43292 , \43413 );
and \U$43072 ( \43415 , \43241 , \43270 , \43288 , \43414 );
not \U$43073 ( \43416 , \36177 );
or \U$43074 ( \43417 , \36171 , \36063 );
not \U$43075 ( \43418 , \43417 );
or \U$43076 ( \43419 , \43416 , \43418 );
nand \U$43077 ( \43420 , \36171 , \36063 );
nand \U$43078 ( \43421 , \43419 , \43420 );
not \U$43079 ( \43422 , \43157 );
and \U$43080 ( \43423 , \43160 , \43422 );
not \U$43081 ( \43424 , \43160 );
and \U$43082 ( \43425 , \43424 , \43157 );
nor \U$43083 ( \43426 , \43423 , \43425 );
not \U$43084 ( \43427 , \43426 );
not \U$43085 ( \43428 , \43427 );
xor \U$43086 ( \43429 , \43332 , \43324 );
xnor \U$43087 ( \43430 , \43429 , \43339 );
not \U$43088 ( \43431 , \43430 );
not \U$43089 ( \43432 , \43431 );
or \U$43090 ( \43433 , \43428 , \43432 );
nand \U$43091 ( \43434 , \43430 , \43426 );
nand \U$43092 ( \43435 , \43433 , \43434 );
xor \U$43093 ( \43436 , \36832 , \36835 );
and \U$43094 ( \43437 , \43436 , \36841 );
and \U$43095 ( \43438 , \36832 , \36835 );
or \U$43096 ( \43439 , \43437 , \43438 );
xnor \U$43097 ( \43440 , \43435 , \43439 );
xor \U$43098 ( \43441 , \43421 , \43440 );
or \U$43099 ( \43442 , \36843 , \36822 );
nand \U$43100 ( \43443 , \43442 , \36845 );
xnor \U$43101 ( \43444 , \43441 , \43443 );
not \U$43102 ( \43445 , \43444 );
not \U$43103 ( \43446 , \36748 );
not \U$43104 ( \43447 , \36821 );
or \U$43105 ( \43448 , \43446 , \43447 );
nand \U$43106 ( \43449 , \43448 , \36747 );
not \U$43107 ( \43450 , \43449 );
not \U$43108 ( \43451 , \43302 );
xnor \U$43109 ( \43452 , \43310 , \43316 );
not \U$43110 ( \43453 , \43452 );
or \U$43111 ( \43454 , \43451 , \43453 );
or \U$43112 ( \43455 , \43452 , \43302 );
nand \U$43113 ( \43456 , \43454 , \43455 );
xor \U$43114 ( \43457 , \43450 , \43456 );
not \U$43115 ( \43458 , \43457 );
xor \U$43116 ( \43459 , \43380 , \43382 );
xnor \U$43117 ( \43460 , \43459 , \43373 );
buf \U$43118 ( \43461 , \43460 );
not \U$43119 ( \43462 , \43461 );
or \U$43120 ( \43463 , \43458 , \43462 );
or \U$43121 ( \43464 , \43461 , \43457 );
nand \U$43122 ( \43465 , \43463 , \43464 );
not \U$43123 ( \43466 , \43465 );
not \U$43124 ( \43467 , \36178 );
not \U$43125 ( \43468 , \35703 );
not \U$43126 ( \43469 , \43468 );
or \U$43127 ( \43470 , \43467 , \43469 );
nand \U$43128 ( \43471 , \43470 , \36058 );
not \U$43129 ( \43472 , \36178 );
nand \U$43130 ( \43473 , \43472 , \35703 );
nand \U$43131 ( \43474 , \43471 , \43473 );
not \U$43132 ( \43475 , \43474 );
or \U$43133 ( \43476 , \43466 , \43475 );
or \U$43134 ( \43477 , \43474 , \43465 );
nand \U$43135 ( \43478 , \43476 , \43477 );
not \U$43136 ( \43479 , \43478 );
or \U$43137 ( \43480 , \43445 , \43479 );
or \U$43138 ( \43481 , \43478 , \43444 );
nand \U$43139 ( \43482 , \43480 , \43481 );
not \U$43140 ( \43483 , \36186 );
not \U$43141 ( \43484 , \36854 );
not \U$43142 ( \43485 , \43484 );
or \U$43143 ( \43486 , \43483 , \43485 );
nand \U$43144 ( \43487 , \36850 , \36641 , \36643 );
nand \U$43145 ( \43488 , \43486 , \43487 );
nand \U$43146 ( \43489 , \43482 , \43488 );
not \U$43147 ( \43490 , \43439 );
not \U$43148 ( \43491 , \43435 );
or \U$43149 ( \43492 , \43490 , \43491 );
nand \U$43150 ( \43493 , \43430 , \43427 );
nand \U$43151 ( \43494 , \43492 , \43493 );
xor \U$43152 ( \43495 , \43297 , \43318 );
xor \U$43153 ( \43496 , \43495 , \43348 );
xor \U$43154 ( \43497 , \43494 , \43496 );
nand \U$43155 ( \43498 , \43456 , \43450 );
not \U$43156 ( \43499 , \43498 );
not \U$43157 ( \43500 , \43460 );
or \U$43158 ( \43501 , \43499 , \43500 );
not \U$43159 ( \43502 , \43456 );
nand \U$43160 ( \43503 , \43502 , \43449 );
nand \U$43161 ( \43504 , \43501 , \43503 );
buf \U$43162 ( \43505 , \43504 );
and \U$43163 ( \43506 , \43497 , \43505 );
not \U$43164 ( \43507 , \43497 );
not \U$43165 ( \43508 , \43505 );
and \U$43166 ( \43509 , \43507 , \43508 );
nor \U$43167 ( \43510 , \43506 , \43509 );
not \U$43168 ( \43511 , \43421 );
not \U$43169 ( \43512 , \43511 );
not \U$43170 ( \43513 , \43440 );
or \U$43171 ( \43514 , \43512 , \43513 );
nand \U$43172 ( \43515 , \43514 , \43443 );
not \U$43173 ( \43516 , \43440 );
nand \U$43174 ( \43517 , \43516 , \43421 );
nand \U$43175 ( \43518 , \43515 , \43517 );
and \U$43176 ( \43519 , \43391 , \43363 );
not \U$43177 ( \43520 , \43391 );
and \U$43178 ( \43521 , \43520 , \43364 );
or \U$43179 ( \43522 , \43519 , \43521 );
and \U$43180 ( \43523 , \43522 , \43359 );
not \U$43181 ( \43524 , \43522 );
and \U$43182 ( \43525 , \43524 , \43360 );
nor \U$43183 ( \43526 , \43523 , \43525 );
xnor \U$43184 ( \43527 , \43518 , \43526 );
xnor \U$43185 ( \43528 , \43510 , \43527 );
not \U$43186 ( \43529 , \43444 );
not \U$43187 ( \43530 , \43529 );
not \U$43188 ( \43531 , \43478 );
or \U$43189 ( \43532 , \43530 , \43531 );
nand \U$43190 ( \43533 , \43471 , \43473 , \43465 );
nand \U$43191 ( \43534 , \43532 , \43533 );
nand \U$43192 ( \43535 , \43528 , \43534 );
not \U$43193 ( \43536 , \43396 );
not \U$43194 ( \43537 , \43355 );
or \U$43195 ( \43538 , \43536 , \43537 );
or \U$43196 ( \43539 , \43355 , \43396 );
nand \U$43197 ( \43540 , \43538 , \43539 );
buf \U$43198 ( \43541 , \43393 );
not \U$43199 ( \43542 , \43541 );
and \U$43200 ( \43543 , \43540 , \43542 );
not \U$43201 ( \43544 , \43540 );
and \U$43202 ( \43545 , \43544 , \43541 );
nor \U$43203 ( \43546 , \43543 , \43545 );
not \U$43204 ( \43547 , \43494 );
not \U$43205 ( \43548 , \43504 );
or \U$43206 ( \43549 , \43547 , \43548 );
or \U$43207 ( \43550 , \43504 , \43494 );
nand \U$43208 ( \43551 , \43550 , \43496 );
nand \U$43209 ( \43552 , \43549 , \43551 );
xor \U$43210 ( \43553 , \43175 , \43221 );
xor \U$43211 ( \43554 , \43553 , \43224 );
nor \U$43212 ( \43555 , \43552 , \43554 );
not \U$43213 ( \43556 , \43555 );
nand \U$43214 ( \43557 , \43552 , \43554 );
nand \U$43215 ( \43558 , \43556 , \43557 );
xnor \U$43216 ( \43559 , \43546 , \43558 );
not \U$43217 ( \43560 , \43510 );
not \U$43218 ( \43561 , \43560 );
not \U$43219 ( \43562 , \43527 );
or \U$43220 ( \43563 , \43561 , \43562 );
nand \U$43221 ( \43564 , \43515 , \43517 , \43526 );
nand \U$43222 ( \43565 , \43563 , \43564 );
nand \U$43223 ( \43566 , \43559 , \43565 );
or \U$43224 ( \43567 , \43555 , \43546 );
nand \U$43225 ( \43568 , \43567 , \43557 );
not \U$43226 ( \43569 , \43568 );
xor \U$43227 ( \43570 , \43409 , \43294 );
nand \U$43228 ( \43571 , \43569 , \43570 );
nand \U$43229 ( \43572 , \43489 , \43535 , \43566 , \43571 );
not \U$43230 ( \43573 , \43572 );
nand \U$43231 ( \43574 , \42648 , \43415 , \43573 );
not \U$43232 ( \43575 , \43288 );
not \U$43233 ( \43576 , \43241 );
nor \U$43234 ( \43577 , \43413 , \43292 );
not \U$43235 ( \43578 , \43577 );
or \U$43236 ( \43579 , \43576 , \43578 );
not \U$43237 ( \43580 , \43105 );
not \U$43238 ( \43581 , \43240 );
nand \U$43239 ( \43582 , \43580 , \43581 );
nand \U$43240 ( \43583 , \43579 , \43582 );
not \U$43241 ( \43584 , \43583 );
or \U$43242 ( \43585 , \43575 , \43584 );
not \U$43243 ( \43586 , \43279 );
not \U$43244 ( \43587 , \43287 );
nand \U$43245 ( \43588 , \43586 , \43587 );
nand \U$43246 ( \43589 , \43585 , \43588 );
buf \U$43247 ( \43590 , \43270 );
nand \U$43248 ( \43591 , \43589 , \43590 );
not \U$43249 ( \43592 , \43570 );
nand \U$43250 ( \43593 , \43592 , \43568 );
not \U$43251 ( \43594 , \43593 );
nand \U$43252 ( \43595 , \43594 , \43415 );
not \U$43253 ( \43596 , \43265 );
not \U$43254 ( \43597 , \43262 );
or \U$43255 ( \43598 , \43596 , \43597 );
not \U$43256 ( \43599 , \43269 );
nand \U$43257 ( \43600 , \43598 , \43599 );
and \U$43258 ( \43601 , \43574 , \43591 , \43595 , \43600 );
not \U$43259 ( \43602 , \37764 );
not \U$43260 ( \43603 , \42618 );
not \U$43261 ( \43604 , \42587 );
or \U$43262 ( \43605 , \43603 , \43604 );
nand \U$43263 ( \43606 , \42625 , \42629 );
nand \U$43264 ( \43607 , \43605 , \43606 );
nand \U$43265 ( \43608 , \43607 , \42585 , \42620 , \42645 );
not \U$43266 ( \43609 , \42584 );
nand \U$43267 ( \43610 , \43609 , \42563 );
not \U$43268 ( \43611 , \42645 );
nor \U$43269 ( \43612 , \43610 , \43611 );
nor \U$43270 ( \43613 , \42640 , \42644 );
nor \U$43271 ( \43614 , \43612 , \43613 );
nand \U$43272 ( \43615 , \43608 , \43614 );
nand \U$43273 ( \43616 , \43602 , \43615 );
or \U$43274 ( \43617 , \37164 , \37309 );
not \U$43275 ( \43618 , \43617 );
nor \U$43276 ( \43619 , \37730 , \37762 );
not \U$43277 ( \43620 , \43619 );
not \U$43278 ( \43621 , \37725 );
or \U$43279 ( \43622 , \43620 , \43621 );
not \U$43280 ( \43623 , \37311 );
not \U$43281 ( \43624 , \37724 );
nand \U$43282 ( \43625 , \43623 , \43624 );
nand \U$43283 ( \43626 , \43622 , \43625 );
nand \U$43284 ( \43627 , \43626 , \37310 );
not \U$43285 ( \43628 , \43627 );
or \U$43286 ( \43629 , \43618 , \43628 );
buf \U$43287 ( \43630 , \37159 );
nand \U$43288 ( \43631 , \43629 , \43630 );
or \U$43289 ( \43632 , \36858 , \37158 );
nand \U$43290 ( \43633 , \43616 , \43631 , \43632 );
nand \U$43291 ( \43634 , \43633 , \43573 );
not \U$43292 ( \43635 , \43634 );
not \U$43293 ( \43636 , \43566 );
nor \U$43294 ( \43637 , \43482 , \43488 );
not \U$43295 ( \43638 , \43637 );
not \U$43296 ( \43639 , \43535 );
or \U$43297 ( \43640 , \43638 , \43639 );
or \U$43298 ( \43641 , \43534 , \43528 );
nand \U$43299 ( \43642 , \43640 , \43641 );
not \U$43300 ( \43643 , \43642 );
or \U$43301 ( \43644 , \43636 , \43643 );
or \U$43302 ( \43645 , \43565 , \43559 );
nand \U$43303 ( \43646 , \43644 , \43645 );
nand \U$43304 ( \43647 , \43646 , \43571 );
not \U$43305 ( \43648 , \43647 );
or \U$43306 ( \43649 , \43635 , \43648 );
buf \U$43307 ( \43650 , \43415 );
nand \U$43308 ( \43651 , \43649 , \43650 );
nand \U$43309 ( \43652 , \43601 , \43651 );
nand \U$43310 ( \43653 , \29091 , \31085 , \34842 , \43652 );
not \U$43311 ( \43654 , \28107 );
nand \U$43312 ( \43655 , \28601 , \28605 );
and \U$43313 ( \43656 , \43654 , \43655 );
buf \U$43314 ( \43657 , \28606 );
nor \U$43315 ( \43658 , \43656 , \43657 );
not \U$43316 ( \43659 , \28106 );
nand \U$43317 ( \43660 , \43659 , \27499 );
and \U$43318 ( \43661 , \43660 , \43655 );
nor \U$43319 ( \43662 , \28609 , \29088 );
nand \U$43320 ( \43663 , \43662 , \28598 );
or \U$43321 ( \43664 , \28597 , \28596 );
nand \U$43322 ( \43665 , \43661 , \43663 , \43664 );
nand \U$43323 ( \43666 , \43658 , \43665 );
nand \U$43324 ( \43667 , \43653 , \43666 );
not \U$43325 ( \43668 , \43667 );
not \U$43326 ( \43669 , \31073 );
not \U$43327 ( \43670 , \43669 );
not \U$43328 ( \43671 , \31082 );
and \U$43329 ( \43672 , \43670 , \43671 );
and \U$43330 ( \43673 , \31052 , \31070 );
nor \U$43331 ( \43674 , \43672 , \43673 );
buf \U$43332 ( \43675 , \30828 );
nor \U$43333 ( \43676 , \30833 , \31048 );
nand \U$43334 ( \43677 , \43675 , \43676 );
or \U$43335 ( \43678 , \29891 , \30827 );
nand \U$43336 ( \43679 , \43677 , \43678 );
and \U$43337 ( \43680 , \43674 , \43679 );
not \U$43338 ( \43681 , \31071 );
nor \U$43339 ( \43682 , \31073 , \31083 );
not \U$43340 ( \43683 , \43682 );
or \U$43341 ( \43684 , \43681 , \43683 );
or \U$43342 ( \43685 , \31052 , \31070 );
nand \U$43343 ( \43686 , \43684 , \43685 );
nor \U$43344 ( \43687 , \43680 , \43686 );
not \U$43345 ( \43688 , \43687 );
nand \U$43346 ( \43689 , \34827 , \34807 );
or \U$43347 ( \43690 , \34840 , \43689 );
nand \U$43348 ( \43691 , \34834 , \34839 );
nand \U$43349 ( \43692 , \43690 , \43691 );
not \U$43350 ( \43693 , \43692 );
nand \U$43351 ( \43694 , \31709 , \32119 );
nand \U$43352 ( \43695 , \43693 , \43694 );
and \U$43353 ( \43696 , \43695 , \32121 );
and \U$43354 ( \43697 , \31704 , \31706 );
nor \U$43355 ( \43698 , \43696 , \43697 );
not \U$43356 ( \43699 , \43698 );
not \U$43357 ( \43700 , \34126 );
not \U$43358 ( \43701 , \33730 );
or \U$43359 ( \43702 , \43700 , \43701 );
nand \U$43360 ( \43703 , \34134 , \34794 );
nand \U$43361 ( \43704 , \43702 , \43703 );
not \U$43362 ( \43705 , \43704 );
nor \U$43363 ( \43706 , \34127 , \33727 );
not \U$43364 ( \43707 , \43706 );
or \U$43365 ( \43708 , \43705 , \43707 );
nand \U$43366 ( \43709 , \33726 , \33721 );
not \U$43367 ( \43710 , \43709 );
nor \U$43368 ( \43711 , \32725 , \33454 );
nor \U$43369 ( \43712 , \43710 , \43711 );
nand \U$43370 ( \43713 , \43708 , \43712 );
buf \U$43371 ( \43714 , \33455 );
nand \U$43372 ( \43715 , \43713 , \32121 , \34841 , \43714 );
not \U$43373 ( \43716 , \43715 );
or \U$43374 ( \43717 , \43699 , \43716 );
nand \U$43375 ( \43718 , \43717 , \31085 );
not \U$43376 ( \43719 , \43718 );
or \U$43377 ( \43720 , \43688 , \43719 );
buf \U$43378 ( \43721 , \29091 );
nand \U$43379 ( \43722 , \43720 , \43721 );
nand \U$43380 ( \43723 , \43668 , \43722 );
or \U$43381 ( \43724 , \25933 , \25137 );
not \U$43382 ( \43725 , \25118 );
not \U$43383 ( \43726 , \25133 );
and \U$43384 ( \43727 , \24044 , \43724 , \43725 , \43726 );
and \U$43385 ( \43728 , \25949 , \25952 , \43727 );
nand \U$43386 ( \43729 , \43723 , \27104 , \43728 );
or \U$43387 ( \43730 , \26801 , \26805 );
not \U$43388 ( \43731 , \26934 );
nand \U$43389 ( \43732 , \43731 , \26939 );
and \U$43390 ( \43733 , \43730 , \43732 );
not \U$43391 ( \43734 , \43733 );
not \U$43392 ( \43735 , \26615 );
not \U$43393 ( \43736 , \26320 );
nand \U$43394 ( \43737 , \43736 , \25961 );
or \U$43395 ( \43738 , \43735 , \43737 );
not \U$43396 ( \43739 , \26614 );
nand \U$43397 ( \43740 , \43739 , \26325 , \26331 );
nand \U$43398 ( \43741 , \43738 , \43740 );
nand \U$43399 ( \43742 , \43741 , \26806 );
not \U$43400 ( \43743 , \43742 );
or \U$43401 ( \43744 , \43734 , \43743 );
not \U$43402 ( \43745 , \27103 );
nand \U$43403 ( \43746 , \43744 , \43745 );
buf \U$43404 ( \43747 , \27030 );
not \U$43405 ( \43748 , \43747 );
not \U$43406 ( \43749 , \27102 );
nand \U$43407 ( \43750 , \27084 , \27092 );
or \U$43408 ( \43751 , \27081 , \43750 );
nand \U$43409 ( \43752 , \27066 , \27080 );
nand \U$43410 ( \43753 , \43751 , \43752 );
not \U$43411 ( \43754 , \43753 );
or \U$43412 ( \43755 , \43749 , \43754 );
or \U$43413 ( \43756 , \27095 , \27101 );
nand \U$43414 ( \43757 , \43755 , \43756 );
not \U$43415 ( \43758 , \43757 );
or \U$43416 ( \43759 , \43748 , \43758 );
not \U$43417 ( \43760 , \27029 );
nand \U$43418 ( \43761 , \43760 , \27014 , \27016 );
nand \U$43419 ( \43762 , \43759 , \43761 );
not \U$43420 ( \43763 , \43762 );
nand \U$43421 ( \43764 , \27105 , \43729 , \43746 , \43763 );
not \U$43422 ( \43765 , \43764 );
or \U$43423 ( \43766 , \16879 , \43765 );
not \U$43424 ( \43767 , \15935 );
not \U$43425 ( \43768 , \13787 );
not \U$43426 ( \43769 , \12928 );
or \U$43427 ( \43770 , \43768 , \43769 );
not \U$43428 ( \43771 , \14265 );
nand \U$43429 ( \43772 , \43771 , \13791 );
nand \U$43430 ( \43773 , \43770 , \43772 );
nand \U$43431 ( \43774 , \43773 , \13789 );
or \U$43432 ( \43775 , \43774 , \14278 );
nand \U$43433 ( \43776 , \14270 , \14277 );
nand \U$43434 ( \43777 , \43775 , \43776 );
nand \U$43435 ( \43778 , \43777 , \12367 );
or \U$43436 ( \43779 , \12366 , \11887 );
nand \U$43437 ( \43780 , \43778 , \43779 );
not \U$43438 ( \43781 , \43780 );
or \U$43439 ( \43782 , \43767 , \43781 );
not \U$43440 ( \43783 , \15527 );
not \U$43441 ( \43784 , \15933 );
nor \U$43442 ( \43785 , \15924 , \43784 );
nand \U$43443 ( \43786 , \43783 , \43785 );
nor \U$43444 ( \43787 , \15122 , \14695 );
and \U$43445 ( \43788 , \43787 , \15526 );
nor \U$43446 ( \43789 , \15519 , \15525 );
nor \U$43447 ( \43790 , \43788 , \43789 );
nand \U$43448 ( \43791 , \43786 , \43790 );
not \U$43449 ( \43792 , \15919 );
and \U$43450 ( \43793 , \43791 , \43792 );
nand \U$43451 ( \43794 , \15918 , \15536 );
not \U$43452 ( \43795 , \43794 );
nor \U$43453 ( \43796 , \43793 , \43795 );
nand \U$43454 ( \43797 , \43782 , \43796 );
not \U$43455 ( \43798 , \43797 );
not \U$43456 ( \43799 , \16877 );
not \U$43457 ( \43800 , \43799 );
or \U$43458 ( \43801 , \43798 , \43800 );
not \U$43459 ( \43802 , \16868 );
not \U$43460 ( \43803 , \16706 );
or \U$43461 ( \43804 , \16708 , \16726 );
not \U$43462 ( \43805 , \43804 );
not \U$43463 ( \43806 , \16731 );
nor \U$43464 ( \43807 , \43806 , \16738 );
nand \U$43465 ( \43808 , \16727 , \43807 );
not \U$43466 ( \43809 , \43808 );
or \U$43467 ( \43810 , \43805 , \43809 );
nand \U$43468 ( \43811 , \43810 , \16586 );
or \U$43469 ( \43812 , \16545 , \16585 );
nand \U$43470 ( \43813 , \43811 , \43812 );
not \U$43471 ( \43814 , \43813 );
or \U$43472 ( \43815 , \43803 , \43814 );
or \U$43473 ( \43816 , \16701 , \16705 );
nand \U$43474 ( \43817 , \43815 , \43816 );
not \U$43475 ( \43818 , \43817 );
or \U$43476 ( \43819 , \43802 , \43818 );
not \U$43477 ( \43820 , \16814 );
not \U$43478 ( \43821 , \16742 );
or \U$43479 ( \43822 , \43820 , \43821 );
not \U$43480 ( \43823 , \16813 );
nand \U$43481 ( \43824 , \43822 , \43823 );
not \U$43482 ( \43825 , \16850 );
or \U$43483 ( \43826 , \43824 , \43825 );
not \U$43484 ( \43827 , \16849 );
nand \U$43485 ( \43828 , \43827 , \16823 );
nand \U$43486 ( \43829 , \43826 , \43828 );
and \U$43487 ( \43830 , \43829 , \16867 );
nor \U$43488 ( \43831 , \16854 , \16866 );
nor \U$43489 ( \43832 , \43830 , \43831 );
nand \U$43490 ( \43833 , \43819 , \43832 );
buf \U$43491 ( \43834 , \16876 );
and \U$43492 ( \43835 , \43833 , \43834 );
not \U$43493 ( \43836 , \16875 );
not \U$43494 ( \43837 , \16870 );
or \U$43495 ( \43838 , \43836 , \43837 );
not \U$43496 ( \43839 , \16874 );
nand \U$43497 ( \43840 , \43838 , \43839 );
not \U$43498 ( \43841 , \43840 );
nor \U$43499 ( \43842 , \43835 , \43841 );
nand \U$43500 ( \43843 , \43801 , \43842 );
not \U$43501 ( \43844 , \43843 );
nand \U$43502 ( \43845 , \43766 , \43844 );
not \U$43503 ( \43846 , \43845 );
or \U$43504 ( \43847 , \8535 , \43846 );
not \U$43505 ( \43848 , \3088 );
not \U$43506 ( \43849 , \5592 );
not \U$43507 ( \43850 , \8532 );
not \U$43508 ( \43851 , \6988 );
not \U$43509 ( \43852 , \7742 );
not \U$43510 ( \43853 , \7423 );
nand \U$43511 ( \43854 , \43852 , \43853 );
not \U$43512 ( \43855 , \43854 );
not \U$43513 ( \43856 , \8430 );
nand \U$43514 ( \43857 , \43856 , \7765 );
not \U$43515 ( \43858 , \43857 );
nand \U$43516 ( \43859 , \43858 , \7743 );
not \U$43517 ( \43860 , \43859 );
or \U$43518 ( \43861 , \43855 , \43860 );
nand \U$43519 ( \43862 , \43861 , \7760 );
not \U$43520 ( \43863 , \7759 );
not \U$43521 ( \43864 , \7755 );
or \U$43522 ( \43865 , \43863 , \43864 );
not \U$43523 ( \43866 , \7754 );
nand \U$43524 ( \43867 , \43865 , \43866 );
nand \U$43525 ( \43868 , \43862 , \43867 );
not \U$43526 ( \43869 , \43868 );
or \U$43527 ( \43870 , \43851 , \43869 );
not \U$43528 ( \43871 , \6987 );
nand \U$43529 ( \43872 , \43871 , \6940 );
nand \U$43530 ( \43873 , \43870 , \43872 );
not \U$43531 ( \43874 , \43873 );
or \U$43532 ( \43875 , \43850 , \43874 );
not \U$43533 ( \43876 , \8493 );
not \U$43534 ( \43877 , \8524 );
not \U$43535 ( \43878 , \8529 );
or \U$43536 ( \43879 , \43877 , \43878 );
nand \U$43537 ( \43880 , \8512 , \8518 );
or \U$43538 ( \43881 , \8530 , \43880 );
nand \U$43539 ( \43882 , \43879 , \43881 );
not \U$43540 ( \43883 , \43882 );
or \U$43541 ( \43884 , \43876 , \43883 );
not \U$43542 ( \43885 , \8492 );
nand \U$43543 ( \43886 , \43885 , \8480 , \8483 );
nand \U$43544 ( \43887 , \43884 , \43886 );
not \U$43545 ( \43888 , \43887 );
nand \U$43546 ( \43889 , \43875 , \43888 );
not \U$43547 ( \43890 , \43889 );
or \U$43548 ( \43891 , \43849 , \43890 );
not \U$43549 ( \43892 , \5588 );
nor \U$43550 ( \43893 , \43892 , \5590 );
not \U$43551 ( \43894 , \43893 );
nor \U$43552 ( \43895 , \4042 , \5303 );
not \U$43553 ( \43896 , \43895 );
or \U$43554 ( \43897 , \43894 , \43896 );
not \U$43555 ( \43898 , \4041 );
or \U$43556 ( \43899 , \3819 , \4028 );
or \U$43557 ( \43900 , \43898 , \43899 );
not \U$43558 ( \43901 , \4040 );
not \U$43559 ( \43902 , \4030 );
or \U$43560 ( \43903 , \43901 , \43902 );
not \U$43561 ( \43904 , \4035 );
nand \U$43562 ( \43905 , \43903 , \43904 );
nand \U$43563 ( \43906 , \43900 , \43905 );
buf \U$43564 ( \43907 , \3345 );
and \U$43565 ( \43908 , \43906 , \43907 );
nor \U$43566 ( \43909 , \3338 , \3344 );
nor \U$43567 ( \43910 , \43908 , \43909 );
nand \U$43568 ( \43911 , \43897 , \43910 );
not \U$43569 ( \43912 , \5297 );
not \U$43570 ( \43913 , \5300 );
or \U$43571 ( \43914 , \43912 , \43913 );
not \U$43572 ( \43915 , \4667 );
nand \U$43573 ( \43916 , \4622 , \43915 );
nand \U$43574 ( \43917 , \43914 , \43916 );
not \U$43575 ( \43918 , \43917 );
not \U$43576 ( \43919 , \4690 );
or \U$43577 ( \43920 , \43918 , \43919 );
nand \U$43578 ( \43921 , \4673 , \4688 );
nand \U$43579 ( \43922 , \43920 , \43921 );
nand \U$43580 ( \43923 , \43922 , \4700 );
or \U$43581 ( \43924 , \4699 , \4695 );
and \U$43582 ( \43925 , \43923 , \43924 );
not \U$43583 ( \43926 , \4043 );
nor \U$43584 ( \43927 , \43925 , \43926 );
nor \U$43585 ( \43928 , \43911 , \43927 );
nand \U$43586 ( \43929 , \43891 , \43928 );
not \U$43587 ( \43930 , \43929 );
or \U$43588 ( \43931 , \43848 , \43930 );
or \U$43589 ( \43932 , \3083 , \3087 );
nand \U$43590 ( \43933 , \43931 , \43932 );
not \U$43591 ( \43934 , \43933 );
nand \U$43592 ( \43935 , \43847 , \43934 );
not \U$43593 ( \43936 , \43935 );
or \U$43594 ( \43937 , \2797 , \43936 );
not \U$43595 ( \43938 , \2728 );
not \U$43596 ( \43939 , \2529 );
not \U$43597 ( \43940 , \43939 );
nand \U$43598 ( \43941 , \2172 , \2015 );
or \U$43599 ( \43942 , \2540 , \43941 );
nand \U$43600 ( \43943 , \2533 , \2539 );
nand \U$43601 ( \43944 , \43942 , \43943 );
not \U$43602 ( \43945 , \43944 );
or \U$43603 ( \43946 , \43940 , \43945 );
nor \U$43604 ( \43947 , \2527 , \2414 );
and \U$43605 ( \43948 , \43947 , \2303 );
and \U$43606 ( \43949 , \2522 , \2526 );
nor \U$43607 ( \43950 , \43948 , \43949 );
nand \U$43608 ( \43951 , \43946 , \43950 );
not \U$43609 ( \43952 , \43951 );
or \U$43610 ( \43953 , \43938 , \43952 );
nor \U$43611 ( \43954 , \2546 , \2643 );
and \U$43612 ( \43955 , \43954 , \2727 );
and \U$43613 ( \43956 , \2648 , \2726 );
nor \U$43614 ( \43957 , \43955 , \43956 );
nand \U$43615 ( \43958 , \43953 , \43957 );
nand \U$43616 ( \43959 , \43958 , \2795 );
or \U$43617 ( \43960 , \2732 , \2794 );
and \U$43618 ( \43961 , \43959 , \43960 );
nand \U$43619 ( \43962 , \43937 , \43961 );
not \U$43620 ( \43963 , \43962 );
and \U$43621 ( \43964 , RI9871e60_141, \1106 );
not \U$43622 ( \43965 , RI9871e60_141);
and \U$43623 ( \43966 , \43965 , \1098 );
nor \U$43624 ( \43967 , \43964 , \43966 );
and \U$43625 ( \43968 , \43967 , \1353 );
and \U$43626 ( \43969 , \2746 , \1382 );
nor \U$43627 ( \43970 , \43968 , \43969 );
not \U$43628 ( \43971 , \43970 );
xor \U$43629 ( \43972 , \2742 , \2744 );
and \U$43630 ( \43973 , \43972 , \2749 );
and \U$43631 ( \43974 , \2742 , \2744 );
nor \U$43632 ( \43975 , \43973 , \43974 );
not \U$43633 ( \43976 , \43975 );
or \U$43634 ( \43977 , \43971 , \43976 );
or \U$43635 ( \43978 , \43975 , \43970 );
nand \U$43636 ( \43979 , \43977 , \43978 );
not \U$43637 ( \43980 , \43979 );
xor \U$43638 ( \43981 , \2757 , \2763 );
and \U$43639 ( \43982 , \43981 , \2773 );
and \U$43640 ( \43983 , \2757 , \2763 );
nor \U$43641 ( \43984 , \43982 , \43983 );
not \U$43642 ( \43985 , \43984 );
not \U$43643 ( \43986 , \1162 );
not \U$43644 ( \43987 , \2755 );
or \U$43645 ( \43988 , \43986 , \43987 );
and \U$43646 ( \43989 , \1834 , \1165 );
and \U$43647 ( \43990 , \1275 , \1166 );
nor \U$43648 ( \43991 , \43989 , \43990 );
or \U$43649 ( \43992 , \43991 , \1719 );
nand \U$43650 ( \43993 , \43988 , \43992 );
not \U$43651 ( \43994 , \43993 );
not \U$43652 ( \43995 , \2711 );
not \U$43653 ( \43996 , \43995 );
and \U$43654 ( \43997 , \2740 , \876 );
and \U$43655 ( \43998 , \924 , RI9872130_147);
nor \U$43656 ( \43999 , \43997 , \43998 );
not \U$43657 ( \44000 , \43999 );
and \U$43658 ( \44001 , \43996 , \44000 );
and \U$43659 ( \44002 , \43995 , \43999 );
nor \U$43660 ( \44003 , \44001 , \44002 );
not \U$43661 ( \44004 , \44003 );
or \U$43662 ( \44005 , \43994 , \44004 );
or \U$43663 ( \44006 , \44003 , \43993 );
nand \U$43664 ( \44007 , \44005 , \44006 );
not \U$43665 ( \44008 , \44007 );
xnor \U$43666 ( \44009 , \1672 , RI9871d70_139);
and \U$43667 ( \44010 , \44009 , \832 );
and \U$43668 ( \44011 , \2761 , \859 );
nor \U$43669 ( \44012 , \44010 , \44011 );
not \U$43670 ( \44013 , \44012 );
or \U$43671 ( \44014 , \2768 , \1612 );
xnor \U$43672 ( \44015 , \1447 , \1758 );
or \U$43673 ( \44016 , \44015 , \1068 );
nand \U$43674 ( \44017 , \44014 , \44016 );
not \U$43675 ( \44018 , \44017 );
and \U$43676 ( \44019 , \44013 , \44018 );
and \U$43677 ( \44020 , \44012 , \44017 );
nor \U$43678 ( \44021 , \44019 , \44020 );
not \U$43679 ( \44022 , \44021 );
and \U$43680 ( \44023 , \44008 , \44022 );
and \U$43681 ( \44024 , \44007 , \44021 );
nor \U$43682 ( \44025 , \44023 , \44024 );
not \U$43683 ( \44026 , \44025 );
and \U$43684 ( \44027 , \43985 , \44026 );
and \U$43685 ( \44028 , \43984 , \44025 );
nor \U$43686 ( \44029 , \44027 , \44028 );
not \U$43687 ( \44030 , \44029 );
or \U$43688 ( \44031 , \43980 , \44030 );
or \U$43689 ( \44032 , \44029 , \43979 );
nand \U$43690 ( \44033 , \44031 , \44032 );
not \U$43691 ( \44034 , \44033 );
xor \U$43692 ( \44035 , \2738 , \2750 );
and \U$43693 ( \44036 , \44035 , \2774 );
and \U$43694 ( \44037 , \2738 , \2750 );
nor \U$43695 ( \44038 , \44036 , \44037 );
not \U$43696 ( \44039 , \44038 );
and \U$43697 ( \44040 , \2782 , \2787 );
and \U$43698 ( \44041 , \2664 , \2783 );
nor \U$43699 ( \44042 , \44040 , \44041 );
not \U$43700 ( \44043 , \44042 );
and \U$43701 ( \44044 , \44039 , \44043 );
and \U$43702 ( \44045 , \44038 , \44042 );
nor \U$43703 ( \44046 , \44044 , \44045 );
not \U$43704 ( \44047 , \44046 );
or \U$43705 ( \44048 , \44034 , \44047 );
or \U$43706 ( \44049 , \44046 , \44033 );
nand \U$43707 ( \44050 , \44048 , \44049 );
not \U$43708 ( \44051 , \44050 );
xor \U$43709 ( \44052 , \2779 , \2788 );
and \U$43710 ( \44053 , \44052 , \2792 );
and \U$43711 ( \44054 , \2779 , \2788 );
or \U$43712 ( \44055 , \44053 , \44054 );
not \U$43713 ( \44056 , \44055 );
or \U$43714 ( \44057 , \44051 , \44056 );
or \U$43715 ( \44058 , \44055 , \44050 );
nand \U$43716 ( \44059 , \44057 , \44058 );
xor \U$43717 ( \44060 , \2735 , \2775 );
and \U$43718 ( \44061 , \44060 , \2793 );
and \U$43719 ( \44062 , \2735 , \2775 );
nor \U$43720 ( \44063 , \44061 , \44062 );
xnor \U$43721 ( \44064 , \44059 , \44063 );
not \U$43722 ( \44065 , \44064 );
and \U$43723 ( \44066 , \43963 , \44065 );
and \U$43724 ( \44067 , \43962 , \44064 );
nor \U$43725 ( \44068 , \44066 , \44067 );
xnor \U$43726 ( \44069 , RI9874020_213, RI9874098_214);
not \U$43727 ( \44070 , \44069 );
xor \U$43728 ( \44071 , RI9875100_249, RI9875178_250);
not \U$43729 ( \44072 , \44071 );
and \U$43730 ( \44073 , \44070 , \44072 );
and \U$43731 ( \44074 , \44069 , \44071 );
nor \U$43732 ( \44075 , \44073 , \44074 );
not \U$43733 ( \44076 , \44075 );
xor \U$43734 ( \44077 , RI98751f0_251, RI9875268_252);
not \U$43735 ( \44078 , \44077 );
xnor \U$43736 ( \44079 , RI9874200_217, RI9874278_218);
not \U$43737 ( \44080 , \44079 );
or \U$43738 ( \44081 , \44078 , \44080 );
or \U$43739 ( \44082 , \44079 , \44077 );
nand \U$43740 ( \44083 , \44081 , \44082 );
not \U$43741 ( \44084 , \44083 );
and \U$43742 ( \44085 , \44076 , \44084 );
and \U$43743 ( \44086 , \44075 , \44083 );
nor \U$43744 ( \44087 , \44085 , \44086 );
not \U$43745 ( \44088 , \44087 );
not \U$43746 ( \44089 , RI9874b60_237);
not \U$43747 ( \44090 , RI9874bd8_238);
and \U$43748 ( \44091 , \44089 , \44090 );
and \U$43749 ( \44092 , RI9874b60_237, RI9874bd8_238);
nor \U$43750 ( \44093 , \44091 , \44092 );
not \U$43751 ( \44094 , \44093 );
xor \U$43752 ( \44095 , RI9874c50_239, RI9874cc8_240);
not \U$43753 ( \44096 , \44095 );
and \U$43754 ( \44097 , \44094 , \44096 );
and \U$43755 ( \44098 , \44093 , \44095 );
nor \U$43756 ( \44099 , \44097 , \44098 );
not \U$43757 ( \44100 , \44099 );
xor \U$43758 ( \44101 , RI9874110_215, RI9874188_216);
not \U$43759 ( \44102 , \44101 );
xnor \U$43760 ( \44103 , RI98736c0_193, RI9873738_194);
not \U$43761 ( \44104 , \44103 );
or \U$43762 ( \44105 , \44102 , \44104 );
or \U$43763 ( \44106 , \44103 , \44101 );
nand \U$43764 ( \44107 , \44105 , \44106 );
not \U$43765 ( \44108 , \44107 );
or \U$43766 ( \44109 , \44100 , \44108 );
or \U$43767 ( \44110 , \44099 , \44107 );
nand \U$43768 ( \44111 , \44109 , \44110 );
not \U$43769 ( \44112 , \44111 );
and \U$43770 ( \44113 , \44088 , \44112 );
and \U$43771 ( \44114 , \44087 , \44111 );
nor \U$43772 ( \44115 , \44113 , \44114 );
not \U$43773 ( \44116 , \44115 );
not \U$43774 ( \44117 , RI9873a08_200);
not \U$43775 ( \44118 , RI9873990_199);
or \U$43776 ( \44119 , \44117 , \44118 );
or \U$43777 ( \44120 , RI9873990_199, RI9873a08_200);
nand \U$43778 ( \44121 , \44119 , \44120 );
not \U$43779 ( \44122 , \44121 );
xor \U$43780 ( \44123 , RI98738a0_197, RI9873918_198);
not \U$43781 ( \44124 , \44123 );
and \U$43782 ( \44125 , \44122 , \44124 );
and \U$43783 ( \44126 , \44121 , \44123 );
nor \U$43784 ( \44127 , \44125 , \44126 );
not \U$43785 ( \44128 , \44127 );
xor \U$43786 ( \44129 , RI9873c60_205, RI9873cd8_206);
not \U$43787 ( \44130 , \44129 );
not \U$43788 ( \44131 , RI9873dc8_208);
not \U$43789 ( \44132 , RI9873d50_207);
or \U$43790 ( \44133 , \44131 , \44132 );
or \U$43791 ( \44134 , RI9873d50_207, RI9873dc8_208);
nand \U$43792 ( \44135 , \44133 , \44134 );
not \U$43793 ( \44136 , \44135 );
or \U$43794 ( \44137 , \44130 , \44136 );
or \U$43795 ( \44138 , \44135 , \44129 );
nand \U$43796 ( \44139 , \44137 , \44138 );
not \U$43797 ( \44140 , \44139 );
and \U$43798 ( \44141 , \44128 , \44140 );
and \U$43799 ( \44142 , \44127 , \44139 );
nor \U$43800 ( \44143 , \44141 , \44142 );
not \U$43801 ( \44144 , \44143 );
not \U$43802 ( \44145 , RI9874f20_245);
not \U$43803 ( \44146 , RI9874f98_246);
and \U$43804 ( \44147 , \44145 , \44146 );
and \U$43805 ( \44148 , RI9874f20_245, RI9874f98_246);
nor \U$43806 ( \44149 , \44147 , \44148 );
not \U$43807 ( \44150 , \44149 );
xor \U$43808 ( \44151 , RI9875010_247, RI9875088_248);
not \U$43809 ( \44152 , \44151 );
and \U$43810 ( \44153 , \44150 , \44152 );
and \U$43811 ( \44154 , \44149 , \44151 );
nor \U$43812 ( \44155 , \44153 , \44154 );
not \U$43813 ( \44156 , \44155 );
xnor \U$43814 ( \44157 , RI9874d40_241, RI9874db8_242);
not \U$43815 ( \44158 , \44157 );
xor \U$43816 ( \44159 , RI9874e30_243, RI9874ea8_244);
not \U$43817 ( \44160 , \44159 );
and \U$43818 ( \44161 , \44158 , \44160 );
and \U$43819 ( \44162 , \44157 , \44159 );
nor \U$43820 ( \44163 , \44161 , \44162 );
not \U$43821 ( \44164 , \44163 );
or \U$43822 ( \44165 , \44156 , \44164 );
or \U$43823 ( \44166 , \44163 , \44155 );
nand \U$43824 ( \44167 , \44165 , \44166 );
not \U$43825 ( \44168 , \44167 );
or \U$43826 ( \44169 , \44144 , \44168 );
or \U$43827 ( \44170 , \44143 , \44167 );
nand \U$43828 ( \44171 , \44169 , \44170 );
not \U$43829 ( \44172 , \44171 );
and \U$43830 ( \44173 , \44116 , \44172 );
and \U$43831 ( \44174 , \44115 , \44171 );
nor \U$43832 ( \44175 , \44173 , \44174 );
not \U$43833 ( \44176 , \44175 );
xnor \U$43834 ( \44177 , RI98742f0_219, RI9874368_220);
not \U$43835 ( \44178 , \44177 );
xor \U$43836 ( \44179 , RI9874890_231, RI9874908_232);
not \U$43837 ( \44180 , \44179 );
and \U$43838 ( \44181 , \44178 , \44180 );
and \U$43839 ( \44182 , \44177 , \44179 );
nor \U$43840 ( \44183 , \44181 , \44182 );
not \U$43841 ( \44184 , \44183 );
xor \U$43842 ( \44185 , RI98752e0_253, RI9875358_254);
not \U$43843 ( \44186 , \44185 );
xnor \U$43844 ( \44187 , RI98747a0_229, RI9874818_230);
not \U$43845 ( \44188 , \44187 );
or \U$43846 ( \44189 , \44186 , \44188 );
or \U$43847 ( \44190 , \44187 , \44185 );
nand \U$43848 ( \44191 , \44189 , \44190 );
not \U$43849 ( \44192 , \44191 );
and \U$43850 ( \44193 , \44184 , \44192 );
and \U$43851 ( \44194 , \44183 , \44191 );
nor \U$43852 ( \44195 , \44193 , \44194 );
not \U$43853 ( \44196 , \44195 );
xor \U$43854 ( \44197 , RI98743e0_221, RI9874458_222);
not \U$43855 ( \44198 , \44197 );
not \U$43856 ( \44199 , RI9874548_224);
not \U$43857 ( \44200 , RI98744d0_223);
or \U$43858 ( \44201 , \44199 , \44200 );
or \U$43859 ( \44202 , RI98744d0_223, RI9874548_224);
nand \U$43860 ( \44203 , \44201 , \44202 );
not \U$43861 ( \44204 , \44203 );
or \U$43862 ( \44205 , \44198 , \44204 );
or \U$43863 ( \44206 , \44203 , \44197 );
nand \U$43864 ( \44207 , \44205 , \44206 );
not \U$43865 ( \44208 , \44207 );
not \U$43866 ( \44209 , RI9873fa8_212);
not \U$43867 ( \44210 , RI9873f30_211);
or \U$43868 ( \44211 , \44209 , \44210 );
or \U$43869 ( \44212 , RI9873f30_211, RI9873fa8_212);
nand \U$43870 ( \44213 , \44211 , \44212 );
not \U$43871 ( \44214 , \44213 );
xor \U$43872 ( \44215 , RI9873e40_209, RI9873eb8_210);
not \U$43873 ( \44216 , \44215 );
and \U$43874 ( \44217 , \44214 , \44216 );
and \U$43875 ( \44218 , \44213 , \44215 );
nor \U$43876 ( \44219 , \44217 , \44218 );
not \U$43877 ( \44220 , \44219 );
or \U$43878 ( \44221 , \44208 , \44220 );
or \U$43879 ( \44222 , \44219 , \44207 );
nand \U$43880 ( \44223 , \44221 , \44222 );
not \U$43881 ( \44224 , \44223 );
and \U$43882 ( \44225 , \44196 , \44224 );
and \U$43883 ( \44226 , \44195 , \44223 );
nor \U$43884 ( \44227 , \44225 , \44226 );
not \U$43885 ( \44228 , \44227 );
xnor \U$43886 ( \44229 , RI98737b0_195, RI9873828_196);
not \U$43887 ( \44230 , \44229 );
xor \U$43888 ( \44231 , RI98753d0_255, RI9875448_256);
not \U$43889 ( \44232 , \44231 );
and \U$43890 ( \44233 , \44230 , \44232 );
and \U$43891 ( \44234 , \44229 , \44231 );
nor \U$43892 ( \44235 , \44233 , \44234 );
not \U$43893 ( \44236 , \44235 );
not \U$43894 ( \44237 , RI9873a80_201);
not \U$43895 ( \44238 , RI9873af8_202);
and \U$43896 ( \44239 , \44237 , \44238 );
and \U$43897 ( \44240 , RI9873a80_201, RI9873af8_202);
nor \U$43898 ( \44241 , \44239 , \44240 );
not \U$43899 ( \44242 , \44241 );
xor \U$43900 ( \44243 , RI9873b70_203, RI9873be8_204);
not \U$43901 ( \44244 , \44243 );
and \U$43902 ( \44245 , \44242 , \44244 );
and \U$43903 ( \44246 , \44241 , \44243 );
nor \U$43904 ( \44247 , \44245 , \44246 );
not \U$43905 ( \44248 , \44247 );
and \U$43906 ( \44249 , \44236 , \44248 );
and \U$43907 ( \44250 , \44235 , \44247 );
nor \U$43908 ( \44251 , \44249 , \44250 );
not \U$43909 ( \44252 , \44251 );
xor \U$43910 ( \44253 , RI9874980_233, RI98749f8_234);
not \U$43911 ( \44254 , \44253 );
not \U$43912 ( \44255 , RI9874ae8_236);
not \U$43913 ( \44256 , RI9874a70_235);
or \U$43914 ( \44257 , \44255 , \44256 );
or \U$43915 ( \44258 , RI9874a70_235, RI9874ae8_236);
nand \U$43916 ( \44259 , \44257 , \44258 );
not \U$43917 ( \44260 , \44259 );
or \U$43918 ( \44261 , \44254 , \44260 );
or \U$43919 ( \44262 , \44259 , \44253 );
nand \U$43920 ( \44263 , \44261 , \44262 );
not \U$43921 ( \44264 , \44263 );
xor \U$43922 ( \44265 , RI98746b0_227, RI9874728_228);
not \U$43923 ( \44266 , \44265 );
xor \U$43924 ( \44267 , RI98745c0_225, RI9874638_226);
not \U$43925 ( \44268 , \44267 );
or \U$43926 ( \44269 , \44266 , \44268 );
or \U$43927 ( \44270 , \44267 , \44265 );
nand \U$43928 ( \44271 , \44269 , \44270 );
not \U$43929 ( \44272 , \44271 );
or \U$43930 ( \44273 , \44264 , \44272 );
or \U$43931 ( \44274 , \44271 , \44263 );
nand \U$43932 ( \44275 , \44273 , \44274 );
not \U$43933 ( \44276 , \44275 );
or \U$43934 ( \44277 , \44252 , \44276 );
or \U$43935 ( \44278 , \44251 , \44275 );
nand \U$43936 ( \44279 , \44277 , \44278 );
not \U$43937 ( \44280 , \44279 );
or \U$43938 ( \44281 , \44228 , \44280 );
or \U$43939 ( \44282 , \44227 , \44279 );
nand \U$43940 ( \44283 , \44281 , \44282 );
not \U$43941 ( \44284 , \44283 );
and \U$43942 ( \44285 , \44176 , \44284 );
and \U$43943 ( \44286 , \44175 , \44283 );
nor \U$43944 ( \44287 , \44285 , \44286 );
not \U$43945 ( \44288 , \44287 );
buf \U$43946 ( \44289 , \44288 );
nor \U$43947 ( \44290 , \44068 , \44289 );
buf \U$43948 ( \44291 , \44290 );
not \U$43949 ( \44292 , \2728 );
not \U$43950 ( \44293 , \8533 );
and \U$43951 ( \44294 , \44293 , \2542 , \3088 );
not \U$43952 ( \44295 , \44294 );
not \U$43953 ( \44296 , \43845 );
or \U$43954 ( \44297 , \44295 , \44296 );
not \U$43955 ( \44298 , \2542 );
not \U$43956 ( \44299 , \43933 );
or \U$43957 ( \44300 , \44298 , \44299 );
not \U$43958 ( \44301 , \43951 );
nand \U$43959 ( \44302 , \44300 , \44301 );
not \U$43960 ( \44303 , \44302 );
nand \U$43961 ( \44304 , \44297 , \44303 );
not \U$43962 ( \44305 , \44304 );
or \U$43963 ( \44306 , \44292 , \44305 );
nand \U$43964 ( \44307 , \44306 , \43957 );
not \U$43965 ( \44308 , \43960 );
not \U$43966 ( \44309 , \2795 );
or \U$43967 ( \44310 , \44308 , \44309 );
not \U$43968 ( \44311 , \44288 );
buf \U$43969 ( \44312 , \44311 );
nand \U$43970 ( \44313 , \44310 , \44312 );
and \U$43971 ( \44314 , \44307 , \44313 );
not \U$43972 ( \44315 , \44307 );
nand \U$43973 ( \44316 , \2795 , \43960 , \44312 );
and \U$43974 ( \44317 , \44315 , \44316 );
nor \U$43975 ( \44318 , \44314 , \44317 );
buf \U$43976 ( \44319 , \44318 );
not \U$43977 ( \44320 , \43954 );
nand \U$43978 ( \44321 , \44320 , \2644 );
not \U$43979 ( \44322 , \44321 );
not \U$43980 ( \44323 , \44304 );
and \U$43981 ( \44324 , \44322 , \44323 );
buf \U$43982 ( \44325 , \44304 );
and \U$43983 ( \44326 , \44325 , \44321 );
nor \U$43984 ( \44327 , \44324 , \44326 );
nor \U$43985 ( \44328 , \44327 , \44289 );
buf \U$43986 ( \44329 , \44328 );
not \U$43987 ( \44330 , \2174 );
not \U$43988 ( \44331 , \43935 );
or \U$43989 ( \44332 , \44330 , \44331 );
nand \U$43990 ( \44333 , \44332 , \43941 );
not \U$43991 ( \44334 , \44333 );
not \U$43992 ( \44335 , \2540 );
nand \U$43993 ( \44336 , \44335 , \43943 );
not \U$43994 ( \44337 , \44336 );
and \U$43995 ( \44338 , \44334 , \44337 );
and \U$43996 ( \44339 , \44333 , \44336 );
nor \U$43997 ( \44340 , \44338 , \44339 );
nor \U$43998 ( \44341 , \44340 , \44289 );
buf \U$43999 ( \44342 , \44341 );
not \U$44000 ( \44343 , \44293 );
buf \U$44001 ( \44344 , \43845 );
not \U$44002 ( \44345 , \44344 );
or \U$44003 ( \44346 , \44343 , \44345 );
not \U$44004 ( \44347 , \43929 );
nand \U$44005 ( \44348 , \44346 , \44347 );
not \U$44006 ( \44349 , \44348 );
nand \U$44007 ( \44350 , \3088 , \43932 );
not \U$44008 ( \44351 , \44350 );
and \U$44009 ( \44352 , \44349 , \44351 );
and \U$44010 ( \44353 , \44348 , \44350 );
nor \U$44011 ( \44354 , \44352 , \44353 );
nor \U$44012 ( \44355 , \44354 , \44289 );
buf \U$44013 ( \44356 , \44355 );
not \U$44014 ( \44357 , \5591 );
nor \U$44015 ( \44358 , \44357 , \43893 );
and \U$44016 ( \44359 , \44358 , \44312 );
nand \U$44017 ( \44360 , \43888 , \44359 );
not \U$44018 ( \44361 , \8432 );
not \U$44019 ( \44362 , \44344 );
or \U$44020 ( \44363 , \44361 , \44362 );
not \U$44021 ( \44364 , \43873 );
nand \U$44022 ( \44365 , \44363 , \44364 );
or \U$44023 ( \44366 , \44360 , \44365 );
not \U$44024 ( \44367 , \44312 );
nor \U$44025 ( \44368 , \44358 , \44367 );
and \U$44026 ( \44369 , \8532 , \44368 );
nand \U$44027 ( \44370 , \44369 , \44365 );
not \U$44028 ( \44371 , \44359 );
nor \U$44029 ( \44372 , \44371 , \8532 );
and \U$44030 ( \44373 , \43888 , \44372 );
not \U$44031 ( \44374 , \43888 );
and \U$44032 ( \44375 , \44374 , \44368 );
nor \U$44033 ( \44376 , \44373 , \44375 );
nand \U$44034 ( \44377 , \44366 , \44370 , \44376 );
buf \U$44035 ( \44378 , \44377 );
not \U$44036 ( \44379 , \44365 );
nand \U$44037 ( \44380 , \43880 , \8519 );
not \U$44038 ( \44381 , \44380 );
and \U$44039 ( \44382 , \44379 , \44381 );
and \U$44040 ( \44383 , \44365 , \44380 );
nor \U$44041 ( \44384 , \44382 , \44383 );
nor \U$44042 ( \44385 , \44384 , \44289 );
buf \U$44043 ( \44386 , \44385 );
and \U$44044 ( \44387 , \7760 , \7744 , \8431 );
not \U$44045 ( \44388 , \44387 );
not \U$44046 ( \44389 , \44344 );
or \U$44047 ( \44390 , \44388 , \44389 );
not \U$44048 ( \44391 , \43868 );
nand \U$44049 ( \44392 , \44390 , \44391 );
not \U$44050 ( \44393 , \44392 );
nand \U$44051 ( \44394 , \6988 , \43872 );
not \U$44052 ( \44395 , \44394 );
and \U$44053 ( \44396 , \44393 , \44395 );
and \U$44054 ( \44397 , \44392 , \44394 );
nor \U$44055 ( \44398 , \44396 , \44397 );
nor \U$44056 ( \44399 , \44398 , \44289 );
buf \U$44057 ( \44400 , \44399 );
not \U$44058 ( \44401 , \8431 );
not \U$44059 ( \44402 , \44344 );
or \U$44060 ( \44403 , \44401 , \44402 );
buf \U$44061 ( \44404 , \43857 );
nand \U$44062 ( \44405 , \44403 , \44404 );
not \U$44063 ( \44406 , \44405 );
nand \U$44064 ( \44407 , \43854 , \7744 );
not \U$44065 ( \44408 , \44407 );
and \U$44066 ( \44409 , \44406 , \44408 );
and \U$44067 ( \44410 , \44405 , \44407 );
nor \U$44068 ( \44411 , \44409 , \44410 );
nor \U$44069 ( \44412 , \44411 , \44289 );
buf \U$44070 ( \44413 , \44412 );
not \U$44071 ( \44414 , \16815 );
nor \U$44072 ( \44415 , \44414 , \43825 );
not \U$44073 ( \44416 , \44415 );
not \U$44074 ( \44417 , \27105 );
not \U$44075 ( \44418 , \43729 );
or \U$44076 ( \44419 , \44417 , \44418 );
buf \U$44077 ( \44420 , \16741 );
and \U$44078 ( \44421 , \15936 , \14280 , \44420 );
nand \U$44079 ( \44422 , \44419 , \44421 );
not \U$44080 ( \44423 , \43763 );
not \U$44081 ( \44424 , \43746 );
or \U$44082 ( \44425 , \44423 , \44424 );
nand \U$44083 ( \44426 , \44425 , \44421 );
buf \U$44084 ( \44427 , \43797 );
nand \U$44085 ( \44428 , \44427 , \44420 );
not \U$44086 ( \44429 , \43817 );
nand \U$44087 ( \44430 , \44422 , \44426 , \44428 , \44429 );
not \U$44088 ( \44431 , \44430 );
or \U$44089 ( \44432 , \44416 , \44431 );
not \U$44090 ( \44433 , \43829 );
nand \U$44091 ( \44434 , \44432 , \44433 );
not \U$44092 ( \44435 , \43831 );
nand \U$44093 ( \44436 , \44435 , \16867 );
and \U$44094 ( \44437 , \44434 , \44436 );
not \U$44095 ( \44438 , \44434 );
not \U$44096 ( \44439 , \44436 );
and \U$44097 ( \44440 , \44438 , \44439 );
nor \U$44098 ( \44441 , \44437 , \44440 );
nor \U$44099 ( \44442 , \44441 , \44367 );
buf \U$44100 ( \44443 , \44442 );
not \U$44101 ( \44444 , \16815 );
not \U$44102 ( \44445 , \44430 );
or \U$44103 ( \44446 , \44444 , \44445 );
buf \U$44104 ( \44447 , \43824 );
nand \U$44105 ( \44448 , \44446 , \44447 );
not \U$44106 ( \44449 , \43825 );
nand \U$44107 ( \44450 , \44449 , \43828 );
and \U$44108 ( \44451 , \44448 , \44450 );
not \U$44109 ( \44452 , \44448 );
not \U$44110 ( \44453 , \44450 );
and \U$44111 ( \44454 , \44452 , \44453 );
nor \U$44112 ( \44455 , \44451 , \44454 );
nor \U$44113 ( \44456 , \44455 , \44367 );
buf \U$44114 ( \44457 , \44456 );
not \U$44115 ( \44458 , \44414 );
nand \U$44116 ( \44459 , \44458 , \44447 );
and \U$44117 ( \44460 , \44459 , \44430 );
not \U$44118 ( \44461 , \44459 );
not \U$44119 ( \44462 , \44430 );
and \U$44120 ( \44463 , \44461 , \44462 );
nor \U$44121 ( \44464 , \44460 , \44463 );
nor \U$44122 ( \44465 , \44464 , \44367 );
buf \U$44123 ( \44466 , \44465 );
and \U$44124 ( \44467 , \16587 , \16740 );
not \U$44125 ( \44468 , \44467 );
not \U$44126 ( \44469 , \15937 );
not \U$44127 ( \44470 , \44469 );
nand \U$44128 ( \44471 , \27105 , \43729 , \43746 , \43763 );
not \U$44129 ( \44472 , \44471 );
or \U$44130 ( \44473 , \44470 , \44472 );
not \U$44131 ( \44474 , \44427 );
nand \U$44132 ( \44475 , \44473 , \44474 );
not \U$44133 ( \44476 , \44475 );
or \U$44134 ( \44477 , \44468 , \44476 );
not \U$44135 ( \44478 , \43813 );
nand \U$44136 ( \44479 , \44477 , \44478 );
not \U$44137 ( \44480 , \44479 );
nand \U$44138 ( \44481 , \43816 , \16706 );
not \U$44139 ( \44482 , \44481 );
and \U$44140 ( \44483 , \44480 , \44482 );
and \U$44141 ( \44484 , \44479 , \44481 );
nor \U$44142 ( \44485 , \44483 , \44484 );
nor \U$44143 ( \44486 , \44485 , \44289 );
buf \U$44144 ( \44487 , \44486 );
not \U$44145 ( \44488 , \16739 );
not \U$44146 ( \44489 , \44475 );
or \U$44147 ( \44490 , \44488 , \44489 );
not \U$44148 ( \44491 , \43807 );
nand \U$44149 ( \44492 , \44490 , \44491 );
not \U$44150 ( \44493 , \44492 );
not \U$44151 ( \44494 , \43804 );
not \U$44152 ( \44495 , \44494 );
nand \U$44153 ( \44496 , \44495 , \16727 );
not \U$44154 ( \44497 , \44496 );
and \U$44155 ( \44498 , \44493 , \44497 );
and \U$44156 ( \44499 , \44492 , \44496 );
nor \U$44157 ( \44500 , \44498 , \44499 );
nor \U$44158 ( \44501 , \44500 , \44289 );
buf \U$44159 ( \44502 , \44501 );
not \U$44160 ( \44503 , \16739 );
not \U$44161 ( \44504 , \44503 );
nand \U$44162 ( \44505 , \44504 , \44491 );
xor \U$44163 ( \44506 , \44475 , \44505 );
nor \U$44164 ( \44507 , \44506 , \44289 );
buf \U$44165 ( \44508 , \44507 );
nor \U$44166 ( \44509 , \15528 , \15934 );
not \U$44167 ( \44510 , \44509 );
not \U$44168 ( \44511 , \14280 );
not \U$44169 ( \44512 , \44471 );
or \U$44170 ( \44513 , \44511 , \44512 );
not \U$44171 ( \44514 , \43780 );
nand \U$44172 ( \44515 , \44513 , \44514 );
not \U$44173 ( \44516 , \44515 );
or \U$44174 ( \44517 , \44510 , \44516 );
not \U$44175 ( \44518 , \43791 );
nand \U$44176 ( \44519 , \44517 , \44518 );
not \U$44177 ( \44520 , \44519 );
not \U$44178 ( \44521 , \15919 );
nand \U$44179 ( \44522 , \44521 , \43794 );
not \U$44180 ( \44523 , \44522 );
and \U$44181 ( \44524 , \44520 , \44523 );
and \U$44182 ( \44525 , \44519 , \44522 );
nor \U$44183 ( \44526 , \44524 , \44525 );
nor \U$44184 ( \44527 , \44526 , \44289 );
buf \U$44185 ( \44528 , \44527 );
not \U$44186 ( \44529 , \15934 );
not \U$44187 ( \44530 , \44529 );
not \U$44188 ( \44531 , \44515 );
or \U$44189 ( \44532 , \44530 , \44531 );
not \U$44190 ( \44533 , \43785 );
nand \U$44191 ( \44534 , \44532 , \44533 );
not \U$44192 ( \44535 , \44534 );
buf \U$44193 ( \44536 , \14695 );
not \U$44194 ( \44537 , \44536 );
buf \U$44195 ( \44538 , \15122 );
not \U$44196 ( \44539 , \44538 );
or \U$44197 ( \44540 , \44537 , \44539 );
or \U$44198 ( \44541 , \44538 , \44536 );
nand \U$44199 ( \44542 , \44540 , \44541 );
not \U$44200 ( \44543 , \44542 );
and \U$44201 ( \44544 , \44535 , \44543 );
and \U$44202 ( \44545 , \44534 , \44542 );
nor \U$44203 ( \44546 , \44544 , \44545 );
nor \U$44204 ( \44547 , \44546 , \44289 );
buf \U$44205 ( \44548 , \44547 );
not \U$44206 ( \44549 , \15934 );
nand \U$44207 ( \44550 , \44549 , \44533 );
xor \U$44208 ( \44551 , \44515 , \44550 );
nor \U$44209 ( \44552 , \44551 , \44289 );
buf \U$44210 ( \44553 , \44552 );
not \U$44211 ( \44554 , \14268 );
nand \U$44212 ( \44555 , \27105 , \43746 , \43763 , \43729 );
not \U$44213 ( \44556 , \44555 );
or \U$44214 ( \44557 , \44554 , \44556 );
buf \U$44215 ( \44558 , \43774 );
nand \U$44216 ( \44559 , \44557 , \44558 );
not \U$44217 ( \44560 , \44559 );
nand \U$44218 ( \44561 , \14279 , \43776 );
not \U$44219 ( \44562 , \44561 );
and \U$44220 ( \44563 , \44560 , \44562 );
and \U$44221 ( \44564 , \44559 , \44561 );
nor \U$44222 ( \44565 , \44563 , \44564 );
nor \U$44223 ( \44566 , \44565 , \44367 );
buf \U$44224 ( \44567 , \44566 );
not \U$44225 ( \44568 , \14266 );
not \U$44226 ( \44569 , \44471 );
or \U$44227 ( \44570 , \44568 , \44569 );
buf \U$44228 ( \44571 , \43772 );
nand \U$44229 ( \44572 , \44570 , \44571 );
not \U$44230 ( \44573 , \44572 );
nor \U$44231 ( \44574 , \13788 , \12929 );
not \U$44232 ( \44575 , \44574 );
nand \U$44233 ( \44576 , \44575 , \13790 );
not \U$44234 ( \44577 , \44576 );
and \U$44235 ( \44578 , \44573 , \44577 );
and \U$44236 ( \44579 , \44572 , \44576 );
nor \U$44237 ( \44580 , \44578 , \44579 );
nor \U$44238 ( \44581 , \44580 , \44367 );
buf \U$44239 ( \44582 , \44581 );
nand \U$44240 ( \44583 , \44571 , \14266 );
xor \U$44241 ( \44584 , \44583 , \44555 );
not \U$44242 ( \44585 , \44312 );
nor \U$44243 ( \44586 , \44584 , \44585 );
buf \U$44244 ( \44587 , \44586 );
buf \U$44245 ( \44588 , \26941 );
not \U$44246 ( \44589 , \44588 );
not \U$44247 ( \44590 , \26807 );
not \U$44248 ( \44591 , \44590 );
not \U$44249 ( \44592 , \43728 );
not \U$44250 ( \44593 , \43723 );
or \U$44251 ( \44594 , \44592 , \44593 );
not \U$44252 ( \44595 , \25956 );
nand \U$44253 ( \44596 , \44594 , \44595 );
not \U$44254 ( \44597 , \44596 );
or \U$44255 ( \44598 , \44591 , \44597 );
buf \U$44256 ( \44599 , \43741 );
and \U$44257 ( \44600 , \44599 , \26806 );
not \U$44258 ( \44601 , \43730 );
nor \U$44259 ( \44602 , \44600 , \44601 );
nand \U$44260 ( \44603 , \44598 , \44602 );
not \U$44261 ( \44604 , \44603 );
or \U$44262 ( \44605 , \44589 , \44604 );
buf \U$44263 ( \44606 , \43732 );
nand \U$44264 ( \44607 , \44605 , \44606 );
and \U$44265 ( \44608 , \27082 , \27094 , \27102 );
nand \U$44266 ( \44609 , \44607 , \44608 );
not \U$44267 ( \44610 , \43757 );
nand \U$44268 ( \44611 , \44609 , \44610 );
not \U$44269 ( \44612 , \44611 );
not \U$44270 ( \44613 , \43761 );
not \U$44271 ( \44614 , \44613 );
nand \U$44272 ( \44615 , \44614 , \43747 );
not \U$44273 ( \44616 , \44615 );
and \U$44274 ( \44617 , \44612 , \44616 );
and \U$44275 ( \44618 , \44611 , \44615 );
nor \U$44276 ( \44619 , \44617 , \44618 );
nor \U$44277 ( \44620 , \44619 , \44289 );
buf \U$44278 ( \44621 , \44620 );
nand \U$44279 ( \44622 , \44606 , \44588 );
and \U$44280 ( \44623 , \44603 , \44622 );
not \U$44281 ( \44624 , \44603 );
not \U$44282 ( \44625 , \44622 );
and \U$44283 ( \44626 , \44624 , \44625 );
nor \U$44284 ( \44627 , \44623 , \44626 );
nor \U$44285 ( \44628 , \44627 , \44289 );
buf \U$44286 ( \44629 , \44628 );
buf \U$44287 ( \44630 , \26321 );
not \U$44288 ( \44631 , \44630 );
nor \U$44289 ( \44632 , \44631 , \43735 );
not \U$44290 ( \44633 , \44632 );
not \U$44291 ( \44634 , \44596 );
or \U$44292 ( \44635 , \44633 , \44634 );
not \U$44293 ( \44636 , \44599 );
nand \U$44294 ( \44637 , \44635 , \44636 );
nand \U$44295 ( \44638 , \26806 , \43730 );
and \U$44296 ( \44639 , \44637 , \44638 );
not \U$44297 ( \44640 , \44637 );
not \U$44298 ( \44641 , \44638 );
and \U$44299 ( \44642 , \44640 , \44641 );
nor \U$44300 ( \44643 , \44639 , \44642 );
nor \U$44301 ( \44644 , \44643 , \44289 );
buf \U$44302 ( \44645 , \44644 );
not \U$44303 ( \44646 , \44630 );
not \U$44304 ( \44647 , \44596 );
or \U$44305 ( \44648 , \44646 , \44647 );
buf \U$44306 ( \44649 , \43737 );
nand \U$44307 ( \44650 , \44648 , \44649 );
not \U$44308 ( \44651 , \44650 );
nand \U$44309 ( \44652 , \43740 , \26615 );
not \U$44310 ( \44653 , \44652 );
and \U$44311 ( \44654 , \44651 , \44653 );
and \U$44312 ( \44655 , \44650 , \44652 );
nor \U$44313 ( \44656 , \44654 , \44655 );
nor \U$44314 ( \44657 , \44656 , \44289 );
buf \U$44315 ( \44658 , \44657 );
nand \U$44316 ( \44659 , \44649 , \44630 );
and \U$44317 ( \44660 , \44596 , \44659 );
not \U$44318 ( \44661 , \44596 );
not \U$44319 ( \44662 , \44659 );
and \U$44320 ( \44663 , \44661 , \44662 );
nor \U$44321 ( \44664 , \44660 , \44663 );
nor \U$44322 ( \44665 , \44664 , \44367 );
buf \U$44323 ( \44666 , \44665 );
not \U$44324 ( \44667 , \25952 );
nor \U$44325 ( \44668 , \44667 , \25948 );
not \U$44326 ( \44669 , \44668 );
not \U$44327 ( \44670 , \43727 );
buf \U$44328 ( \44671 , \43723 );
not \U$44329 ( \44672 , \44671 );
or \U$44330 ( \44673 , \44670 , \44672 );
not \U$44331 ( \44674 , \25947 );
nand \U$44332 ( \44675 , \44673 , \44674 );
not \U$44333 ( \44676 , \44675 );
or \U$44334 ( \44677 , \44669 , \44676 );
not \U$44335 ( \44678 , \23239 );
nand \U$44336 ( \44679 , \44677 , \44678 );
nand \U$44337 ( \44680 , \23813 , \25955 );
and \U$44338 ( \44681 , \44679 , \44680 );
not \U$44339 ( \44682 , \44679 );
not \U$44340 ( \44683 , \44680 );
and \U$44341 ( \44684 , \44682 , \44683 );
nor \U$44342 ( \44685 , \44681 , \44684 );
nor \U$44343 ( \44686 , \44685 , \44367 );
buf \U$44344 ( \44687 , \44686 );
not \U$44345 ( \44688 , \25951 );
not \U$44346 ( \44689 , \44688 );
not \U$44347 ( \44690 , \44675 );
or \U$44348 ( \44691 , \44689 , \44690 );
buf \U$44349 ( \44692 , \23233 );
nand \U$44350 ( \44693 , \44691 , \44692 );
not \U$44351 ( \44694 , \22236 );
not \U$44352 ( \44695 , \21481 );
or \U$44353 ( \44696 , \44694 , \44695 );
or \U$44354 ( \44697 , \21481 , \22236 );
nand \U$44355 ( \44698 , \44696 , \44697 );
and \U$44356 ( \44699 , \44693 , \44698 );
not \U$44357 ( \44700 , \44693 );
not \U$44358 ( \44701 , \44698 );
and \U$44359 ( \44702 , \44700 , \44701 );
nor \U$44360 ( \44703 , \44699 , \44702 );
nor \U$44361 ( \44704 , \44703 , \44367 );
buf \U$44362 ( \44705 , \44704 );
not \U$44363 ( \44706 , \25936 );
not \U$44364 ( \44707 , \44706 );
nand \U$44365 ( \44708 , \43722 , \43666 , \43653 );
nand \U$44366 ( \44709 , \44708 , \43724 );
not \U$44367 ( \44710 , \44709 );
or \U$44368 ( \44711 , \44707 , \44710 );
nand \U$44369 ( \44712 , \44711 , \43725 );
not \U$44370 ( \44713 , \43726 );
or \U$44371 ( \44714 , \44712 , \44713 );
nand \U$44372 ( \44715 , \44714 , \25940 );
not \U$44373 ( \44716 , \44715 );
not \U$44374 ( \44717 , \25945 );
not \U$44375 ( \44718 , \25944 );
or \U$44376 ( \44719 , \44717 , \44718 );
or \U$44377 ( \44720 , \25944 , \25945 );
nand \U$44378 ( \44721 , \44719 , \44720 );
not \U$44379 ( \44722 , \44721 );
and \U$44380 ( \44723 , \44716 , \44722 );
and \U$44381 ( \44724 , \44715 , \44721 );
nor \U$44382 ( \44725 , \44723 , \44724 );
nor \U$44383 ( \44726 , \44725 , \44367 );
buf \U$44384 ( \44727 , \44726 );
and \U$44385 ( \44728 , \43726 , \25940 );
xor \U$44386 ( \44729 , \44712 , \44728 );
nor \U$44387 ( \44730 , \44729 , \44367 );
buf \U$44388 ( \44731 , \44730 );
buf \U$44389 ( \44732 , \25934 );
nand \U$44390 ( \44733 , \44709 , \44732 );
nand \U$44391 ( \44734 , \43725 , \25935 );
and \U$44392 ( \44735 , \44733 , \44734 );
not \U$44393 ( \44736 , \44733 );
not \U$44394 ( \44737 , \44734 );
and \U$44395 ( \44738 , \44736 , \44737 );
nor \U$44396 ( \44739 , \44735 , \44738 );
nor \U$44397 ( \44740 , \44739 , \44367 );
buf \U$44398 ( \44741 , \44740 );
nand \U$44399 ( \44742 , \44732 , \43724 );
and \U$44400 ( \44743 , \44671 , \44742 );
not \U$44401 ( \44744 , \44671 );
not \U$44402 ( \44745 , \44742 );
and \U$44403 ( \44746 , \44744 , \44745 );
nor \U$44404 ( \44747 , \44743 , \44746 );
nor \U$44405 ( \44748 , \44747 , \44585 );
buf \U$44406 ( \44749 , \44748 );
buf \U$44407 ( \44750 , \29089 );
not \U$44408 ( \44751 , \44750 );
buf \U$44409 ( \44752 , \28599 );
nor \U$44410 ( \44753 , \44751 , \44752 );
not \U$44411 ( \44754 , \44753 );
not \U$44412 ( \44755 , \31085 );
nand \U$44413 ( \44756 , \43601 , \43651 );
not \U$44414 ( \44757 , \44756 );
not \U$44415 ( \44758 , \34842 );
or \U$44416 ( \44759 , \44757 , \44758 );
nand \U$44417 ( \44760 , \32121 , \43695 );
not \U$44418 ( \44761 , \43697 );
and \U$44419 ( \44762 , \43715 , \44760 , \44761 );
nand \U$44420 ( \44763 , \44759 , \44762 );
not \U$44421 ( \44764 , \44763 );
or \U$44422 ( \44765 , \44755 , \44764 );
buf \U$44423 ( \44766 , \43687 );
nand \U$44424 ( \44767 , \44765 , \44766 );
not \U$44425 ( \44768 , \44767 );
or \U$44426 ( \44769 , \44754 , \44768 );
not \U$44427 ( \44770 , \44752 );
buf \U$44428 ( \44771 , \43662 );
not \U$44429 ( \44772 , \44771 );
not \U$44430 ( \44773 , \44772 );
and \U$44431 ( \44774 , \44770 , \44773 );
or \U$44432 ( \44775 , \43654 , \43664 );
nand \U$44433 ( \44776 , \44775 , \43660 );
nor \U$44434 ( \44777 , \44774 , \44776 );
nand \U$44435 ( \44778 , \44769 , \44777 );
not \U$44436 ( \44779 , \44778 );
not \U$44437 ( \44780 , \43657 );
nand \U$44438 ( \44781 , \44780 , \43655 );
not \U$44439 ( \44782 , \44781 );
and \U$44440 ( \44783 , \44779 , \44782 );
and \U$44441 ( \44784 , \44778 , \44781 );
nor \U$44442 ( \44785 , \44783 , \44784 );
or \U$44443 ( \44786 , \44785 , \44367 );
not \U$44444 ( \44787 , RI9871fc8_144);
or \U$44445 ( \44788 , \44312 , \44787 );
nand \U$44446 ( \44789 , \44786 , \44788 );
buf \U$44447 ( \44790 , \44789 );
not \U$44448 ( \44791 , \44750 );
not \U$44449 ( \44792 , \44767 );
or \U$44450 ( \44793 , \44791 , \44792 );
not \U$44451 ( \44794 , \44771 );
nand \U$44452 ( \44795 , \44793 , \44794 );
not \U$44453 ( \44796 , \44795 );
nand \U$44454 ( \44797 , \28598 , \43664 );
not \U$44455 ( \44798 , \44797 );
and \U$44456 ( \44799 , \44796 , \44798 );
and \U$44457 ( \44800 , \44795 , \44797 );
nor \U$44458 ( \44801 , \44799 , \44800 );
or \U$44459 ( \44802 , \44801 , \44367 );
not \U$44460 ( \44803 , RI9871ed8_142);
or \U$44461 ( \44804 , \44312 , \44803 );
nand \U$44462 ( \44805 , \44802 , \44804 );
buf \U$44463 ( \44806 , \44805 );
not \U$44464 ( \44807 , \44767 );
not \U$44465 ( \44808 , \44771 );
nand \U$44466 ( \44809 , \44808 , \44750 );
not \U$44467 ( \44810 , \44809 );
and \U$44468 ( \44811 , \44807 , \44810 );
and \U$44469 ( \44812 , \44767 , \44809 );
nor \U$44470 ( \44813 , \44811 , \44812 );
or \U$44471 ( \44814 , \44813 , \44289 );
or \U$44472 ( \44815 , \44312 , \1009 );
nand \U$44473 ( \44816 , \44814 , \44815 );
buf \U$44474 ( \44817 , \44816 );
not \U$44475 ( \44818 , \31084 );
not \U$44476 ( \44819 , \31050 );
not \U$44477 ( \44820 , \44763 );
or \U$44478 ( \44821 , \44819 , \44820 );
not \U$44479 ( \44822 , \43679 );
nand \U$44480 ( \44823 , \44821 , \44822 );
not \U$44481 ( \44824 , \44823 );
or \U$44482 ( \44825 , \44818 , \44824 );
not \U$44483 ( \44826 , \43682 );
nand \U$44484 ( \44827 , \44825 , \44826 );
not \U$44485 ( \44828 , \44827 );
nand \U$44486 ( \44829 , \43685 , \31071 );
not \U$44487 ( \44830 , \44829 );
and \U$44488 ( \44831 , \44828 , \44830 );
and \U$44489 ( \44832 , \44827 , \44829 );
nor \U$44490 ( \44833 , \44831 , \44832 );
or \U$44491 ( \44834 , \44833 , \44289 );
or \U$44492 ( \44835 , \44312 , \1367 );
nand \U$44493 ( \44836 , \44834 , \44835 );
buf \U$44494 ( \44837 , \44836 );
nand \U$44495 ( \44838 , \44826 , \31084 );
and \U$44496 ( \44839 , \44823 , \44838 );
not \U$44497 ( \44840 , \44823 );
not \U$44498 ( \44841 , \44838 );
and \U$44499 ( \44842 , \44840 , \44841 );
nor \U$44500 ( \44843 , \44839 , \44842 );
or \U$44501 ( \44844 , \44843 , \44585 );
or \U$44502 ( \44845 , \44312 , \1348 );
nand \U$44503 ( \44846 , \44844 , \44845 );
buf \U$44504 ( \44847 , \44846 );
not \U$44505 ( \44848 , \31049 );
not \U$44506 ( \44849 , \44763 );
or \U$44507 ( \44850 , \44848 , \44849 );
not \U$44508 ( \44851 , \43676 );
nand \U$44509 ( \44852 , \44850 , \44851 );
nand \U$44510 ( \44853 , \43675 , \43678 );
and \U$44511 ( \44854 , \44852 , \44853 );
not \U$44512 ( \44855 , \44852 );
not \U$44513 ( \44856 , \44853 );
and \U$44514 ( \44857 , \44855 , \44856 );
nor \U$44515 ( \44858 , \44854 , \44857 );
or \U$44516 ( \44859 , \44858 , \44585 );
or \U$44517 ( \44860 , \44312 , \1347 );
nand \U$44518 ( \44861 , \44859 , \44860 );
buf \U$44519 ( \44862 , \44861 );
nand \U$44520 ( \44863 , \31049 , \44851 );
and \U$44521 ( \44864 , \44763 , \44863 );
not \U$44522 ( \44865 , \44763 );
not \U$44523 ( \44866 , \44863 );
and \U$44524 ( \44867 , \44865 , \44866 );
nor \U$44525 ( \44868 , \44864 , \44867 );
or \U$44526 ( \44869 , \44868 , \44367 );
or \U$44527 ( \44870 , \44312 , \829 );
nand \U$44528 ( \44871 , \44869 , \44870 );
buf \U$44529 ( \44872 , \44871 );
not \U$44530 ( \44873 , \32120 );
not \U$44531 ( \44874 , \44873 );
not \U$44532 ( \44875 , \34841 );
not \U$44533 ( \44876 , \34796 );
not \U$44534 ( \44877 , \43652 );
or \U$44535 ( \44878 , \44876 , \44877 );
nand \U$44536 ( \44879 , \43714 , \43713 );
nand \U$44537 ( \44880 , \44878 , \44879 );
not \U$44538 ( \44881 , \44880 );
or \U$44539 ( \44882 , \44875 , \44881 );
nand \U$44540 ( \44883 , \44882 , \43693 );
not \U$44541 ( \44884 , \44883 );
or \U$44542 ( \44885 , \44874 , \44884 );
buf \U$44543 ( \44886 , \43694 );
nand \U$44544 ( \44887 , \44885 , \44886 );
not \U$44545 ( \44888 , \44887 );
not \U$44546 ( \44889 , \31707 );
nand \U$44547 ( \44890 , \44889 , \44761 );
not \U$44548 ( \44891 , \44890 );
and \U$44549 ( \44892 , \44888 , \44891 );
and \U$44550 ( \44893 , \44887 , \44890 );
nor \U$44551 ( \44894 , \44892 , \44893 );
or \U$44552 ( \44895 , \44894 , \44367 );
or \U$44553 ( \44896 , \44312 , \919 );
nand \U$44554 ( \44897 , \44895 , \44896 );
buf \U$44555 ( \44898 , \44897 );
and \U$44556 ( \44899 , \44288 , \866 );
not \U$44557 ( \44900 , \44288 );
not \U$44558 ( \44901 , \44883 );
not \U$44559 ( \44902 , \32120 );
nand \U$44560 ( \44903 , \44902 , \44886 );
not \U$44561 ( \44904 , \44903 );
and \U$44562 ( \44905 , \44901 , \44904 );
and \U$44563 ( \44906 , \44883 , \44903 );
nor \U$44564 ( \44907 , \44905 , \44906 );
and \U$44565 ( \44908 , \44900 , \44907 );
nor \U$44566 ( \44909 , \44899 , \44908 );
buf \U$44567 ( \44910 , \44909 );
buf \U$44568 ( \44911 , \34829 );
not \U$44569 ( \44912 , \44911 );
not \U$44570 ( \44913 , \44912 );
not \U$44571 ( \44914 , \44880 );
or \U$44572 ( \44915 , \44913 , \44914 );
buf \U$44573 ( \44916 , \43689 );
nand \U$44574 ( \44917 , \44915 , \44916 );
not \U$44575 ( \44918 , \34840 );
nand \U$44576 ( \44919 , \44918 , \43691 );
xor \U$44577 ( \44920 , \44917 , \44919 );
or \U$44578 ( \44921 , \44920 , \44289 );
or \U$44579 ( \44922 , \44312 , \1584 );
nand \U$44580 ( \44923 , \44921 , \44922 );
buf \U$44581 ( \44924 , \44923 );
and \U$44582 ( \44925 , \44288 , \1491 );
not \U$44583 ( \44926 , \44288 );
not \U$44584 ( \44927 , \44880 );
not \U$44585 ( \44928 , \44911 );
nand \U$44586 ( \44929 , \44928 , \44916 );
not \U$44587 ( \44930 , \44929 );
and \U$44588 ( \44931 , \44927 , \44930 );
and \U$44589 ( \44932 , \44880 , \44929 );
nor \U$44590 ( \44933 , \44931 , \44932 );
and \U$44591 ( \44934 , \44926 , \44933 );
nor \U$44592 ( \44935 , \44925 , \44934 );
buf \U$44593 ( \44936 , \44935 );
not \U$44594 ( \44937 , \43704 );
not \U$44595 ( \44938 , \44937 );
nand \U$44596 ( \44939 , \44756 , \34795 );
not \U$44597 ( \44940 , \44939 );
or \U$44598 ( \44941 , \44938 , \44940 );
buf \U$44599 ( \44942 , \34128 );
nand \U$44600 ( \44943 , \44941 , \44942 );
not \U$44601 ( \44944 , \33728 );
or \U$44602 ( \44945 , \44943 , \44944 );
buf \U$44603 ( \44946 , \43709 );
nand \U$44604 ( \44947 , \44945 , \44946 );
not \U$44605 ( \44948 , \44947 );
not \U$44606 ( \44949 , \43711 );
nand \U$44607 ( \44950 , \44949 , \43714 );
not \U$44608 ( \44951 , \44950 );
and \U$44609 ( \44952 , \44948 , \44951 );
and \U$44610 ( \44953 , \44947 , \44950 );
nor \U$44611 ( \44954 , \44952 , \44953 );
or \U$44612 ( \44955 , \44954 , \44289 );
or \U$44613 ( \44956 , \44312 , \2479 );
nand \U$44614 ( \44957 , \44955 , \44956 );
buf \U$44615 ( \44958 , \44957 );
nand \U$44616 ( \44959 , \33728 , \44946 );
not \U$44617 ( \44960 , \44959 );
and \U$44618 ( \44961 , \44943 , \44960 );
not \U$44619 ( \44962 , \44943 );
and \U$44620 ( \44963 , \44962 , \44959 );
nor \U$44621 ( \44964 , \44961 , \44963 );
or \U$44622 ( \44965 , \44964 , \44367 );
or \U$44623 ( \44966 , \44312 , \1284 );
nand \U$44624 ( \44967 , \44965 , \44966 );
buf \U$44625 ( \44968 , \44967 );
nand \U$44626 ( \44969 , \44939 , \43703 );
nand \U$44627 ( \44970 , \33730 , \34126 );
nand \U$44628 ( \44971 , \44970 , \44942 );
and \U$44629 ( \44972 , \44969 , \44971 );
not \U$44630 ( \44973 , \44969 );
not \U$44631 ( \44974 , \44971 );
and \U$44632 ( \44975 , \44973 , \44974 );
nor \U$44633 ( \44976 , \44972 , \44975 );
or \U$44634 ( \44977 , \44976 , \44288 );
or \U$44635 ( \44978 , \44311 , \1850 );
nand \U$44636 ( \44979 , \44977 , \44978 );
buf \U$44637 ( \44980 , \44979 );
not \U$44638 ( \44981 , \44756 );
not \U$44639 ( \44982 , \34795 );
not \U$44640 ( \44983 , \44982 );
nand \U$44641 ( \44984 , \44983 , \43703 );
not \U$44642 ( \44985 , \44984 );
and \U$44643 ( \44986 , \44981 , \44985 );
and \U$44644 ( \44987 , \44756 , \44984 );
nor \U$44645 ( \44988 , \44986 , \44987 );
and \U$44646 ( \44989 , \44312 , \44988 );
not \U$44647 ( \44990 , \44312 );
and \U$44648 ( \44991 , \44990 , \1425 );
nor \U$44649 ( \44992 , \44989 , \44991 );
buf \U$44650 ( \44993 , \44992 );
buf \U$44651 ( \44994 , \43288 );
not \U$44652 ( \44995 , \44994 );
buf \U$44653 ( \44996 , \43241 );
buf \U$44654 ( \44997 , \43414 );
and \U$44655 ( \44998 , \44996 , \44997 );
not \U$44656 ( \44999 , \44998 );
and \U$44657 ( \45000 , \42647 , \43616 , \43631 , \43632 );
not \U$44658 ( \45001 , \45000 );
nand \U$44659 ( \45002 , \45001 , \43573 );
buf \U$44660 ( \45003 , \43647 );
buf \U$44661 ( \45004 , \43593 );
nand \U$44662 ( \45005 , \45002 , \45003 , \45004 );
not \U$44663 ( \45006 , \45005 );
or \U$44664 ( \45007 , \44999 , \45006 );
not \U$44665 ( \45008 , \43583 );
nand \U$44666 ( \45009 , \45007 , \45008 );
not \U$44667 ( \45010 , \45009 );
or \U$44668 ( \45011 , \44995 , \45010 );
nand \U$44669 ( \45012 , \45011 , \43588 );
nand \U$44670 ( \45013 , \43590 , \43600 );
and \U$44671 ( \45014 , \45012 , \45013 );
not \U$44672 ( \45015 , \45012 );
not \U$44673 ( \45016 , \45013 );
and \U$44674 ( \45017 , \45015 , \45016 );
nor \U$44675 ( \45018 , \45014 , \45017 );
or \U$44676 ( \45019 , \45018 , \44367 );
or \U$44677 ( \45020 , \44312 , \1111 );
nand \U$44678 ( \45021 , \45019 , \45020 );
buf \U$44679 ( \45022 , \45021 );
nand \U$44680 ( \45023 , \44994 , \43588 );
and \U$44681 ( \45024 , \45009 , \45023 );
not \U$44682 ( \45025 , \45009 );
not \U$44683 ( \45026 , \45023 );
and \U$44684 ( \45027 , \45025 , \45026 );
nor \U$44685 ( \45028 , \45024 , \45027 );
or \U$44686 ( \45029 , \45028 , \44585 );
or \U$44687 ( \45030 , \44312 , \1074 );
nand \U$44688 ( \45031 , \45029 , \45030 );
buf \U$44689 ( \45032 , \45031 );
not \U$44690 ( \45033 , \44997 );
not \U$44691 ( \45034 , \45005 );
or \U$44692 ( \45035 , \45033 , \45034 );
not \U$44693 ( \45036 , \43577 );
nand \U$44694 ( \45037 , \45035 , \45036 );
nand \U$44695 ( \45038 , \44996 , \43582 );
and \U$44696 ( \45039 , \45037 , \45038 );
not \U$44697 ( \45040 , \45037 );
not \U$44698 ( \45041 , \45038 );
and \U$44699 ( \45042 , \45040 , \45041 );
nor \U$44700 ( \45043 , \45039 , \45042 );
or \U$44701 ( \45044 , \45043 , \44585 );
or \U$44702 ( \45045 , \44312 , \1078 );
nand \U$44703 ( \45046 , \45044 , \45045 );
buf \U$44704 ( \45047 , \45046 );
nand \U$44705 ( \45048 , \45036 , \44997 );
and \U$44706 ( \45049 , \45005 , \45048 );
not \U$44707 ( \45050 , \45005 );
not \U$44708 ( \45051 , \45048 );
and \U$44709 ( \45052 , \45050 , \45051 );
nor \U$44710 ( \45053 , \45049 , \45052 );
or \U$44711 ( \45054 , \45053 , \44367 );
or \U$44712 ( \45055 , \44312 , \784 );
nand \U$44713 ( \45056 , \45054 , \45055 );
buf \U$44714 ( \45057 , \45056 );
buf \U$44715 ( \45058 , \43566 );
not \U$44716 ( \45059 , \45058 );
buf \U$44717 ( \45060 , \43535 );
not \U$44718 ( \45061 , \45060 );
not \U$44719 ( \45062 , \43489 );
nor \U$44720 ( \45063 , \45000 , \45062 );
not \U$44721 ( \45064 , \45063 );
or \U$44722 ( \45065 , \45061 , \45064 );
not \U$44723 ( \45066 , \43642 );
nand \U$44724 ( \45067 , \45065 , \45066 );
not \U$44725 ( \45068 , \45067 );
or \U$44726 ( \45069 , \45059 , \45068 );
nand \U$44727 ( \45070 , \45069 , \43645 );
nand \U$44728 ( \45071 , \43571 , \45004 );
and \U$44729 ( \45072 , \45070 , \45071 );
not \U$44730 ( \45073 , \45070 );
not \U$44731 ( \45074 , \45071 );
and \U$44732 ( \45075 , \45073 , \45074 );
nor \U$44733 ( \45076 , \45072 , \45075 );
or \U$44734 ( \45077 , \45076 , \44367 );
or \U$44735 ( \45078 , \44312 , \2080 );
nand \U$44736 ( \45079 , \45077 , \45078 );
buf \U$44737 ( \45080 , \45079 );
nand \U$44738 ( \45081 , \43645 , \45058 );
and \U$44739 ( \45082 , \45067 , \45081 );
not \U$44740 ( \45083 , \45067 );
not \U$44741 ( \45084 , \45081 );
and \U$44742 ( \45085 , \45083 , \45084 );
nor \U$44743 ( \45086 , \45082 , \45085 );
or \U$44744 ( \45087 , \45086 , \44367 );
or \U$44745 ( \45088 , \44312 , \2067 );
nand \U$44746 ( \45089 , \45087 , \45088 );
buf \U$44747 ( \45090 , \45089 );
not \U$44748 ( \45091 , \43489 );
not \U$44749 ( \45092 , \45001 );
or \U$44750 ( \45093 , \45091 , \45092 );
not \U$44751 ( \45094 , \43637 );
nand \U$44752 ( \45095 , \45093 , \45094 );
nand \U$44753 ( \45096 , \43641 , \45060 );
and \U$44754 ( \45097 , \45095 , \45096 );
not \U$44755 ( \45098 , \45095 );
not \U$44756 ( \45099 , \45096 );
and \U$44757 ( \45100 , \45098 , \45099 );
nor \U$44758 ( \45101 , \45097 , \45100 );
or \U$44759 ( \45102 , \45101 , \44585 );
or \U$44760 ( \45103 , \44312 , \3154 );
nand \U$44761 ( \45104 , \45102 , \45103 );
buf \U$44762 ( \45105 , \45104 );
not \U$44763 ( \45106 , \45094 );
nor \U$44764 ( \45107 , \45106 , \45062 );
and \U$44765 ( \45108 , \45107 , \45000 );
not \U$44766 ( \45109 , \45107 );
and \U$44767 ( \45110 , \45109 , \45001 );
nor \U$44768 ( \45111 , \45108 , \45110 );
or \U$44769 ( \45112 , \45111 , \44288 );
or \U$44770 ( \45113 , \44312 , \3155 );
nand \U$44771 ( \45114 , \45112 , \45113 );
buf \U$44772 ( \45115 , \45114 );
not \U$44773 ( \45116 , \37310 );
not \U$44774 ( \45117 , \43615 );
nand \U$44775 ( \45118 , \42448 , \42646 );
nand \U$44776 ( \45119 , \45117 , \45118 );
buf \U$44777 ( \45120 , \37763 );
nand \U$44778 ( \45121 , \45119 , \45120 );
buf \U$44779 ( \45122 , \37725 );
not \U$44780 ( \45123 , \45122 );
or \U$44781 ( \45124 , \45121 , \45123 );
not \U$44782 ( \45125 , \43626 );
nand \U$44783 ( \45126 , \45124 , \45125 );
not \U$44784 ( \45127 , \45126 );
or \U$44785 ( \45128 , \45116 , \45127 );
nand \U$44786 ( \45129 , \45128 , \43617 );
not \U$44787 ( \45130 , \45129 );
not \U$44788 ( \45131 , \43632 );
not \U$44789 ( \45132 , \45131 );
nand \U$44790 ( \45133 , \45132 , \43630 );
not \U$44791 ( \45134 , \45133 );
and \U$44792 ( \45135 , \45130 , \45134 );
and \U$44793 ( \45136 , \45129 , \45133 );
nor \U$44794 ( \45137 , \45135 , \45136 );
or \U$44795 ( \45138 , \45137 , \44288 );
or \U$44796 ( \45139 , \44312 , \3593 );
nand \U$44797 ( \45140 , \45138 , \45139 );
buf \U$44798 ( \45141 , \45140 );
not \U$44799 ( \45142 , \45126 );
nand \U$44800 ( \45143 , \43617 , \37310 );
not \U$44801 ( \45144 , \45143 );
and \U$44802 ( \45145 , \45142 , \45144 );
and \U$44803 ( \45146 , \45126 , \45143 );
nor \U$44804 ( \45147 , \45145 , \45146 );
or \U$44805 ( \45148 , \45147 , \44367 );
or \U$44806 ( \45149 , \44311 , \3455 );
nand \U$44807 ( \45150 , \45148 , \45149 );
buf \U$44808 ( \45151 , \45150 );
not \U$44809 ( \45152 , \43619 );
nand \U$44810 ( \45153 , \45121 , \45152 );
nand \U$44811 ( \45154 , \43625 , \45122 );
and \U$44812 ( \45155 , \45153 , \45154 );
not \U$44813 ( \45156 , \45153 );
not \U$44814 ( \45157 , \45154 );
and \U$44815 ( \45158 , \45156 , \45157 );
nor \U$44816 ( \45159 , \45155 , \45158 );
not \U$44817 ( \45160 , \44312 );
or \U$44818 ( \45161 , \45159 , \45160 );
or \U$44819 ( \45162 , \44311 , \4088 );
nand \U$44820 ( \45163 , \45161 , \45162 );
buf \U$44821 ( \45164 , \45163 );
nand \U$44822 ( \45165 , \45120 , \45152 );
and \U$44823 ( \45166 , \45119 , \45165 );
not \U$44824 ( \45167 , \45119 );
not \U$44825 ( \45168 , \45165 );
and \U$44826 ( \45169 , \45167 , \45168 );
nor \U$44827 ( \45170 , \45166 , \45169 );
or \U$44828 ( \45171 , \45170 , \44288 );
or \U$44829 ( \45172 , \44311 , \4081 );
nand \U$44830 ( \45173 , \45171 , \45172 );
buf \U$44831 ( \45174 , \45173 );
not \U$44832 ( \45175 , \42585 );
nand \U$44833 ( \45176 , \42448 , \42630 );
buf \U$44834 ( \45177 , \42620 );
not \U$44835 ( \45178 , \45177 );
or \U$44836 ( \45179 , \45176 , \45178 );
nand \U$44837 ( \45180 , \43607 , \45177 );
nand \U$44838 ( \45181 , \45179 , \45180 );
not \U$44839 ( \45182 , \45181 );
or \U$44840 ( \45183 , \45175 , \45182 );
nand \U$44841 ( \45184 , \45183 , \43610 );
not \U$44842 ( \45185 , \45184 );
not \U$44843 ( \45186 , \43613 );
nand \U$44844 ( \45187 , \45186 , \42645 );
not \U$44845 ( \45188 , \45187 );
and \U$44846 ( \45189 , \45185 , \45188 );
and \U$44847 ( \45190 , \45184 , \45187 );
nor \U$44848 ( \45191 , \45189 , \45190 );
or \U$44849 ( \45192 , \45191 , \45160 );
or \U$44850 ( \45193 , \44312 , \4902 );
nand \U$44851 ( \45194 , \45192 , \45193 );
buf \U$44852 ( \45195 , \45194 );
not \U$44853 ( \45196 , \45181 );
nand \U$44854 ( \45197 , \42585 , \43610 );
not \U$44855 ( \45198 , \45197 );
and \U$44856 ( \45199 , \45196 , \45198 );
and \U$44857 ( \45200 , \45181 , \45197 );
nor \U$44858 ( \45201 , \45199 , \45200 );
or \U$44859 ( \45202 , \45201 , \44288 );
or \U$44860 ( \45203 , \44311 , \4908 );
nand \U$44861 ( \45204 , \45202 , \45203 );
buf \U$44862 ( \45205 , \45204 );
nand \U$44863 ( \45206 , \45176 , \43606 );
not \U$44864 ( \45207 , \42618 );
not \U$44865 ( \45208 , \42587 );
or \U$44866 ( \45209 , \45207 , \45208 );
nand \U$44867 ( \45210 , \45209 , \45177 );
and \U$44868 ( \45211 , \45206 , \45210 );
not \U$44869 ( \45212 , \45206 );
not \U$44870 ( \45213 , \45210 );
and \U$44871 ( \45214 , \45212 , \45213 );
nor \U$44872 ( \45215 , \45211 , \45214 );
or \U$44873 ( \45216 , \45215 , \44288 );
or \U$44874 ( \45217 , \44311 , \5025 );
nand \U$44875 ( \45218 , \45216 , \45217 );
buf \U$44876 ( \45219 , \45218 );
nand \U$44877 ( \45220 , \43606 , \42630 );
xor \U$44878 ( \45221 , \42448 , \45220 );
or \U$44879 ( \45222 , \45221 , \44288 );
not \U$44880 ( \45223 , \44288 );
or \U$44881 ( \45224 , \45223 , \5026 );
nand \U$44882 ( \45225 , \45222 , \45224 );
buf \U$44883 ( \45226 , \45225 );
not \U$44884 ( \45227 , \39720 );
not \U$44885 ( \45228 , \42445 );
buf \U$44886 ( \45229 , \42443 );
not \U$44887 ( \45230 , \45229 );
or \U$44888 ( \45231 , \45228 , \45230 );
not \U$44889 ( \45232 , \39710 );
nand \U$44890 ( \45233 , \45231 , \45232 );
not \U$44891 ( \45234 , \45233 );
or \U$44892 ( \45235 , \45227 , \45234 );
buf \U$44893 ( \45236 , \39723 );
nand \U$44894 ( \45237 , \45235 , \45236 );
not \U$44895 ( \45238 , \45237 );
nand \U$44896 ( \45239 , \39727 , \38887 );
not \U$44897 ( \45240 , \45239 );
and \U$44898 ( \45241 , \45238 , \45240 );
and \U$44899 ( \45242 , \45237 , \45239 );
nor \U$44900 ( \45243 , \45241 , \45242 );
or \U$44901 ( \45244 , \45243 , \44288 );
or \U$44902 ( \45245 , \44311 , \5644 );
nand \U$44903 ( \45246 , \45244 , \45245 );
buf \U$44904 ( \45247 , \45246 );
and \U$44905 ( \45248 , \44288 , \5631 );
not \U$44906 ( \45249 , \44288 );
not \U$44907 ( \45250 , \45233 );
nand \U$44908 ( \45251 , \39720 , \45236 );
not \U$44909 ( \45252 , \45251 );
and \U$44910 ( \45253 , \45250 , \45252 );
and \U$44911 ( \45254 , \45233 , \45251 );
nor \U$44912 ( \45255 , \45253 , \45254 );
and \U$44913 ( \45256 , \45249 , \45255 );
nor \U$44914 ( \45257 , \45248 , \45256 );
buf \U$44915 ( \45258 , \45257 );
buf \U$44916 ( \45259 , \42444 );
not \U$44917 ( \45260 , \45259 );
not \U$44918 ( \45261 , \45229 );
or \U$44919 ( \45262 , \45260 , \45261 );
not \U$44920 ( \45263 , \39671 );
nand \U$44921 ( \45264 , \45262 , \45263 );
nand \U$44922 ( \45265 , \39709 , \39704 );
and \U$44923 ( \45266 , \45264 , \45265 );
not \U$44924 ( \45267 , \45264 );
not \U$44925 ( \45268 , \45265 );
and \U$44926 ( \45269 , \45267 , \45268 );
nor \U$44927 ( \45270 , \45266 , \45269 );
or \U$44928 ( \45271 , \45270 , \44288 );
or \U$44929 ( \45272 , \45223 , \5632 );
nand \U$44930 ( \45273 , \45271 , \45272 );
buf \U$44931 ( \45274 , \45273 );
and \U$44932 ( \45275 , \44288 , \6279 );
not \U$44933 ( \45276 , \44288 );
nand \U$44934 ( \45277 , \45263 , \45259 );
and \U$44935 ( \45278 , \45229 , \45277 );
not \U$44936 ( \45279 , \45229 );
not \U$44937 ( \45280 , \45277 );
and \U$44938 ( \45281 , \45279 , \45280 );
nor \U$44939 ( \45282 , \45278 , \45281 );
and \U$44940 ( \45283 , \45276 , \45282 );
nor \U$44941 ( \45284 , \45275 , \45283 );
buf \U$44942 ( \45285 , \45284 );
not \U$44943 ( \45286 , \40112 );
not \U$44944 ( \45287 , \42440 );
buf \U$44945 ( \45288 , \42438 );
not \U$44946 ( \45289 , \45288 );
or \U$44947 ( \45290 , \45287 , \45289 );
not \U$44948 ( \45291 , \40398 );
nand \U$44949 ( \45292 , \45290 , \45291 );
not \U$44950 ( \45293 , \45292 );
or \U$44951 ( \45294 , \45286 , \45293 );
buf \U$44952 ( \45295 , \40401 );
nand \U$44953 ( \45296 , \45294 , \45295 );
not \U$44954 ( \45297 , \42442 );
not \U$44955 ( \45298 , \45297 );
nand \U$44956 ( \45299 , \45298 , \40412 );
xor \U$44957 ( \45300 , \45296 , \45299 );
or \U$44958 ( \45301 , \45300 , \44288 );
or \U$44959 ( \45302 , \45223 , \7333 );
nand \U$44960 ( \45303 , \45301 , \45302 );
buf \U$44961 ( \45304 , \45303 );
not \U$44962 ( \45305 , \45292 );
nand \U$44963 ( \45306 , \45295 , \40112 );
not \U$44964 ( \45307 , \45306 );
and \U$44965 ( \45308 , \45305 , \45307 );
and \U$44966 ( \45309 , \45292 , \45306 );
nor \U$44967 ( \45310 , \45308 , \45309 );
or \U$44968 ( \45311 , \45310 , \44288 );
or \U$44969 ( \45312 , \44311 , \7316 );
nand \U$44970 ( \45313 , \45311 , \45312 );
buf \U$44971 ( \45314 , \45313 );
not \U$44972 ( \45315 , \42439 );
not \U$44973 ( \45316 , \45288 );
or \U$44974 ( \45317 , \45315 , \45316 );
not \U$44975 ( \45318 , \40394 );
nand \U$44976 ( \45319 , \45317 , \45318 );
nand \U$44977 ( \45320 , \40397 , \40302 );
xor \U$44978 ( \45321 , \45319 , \45320 );
or \U$44979 ( \45322 , \45321 , \44288 );
or \U$44980 ( \45323 , \45223 , \8031 );
nand \U$44981 ( \45324 , \45322 , \45323 );
buf \U$44982 ( \45325 , \45324 );
and \U$44983 ( \45326 , \44288 , \8017 );
not \U$44984 ( \45327 , \44288 );
not \U$44985 ( \45328 , \40394 );
nand \U$44986 ( \45329 , \45328 , \42439 );
xor \U$44987 ( \45330 , \45288 , \45329 );
and \U$44988 ( \45331 , \45327 , \45330 );
nor \U$44989 ( \45332 , \45326 , \45331 );
buf \U$44990 ( \45333 , \45332 );
not \U$44991 ( \45334 , \41111 );
not \U$44992 ( \45335 , \41084 );
buf \U$44993 ( \45336 , \42422 );
not \U$44994 ( \45337 , \45336 );
or \U$44995 ( \45338 , \45335 , \45337 );
not \U$44996 ( \45339 , \42429 );
nand \U$44997 ( \45340 , \45338 , \45339 );
not \U$44998 ( \45341 , \45340 );
or \U$44999 ( \45342 , \45334 , \45341 );
nand \U$45000 ( \45343 , \45342 , \42433 );
not \U$45001 ( \45344 , \45343 );
nand \U$45002 ( \45345 , \41118 , \42437 );
not \U$45003 ( \45346 , \45345 );
and \U$45004 ( \45347 , \45344 , \45346 );
and \U$45005 ( \45348 , \45343 , \45345 );
nor \U$45006 ( \45349 , \45347 , \45348 );
or \U$45007 ( \45350 , \45349 , \44288 );
or \U$45008 ( \45351 , \45223 , \9198 );
nand \U$45009 ( \45352 , \45350 , \45351 );
buf \U$45010 ( \45353 , \45352 );
not \U$45011 ( \45354 , \45340 );
not \U$45012 ( \45355 , \42433 );
not \U$45013 ( \45356 , \45355 );
nand \U$45014 ( \45357 , \45356 , \41111 );
not \U$45015 ( \45358 , \45357 );
and \U$45016 ( \45359 , \45354 , \45358 );
and \U$45017 ( \45360 , \45340 , \45357 );
nor \U$45018 ( \45361 , \45359 , \45360 );
or \U$45019 ( \45362 , \45361 , \44288 );
or \U$45020 ( \45363 , \44311 , \9186 );
nand \U$45021 ( \45364 , \45362 , \45363 );
buf \U$45022 ( \45365 , \45364 );
not \U$45023 ( \45366 , \41083 );
not \U$45024 ( \45367 , \45336 );
or \U$45025 ( \45368 , \45366 , \45367 );
not \U$45026 ( \45369 , \42424 );
nand \U$45027 ( \45370 , \45368 , \45369 );
not \U$45028 ( \45371 , \45370 );
not \U$45029 ( \45372 , \40955 );
not \U$45030 ( \45373 , \45372 );
nand \U$45031 ( \45374 , \45373 , \42428 );
not \U$45032 ( \45375 , \45374 );
and \U$45033 ( \45376 , \45371 , \45375 );
and \U$45034 ( \45377 , \45370 , \45374 );
nor \U$45035 ( \45378 , \45376 , \45377 );
or \U$45036 ( \45379 , \45378 , \44288 );
or \U$45037 ( \45380 , \45223 , \9185 );
nand \U$45038 ( \45381 , \45379 , \45380 );
buf \U$45039 ( \45382 , \45381 );
not \U$45040 ( \45383 , \42424 );
nand \U$45041 ( \45384 , \45383 , \41083 );
xor \U$45042 ( \45385 , \45336 , \45384 );
or \U$45043 ( \45386 , \45385 , \44288 );
or \U$45044 ( \45387 , \44287 , \9243 );
nand \U$45045 ( \45388 , \45386 , \45387 );
buf \U$45046 ( \45389 , \45388 );
not \U$45047 ( \45390 , \41573 );
not \U$45048 ( \45391 , \42418 );
not \U$45049 ( \45392 , \45391 );
not \U$45050 ( \45393 , \42415 );
or \U$45051 ( \45394 , \45392 , \45393 );
not \U$45052 ( \45395 , \41572 );
nand \U$45053 ( \45396 , \45394 , \45395 );
not \U$45054 ( \45397 , \45396 );
or \U$45055 ( \45398 , \45390 , \45397 );
nand \U$45056 ( \45399 , \45398 , \41359 );
not \U$45057 ( \45400 , \45399 );
not \U$45058 ( \45401 , \42421 );
not \U$45059 ( \45402 , \45401 );
nand \U$45060 ( \45403 , \45402 , \41588 );
not \U$45061 ( \45404 , \45403 );
and \U$45062 ( \45405 , \45400 , \45404 );
and \U$45063 ( \45406 , \45399 , \45403 );
nor \U$45064 ( \45407 , \45405 , \45406 );
or \U$45065 ( \45408 , \45407 , \44288 );
or \U$45066 ( \45409 , \45223 , \8807 );
nand \U$45067 ( \45410 , \45408 , \45409 );
buf \U$45068 ( \45411 , \45410 );
not \U$45069 ( \45412 , \45396 );
not \U$45070 ( \45413 , \42416 );
nand \U$45071 ( \45414 , \45413 , \41359 );
not \U$45072 ( \45415 , \45414 );
and \U$45073 ( \45416 , \45412 , \45415 );
and \U$45074 ( \45417 , \45396 , \45414 );
nor \U$45075 ( \45418 , \45416 , \45417 );
or \U$45076 ( \45419 , \45418 , \44288 );
or \U$45077 ( \45420 , \44287 , \8797 );
nand \U$45078 ( \45421 , \45419 , \45420 );
buf \U$45079 ( \45422 , \45421 );
not \U$45080 ( \45423 , \42417 );
not \U$45081 ( \45424 , \42415 );
or \U$45082 ( \45425 , \45423 , \45424 );
not \U$45083 ( \45426 , \41558 );
nand \U$45084 ( \45427 , \45425 , \45426 );
not \U$45085 ( \45428 , \45427 );
nand \U$45086 ( \45429 , \41571 , \41568 );
not \U$45087 ( \45430 , \45429 );
and \U$45088 ( \45431 , \45428 , \45430 );
and \U$45089 ( \45432 , \45427 , \45429 );
nor \U$45090 ( \45433 , \45431 , \45432 );
or \U$45091 ( \45434 , \45433 , \44288 );
or \U$45092 ( \45435 , \44287 , \9690 );
nand \U$45093 ( \45436 , \45434 , \45435 );
buf \U$45094 ( \45437 , \45436 );
not \U$45095 ( \45438 , \41558 );
nand \U$45096 ( \45439 , \45438 , \42417 );
xor \U$45097 ( \45440 , \42415 , \45439 );
or \U$45098 ( \45441 , \45440 , \44288 );
or \U$45099 ( \45442 , \44287 , \9290 );
nand \U$45100 ( \45443 , \45441 , \45442 );
buf \U$45101 ( \45444 , \45443 );
buf \U$45102 ( \45445 , \42410 );
not \U$45103 ( \45446 , \45445 );
not \U$45104 ( \45447 , \42413 );
nand \U$45105 ( \45448 , \45447 , \41678 );
not \U$45106 ( \45449 , \45448 );
and \U$45107 ( \45450 , \45446 , \45449 );
and \U$45108 ( \45451 , \45445 , \45448 );
nor \U$45109 ( \45452 , \45450 , \45451 );
or \U$45110 ( \45453 , \45452 , \44288 );
or \U$45111 ( \45454 , \44287 , \8732 );
nand \U$45112 ( \45455 , \45453 , \45454 );
buf \U$45113 ( \45456 , \45455 );
nand \U$45114 ( \45457 , \42409 , \41782 );
xor \U$45115 ( \45458 , \45457 , \42404 );
or \U$45116 ( \45459 , \45458 , \44288 );
or \U$45117 ( \45460 , \44287 , \8733 );
nand \U$45118 ( \45461 , \45459 , \45460 );
buf \U$45119 ( \45462 , \45461 );
nand \U$45120 ( \45463 , \42403 , \41859 );
xor \U$45121 ( \45464 , \45463 , \42399 );
or \U$45122 ( \45465 , \45464 , \44288 );
or \U$45123 ( \45466 , \44287 , \17560 );
nand \U$45124 ( \45467 , \45465 , \45466 );
buf \U$45125 ( \45468 , \45467 );
nand \U$45126 ( \45469 , \42398 , \42393 );
xor \U$45127 ( \45470 , \45469 , \42373 );
or \U$45128 ( \45471 , \45470 , \44288 );
or \U$45129 ( \45472 , \44287 , \9947 );
nand \U$45130 ( \45473 , \45471 , \45472 );
buf \U$45131 ( \45474 , \45473 );
nand \U$45132 ( \45475 , \42372 , \41995 );
xor \U$45133 ( \45476 , \45475 , \42368 );
or \U$45134 ( \45477 , \45476 , \44288 );
or \U$45135 ( \45478 , \44287 , \13022 );
nand \U$45136 ( \45479 , \45477 , \45478 );
buf \U$45137 ( \45480 , \45479 );
not \U$45138 ( \45481 , RI9873198_182);
not \U$45139 ( \45482 , \44288 );
or \U$45140 ( \45483 , \45481 , \45482 );
nand \U$45141 ( \45484 , \42060 , \42367 );
not \U$45142 ( \45485 , \45484 );
not \U$45143 ( \45486 , \42364 );
and \U$45144 ( \45487 , \45485 , \45486 );
and \U$45145 ( \45488 , \42364 , \45484 );
nor \U$45146 ( \45489 , \45487 , \45488 );
or \U$45147 ( \45490 , \45489 , \44288 );
nand \U$45148 ( \45491 , \45483 , \45490 );
buf \U$45149 ( \45492 , \45491 );
endmodule

