//
// Conformal-LEC Version 20.10-d214 (03-Sep-2020)
//
module top(RIaa97c98_14,RIaa9e7f0_243,RIaa9e868_244,RIaa9e778_242,RIaa9e9d0_247,RIaa97d88_16,RIaa97d10_15,RIaa97e00_17,RIaa97c20_13,
        RIaa9e688_240,RIaa9e700_241,RIaa9e8e0_245,RIaa9e958_246,RIaa9cf90_191,RIaa9d170_195,RIaa9cea0_189,RIaa9d1e8_196,RIaa9d080_193,RIaa9d0f8_194,
        RIaa9d5a8_204,RIaa9d620_205,RIaa9d2d8_198,RIaa9d008_192,RIaa9d3c8_200,RIaa9d4b8_202,RIaa9d260_197,RIaa9d350_199,RIaa9cf18_190,RIaa9d530_203,
        RIaa9d440_201,RIaa97860_5,RIaa976f8_2,RIaa97770_3,RIaa977e8_4,RIaa9ba00_145,RIaa9b640_137,RIaa9b910_143,RIaa9bd48_152,RIaa9ba78_146,
        RIaa9bb68_148,RIaa9b7a8_140,RIaa9bdc0_153,RIaa9baf0_147,RIaa9b730_139,RIaa9bc58_150,RIaa9b6b8_138,RIaa9b898_142,RIaa9bcd0_151,RIaa9b988_144,
        RIaa9b820_141,RIaa9bbe0_149,RIaa9b370_131,RIaa9b0a0_125,RIaa9b5c8_136,RIaa9b3e8_132,RIaa9ae48_120,RIaa9b460_133,RIaa9b190_127,RIaa9b118_126,
        RIaa9b4d8_134,RIaa9b280_129,RIaa9b028_124,RIaa9af38_122,RIaa9b2f8_130,RIaa9aec0_121,RIaa9b550_135,RIaa9afb0_123,RIaa9b208_128,RIaa9c2e8_164,
        RIaa9c4c8_168,RIaa9c018_158,RIaa9c3d8_166,RIaa9c450_167,RIaa9be38_154,RIaa9bfa0_157,RIaa9beb0_155,RIaa9c270_163,RIaa9c090_159,RIaa9c108_160,
        RIaa9c180_161,RIaa9bf28_156,RIaa9c5b8_170,RIaa9c1f8_162,RIaa9c360_165,RIaa9c540_169,RIaa9ce28_188,RIaa9c978_178,RIaa9c9f0_179,RIaa9c900_177,
        RIaa9cdb0_187,RIaa9c810_175,RIaa9c720_173,RIaa9cb58_182,RIaa9cae0_181,RIaa9c630_171,RIaa9ca68_180,RIaa9cc48_184,RIaa9ccc0_185,RIaa9c888_176,
        RIaa9c6a8_172,RIaa9c798_174,RIaa9cbd0_183,RIaa9cd38_186,RIaa9ab78_114,RIaa9aa10_111,RIaa9ac68_116,RIaa9a7b8_106,RIaa9a6c8_104,RIaa9add0_119,
        RIaa9abf0_115,RIaa9a8a8_108,RIaa9a998_110,RIaa9a920_109,RIaa9a830_107,RIaa9ad58_118,RIaa9a740_105,RIaa9ab00_113,RIaa9aa88_112,RIaa9a650_103,
        RIaa9ace0_117,RIaa978d8_6,RIaa9a308_96,RIaa9a218_94,RIaa9a380_97,RIaa9a038_90,RIaa99ed0_87,RIaa9a290_95,RIaa9a0b0_91,RIaa99fc0_89,
        RIaa9a470_99,RIaa99f48_88,RIaa9a4e8_100,RIaa9a1a0_93,RIaa9a3f8_98,RIaa99e58_86,RIaa9a560_101,RIaa9a128_92,RIaa9a5d8_102,RIaa97950_7,
        RIaa99b10_79,RIaa999a8_76,RIaa99a20_77,RIaa996d8_70,RIaa99930_75,RIaa99d68_84,RIaa99b88_80,RIaa99660_69,RIaa99cf0_83,RIaa99c00_81,
        RIaa998b8_74,RIaa99de0_85,RIaa99a98_78,RIaa99c78_82,RIaa997c8_72,RIaa99840_73,RIaa99750_71,RIaa979c8_8,RIaa9f6f0_275,RIaa9f768_276,
        RIaa9f3a8_268,RIaa9f600_273,RIaa9f2b8_266,RIaa9f330_267,RIaa9f420_269,RIaa9f9c0_281,RIaa9f948_280,RIaa9f678_274,RIaa9f8d0_279,RIaa9f588_272,
        RIaa9f240_265,RIaa9f510_271,RIaa9f7e0_277,RIaa9f858_278,RIaa9f498_270,RIaa9eca0_253,RIaa9ee08_256,RIaa9eef8_258,RIaa9ed90_255,RIaa9f1c8_264,
        RIaa9efe8_260,RIaa9ef70_259,RIaa9ed18_254,RIaa9eb38_250,RIaa9ebb0_251,RIaa9ea48_248,RIaa9f0d8_262,RIaa9ee80_257,RIaa9eac0_249,RIaa9f150_263,
        RIaa9f060_261,RIaa9ec28_252,RIaa97b30_11,RIaa97ba8_12,RIaa9de18_222,RIaa9db48_216,RIaa9d968_212,RIaa9dbc0_217,RIaa9dda0_221,RIaa9dd28_220,
        RIaa9dad0_215,RIaa9d800_209,RIaa9dc38_218,RIaa9d710_207,RIaa9dcb0_219,RIaa9d788_208,RIaa9d698_206,RIaa9da58_214,RIaa9d9e0_213,RIaa9d878_210,
        RIaa9d8f0_211,RIaa994f8_66,RIaa99048_56,RIaa98f58_54,RIaa99570_67,RIaa990c0_57,RIaa99138_58,RIaa99390_63,RIaa98ee0_53,RIaa99480_65,
        RIaa98fd0_55,RIaa995e8_68,RIaa99318_62,RIaa991b0_59,RIaa99408_64,RIaa992a0_61,RIaa98e68_52,RIaa99228_60,RIaa9e160_229,RIaa9df80_225,
        RIaa9e3b8_234,RIaa9de90_223,RIaa9e610_239,RIaa9e2c8_232,RIaa9e598_238,RIaa9e1d8_230,RIaa9df08_224,RIaa9e520_237,RIaa9e340_233,RIaa9e250_231,
        RIaa9e430_235,RIaa9e0e8_228,RIaa9dff8_226,RIaa9e4a8_236,RIaa9e070_227,RIaa97ab8_10,RIaa97a40_9,RIaa98b20_45,RIaa989b8_42,RIaa98c88_48,
        RIaa98a30_43,RIaa98aa8_44,RIaa98df0_51,RIaa98940_41,RIaa98c10_47,RIaa98670_35,RIaa98850_39,RIaa98760_37,RIaa986e8_36,RIaa98d00_49,
        RIaa98b98_46,RIaa987d8_38,RIaa988c8_40,RIaa98d78_50,RIaaa1ce8_356,RIaaa1e50_359,RIaaa2030_363,RIaaa1fb8_362,RIaaa1f40_361,RIaaa1c70_355,
        RIaaa1d60_357,RIaaa1ec8_360,RIaaa1b80_353,RIaaa1bf8_354,RIaaa20a8_364,RIaaa1a90_351,RIaaa2120_365,RIaaa1dd8_358,RIaaa2198_366,RIaaa1b08_352,
        RIaaa1a18_350,RIaaa1130_331,RIaaa0f50_327,RIaaa0a28_316,RIaaa0b90_319,RIaaa0b18_318,RIaaa1040_329,RIaaa0c80_321,RIaaa0cf8_322,RIaaa0c08_320,
        RIaaa0ed8_326,RIaaa0d70_323,RIaaa0aa0_317,RIaaa0fc8_328,RIaaa11a8_332,RIaaa10b8_330,RIaaa0e60_325,RIaaa0de8_324,RIaa97680_1,RIaa98508_32,
        RIaa98328_28,RIaa98238_26,RIaa98418_30,RIaa97e78_18,RIaa981c0_25,RIaa985f8_34,RIaa982b0_27,RIaa98580_33,RIaa97ef0_19,RIaa98058_22,
        RIaa98148_24,RIaa97f68_20,RIaa97fe0_21,RIaa983a0_29,RIaa980d0_23,RIaa98490_31,RIaaa2cd8_390,RIaaa2af8_386,RIaaa3110_399,RIaaa3188_400,
        RIaaa2f30_395,RIaaa2c60_389,RIaaa2eb8_394,RIaaa2dc8_392,RIaaa2e40_393,RIaaa2fa8_396,RIaaa3020_397,RIaaa2a08_384,RIaaa3098_398,RIaaa2be8_388,
        RIaaa2b70_387,RIaaa2a80_385,RIaaa2d50_391,RIaaa1298_334,RIaaa16d0_343,RIaaa1928_348,RIaaa1658_342,RIaaa1838_346,RIaaa14f0_339,RIaaa1388_336,
        RIaaa1400_337,RIaaa19a0_349,RIaaa1748_344,RIaaa15e0_341,RIaaa1310_335,RIaaa1220_333,RIaaa1478_338,RIaaa1568_340,RIaaa17c0_345,RIaaa18b0_347,
        RIaa9ff60_293,RIaa9fba0_285,RIaa9fa38_282,RIaaa0050_295,RIaa9ffd8_294,RIaa9fe70_291,RIaa9fc90_287,RIaaa01b8_298,RIaaa0140_297,RIaa9fdf8_290,
        RIaa9fab0_283,RIaa9fc18_286,RIaa9fb28_284,RIaa9fd08_288,RIaaa00c8_296,RIaa9fee8_292,RIaa9fd80_289,RIaaa05f0_307,RIaaa0938_314,RIaaa0758_310,
        RIaaa0488_304,RIaaa0578_306,RIaaa0230_299,RIaaa06e0_309,RIaaa0848_312,RIaaa0398_302,RIaaa0320_301,RIaaa0668_308,RIaaa0410_303,RIaaa02a8_300,
        RIaaa08c0_313,RIaaa0500_305,RIaaa07d0_311,RIaaa09b0_315,RIaaa24e0_373,RIaaa2558_374,RIaaa2738_378,RIaaa2828_380,RIaaa2300_369,RIaaa26c0_377,
        RIaaa2918_382,RIaaa2468_372,RIaaa2378_370,RIaaa2288_368,RIaaa2648_376,RIaaa23f0_371,RIaaa2210_367,RIaaa25d0_375,RIaaa27b0_379,RIaaa28a0_381,
        RIaaa2990_383,RIaaa3f20_429,RIaaa3f98_430,RIaaa3cc8_424,RIaaa3c50_423,RIaaa4010_431,RIaaa4100_433,RIaaa3db8_426,RIaaa3b60_421,RIaaa3d40_425,
        RIaaa3ae8_420,RIaaa3a70_419,RIaaa39f8_418,RIaaa4178_434,RIaaa3e30_427,RIaaa3bd8_422,RIaaa4088_432,RIaaa3ea8_428,RIaaa32f0_403,RIaaa3890_415,
        RIaaa34d0_407,RIaaa3638_410,RIaaa3728_412,RIaaa35c0_409,RIaaa3278_402,RIaaa3818_414,RIaaa33e0_405,RIaaa3368_404,RIaaa37a0_413,RIaaa3980_417,
        RIaaa3908_416,RIaaa36b0_411,RIaaa3458_406,RIaaa3548_408,RIaaa3200_401,RIaaa4448_440,RIaaa4538_442,RIaaa4268_436,RIaaa43d0_439,RIaaa42e0_437,
        RIaaa41f0_435,RIaaa4628_444,RIaaa4808_448,RIaaa45b0_443,RIaaa4718_446,RIaaa44c0_441,RIaaa48f8_450,RIaaa4358_438,RIaaa4970_451,RIaaa4880_449,
        RIaaa4790_447,RIaaa46a0_445,RIaaa6248_504,RIaaa66f8_514,RIaaa6860_517,RIaaa67e8_516,RIaaa6680_513,RIaaa64a0_509,RIaaa6338_506,RIaaa63b0_507,
        RIaaa6950_519,RIaaa6608_512,RIaaa6590_511,RIaaa6428_508,RIaaa6770_515,RIaaa68d8_518,RIaaa6518_510,RIaaa62c0_505,RIaaa61d0_503,RIaaa57f8_482,
        RIaaa54b0_475,RIaaa5618_478,RIaaa52d0_471,RIaaa5528_476,RIaaa5258_470,RIaaa5708_480,RIaaa5690_479,RIaaa5348_472,RIaaa53c0_473,RIaaa58e8_484,
        RIaaa5960_485,RIaaa5780_481,RIaaa5438_474,RIaaa5870_483,RIaaa55a0_477,RIaaa51e0_469,RIaaa4e98_462,RIaaa49e8_452,RIaaa4b50_455,RIaaa4e20_461,
        RIaaa50f0_467,RIaaa4f88_464,RIaaa5000_465,RIaaa4c40_457,RIaaa4cb8_458,RIaaa4a60_453,RIaaa4f10_463,RIaaa4bc8_456,RIaaa4ad8_454,RIaaa5168_468,
        RIaaa4d30_459,RIaaa4da8_460,RIaaa5078_466,RIaaa5e10_495,RIaaa5ca8_492,RIaaa59d8_486,RIaaa60e0_501,RIaaa5b40_489,RIaaa5a50_487,RIaaa5f00_497,
        RIaaa5bb8_490,RIaaa6158_502,RIaaa5f78_498,RIaaa5ac8_488,RIaaa5e88_496,RIaaa5d98_494,RIaaa5ff0_499,RIaaa5d20_493,RIaaa6068_500,RIaaa5c30_491,
        RIaaa6d10_527,RIaaa6a40_521,RIaaa7058_534,RIaaa7148_536,RIaaa6e00_529,RIaaa6ba8_524,RIaaa6e78_530,RIaaa6c98_526,RIaaa6f68_532,RIaaa6ab8_522,
        RIaaa70d0_535,RIaaa6c20_525,RIaaa69c8_520,RIaaa6d88_528,RIaaa6fe0_533,RIaaa6ef0_531,RIaaa6b30_523,RIaaa8408_576,RIaaa87c8_584,RIaaa84f8_578,
        RIaaa8390_575,RIaaa8318_574,RIaaa8660_581,RIaaa8228_572,RIaaa88b8_586,RIaaa8930_587,RIaaa8750_583,RIaaa8480_577,RIaaa8840_585,RIaaa86d8_582,
        RIaaa85e8_580,RIaaa8570_579,RIaaa82a0_573,RIaaa81b0_571,RIaaa7670_547,RIaaa7238_538,RIaaa7490_543,RIaaa75f8_546,RIaaa78c8_552,RIaaa7328_540,
        RIaaa73a0_541,RIaaa77d8_550,RIaaa7850_551,RIaaa76e8_548,RIaaa7580_545,RIaaa72b0_539,RIaaa71c0_537,RIaaa7508_544,RIaaa7418_542,RIaaa7940_553,
        RIaaa7760_549,RIaaa7d00_561,RIaaa7f58_566,RIaaa7fd0_567,RIaaa7b98_558,RIaaa7b20_557,RIaaa7df0_563,RIaaa7c88_560,RIaaa7e68_564,RIaaa7ee0_565,
        RIaaa7d78_562,RIaaa8048_568,RIaaa7c10_559,RIaaa8138_570,RIaaa80c0_569,RIaaa7aa8_556,RIaaa7a30_555,RIaaa79b8_554,RIaaa89a8_588,RIaaa95d8_614,
        RIaaa9218_606,RIaaa90b0_603,RIaaa9128_604,RIaaa91a0_605,RIaaa9380_609,RIaaa9308_608,RIaaa9290_607,RIaaa9038_602,RIaaa93f8_610,RIaaa9470_611,
        RIaaa94e8_612,RIaaa8c78_594,RIaaa8cf0_595,RIaaa8a98_590,RIaaa8b10_591,RIaaa8a20_589,RIaaa8b88_592,RIaaa8c00_593,RIaaa8d68_596,RIaaa8de0_597,
        RIaaa8e58_598,RIaaa8ed0_599,RIaaa8f48_600,RIaaa8fc0_601,RIaaa9560_613,R_267_b0ecd58,R_268_b0ece00,R_269_b0ecea8,R_26a_b0ecf50,R_26b_b0ecff8,
        R_26c_b0ed0a0,R_26d_b0ed148,R_26e_b0ed1f0,R_26f_b0ed298,R_270_b0ed340,R_271_b0ed3e8,R_272_b0ed490,R_273_b0ed538,R_274_b0ed5e0,R_275_b0ed688,
        R_276_b0ed730,R_277_b0ed7d8,R_278_b0ed880,R_279_b0ed928,R_27a_b0ed9d0,R_27b_b0eda78,R_27c_b0edb20,R_27d_b0edbc8,R_27e_b0edc70,R_27f_b0edd18,
        R_280_b0eddc0,R_281_b0ede68,R_282_b0edf10,R_283_b0edfb8,R_284_b0ee060,R_285_b0ee108,R_286_b0ee1b0,R_287_b0ee258,R_288_b0ee300,R_289_b0ee3a8,
        R_28a_b0ee450,R_28b_b0ee4f8,R_28c_b0ee5a0,R_28d_b0ee648,R_28e_b0ee6f0,R_28f_b0ee798,R_290_b0ee840,R_291_b0ee8e8,R_292_b0ee990,R_293_b0eea38,
        R_294_b0eeae0,R_295_b0eeb88,R_296_b0eec30,R_297_b0eecd8,R_298_b0eed80,R_299_b0eee28,R_29a_b0eeed0,R_29b_b0eef78,R_29c_b0ef020);
input RIaa97c98_14,RIaa9e7f0_243,RIaa9e868_244,RIaa9e778_242,RIaa9e9d0_247,RIaa97d88_16,RIaa97d10_15,RIaa97e00_17,RIaa97c20_13,
        RIaa9e688_240,RIaa9e700_241,RIaa9e8e0_245,RIaa9e958_246,RIaa9cf90_191,RIaa9d170_195,RIaa9cea0_189,RIaa9d1e8_196,RIaa9d080_193,RIaa9d0f8_194,
        RIaa9d5a8_204,RIaa9d620_205,RIaa9d2d8_198,RIaa9d008_192,RIaa9d3c8_200,RIaa9d4b8_202,RIaa9d260_197,RIaa9d350_199,RIaa9cf18_190,RIaa9d530_203,
        RIaa9d440_201,RIaa97860_5,RIaa976f8_2,RIaa97770_3,RIaa977e8_4,RIaa9ba00_145,RIaa9b640_137,RIaa9b910_143,RIaa9bd48_152,RIaa9ba78_146,
        RIaa9bb68_148,RIaa9b7a8_140,RIaa9bdc0_153,RIaa9baf0_147,RIaa9b730_139,RIaa9bc58_150,RIaa9b6b8_138,RIaa9b898_142,RIaa9bcd0_151,RIaa9b988_144,
        RIaa9b820_141,RIaa9bbe0_149,RIaa9b370_131,RIaa9b0a0_125,RIaa9b5c8_136,RIaa9b3e8_132,RIaa9ae48_120,RIaa9b460_133,RIaa9b190_127,RIaa9b118_126,
        RIaa9b4d8_134,RIaa9b280_129,RIaa9b028_124,RIaa9af38_122,RIaa9b2f8_130,RIaa9aec0_121,RIaa9b550_135,RIaa9afb0_123,RIaa9b208_128,RIaa9c2e8_164,
        RIaa9c4c8_168,RIaa9c018_158,RIaa9c3d8_166,RIaa9c450_167,RIaa9be38_154,RIaa9bfa0_157,RIaa9beb0_155,RIaa9c270_163,RIaa9c090_159,RIaa9c108_160,
        RIaa9c180_161,RIaa9bf28_156,RIaa9c5b8_170,RIaa9c1f8_162,RIaa9c360_165,RIaa9c540_169,RIaa9ce28_188,RIaa9c978_178,RIaa9c9f0_179,RIaa9c900_177,
        RIaa9cdb0_187,RIaa9c810_175,RIaa9c720_173,RIaa9cb58_182,RIaa9cae0_181,RIaa9c630_171,RIaa9ca68_180,RIaa9cc48_184,RIaa9ccc0_185,RIaa9c888_176,
        RIaa9c6a8_172,RIaa9c798_174,RIaa9cbd0_183,RIaa9cd38_186,RIaa9ab78_114,RIaa9aa10_111,RIaa9ac68_116,RIaa9a7b8_106,RIaa9a6c8_104,RIaa9add0_119,
        RIaa9abf0_115,RIaa9a8a8_108,RIaa9a998_110,RIaa9a920_109,RIaa9a830_107,RIaa9ad58_118,RIaa9a740_105,RIaa9ab00_113,RIaa9aa88_112,RIaa9a650_103,
        RIaa9ace0_117,RIaa978d8_6,RIaa9a308_96,RIaa9a218_94,RIaa9a380_97,RIaa9a038_90,RIaa99ed0_87,RIaa9a290_95,RIaa9a0b0_91,RIaa99fc0_89,
        RIaa9a470_99,RIaa99f48_88,RIaa9a4e8_100,RIaa9a1a0_93,RIaa9a3f8_98,RIaa99e58_86,RIaa9a560_101,RIaa9a128_92,RIaa9a5d8_102,RIaa97950_7,
        RIaa99b10_79,RIaa999a8_76,RIaa99a20_77,RIaa996d8_70,RIaa99930_75,RIaa99d68_84,RIaa99b88_80,RIaa99660_69,RIaa99cf0_83,RIaa99c00_81,
        RIaa998b8_74,RIaa99de0_85,RIaa99a98_78,RIaa99c78_82,RIaa997c8_72,RIaa99840_73,RIaa99750_71,RIaa979c8_8,RIaa9f6f0_275,RIaa9f768_276,
        RIaa9f3a8_268,RIaa9f600_273,RIaa9f2b8_266,RIaa9f330_267,RIaa9f420_269,RIaa9f9c0_281,RIaa9f948_280,RIaa9f678_274,RIaa9f8d0_279,RIaa9f588_272,
        RIaa9f240_265,RIaa9f510_271,RIaa9f7e0_277,RIaa9f858_278,RIaa9f498_270,RIaa9eca0_253,RIaa9ee08_256,RIaa9eef8_258,RIaa9ed90_255,RIaa9f1c8_264,
        RIaa9efe8_260,RIaa9ef70_259,RIaa9ed18_254,RIaa9eb38_250,RIaa9ebb0_251,RIaa9ea48_248,RIaa9f0d8_262,RIaa9ee80_257,RIaa9eac0_249,RIaa9f150_263,
        RIaa9f060_261,RIaa9ec28_252,RIaa97b30_11,RIaa97ba8_12,RIaa9de18_222,RIaa9db48_216,RIaa9d968_212,RIaa9dbc0_217,RIaa9dda0_221,RIaa9dd28_220,
        RIaa9dad0_215,RIaa9d800_209,RIaa9dc38_218,RIaa9d710_207,RIaa9dcb0_219,RIaa9d788_208,RIaa9d698_206,RIaa9da58_214,RIaa9d9e0_213,RIaa9d878_210,
        RIaa9d8f0_211,RIaa994f8_66,RIaa99048_56,RIaa98f58_54,RIaa99570_67,RIaa990c0_57,RIaa99138_58,RIaa99390_63,RIaa98ee0_53,RIaa99480_65,
        RIaa98fd0_55,RIaa995e8_68,RIaa99318_62,RIaa991b0_59,RIaa99408_64,RIaa992a0_61,RIaa98e68_52,RIaa99228_60,RIaa9e160_229,RIaa9df80_225,
        RIaa9e3b8_234,RIaa9de90_223,RIaa9e610_239,RIaa9e2c8_232,RIaa9e598_238,RIaa9e1d8_230,RIaa9df08_224,RIaa9e520_237,RIaa9e340_233,RIaa9e250_231,
        RIaa9e430_235,RIaa9e0e8_228,RIaa9dff8_226,RIaa9e4a8_236,RIaa9e070_227,RIaa97ab8_10,RIaa97a40_9,RIaa98b20_45,RIaa989b8_42,RIaa98c88_48,
        RIaa98a30_43,RIaa98aa8_44,RIaa98df0_51,RIaa98940_41,RIaa98c10_47,RIaa98670_35,RIaa98850_39,RIaa98760_37,RIaa986e8_36,RIaa98d00_49,
        RIaa98b98_46,RIaa987d8_38,RIaa988c8_40,RIaa98d78_50,RIaaa1ce8_356,RIaaa1e50_359,RIaaa2030_363,RIaaa1fb8_362,RIaaa1f40_361,RIaaa1c70_355,
        RIaaa1d60_357,RIaaa1ec8_360,RIaaa1b80_353,RIaaa1bf8_354,RIaaa20a8_364,RIaaa1a90_351,RIaaa2120_365,RIaaa1dd8_358,RIaaa2198_366,RIaaa1b08_352,
        RIaaa1a18_350,RIaaa1130_331,RIaaa0f50_327,RIaaa0a28_316,RIaaa0b90_319,RIaaa0b18_318,RIaaa1040_329,RIaaa0c80_321,RIaaa0cf8_322,RIaaa0c08_320,
        RIaaa0ed8_326,RIaaa0d70_323,RIaaa0aa0_317,RIaaa0fc8_328,RIaaa11a8_332,RIaaa10b8_330,RIaaa0e60_325,RIaaa0de8_324,RIaa97680_1,RIaa98508_32,
        RIaa98328_28,RIaa98238_26,RIaa98418_30,RIaa97e78_18,RIaa981c0_25,RIaa985f8_34,RIaa982b0_27,RIaa98580_33,RIaa97ef0_19,RIaa98058_22,
        RIaa98148_24,RIaa97f68_20,RIaa97fe0_21,RIaa983a0_29,RIaa980d0_23,RIaa98490_31,RIaaa2cd8_390,RIaaa2af8_386,RIaaa3110_399,RIaaa3188_400,
        RIaaa2f30_395,RIaaa2c60_389,RIaaa2eb8_394,RIaaa2dc8_392,RIaaa2e40_393,RIaaa2fa8_396,RIaaa3020_397,RIaaa2a08_384,RIaaa3098_398,RIaaa2be8_388,
        RIaaa2b70_387,RIaaa2a80_385,RIaaa2d50_391,RIaaa1298_334,RIaaa16d0_343,RIaaa1928_348,RIaaa1658_342,RIaaa1838_346,RIaaa14f0_339,RIaaa1388_336,
        RIaaa1400_337,RIaaa19a0_349,RIaaa1748_344,RIaaa15e0_341,RIaaa1310_335,RIaaa1220_333,RIaaa1478_338,RIaaa1568_340,RIaaa17c0_345,RIaaa18b0_347,
        RIaa9ff60_293,RIaa9fba0_285,RIaa9fa38_282,RIaaa0050_295,RIaa9ffd8_294,RIaa9fe70_291,RIaa9fc90_287,RIaaa01b8_298,RIaaa0140_297,RIaa9fdf8_290,
        RIaa9fab0_283,RIaa9fc18_286,RIaa9fb28_284,RIaa9fd08_288,RIaaa00c8_296,RIaa9fee8_292,RIaa9fd80_289,RIaaa05f0_307,RIaaa0938_314,RIaaa0758_310,
        RIaaa0488_304,RIaaa0578_306,RIaaa0230_299,RIaaa06e0_309,RIaaa0848_312,RIaaa0398_302,RIaaa0320_301,RIaaa0668_308,RIaaa0410_303,RIaaa02a8_300,
        RIaaa08c0_313,RIaaa0500_305,RIaaa07d0_311,RIaaa09b0_315,RIaaa24e0_373,RIaaa2558_374,RIaaa2738_378,RIaaa2828_380,RIaaa2300_369,RIaaa26c0_377,
        RIaaa2918_382,RIaaa2468_372,RIaaa2378_370,RIaaa2288_368,RIaaa2648_376,RIaaa23f0_371,RIaaa2210_367,RIaaa25d0_375,RIaaa27b0_379,RIaaa28a0_381,
        RIaaa2990_383,RIaaa3f20_429,RIaaa3f98_430,RIaaa3cc8_424,RIaaa3c50_423,RIaaa4010_431,RIaaa4100_433,RIaaa3db8_426,RIaaa3b60_421,RIaaa3d40_425,
        RIaaa3ae8_420,RIaaa3a70_419,RIaaa39f8_418,RIaaa4178_434,RIaaa3e30_427,RIaaa3bd8_422,RIaaa4088_432,RIaaa3ea8_428,RIaaa32f0_403,RIaaa3890_415,
        RIaaa34d0_407,RIaaa3638_410,RIaaa3728_412,RIaaa35c0_409,RIaaa3278_402,RIaaa3818_414,RIaaa33e0_405,RIaaa3368_404,RIaaa37a0_413,RIaaa3980_417,
        RIaaa3908_416,RIaaa36b0_411,RIaaa3458_406,RIaaa3548_408,RIaaa3200_401,RIaaa4448_440,RIaaa4538_442,RIaaa4268_436,RIaaa43d0_439,RIaaa42e0_437,
        RIaaa41f0_435,RIaaa4628_444,RIaaa4808_448,RIaaa45b0_443,RIaaa4718_446,RIaaa44c0_441,RIaaa48f8_450,RIaaa4358_438,RIaaa4970_451,RIaaa4880_449,
        RIaaa4790_447,RIaaa46a0_445,RIaaa6248_504,RIaaa66f8_514,RIaaa6860_517,RIaaa67e8_516,RIaaa6680_513,RIaaa64a0_509,RIaaa6338_506,RIaaa63b0_507,
        RIaaa6950_519,RIaaa6608_512,RIaaa6590_511,RIaaa6428_508,RIaaa6770_515,RIaaa68d8_518,RIaaa6518_510,RIaaa62c0_505,RIaaa61d0_503,RIaaa57f8_482,
        RIaaa54b0_475,RIaaa5618_478,RIaaa52d0_471,RIaaa5528_476,RIaaa5258_470,RIaaa5708_480,RIaaa5690_479,RIaaa5348_472,RIaaa53c0_473,RIaaa58e8_484,
        RIaaa5960_485,RIaaa5780_481,RIaaa5438_474,RIaaa5870_483,RIaaa55a0_477,RIaaa51e0_469,RIaaa4e98_462,RIaaa49e8_452,RIaaa4b50_455,RIaaa4e20_461,
        RIaaa50f0_467,RIaaa4f88_464,RIaaa5000_465,RIaaa4c40_457,RIaaa4cb8_458,RIaaa4a60_453,RIaaa4f10_463,RIaaa4bc8_456,RIaaa4ad8_454,RIaaa5168_468,
        RIaaa4d30_459,RIaaa4da8_460,RIaaa5078_466,RIaaa5e10_495,RIaaa5ca8_492,RIaaa59d8_486,RIaaa60e0_501,RIaaa5b40_489,RIaaa5a50_487,RIaaa5f00_497,
        RIaaa5bb8_490,RIaaa6158_502,RIaaa5f78_498,RIaaa5ac8_488,RIaaa5e88_496,RIaaa5d98_494,RIaaa5ff0_499,RIaaa5d20_493,RIaaa6068_500,RIaaa5c30_491,
        RIaaa6d10_527,RIaaa6a40_521,RIaaa7058_534,RIaaa7148_536,RIaaa6e00_529,RIaaa6ba8_524,RIaaa6e78_530,RIaaa6c98_526,RIaaa6f68_532,RIaaa6ab8_522,
        RIaaa70d0_535,RIaaa6c20_525,RIaaa69c8_520,RIaaa6d88_528,RIaaa6fe0_533,RIaaa6ef0_531,RIaaa6b30_523,RIaaa8408_576,RIaaa87c8_584,RIaaa84f8_578,
        RIaaa8390_575,RIaaa8318_574,RIaaa8660_581,RIaaa8228_572,RIaaa88b8_586,RIaaa8930_587,RIaaa8750_583,RIaaa8480_577,RIaaa8840_585,RIaaa86d8_582,
        RIaaa85e8_580,RIaaa8570_579,RIaaa82a0_573,RIaaa81b0_571,RIaaa7670_547,RIaaa7238_538,RIaaa7490_543,RIaaa75f8_546,RIaaa78c8_552,RIaaa7328_540,
        RIaaa73a0_541,RIaaa77d8_550,RIaaa7850_551,RIaaa76e8_548,RIaaa7580_545,RIaaa72b0_539,RIaaa71c0_537,RIaaa7508_544,RIaaa7418_542,RIaaa7940_553,
        RIaaa7760_549,RIaaa7d00_561,RIaaa7f58_566,RIaaa7fd0_567,RIaaa7b98_558,RIaaa7b20_557,RIaaa7df0_563,RIaaa7c88_560,RIaaa7e68_564,RIaaa7ee0_565,
        RIaaa7d78_562,RIaaa8048_568,RIaaa7c10_559,RIaaa8138_570,RIaaa80c0_569,RIaaa7aa8_556,RIaaa7a30_555,RIaaa79b8_554,RIaaa89a8_588,RIaaa95d8_614,
        RIaaa9218_606,RIaaa90b0_603,RIaaa9128_604,RIaaa91a0_605,RIaaa9380_609,RIaaa9308_608,RIaaa9290_607,RIaaa9038_602,RIaaa93f8_610,RIaaa9470_611,
        RIaaa94e8_612,RIaaa8c78_594,RIaaa8cf0_595,RIaaa8a98_590,RIaaa8b10_591,RIaaa8a20_589,RIaaa8b88_592,RIaaa8c00_593,RIaaa8d68_596,RIaaa8de0_597,
        RIaaa8e58_598,RIaaa8ed0_599,RIaaa8f48_600,RIaaa8fc0_601,RIaaa9560_613;
output R_267_b0ecd58,R_268_b0ece00,R_269_b0ecea8,R_26a_b0ecf50,R_26b_b0ecff8,R_26c_b0ed0a0,R_26d_b0ed148,R_26e_b0ed1f0,R_26f_b0ed298,
        R_270_b0ed340,R_271_b0ed3e8,R_272_b0ed490,R_273_b0ed538,R_274_b0ed5e0,R_275_b0ed688,R_276_b0ed730,R_277_b0ed7d8,R_278_b0ed880,R_279_b0ed928,
        R_27a_b0ed9d0,R_27b_b0eda78,R_27c_b0edb20,R_27d_b0edbc8,R_27e_b0edc70,R_27f_b0edd18,R_280_b0eddc0,R_281_b0ede68,R_282_b0edf10,R_283_b0edfb8,
        R_284_b0ee060,R_285_b0ee108,R_286_b0ee1b0,R_287_b0ee258,R_288_b0ee300,R_289_b0ee3a8,R_28a_b0ee450,R_28b_b0ee4f8,R_28c_b0ee5a0,R_28d_b0ee648,
        R_28e_b0ee6f0,R_28f_b0ee798,R_290_b0ee840,R_291_b0ee8e8,R_292_b0ee990,R_293_b0eea38,R_294_b0eeae0,R_295_b0eeb88,R_296_b0eec30,R_297_b0eecd8,
        R_298_b0eed80,R_299_b0eee28,R_29a_b0eeed0,R_29b_b0eef78,R_29c_b0ef020;

wire \669_ZERO , \670_ONE , \671 , \672 , \673 , \674 , \675 , \676 , \677 ,
         \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 ,
         \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 ,
         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,
         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,
         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,
         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,
         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,
         \748 , \749 , \750 , \751 , \752 , \753 , \754 , \755 , \756 , \757 ,
         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,
         \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,
         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787 ,
         \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,
         \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 ,
         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,
         \818 , \819 , \820 , \821 , \822 , \823 , \824 , \825 , \826 , \827 ,
         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,
         \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,
         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,
         \858 , \859 , \860 , \861 , \862 , \863 , \864 , \865 , \866 , \867 ,
         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 ,
         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,
         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,
         \898 , \899 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,
         \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 ,
         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,
         \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937 ,
         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,
         \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,
         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,
         \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975 , \976 , \977 ,
         \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 ,
         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,
         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,
         \1008 , \1009 , \1010 , \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,
         \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,
         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,
         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 ,
         \1048 , \1049 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 ,
         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,
         \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 ,
         \1078 , \1079 , \1080 , \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 ,
         \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 ,
         \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 ,
         \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 ,
         \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 ,
         \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 ,
         \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 ,
         \1148 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 ,
         \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 ,
         \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 ,
         \1178 , \1179 , \1180 , \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 ,
         \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 ,
         \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 ,
         \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 ,
         \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 ,
         \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 ,
         \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 ,
         \1248 , \1249 , \1250 , \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 ,
         \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 ,
         \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 ,
         \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 ,
         \1288 , \1289 , \1290 , \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 ,
         \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 ,
         \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 ,
         \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 ,
         \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 ,
         \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 ,
         \1348 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 ,
         \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 ,
         \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 ,
         \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 ,
         \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 ,
         \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 ,
         \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 ,
         \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 ,
         \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 ,
         \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 ,
         \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 ,
         \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 ,
         \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 ,
         \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 ,
         \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 ,
         \1498 , \1499 , \1500 , \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 ,
         \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 ,
         \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 ,
         \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 ,
         \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 ,
         \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 ,
         \1558 , \1559 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 ,
         \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 ,
         \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 ,
         \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 ,
         \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 ,
         \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 ,
         \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 ,
         \1628 , \1629 , \1630 , \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 ,
         \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 ,
         \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 ,
         \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 ,
         \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 ,
         \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 ,
         \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 ,
         \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 ,
         \1708 , \1709 , \1710 , \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 ,
         \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 ,
         \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 ,
         \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 ,
         \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 ,
         \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 ,
         \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 ,
         \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 ,
         \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 ,
         \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 ,
         \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 ,
         \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 ,
         \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 ,
         \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 ,
         \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 ,
         \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 ,
         \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 ,
         \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 ,
         \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 ,
         \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 ,
         \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 ,
         \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 ,
         \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 ,
         \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 ,
         \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 ,
         \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 ,
         \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 ,
         \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 ,
         \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 ,
         \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 ,
         \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 ,
         \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 ,
         \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 ,
         \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 ,
         \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 ,
         \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 ,
         \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 ,
         \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 ,
         \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 ,
         \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 ,
         \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 ,
         \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 ,
         \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 ,
         \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 ,
         \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 ,
         \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 ,
         \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 ,
         \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 ,
         \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 ,
         \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 ,
         \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 ,
         \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 ,
         \2228 , \2229 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 ,
         \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 ,
         \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 ,
         \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 ,
         \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 ,
         \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 ,
         \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 ,
         \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 ,
         \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 ,
         \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 ,
         \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 ,
         \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 ,
         \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 ,
         \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 ,
         \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 ,
         \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 ,
         \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 ,
         \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 ,
         \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 ,
         \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 ,
         \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 ,
         \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 ,
         \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 ,
         \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 ,
         \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 ,
         \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 ,
         \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 ,
         \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 ,
         \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 ,
         \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 ,
         \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 ,
         \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 ,
         \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 ,
         \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 ,
         \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 ,
         \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 ,
         \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 ,
         \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 ,
         \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 ,
         \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 ,
         \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 ,
         \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 ,
         \2648 , \2649 , \2650 , \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 ,
         \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 ,
         \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 ,
         \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 ,
         \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 ,
         \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 ,
         \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 ,
         \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 ,
         \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 ,
         \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 ,
         \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 ,
         \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 ,
         \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 ,
         \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 ,
         \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 ,
         \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 ,
         \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 ,
         \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 ,
         \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 ,
         \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 ,
         \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 ,
         \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 ,
         \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 ,
         \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 ,
         \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 ,
         \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 ,
         \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 ,
         \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 ,
         \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 ,
         \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 ,
         \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 ,
         \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 ,
         \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 ,
         \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 ,
         \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 ,
         \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 ,
         \3008 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 ,
         \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 ,
         \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 ,
         \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 ,
         \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 ,
         \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 ,
         \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 ,
         \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 ,
         \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 ,
         \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 ,
         \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 ,
         \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 ,
         \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 ,
         \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 ,
         \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 ,
         \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 ,
         \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 ,
         \3178 , \3179 , \3180 , \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 ,
         \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 ,
         \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 ,
         \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 ,
         \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 ,
         \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 ,
         \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 ,
         \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 ,
         \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 ,
         \3268 , \3269 , \3270 , \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 ,
         \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 ,
         \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 ,
         \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 ,
         \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 ,
         \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 ,
         \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 ,
         \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 ,
         \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 ,
         \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 ,
         \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 ,
         \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 ,
         \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 ,
         \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 ,
         \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 ,
         \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 ,
         \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 ,
         \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 ,
         \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 ,
         \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 ,
         \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 ,
         \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 ,
         \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 ,
         \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 ,
         \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 ,
         \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 ,
         \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 ,
         \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 ,
         \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 ,
         \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 ,
         \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 ,
         \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 ,
         \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 ,
         \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 ,
         \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 ,
         \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 ,
         \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 ,
         \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 ,
         \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 ,
         \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 ,
         \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 ,
         \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 ,
         \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 ,
         \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 ,
         \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 ,
         \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 ,
         \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 ,
         \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 ,
         \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 ,
         \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 ,
         \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 ,
         \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 ,
         \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 ,
         \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 ,
         \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 ,
         \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 ,
         \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 ,
         \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 ,
         \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 ,
         \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 ,
         \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 ,
         \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 ,
         \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 ,
         \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 ,
         \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 ,
         \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 ,
         \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 ,
         \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 ,
         \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 ,
         \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 ,
         \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 ,
         \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 ,
         \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 ,
         \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 ,
         \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 ,
         \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 ,
         \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 ,
         \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 ,
         \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 ,
         \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 ,
         \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 ,
         \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 ,
         \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 ,
         \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 ,
         \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 ,
         \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 ,
         \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 ,
         \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 ,
         \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 ,
         \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 ,
         \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 ,
         \4178 , \4179 , \4180 , \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 ,
         \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 ,
         \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 ,
         \4208 , \4209 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 ,
         \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 ,
         \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 ,
         \4238 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 ,
         \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 ,
         \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 ,
         \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 ,
         \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 ,
         \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 ,
         \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 ,
         \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 ,
         \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 ,
         \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 ,
         \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 ,
         \4348 , \4349 , \4350 , \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 ,
         \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 ,
         \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 ,
         \4378 , \4379 , \4380 , \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 ,
         \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 ,
         \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 ,
         \4408 , \4409 , \4410 , \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 ,
         \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 ,
         \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 ,
         \4438 , \4439 , \4440 , \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 ,
         \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 ,
         \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 ,
         \4468 , \4469 , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 ,
         \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 ,
         \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 ,
         \4498 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 ,
         \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 ,
         \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 ,
         \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 ,
         \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 ,
         \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 ,
         \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 ,
         \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 ,
         \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 ,
         \4588 , \4589 , \4590 , \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 ,
         \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 ,
         \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 ,
         \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 ,
         \4628 , \4629 , \4630 , \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 ,
         \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 ,
         \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 ,
         \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 ,
         \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 ,
         \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 ,
         \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 ,
         \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 ,
         \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 ,
         \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 ,
         \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 ,
         \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 ,
         \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 ,
         \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 ,
         \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 ,
         \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 ,
         \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 ,
         \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 ,
         \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 ,
         \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 ,
         \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 ,
         \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 ,
         \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 ,
         \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 ,
         \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 ,
         \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 ,
         \4888 , \4889 , \4890 , \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 ,
         \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 ,
         \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 ,
         \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 ,
         \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 ,
         \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 ,
         \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 ,
         \4958 , \4959 , \4960 , \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 ,
         \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 ,
         \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 ,
         \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 ,
         \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 ,
         \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 ,
         \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 ,
         \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 ,
         \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 ,
         \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 ,
         \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 ,
         \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 ,
         \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 ,
         \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 ,
         \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 ,
         \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 ,
         \5118 , \5119 , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 ,
         \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 ,
         \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 ,
         \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 ,
         \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 ,
         \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 ,
         \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 ,
         \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 ,
         \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 ,
         \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 ,
         \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 ,
         \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 ,
         \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 ,
         \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 ,
         \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 ,
         \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 ,
         \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 ,
         \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 ,
         \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 ,
         \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 ,
         \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 ,
         \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 ,
         \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 ,
         \5348 , \5349 , \5350 , \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 ,
         \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 ,
         \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 ,
         \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 ,
         \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 ,
         \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 ,
         \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 ,
         \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 ,
         \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 ,
         \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 ,
         \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 ,
         \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 ,
         \5468 , \5469 , \5470 , \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 ,
         \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 ,
         \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 ,
         \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 ,
         \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 ,
         \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 ,
         \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 ,
         \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 ,
         \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 ,
         \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 ,
         \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 ,
         \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 ,
         \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 ,
         \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 ,
         \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 ,
         \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 ,
         \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 ,
         \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 ,
         \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 ,
         \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 ,
         \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 ,
         \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 ,
         \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 ,
         \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 ,
         \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 ,
         \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 ,
         \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 ,
         \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 ,
         \5748 , \5749 , \5750 , \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 ,
         \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 ,
         \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 ,
         \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 ,
         \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 ,
         \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 ,
         \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 ,
         \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 ,
         \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 ,
         \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 ,
         \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 ,
         \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 ,
         \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 ,
         \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 ,
         \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 ,
         \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 ,
         \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 ,
         \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 ,
         \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 ,
         \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 ,
         \5948 , \5949 , \5950 , \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 ,
         \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 ,
         \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 ,
         \5978 , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 ,
         \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 ,
         \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 ,
         \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 ,
         \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 ,
         \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 ,
         \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 ,
         \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 ,
         \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 ,
         \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 ,
         \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 ,
         \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 ,
         \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 ,
         \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 ,
         \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 ,
         \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 ,
         \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 ,
         \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 ,
         \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 ,
         \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 ,
         \6178 , \6179 , \6180 , \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 ,
         \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 ,
         \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 ,
         \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 ,
         \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 ,
         \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 ,
         \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 ,
         \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 ,
         \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 ,
         \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 ,
         \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 ,
         \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 ,
         \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 ,
         \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 ,
         \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 ,
         \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 ,
         \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 ,
         \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 ,
         \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 ,
         \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 ,
         \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 ,
         \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 ,
         \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 ,
         \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 ,
         \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 ,
         \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 ,
         \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 ,
         \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 ,
         \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 ,
         \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 ,
         \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 ,
         \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 ,
         \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 ,
         \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 ,
         \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 ,
         \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 ,
         \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 ,
         \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 ,
         \6558 , \6559 , \6560 , \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 ,
         \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 ,
         \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 ,
         \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 ,
         \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 ,
         \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 ,
         \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 ,
         \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 ,
         \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 ,
         \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 ,
         \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 ,
         \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 ,
         \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 ,
         \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 ,
         \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 ,
         \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 ,
         \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 ,
         \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 ,
         \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 ,
         \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 ,
         \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 ,
         \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 ,
         \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 ,
         \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 ,
         \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 ,
         \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 ,
         \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 ,
         \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 ,
         \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 ,
         \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 ,
         \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 ,
         \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 ,
         \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 ,
         \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 ,
         \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 ,
         \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 ,
         \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 ,
         \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 ,
         \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 ,
         \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 ,
         \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 ,
         \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 ,
         \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 ,
         \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 ,
         \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 ,
         \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 ,
         \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 ,
         \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 ,
         \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 ,
         \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 ,
         \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 ,
         \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 ,
         \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 ,
         \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 ,
         \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 ,
         \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 ,
         \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 ,
         \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 ,
         \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 ,
         \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 ,
         \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 ,
         \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 ,
         \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 ,
         \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 ,
         \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 ,
         \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 ,
         \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 ,
         \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 ,
         \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 ,
         \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 ,
         \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 ,
         \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 ,
         \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 ,
         \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 ,
         \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 ,
         \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 ,
         \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 ,
         \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 ,
         \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 ,
         \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 ,
         \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 ,
         \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 ,
         \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 ,
         \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 ,
         \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 ,
         \7408 , \7409 , \7410 , \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 ,
         \7418 , \7419 , \7420 , \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 ,
         \7428 , \7429 , \7430 , \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 ,
         \7438 , \7439 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 ,
         \7448 , \7449 , \7450 , \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 ,
         \7458 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 ,
         \7468 , \7469 , \7470 , \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 ,
         \7478 , \7479 , \7480 , \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 ,
         \7488 , \7489 , \7490 , \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 ,
         \7498 , \7499 , \7500 , \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 ,
         \7508 , \7509 , \7510 , \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 ,
         \7518 , \7519 , \7520 , \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 ,
         \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 ,
         \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 ,
         \7548 , \7549 , \7550 , \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 ,
         \7558 , \7559 , \7560 , \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 ,
         \7568 , \7569 , \7570 , \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 ,
         \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 ,
         \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 ,
         \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
         \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 ,
         \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 ,
         \7628 , \7629 , \7630 , \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 ,
         \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 ,
         \7648 , \7649 , \7650 , \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 ,
         \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 ,
         \7668 , \7669 , \7670 , \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 ,
         \7678 , \7679 , \7680 , \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 ,
         \7688 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 ,
         \7698 , \7699 , \7700 , \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 ,
         \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 ,
         \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 ,
         \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 ,
         \7738 , \7739 , \7740 , \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 ,
         \7748 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 ,
         \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 ,
         \7768 , \7769 , \7770 , \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 ,
         \7778 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 ,
         \7788 , \7789 , \7790 , \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 ,
         \7798 , \7799 , \7800 , \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 ,
         \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 ,
         \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 ,
         \7828 , \7829 , \7830 , \7831 , \7832 , \7833 , \7834 , \7835 , \7836 , \7837 ,
         \7838 , \7839 , \7840 , \7841 , \7842 , \7843 , \7844 , \7845 , \7846 , \7847 ,
         \7848 , \7849 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855 , \7856 , \7857 ,
         \7858 , \7859 , \7860 , \7861 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867 ,
         \7868 , \7869 , \7870 , \7871 , \7872 , \7873 , \7874 , \7875 , \7876 , \7877 ,
         \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 ,
         \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 ,
         \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 ,
         \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 ,
         \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 ,
         \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 ,
         \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 ,
         \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 ,
         \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 ,
         \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974 , \7975 , \7976 , \7977 ,
         \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 ,
         \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 ,
         \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 ,
         \8008 , \8009 , \8010 , \8011 , \8012 , \8013 , \8014 , \8015 , \8016 , \8017 ,
         \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 ,
         \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 ,
         \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 ,
         \8048 , \8049 , \8050 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 ,
         \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 ,
         \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 ,
         \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 ,
         \8088 , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 ,
         \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 ,
         \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 ,
         \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124 , \8125 , \8126 , \8127 ,
         \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 ,
         \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 ,
         \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 ,
         \8158 , \8159 , \8160 , \8161 , \8162 , \8163 , \8164 , \8165 , \8166 , \8167 ,
         \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 ,
         \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 ,
         \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 ,
         \8198 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 ,
         \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 ,
         \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 ,
         \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234 , \8235 , \8236 , \8237 ,
         \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 ,
         \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 ,
         \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 ,
         \8268 , \8269 , \8270 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 ,
         \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 ,
         \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 ,
         \8298 , \8299 , \8300 , \8301 , \8302 , \8303 , \8304 , \8305 , \8306 , \8307 ,
         \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 ,
         \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 ,
         \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 ,
         \8338 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 ,
         \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 ,
         \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 ,
         \8368 , \8369 , \8370 , \8371 , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 ,
         \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 ,
         \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 ,
         \8398 , \8399 , \8400 , \8401 , \8402 , \8403 , \8404 , \8405 , \8406 , \8407 ,
         \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 ,
         \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 ,
         \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 ,
         \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 ,
         \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 ,
         \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 ,
         \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474 , \8475 , \8476 , \8477 ,
         \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 ,
         \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 ,
         \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 ,
         \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514 , \8515 , \8516 , \8517 ,
         \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 ,
         \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 ,
         \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 ,
         \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 ,
         \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 ,
         \8568 , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 ,
         \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 ,
         \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 ,
         \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 ,
         \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 ,
         \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 ,
         \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 ,
         \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 ,
         \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657 ,
         \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 ,
         \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 ,
         \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 ,
         \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 ,
         \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 ,
         \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 ,
         \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 ,
         \8728 , \8729 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 ,
         \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 ,
         \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 ,
         \8758 , \8759 , \8760 , \8761 , \8762 , \8763 , \8764 , \8765 , \8766 , \8767 ,
         \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 ,
         \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 ,
         \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 ,
         \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 ,
         \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 ,
         \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 ,
         \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 ,
         \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 ,
         \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 ,
         \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 ,
         \8868 , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 ,
         \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 ,
         \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 ,
         \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 ,
         \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 ,
         \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 ,
         \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 ,
         \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947 ,
         \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 ,
         \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 ,
         \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 ,
         \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 ,
         \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 ,
         \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 ,
         \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 ,
         \9018 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 ,
         \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 ,
         \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 ,
         \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 ,
         \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 ,
         \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 ,
         \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 ,
         \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 ,
         \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 ,
         \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 ,
         \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 ,
         \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 ,
         \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 ,
         \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 ,
         \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 ,
         \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 ,
         \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 ,
         \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 ,
         \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 ,
         \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 ,
         \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 ,
         \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 ,
         \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 ,
         \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 ,
         \9258 , \9259 , \9260 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 ,
         \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 ,
         \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 ,
         \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 ,
         \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 ,
         \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317 ,
         \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 ,
         \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 ,
         \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 ,
         \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 ,
         \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 ,
         \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 ,
         \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 ,
         \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 ,
         \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 ,
         \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 ,
         \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 ,
         \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 ,
         \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 ,
         \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 ,
         \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 ,
         \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 ,
         \9478 , \9479 , \9480 , \9481 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 ,
         \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 ,
         \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 ,
         \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 ,
         \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 ,
         \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 ,
         \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 ,
         \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 ,
         \9558 , \9559 , \9560 , \9561 , \9562 , \9563 , \9564 , \9565 , \9566 , \9567 ,
         \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 ,
         \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 ,
         \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 ,
         \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 ,
         \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 ,
         \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 ,
         \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 ,
         \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 ,
         \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 ,
         \9658 , \9659 , \9660 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 ,
         \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 ,
         \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 ,
         \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 ,
         \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 ,
         \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 ,
         \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 ,
         \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 ,
         \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 ,
         \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 ,
         \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 ,
         \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 ,
         \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 ,
         \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 ,
         \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 ,
         \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 ,
         \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 ,
         \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 ,
         \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 ,
         \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 ,
         \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 ,
         \9868 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 ,
         \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 ,
         \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 ,
         \9898 , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 ,
         \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 ,
         \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 ,
         \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 ,
         \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 ,
         \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 ,
         \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 ,
         \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 ,
         \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 ,
         \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 ,
         \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 ,
         \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 ,
         \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 ,
         \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 ,
         \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 ,
         \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 ,
         \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 ,
         \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 ,
         \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 ,
         \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 ,
         \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 ,
         \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 ,
         \10118 , \10119 , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 ,
         \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 ,
         \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 ,
         \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 ,
         \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 ,
         \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 ,
         \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 ,
         \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 ,
         \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 ,
         \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 ,
         \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 ,
         \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235 , \10236 , \10237 ,
         \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 ,
         \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 ,
         \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 ,
         \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 ,
         \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 ,
         \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 ,
         \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 ,
         \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 ,
         \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 ,
         \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 ,
         \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 ,
         \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 ,
         \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 ,
         \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 ,
         \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 ,
         \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 ,
         \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 ,
         \10408 , \10409 , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 ,
         \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 ,
         \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 ,
         \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 ,
         \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 ,
         \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 ,
         \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 ,
         \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 ,
         \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 ,
         \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506 , \10507 ,
         \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 ,
         \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 ,
         \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 ,
         \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 ,
         \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 ,
         \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 ,
         \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 ,
         \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 ,
         \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 ,
         \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 ,
         \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 ,
         \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 ,
         \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 ,
         \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 ,
         \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 ,
         \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 ,
         \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 ,
         \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 ,
         \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 ,
         \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 ,
         \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 ,
         \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 ,
         \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 ,
         \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 ,
         \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 ,
         \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 ,
         \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 ,
         \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 ,
         \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 ,
         \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 ,
         \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 ,
         \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 ,
         \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 ,
         \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 ,
         \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 ,
         \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 ,
         \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 ,
         \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 ,
         \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 ,
         \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 ,
         \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 ,
         \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 ,
         \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 ,
         \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 ,
         \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 ,
         \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 ,
         \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 ,
         \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 ,
         \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 ,
         \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 ,
         \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 ,
         \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 ,
         \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 ,
         \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 ,
         \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 ,
         \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 ,
         \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 ,
         \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 ,
         \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 ,
         \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 ,
         \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 ,
         \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 ,
         \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 ,
         \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 ,
         \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 ,
         \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 ,
         \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 ,
         \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 ,
         \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 ,
         \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 ,
         \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 ,
         \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 ,
         \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 ,
         \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 ,
         \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 ,
         \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 ,
         \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 ,
         \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 ,
         \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 ,
         \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 ,
         \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 ,
         \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 ,
         \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 ,
         \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 ,
         \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 ,
         \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 ,
         \11368 , \11369 , \11370 , \11371 , \11372 , \11373 , \11374 , \11375 , \11376 , \11377 ,
         \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 ,
         \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 ,
         \11398 , \11399 , \11400 , \11401 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 ,
         \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 ,
         \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 ,
         \11428 , \11429 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 ,
         \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 ,
         \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 ,
         \11458 , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 ,
         \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 ,
         \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487 ,
         \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 ,
         \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 ,
         \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516 , \11517 ,
         \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 ,
         \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 ,
         \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545 , \11546 , \11547 ,
         \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 ,
         \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 ,
         \11568 , \11569 , \11570 , \11571 , \11572 , \11573 , \11574 , \11575 , \11576 , \11577 ,
         \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 ,
         \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 ,
         \11598 , \11599 , \11600 , \11601 , \11602 , \11603 , \11604 , \11605 , \11606 , \11607 ,
         \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 ,
         \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 ,
         \11628 , \11629 , \11630 , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 ,
         \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 ,
         \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 ,
         \11658 , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 ,
         \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 ,
         \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687 ,
         \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 ,
         \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 ,
         \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715 , \11716 , \11717 ,
         \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 ,
         \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 ,
         \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 ,
         \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 ,
         \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 ,
         \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 ,
         \11778 , \11779 , \11780 , \11781 , \11782 , \11783 , \11784 , \11785 , \11786 , \11787 ,
         \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 ,
         \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 ,
         \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 ,
         \11818 , \11819 , \11820 , \11821 , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 ,
         \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 ,
         \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 ,
         \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 ,
         \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 ,
         \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874 , \11875 , \11876 , \11877 ,
         \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 ,
         \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 ,
         \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 ,
         \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 ,
         \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 ,
         \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 ,
         \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 ,
         \11948 , \11949 , \11950 , \11951 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 ,
         \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 ,
         \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 ,
         \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 ,
         \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 ,
         \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 ,
         \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 ,
         \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 ,
         \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 ,
         \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 ,
         \12048 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 ,
         \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 ,
         \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076 , \12077 ,
         \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 ,
         \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 ,
         \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 ,
         \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 ,
         \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 ,
         \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 ,
         \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 ,
         \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 ,
         \12158 , \12159 , \12160 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 ,
         \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 ,
         \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 ,
         \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 ,
         \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 ,
         \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 ,
         \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 ,
         \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237 ,
         \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 ,
         \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 ,
         \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 ,
         \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 ,
         \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 ,
         \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 ,
         \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307 ,
         \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 ,
         \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 ,
         \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 ,
         \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 ,
         \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 ,
         \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 ,
         \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 ,
         \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 ,
         \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 ,
         \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 ,
         \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 ,
         \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 ,
         \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 ,
         \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 ,
         \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 ,
         \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 ,
         \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 ,
         \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 ,
         \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 ,
         \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 ,
         \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515 , \12516 , \12517 ,
         \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 ,
         \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 ,
         \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 ,
         \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 ,
         \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 ,
         \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 ,
         \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 ,
         \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 ,
         \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 ,
         \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 ,
         \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 ,
         \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 ,
         \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 ,
         \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 ,
         \12658 , \12659 , \12660 , \12661 , \12662 , \12663 , \12664 , \12665 , \12666 , \12667 ,
         \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 ,
         \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 ,
         \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 ,
         \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706 , \12707 ,
         \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 ,
         \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 ,
         \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 ,
         \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 ,
         \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 ,
         \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 ,
         \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 ,
         \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 ,
         \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 ,
         \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 ,
         \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 ,
         \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 ,
         \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 ,
         \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 ,
         \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 ,
         \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 ,
         \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 ,
         \12878 , \12879 , \12880 , \12881 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 ,
         \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 ,
         \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 ,
         \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 ,
         \12918 , \12919 , \12920 , \12921 , \12922 , \12923 , \12924 , \12925 , \12926 , \12927 ,
         \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 ,
         \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 ,
         \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 ,
         \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 ,
         \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 ,
         \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 ,
         \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 ,
         \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 ,
         \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 ,
         \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 ,
         \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 ,
         \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 ,
         \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 ,
         \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 ,
         \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 ,
         \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 ,
         \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 ,
         \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 ,
         \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 ,
         \13118 , \13119 , \13120 , \13121 , \13122 , \13123 , \13124 , \13125 , \13126 , \13127 ,
         \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 ,
         \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 ,
         \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 ,
         \13158 , \13159 , \13160 , \13161 , \13162 , \13163 , \13164 , \13165 , \13166 , \13167 ,
         \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 ,
         \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 ,
         \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 ,
         \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 ,
         \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 ,
         \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 ,
         \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 ,
         \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 ,
         \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 ,
         \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 ,
         \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 ,
         \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 ,
         \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 ,
         \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 ,
         \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 ,
         \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 ,
         \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 ,
         \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 ,
         \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 ,
         \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364 , \13365 , \13366 , \13367 ,
         \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 ,
         \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 ,
         \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 ,
         \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 ,
         \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 ,
         \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 ,
         \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 ,
         \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 ,
         \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 ,
         \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 ,
         \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 ,
         \13478 , \13479 , \13480 , \13481 , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 ,
         \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 ,
         \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 ,
         \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 ,
         \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 ,
         \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 ,
         \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 ,
         \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 ,
         \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 ,
         \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 ,
         \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 ,
         \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 ,
         \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 ,
         \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 ,
         \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 ,
         \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637 ,
         \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 ,
         \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 ,
         \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 ,
         \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 ,
         \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 ,
         \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 ,
         \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 ,
         \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 ,
         \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726 , \13727 ,
         \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 ,
         \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 ,
         \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 ,
         \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 ,
         \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 ,
         \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 ,
         \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 ,
         \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 ,
         \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 ,
         \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 ,
         \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 ,
         \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 ,
         \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 ,
         \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 ,
         \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 ,
         \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 ,
         \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 ,
         \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 ,
         \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 ,
         \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 ,
         \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 ,
         \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 ,
         \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 ,
         \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 ,
         \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 ,
         \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 ,
         \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 ,
         \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 ,
         \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 ,
         \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 ,
         \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 ,
         \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 ,
         \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 ,
         \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 ,
         \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 ,
         \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 ,
         \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 ,
         \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 ,
         \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 ,
         \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 ,
         \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 ,
         \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 ,
         \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 ,
         \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 ,
         \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 ,
         \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 ,
         \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 ,
         \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 ,
         \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 ,
         \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 ,
         \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 ,
         \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 ,
         \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 ,
         \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 ,
         \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 ,
         \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 ,
         \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 ,
         \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 ,
         \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 ,
         \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 ,
         \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 ,
         \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 ,
         \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 ,
         \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 ,
         \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 ,
         \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 ,
         \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 ,
         \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 ,
         \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 ,
         \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 ,
         \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 ,
         \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 ,
         \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 ,
         \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 ,
         \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 ,
         \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 ,
         \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 ,
         \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 ,
         \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 ,
         \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 ,
         \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 ,
         \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 ,
         \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 ,
         \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567 ,
         \14568 , \14569 , \14570 , \14571 , \14572 , \14573 , \14574 , \14575 , \14576 , \14577 ,
         \14578 , \14579 , \14580 , \14581 , \14582 , \14583 , \14584 , \14585 , \14586 , \14587 ,
         \14588 , \14589 , \14590 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596 , \14597 ,
         \14598 , \14599 , \14600 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606 , \14607 ,
         \14608 , \14609 , \14610 , \14611 , \14612 , \14613 , \14614 , \14615 , \14616 , \14617 ,
         \14618 , \14619 , \14620 , \14621 , \14622 , \14623 , \14624 , \14625 , \14626 , \14627 ,
         \14628 , \14629 , \14630 , \14631 , \14632 , \14633 , \14634 , \14635 , \14636 , \14637 ,
         \14638 , \14639 , \14640 , \14641 , \14642 , \14643 , \14644 , \14645 , \14646 , \14647 ,
         \14648 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654 , \14655 , \14656 , \14657 ,
         \14658 , \14659 , \14660 , \14661 , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 ,
         \14668 , \14669 , \14670 , \14671 , \14672 , \14673 , \14674 , \14675 , \14676 , \14677 ,
         \14678 , \14679 , \14680 , \14681 , \14682 , \14683 , \14684 , \14685 , \14686 , \14687 ,
         \14688 , \14689 , \14690 , \14691 , \14692 , \14693 , \14694 , \14695 , \14696 , \14697 ,
         \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 ,
         \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 ,
         \14718 , \14719 , \14720 , \14721 , \14722 , \14723 , \14724 , \14725 , \14726 , \14727 ,
         \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737 ,
         \14738 , \14739 , \14740 , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 ,
         \14748 , \14749 , \14750 , \14751 , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 ,
         \14758 , \14759 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 ,
         \14768 , \14769 , \14770 , \14771 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 ,
         \14778 , \14779 , \14780 , \14781 , \14782 , \14783 , \14784 , \14785 , \14786 , \14787 ,
         \14788 , \14789 , \14790 , \14791 , \14792 , \14793 , \14794 , \14795 , \14796 , \14797 ,
         \14798 , \14799 , \14800 , \14801 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 ,
         \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 ,
         \14818 , \14819 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827 ,
         \14828 , \14829 , \14830 , \14831 , \14832 , \14833 , \14834 , \14835 , \14836 , \14837 ,
         \14838 , \14839 , \14840 , \14841 , \14842 , \14843 , \14844 , \14845 , \14846 , \14847 ,
         \14848 , \14849 , \14850 , \14851 , \14852 , \14853 , \14854 , \14855 , \14856 , \14857 ,
         \14858 , \14859 , \14860 , \14861 , \14862 , \14863 , \14864 , \14865 , \14866 , \14867 ,
         \14868 , \14869 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876 , \14877 ,
         \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885 , \14886 , \14887 ,
         \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896 , \14897 ,
         \14898 , \14899 , \14900 , \14901 , \14902 , \14903 , \14904 , \14905 , \14906 , \14907 ,
         \14908 , \14909 , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 ,
         \14918 , \14919 , \14920 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926 , \14927 ,
         \14928 , \14929 , \14930 , \14931 , \14932 , \14933 , \14934 , \14935 , \14936 , \14937 ,
         \14938 , \14939 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 ,
         \14948 , \14949 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 ,
         \14958 , \14959 , \14960 , \14961 , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 ,
         \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977 ,
         \14978 , \14979 , \14980 , \14981 , \14982 , \14983 , \14984 , \14985 , \14986 , \14987 ,
         \14988 , \14989 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995 , \14996 , \14997 ,
         \14998 , \14999 , \15000 , \15001 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007 ,
         \15008 , \15009 , \15010 , \15011 , \15012 , \15013 , \15014 , \15015 , \15016 , \15017 ,
         \15018 , \15019 , \15020 , \15021 , \15022 , \15023 , \15024 , \15025 , \15026 , \15027 ,
         \15028 , \15029 , \15030 , \15031 , \15032 , \15033 , \15034 , \15035 , \15036 , \15037 ,
         \15038 , \15039 , \15040 , \15041 , \15042 , \15043 , \15044 , \15045 , \15046 , \15047 ,
         \15048 , \15049 , \15050 , \15051 , \15052 , \15053 , \15054 , \15055 , \15056 , \15057 ,
         \15058 , \15059 , \15060 , \15061 , \15062 , \15063 , \15064 , \15065 , \15066 , \15067 ,
         \15068 , \15069 , \15070 , \15071 , \15072 , \15073 , \15074 , \15075 , \15076 , \15077 ,
         \15078 , \15079 , \15080 , \15081 , \15082 , \15083 , \15084 , \15085 , \15086 , \15087 ,
         \15088 , \15089 , \15090 , \15091 , \15092 , \15093 , \15094 , \15095 , \15096 , \15097 ,
         \15098 , \15099 , \15100 , \15101 , \15102 , \15103 , \15104 , \15105 , \15106 , \15107 ,
         \15108 , \15109 , \15110 , \15111 , \15112 , \15113 , \15114 , \15115 , \15116 , \15117 ,
         \15118 , \15119 , \15120 , \15121 , \15122 , \15123 , \15124 , \15125 , \15126 , \15127 ,
         \15128 , \15129 , \15130 , \15131 , \15132 , \15133 , \15134 , \15135 , \15136 , \15137 ,
         \15138 , \15139 , \15140 , \15141 , \15142 , \15143 , \15144 , \15145 , \15146 , \15147 ,
         \15148 , \15149 , \15150 , \15151 , \15152 , \15153 , \15154 , \15155 , \15156 , \15157 ,
         \15158 , \15159 , \15160 , \15161 , \15162 , \15163 , \15164 , \15165 , \15166 , \15167 ,
         \15168 , \15169 , \15170 , \15171 , \15172 , \15173 , \15174 , \15175 , \15176 , \15177 ,
         \15178 , \15179 , \15180 , \15181 , \15182 , \15183 , \15184 , \15185 , \15186 , \15187 ,
         \15188 , \15189 , \15190 , \15191 , \15192 , \15193 , \15194 , \15195 , \15196 , \15197 ,
         \15198 , \15199 , \15200 , \15201 , \15202 , \15203 , \15204 , \15205 , \15206 , \15207 ,
         \15208 , \15209 , \15210 , \15211 , \15212 , \15213 , \15214 , \15215 , \15216 , \15217 ,
         \15218 , \15219 , \15220 , \15221 , \15222 , \15223 , \15224 , \15225 , \15226 , \15227 ,
         \15228 , \15229 , \15230 , \15231 , \15232 , \15233 , \15234 , \15235 , \15236 , \15237 ,
         \15238 , \15239 , \15240 , \15241 , \15242 , \15243 , \15244 , \15245 , \15246 , \15247 ,
         \15248 , \15249 , \15250 , \15251 , \15252 , \15253 , \15254 , \15255 , \15256 , \15257 ,
         \15258 , \15259 , \15260 , \15261 , \15262 , \15263 , \15264 , \15265 , \15266 , \15267 ,
         \15268 , \15269 , \15270 , \15271 , \15272 , \15273 , \15274 , \15275 , \15276 , \15277 ,
         \15278 , \15279 , \15280 , \15281 , \15282 , \15283 , \15284 , \15285 , \15286 , \15287 ,
         \15288 , \15289 , \15290 , \15291 , \15292 , \15293 , \15294 , \15295 , \15296 , \15297 ,
         \15298 , \15299 , \15300 , \15301 , \15302 , \15303 , \15304 , \15305 , \15306 , \15307 ,
         \15308 , \15309 , \15310 , \15311 , \15312 , \15313 , \15314 , \15315 , \15316 , \15317 ,
         \15318 , \15319 , \15320 , \15321 , \15322 , \15323 , \15324 , \15325 , \15326 , \15327 ,
         \15328 , \15329 , \15330 , \15331 , \15332 , \15333 , \15334 , \15335 , \15336 , \15337 ,
         \15338 , \15339 , \15340 , \15341 , \15342 , \15343 , \15344 , \15345 , \15346 , \15347 ,
         \15348 , \15349 , \15350 , \15351 , \15352 , \15353 , \15354 , \15355 , \15356 , \15357 ,
         \15358 , \15359 , \15360 , \15361 , \15362 , \15363 , \15364 , \15365 , \15366 , \15367 ,
         \15368 , \15369 , \15370 , \15371 , \15372 , \15373 , \15374 , \15375 , \15376 , \15377 ,
         \15378 , \15379 , \15380 , \15381 , \15382 , \15383 , \15384 , \15385 , \15386 , \15387 ,
         \15388 , \15389 , \15390 , \15391 , \15392 , \15393 , \15394 , \15395 , \15396 , \15397 ,
         \15398 , \15399 , \15400 , \15401 , \15402 , \15403 , \15404 , \15405 , \15406 , \15407 ,
         \15408 , \15409 , \15410 , \15411 , \15412 , \15413 , \15414 , \15415 , \15416 , \15417 ,
         \15418 , \15419 , \15420 , \15421 , \15422 , \15423 , \15424 , \15425 , \15426 , \15427 ,
         \15428 , \15429 , \15430 , \15431 , \15432 , \15433 , \15434 , \15435 , \15436 , \15437 ,
         \15438 , \15439 , \15440 , \15441 , \15442 , \15443 , \15444 , \15445 , \15446 , \15447 ,
         \15448 , \15449 , \15450 , \15451 , \15452 , \15453 , \15454 , \15455 , \15456 , \15457 ,
         \15458 , \15459 , \15460 , \15461 , \15462 , \15463 , \15464 , \15465 , \15466 , \15467 ,
         \15468 , \15469 , \15470 , \15471 , \15472 , \15473 , \15474 , \15475 , \15476 , \15477 ,
         \15478 , \15479 , \15480 , \15481 , \15482 , \15483 , \15484 , \15485 , \15486 , \15487 ,
         \15488 , \15489 , \15490 , \15491 , \15492 , \15493 , \15494 , \15495 , \15496 , \15497 ,
         \15498 , \15499 , \15500 , \15501 , \15502 , \15503 , \15504 , \15505 , \15506 , \15507 ,
         \15508 , \15509 , \15510 , \15511 , \15512 , \15513 , \15514 , \15515 , \15516 , \15517 ,
         \15518 , \15519 , \15520 , \15521 , \15522 , \15523 , \15524 , \15525 , \15526 , \15527 ,
         \15528 , \15529 , \15530 , \15531 , \15532 , \15533 , \15534 , \15535 , \15536 , \15537 ,
         \15538 , \15539 , \15540 , \15541 , \15542 , \15543 , \15544 , \15545 , \15546 , \15547 ,
         \15548 , \15549 , \15550 , \15551 , \15552 , \15553 , \15554 , \15555 , \15556 , \15557 ,
         \15558 , \15559 , \15560 , \15561 , \15562 , \15563 , \15564 , \15565 , \15566 , \15567 ,
         \15568 , \15569 , \15570 , \15571 , \15572 , \15573 , \15574 , \15575 , \15576 , \15577 ,
         \15578 , \15579 , \15580 , \15581 , \15582 , \15583 , \15584 , \15585 , \15586 , \15587 ,
         \15588 , \15589 , \15590 , \15591 , \15592 , \15593 , \15594 , \15595 , \15596 , \15597 ,
         \15598 , \15599 , \15600 , \15601 , \15602 , \15603 , \15604 , \15605 , \15606 , \15607 ,
         \15608 , \15609 , \15610 , \15611 , \15612 , \15613 , \15614 , \15615 , \15616 , \15617 ,
         \15618 , \15619 , \15620 , \15621 , \15622 , \15623 , \15624 , \15625 , \15626 , \15627 ,
         \15628 , \15629 , \15630 , \15631 , \15632 , \15633 , \15634 , \15635 , \15636 , \15637 ,
         \15638 , \15639 , \15640 , \15641 , \15642 , \15643 , \15644 , \15645 , \15646 , \15647 ,
         \15648 , \15649 , \15650 , \15651 , \15652 , \15653 , \15654 , \15655 , \15656 , \15657 ,
         \15658 , \15659 , \15660 , \15661 , \15662 , \15663 , \15664 , \15665 , \15666 , \15667 ,
         \15668 , \15669 , \15670 , \15671 , \15672 , \15673 , \15674 , \15675 , \15676 , \15677 ,
         \15678 , \15679 , \15680 , \15681 , \15682 , \15683 , \15684 , \15685 , \15686 , \15687 ,
         \15688 , \15689 , \15690 , \15691 , \15692 , \15693 , \15694 , \15695 , \15696 , \15697 ,
         \15698 , \15699 , \15700 , \15701 , \15702 , \15703 , \15704 , \15705 , \15706 , \15707 ,
         \15708 , \15709 , \15710 , \15711 , \15712 , \15713 , \15714 , \15715 , \15716 , \15717 ,
         \15718 , \15719 , \15720 , \15721 , \15722 , \15723 , \15724 , \15725 , \15726 , \15727 ,
         \15728 , \15729 , \15730 , \15731 , \15732 , \15733 , \15734 , \15735 , \15736 , \15737 ,
         \15738 , \15739 , \15740 , \15741 , \15742 , \15743 , \15744 , \15745 , \15746 , \15747 ,
         \15748 , \15749 , \15750 , \15751 , \15752 , \15753 , \15754 , \15755 , \15756 , \15757 ,
         \15758 , \15759 , \15760 , \15761 , \15762 , \15763 , \15764 , \15765 , \15766 , \15767 ,
         \15768 , \15769 , \15770 , \15771 , \15772 , \15773 , \15774 , \15775 , \15776 , \15777 ,
         \15778 , \15779 , \15780 , \15781 , \15782 , \15783 , \15784 , \15785 , \15786 , \15787 ,
         \15788 , \15789 , \15790 , \15791 , \15792 , \15793 , \15794 , \15795 , \15796 , \15797 ,
         \15798 , \15799 , \15800 , \15801 , \15802 , \15803 , \15804 , \15805 , \15806 , \15807 ,
         \15808 , \15809 , \15810 , \15811 , \15812 , \15813 , \15814 , \15815 , \15816 , \15817 ,
         \15818 , \15819 , \15820 , \15821 , \15822 , \15823 , \15824 , \15825 , \15826 , \15827 ,
         \15828 , \15829 , \15830 , \15831 , \15832 , \15833 , \15834 , \15835 , \15836 , \15837 ,
         \15838 , \15839 , \15840 , \15841 , \15842 , \15843 , \15844 , \15845 , \15846 , \15847 ,
         \15848 , \15849 , \15850 , \15851 , \15852 , \15853 , \15854 , \15855 , \15856 , \15857 ,
         \15858 , \15859 , \15860 , \15861 , \15862 , \15863 , \15864 , \15865 , \15866 , \15867 ,
         \15868 , \15869 , \15870 , \15871 , \15872 , \15873 , \15874 , \15875 , \15876 , \15877 ,
         \15878 , \15879 , \15880 , \15881 , \15882 , \15883 , \15884 , \15885 , \15886 , \15887 ,
         \15888 , \15889 , \15890 , \15891 , \15892 , \15893 , \15894 , \15895 , \15896 , \15897 ,
         \15898 , \15899 , \15900 , \15901 , \15902 , \15903 , \15904 , \15905 , \15906 , \15907 ,
         \15908 , \15909 , \15910 , \15911 , \15912 , \15913 , \15914 , \15915 , \15916 , \15917 ,
         \15918 , \15919 , \15920 , \15921 , \15922 , \15923 , \15924 , \15925 , \15926 , \15927 ,
         \15928 , \15929 , \15930 , \15931 , \15932 , \15933 , \15934 , \15935 , \15936 , \15937 ,
         \15938 , \15939 , \15940 , \15941 , \15942 , \15943 , \15944 , \15945 , \15946 , \15947 ,
         \15948 , \15949 , \15950 , \15951 , \15952 , \15953 , \15954 , \15955 , \15956 , \15957 ,
         \15958 , \15959 , \15960 , \15961 , \15962 , \15963 , \15964 , \15965 , \15966 , \15967 ,
         \15968 , \15969 , \15970 , \15971 , \15972 , \15973 , \15974 , \15975 , \15976 , \15977 ,
         \15978 , \15979 , \15980 , \15981 , \15982 , \15983 , \15984 , \15985 , \15986 , \15987 ,
         \15988 , \15989 , \15990 , \15991 , \15992 , \15993 , \15994 , \15995 , \15996 , \15997 ,
         \15998 , \15999 , \16000 , \16001 , \16002 , \16003 , \16004 , \16005 , \16006 , \16007 ,
         \16008 , \16009 , \16010 , \16011 , \16012 , \16013 , \16014 , \16015 , \16016 , \16017 ,
         \16018 , \16019 , \16020 , \16021 , \16022 , \16023 , \16024 , \16025 , \16026 , \16027 ,
         \16028 , \16029 , \16030 , \16031 , \16032 , \16033 , \16034 , \16035 , \16036 , \16037 ,
         \16038 , \16039 , \16040 , \16041 , \16042 , \16043 , \16044 , \16045 , \16046 , \16047 ,
         \16048 , \16049 , \16050 , \16051 , \16052 , \16053 , \16054 , \16055 , \16056 , \16057 ,
         \16058 , \16059 , \16060 , \16061 , \16062 , \16063 , \16064 , \16065 , \16066 , \16067 ,
         \16068 , \16069 , \16070 , \16071 , \16072 , \16073 , \16074 , \16075 , \16076 , \16077 ,
         \16078 , \16079 , \16080 , \16081 , \16082 , \16083 , \16084 , \16085 , \16086 , \16087 ,
         \16088 , \16089 , \16090 , \16091 , \16092 , \16093 , \16094 , \16095 , \16096 , \16097 ,
         \16098 , \16099 , \16100 , \16101 , \16102 , \16103 , \16104 , \16105 , \16106 , \16107 ,
         \16108 , \16109 , \16110 , \16111 , \16112 , \16113 , \16114 , \16115 , \16116 , \16117 ,
         \16118 , \16119 , \16120 , \16121 , \16122 , \16123 , \16124 , \16125 , \16126 , \16127 ,
         \16128 , \16129 , \16130 , \16131 , \16132 , \16133 , \16134 , \16135 , \16136 , \16137 ,
         \16138 , \16139 , \16140 , \16141 , \16142 , \16143 , \16144 , \16145 , \16146 , \16147 ,
         \16148 , \16149 , \16150 , \16151 , \16152 , \16153 , \16154 , \16155 , \16156 , \16157 ,
         \16158 , \16159 , \16160 , \16161 , \16162 , \16163 , \16164 , \16165 , \16166 , \16167 ,
         \16168 , \16169 , \16170 , \16171 , \16172 , \16173 , \16174 , \16175 , \16176 , \16177 ,
         \16178 , \16179 , \16180 , \16181 , \16182 , \16183 , \16184 , \16185 , \16186 , \16187 ,
         \16188 , \16189 , \16190 , \16191 , \16192 , \16193 , \16194 , \16195 , \16196 , \16197 ,
         \16198 , \16199 , \16200 , \16201 , \16202 , \16203 , \16204 , \16205 , \16206 , \16207 ,
         \16208 , \16209 , \16210 , \16211 , \16212 , \16213 , \16214 , \16215 , \16216 , \16217 ,
         \16218 , \16219 , \16220 , \16221 , \16222 , \16223 , \16224 , \16225 , \16226 , \16227 ,
         \16228 , \16229 , \16230 , \16231 , \16232 , \16233 , \16234 , \16235 , \16236 , \16237 ,
         \16238 , \16239 , \16240 , \16241 , \16242 , \16243 , \16244 , \16245 , \16246 , \16247 ,
         \16248 , \16249 , \16250 , \16251 , \16252 , \16253 , \16254 , \16255 , \16256 , \16257 ,
         \16258 , \16259 , \16260 , \16261 , \16262 , \16263 , \16264 , \16265 , \16266 , \16267 ,
         \16268 , \16269 , \16270 , \16271 , \16272 , \16273 , \16274 , \16275 , \16276 , \16277 ,
         \16278 , \16279 , \16280 , \16281 , \16282 , \16283 , \16284 , \16285 , \16286 , \16287 ,
         \16288 , \16289 , \16290 , \16291 , \16292 , \16293 , \16294 , \16295 , \16296 , \16297 ,
         \16298 , \16299 , \16300 , \16301 , \16302 , \16303 , \16304 , \16305 , \16306 , \16307 ,
         \16308 , \16309 , \16310 , \16311 , \16312 , \16313 , \16314 , \16315 , \16316 , \16317 ,
         \16318 , \16319 , \16320 , \16321 , \16322 , \16323 , \16324 , \16325 , \16326 , \16327 ,
         \16328 , \16329 , \16330 , \16331 , \16332 , \16333 , \16334 , \16335 , \16336 , \16337 ,
         \16338 , \16339 , \16340 , \16341 , \16342 , \16343 , \16344 , \16345 , \16346 , \16347 ,
         \16348 , \16349 , \16350 , \16351 , \16352 , \16353 , \16354 , \16355 , \16356 , \16357 ,
         \16358 , \16359 , \16360 , \16361 , \16362 , \16363 , \16364 , \16365 , \16366 , \16367 ,
         \16368 , \16369 , \16370 , \16371 , \16372 , \16373 , \16374 , \16375 , \16376 , \16377 ,
         \16378 , \16379 , \16380 , \16381 , \16382 , \16383 , \16384 , \16385 , \16386 , \16387 ,
         \16388 , \16389 , \16390 , \16391 , \16392 , \16393 , \16394 , \16395 , \16396 , \16397 ,
         \16398 , \16399 , \16400 , \16401 , \16402 , \16403 , \16404 , \16405 , \16406 , \16407 ,
         \16408 , \16409 , \16410 , \16411 , \16412 , \16413 , \16414 , \16415 , \16416 , \16417 ,
         \16418 , \16419 , \16420 , \16421 , \16422 , \16423 , \16424 , \16425 , \16426 , \16427 ,
         \16428 , \16429 , \16430 , \16431 , \16432 , \16433 , \16434 , \16435 , \16436 , \16437 ,
         \16438 , \16439 , \16440 , \16441 , \16442 , \16443 , \16444 , \16445 , \16446 , \16447 ,
         \16448 , \16449 , \16450 , \16451 , \16452 , \16453 , \16454 , \16455 , \16456 , \16457 ,
         \16458 , \16459 , \16460 , \16461 , \16462 , \16463 , \16464 , \16465 , \16466 , \16467 ,
         \16468 , \16469 , \16470 , \16471 , \16472 , \16473 , \16474 , \16475 , \16476 , \16477 ,
         \16478 , \16479 , \16480 , \16481 , \16482 , \16483 , \16484 , \16485 , \16486 , \16487 ,
         \16488 , \16489 , \16490 , \16491 , \16492 , \16493 , \16494 , \16495 , \16496 , \16497 ,
         \16498 , \16499 , \16500 , \16501 , \16502 , \16503 , \16504 , \16505 , \16506 , \16507 ,
         \16508 , \16509 , \16510 , \16511 , \16512 , \16513 , \16514 , \16515 , \16516 , \16517 ,
         \16518 , \16519 , \16520 , \16521 , \16522 , \16523 , \16524 , \16525 , \16526 , \16527 ,
         \16528 , \16529 , \16530 , \16531 , \16532 , \16533 , \16534 , \16535 , \16536 , \16537 ,
         \16538 , \16539 , \16540 , \16541 , \16542 , \16543 , \16544 , \16545 , \16546 , \16547 ,
         \16548 , \16549 , \16550 , \16551 , \16552 , \16553 , \16554 , \16555 , \16556 , \16557 ,
         \16558 , \16559 , \16560 , \16561 , \16562 , \16563 , \16564 , \16565 , \16566 , \16567 ,
         \16568 , \16569 , \16570 , \16571 , \16572 , \16573 , \16574 , \16575 , \16576 , \16577 ,
         \16578 , \16579 , \16580 , \16581 , \16582 , \16583 , \16584 , \16585 , \16586 , \16587 ,
         \16588 , \16589 , \16590 , \16591 , \16592 , \16593 , \16594 , \16595 , \16596 , \16597 ,
         \16598 , \16599 , \16600 , \16601 , \16602 , \16603 , \16604 , \16605 , \16606 , \16607 ,
         \16608 , \16609 , \16610 , \16611 , \16612 , \16613 , \16614 , \16615 , \16616 , \16617 ,
         \16618 , \16619 , \16620 , \16621 , \16622 , \16623 , \16624 , \16625 , \16626 , \16627 ,
         \16628 , \16629 , \16630 , \16631 , \16632 , \16633 , \16634 , \16635 , \16636 , \16637 ,
         \16638 , \16639 , \16640 , \16641 , \16642 , \16643 , \16644 , \16645 , \16646 , \16647 ,
         \16648 , \16649 , \16650 , \16651 , \16652 , \16653 , \16654 , \16655 , \16656 , \16657 ,
         \16658 , \16659 , \16660 , \16661 , \16662 , \16663 , \16664 , \16665 , \16666 , \16667 ,
         \16668 , \16669 , \16670 , \16671 , \16672 , \16673 , \16674 , \16675 , \16676 , \16677 ,
         \16678 , \16679 , \16680 , \16681 , \16682 , \16683 , \16684 , \16685 , \16686 , \16687 ,
         \16688 , \16689 , \16690 , \16691 , \16692 , \16693 , \16694 , \16695 , \16696 , \16697 ,
         \16698 , \16699 , \16700 , \16701 , \16702 , \16703 , \16704 , \16705 , \16706 , \16707 ,
         \16708 , \16709 , \16710 , \16711 , \16712 , \16713 , \16714 , \16715 , \16716 , \16717 ,
         \16718 , \16719 , \16720 , \16721 , \16722 , \16723 , \16724 , \16725 , \16726 , \16727 ,
         \16728 , \16729 , \16730 , \16731 , \16732 , \16733 , \16734 , \16735 , \16736 , \16737 ,
         \16738 , \16739 , \16740 , \16741 , \16742 , \16743 , \16744 , \16745 , \16746 , \16747 ,
         \16748 , \16749 , \16750 , \16751 , \16752 , \16753 , \16754 , \16755 , \16756 , \16757 ,
         \16758 , \16759 , \16760 , \16761 , \16762 , \16763 , \16764 , \16765 , \16766 , \16767 ,
         \16768 , \16769 , \16770 , \16771 , \16772 , \16773 , \16774 , \16775 , \16776 , \16777 ,
         \16778 , \16779 , \16780 , \16781 , \16782 , \16783 , \16784 , \16785 , \16786 , \16787 ,
         \16788 , \16789 , \16790 , \16791 , \16792 , \16793 , \16794 , \16795 , \16796 , \16797 ,
         \16798 , \16799 , \16800 , \16801 , \16802 , \16803 , \16804 , \16805 , \16806 , \16807 ,
         \16808 , \16809 , \16810 , \16811 , \16812 , \16813 , \16814 , \16815 , \16816 , \16817 ,
         \16818 , \16819 , \16820 , \16821 , \16822 , \16823 , \16824 , \16825 , \16826 , \16827 ,
         \16828 , \16829 , \16830 , \16831 , \16832 , \16833 , \16834 , \16835 , \16836 , \16837 ,
         \16838 , \16839 , \16840 , \16841 , \16842 , \16843 , \16844 , \16845 , \16846 , \16847 ,
         \16848 , \16849 , \16850 , \16851 , \16852 , \16853 , \16854 , \16855 , \16856 , \16857 ,
         \16858 , \16859 , \16860 , \16861 , \16862 , \16863 , \16864 , \16865 , \16866 , \16867 ,
         \16868 , \16869 , \16870 , \16871 , \16872 , \16873 , \16874 , \16875 , \16876 , \16877 ,
         \16878 , \16879 , \16880 , \16881 , \16882 , \16883 , \16884 , \16885 , \16886 , \16887 ,
         \16888 , \16889 , \16890 , \16891 , \16892 , \16893 , \16894 , \16895 , \16896 , \16897 ,
         \16898 , \16899 , \16900 , \16901 , \16902 , \16903 , \16904 , \16905 , \16906 , \16907 ,
         \16908 , \16909 , \16910 , \16911 , \16912 , \16913 , \16914 , \16915 , \16916 , \16917 ,
         \16918 , \16919 , \16920 , \16921 , \16922 , \16923 , \16924 , \16925 , \16926 , \16927 ,
         \16928 , \16929 , \16930 , \16931 , \16932 , \16933 , \16934 , \16935 , \16936 , \16937 ,
         \16938 , \16939 , \16940 , \16941 , \16942 , \16943 , \16944 , \16945 , \16946 , \16947 ,
         \16948 , \16949 , \16950 , \16951 , \16952 , \16953 , \16954 , \16955 , \16956 , \16957 ,
         \16958 , \16959 , \16960 , \16961 , \16962 , \16963 , \16964 , \16965 , \16966 , \16967 ,
         \16968 , \16969 , \16970 , \16971 , \16972 , \16973 , \16974 , \16975 , \16976 , \16977 ,
         \16978 , \16979 , \16980 , \16981 , \16982 , \16983 , \16984 , \16985 , \16986 , \16987 ,
         \16988 , \16989 , \16990 , \16991 , \16992 , \16993 , \16994 , \16995 , \16996 , \16997 ,
         \16998 , \16999 , \17000 , \17001 , \17002 , \17003 , \17004 , \17005 , \17006 , \17007 ,
         \17008 , \17009 , \17010 , \17011 , \17012 , \17013 , \17014 , \17015 , \17016 , \17017 ,
         \17018 , \17019 , \17020 , \17021 , \17022 , \17023 , \17024 , \17025 , \17026 , \17027 ,
         \17028 , \17029 , \17030 , \17031 , \17032 , \17033 , \17034 , \17035 , \17036 , \17037 ,
         \17038 , \17039 , \17040 , \17041 , \17042 , \17043 , \17044 , \17045 , \17046 , \17047 ,
         \17048 , \17049 , \17050 , \17051 , \17052 , \17053 , \17054 , \17055 , \17056 , \17057 ,
         \17058 , \17059 , \17060 , \17061 , \17062 , \17063 , \17064 , \17065 , \17066 , \17067 ,
         \17068 , \17069 , \17070 , \17071 , \17072 , \17073 , \17074 , \17075 , \17076 , \17077 ,
         \17078 , \17079 , \17080 , \17081 , \17082 , \17083 , \17084 , \17085 , \17086 , \17087 ,
         \17088 , \17089 , \17090 , \17091 , \17092 , \17093 , \17094 , \17095 , \17096 , \17097 ,
         \17098 , \17099 , \17100 , \17101 , \17102 , \17103 , \17104 , \17105 , \17106 , \17107 ,
         \17108 , \17109 , \17110 , \17111 , \17112 , \17113 , \17114 , \17115 , \17116 , \17117 ,
         \17118 , \17119 , \17120 , \17121 , \17122 , \17123 , \17124 , \17125 , \17126 , \17127 ,
         \17128 , \17129 , \17130 , \17131 , \17132 , \17133 , \17134 , \17135 , \17136 , \17137 ,
         \17138 , \17139 , \17140 , \17141 , \17142 , \17143 , \17144 , \17145 , \17146 , \17147 ,
         \17148 , \17149 , \17150 , \17151 , \17152 , \17153 , \17154 , \17155 , \17156 , \17157 ,
         \17158 , \17159 , \17160 , \17161 , \17162 , \17163 , \17164 , \17165 , \17166 , \17167 ,
         \17168 , \17169 , \17170 , \17171 , \17172 , \17173 , \17174 , \17175 , \17176 , \17177 ,
         \17178 , \17179 , \17180 , \17181 , \17182 , \17183 , \17184 , \17185 , \17186 , \17187 ,
         \17188 , \17189 , \17190 , \17191 , \17192 , \17193 , \17194 , \17195 , \17196 , \17197 ,
         \17198 , \17199 , \17200 , \17201 , \17202 , \17203 , \17204 , \17205 , \17206 , \17207 ,
         \17208 , \17209 , \17210 , \17211 , \17212 , \17213 , \17214 , \17215 , \17216 , \17217 ,
         \17218 , \17219 , \17220 , \17221 , \17222 , \17223 , \17224 , \17225 , \17226 , \17227 ,
         \17228 , \17229 , \17230 , \17231 , \17232 , \17233 , \17234 , \17235 , \17236 , \17237 ,
         \17238 , \17239 , \17240 , \17241 , \17242 , \17243 , \17244 , \17245 , \17246 , \17247 ,
         \17248 , \17249 , \17250 , \17251 , \17252 , \17253 , \17254 , \17255 , \17256 , \17257 ,
         \17258 , \17259 , \17260 , \17261 , \17262 , \17263 , \17264 , \17265 , \17266 , \17267 ,
         \17268 , \17269 , \17270 , \17271 , \17272 , \17273 , \17274 , \17275 , \17276 , \17277 ,
         \17278 , \17279 , \17280 , \17281 , \17282 , \17283 , \17284 , \17285 , \17286 , \17287 ,
         \17288 , \17289 , \17290 , \17291 , \17292 , \17293 , \17294 , \17295 , \17296 , \17297 ,
         \17298 , \17299 , \17300 , \17301 , \17302 , \17303 , \17304 , \17305 , \17306 , \17307 ,
         \17308 , \17309 , \17310 , \17311 , \17312 , \17313 , \17314 , \17315 , \17316 , \17317 ,
         \17318 , \17319 , \17320 , \17321 , \17322 , \17323 , \17324 , \17325 , \17326 , \17327 ,
         \17328 , \17329 , \17330 , \17331 , \17332 , \17333 , \17334 , \17335 , \17336 , \17337 ,
         \17338 , \17339 , \17340 , \17341 , \17342 , \17343 , \17344 , \17345 , \17346 , \17347 ,
         \17348 , \17349 , \17350 , \17351 , \17352 , \17353 , \17354 , \17355 , \17356 , \17357 ,
         \17358 , \17359 , \17360 , \17361 , \17362 , \17363 , \17364 , \17365 , \17366 , \17367 ,
         \17368 , \17369 , \17370 , \17371 , \17372 , \17373 , \17374 , \17375 , \17376 , \17377 ,
         \17378 , \17379 , \17380 , \17381 , \17382 , \17383 , \17384 , \17385 , \17386 , \17387 ,
         \17388 , \17389 , \17390 , \17391 , \17392 , \17393 , \17394 , \17395 , \17396 , \17397 ,
         \17398 , \17399 , \17400 , \17401 , \17402 , \17403 , \17404 , \17405 , \17406 , \17407 ,
         \17408 , \17409 , \17410 , \17411 , \17412 , \17413 , \17414 , \17415 , \17416 , \17417 ,
         \17418 , \17419 , \17420 , \17421 , \17422 , \17423 , \17424 , \17425 , \17426 , \17427 ,
         \17428 , \17429 , \17430 , \17431 , \17432 , \17433 , \17434 , \17435 , \17436 , \17437 ,
         \17438 , \17439 , \17440 , \17441 , \17442 , \17443 , \17444 , \17445 , \17446 , \17447 ,
         \17448 , \17449 , \17450 , \17451 , \17452 , \17453 , \17454 , \17455 , \17456 , \17457 ,
         \17458 , \17459 , \17460 , \17461 , \17462 , \17463 , \17464 , \17465 , \17466 , \17467 ,
         \17468 , \17469 , \17470 , \17471 , \17472 , \17473 , \17474 , \17475 , \17476 , \17477 ,
         \17478 , \17479 , \17480 , \17481 , \17482 , \17483 , \17484 , \17485 , \17486 , \17487 ,
         \17488 , \17489 , \17490 , \17491 , \17492 , \17493 , \17494 , \17495 , \17496 , \17497 ,
         \17498 , \17499 , \17500 , \17501 , \17502 , \17503 , \17504 , \17505 , \17506 , \17507 ,
         \17508 , \17509 , \17510 , \17511 , \17512 , \17513 , \17514 , \17515 , \17516 , \17517 ,
         \17518 , \17519 , \17520 , \17521 , \17522 , \17523 , \17524 , \17525 , \17526 , \17527 ,
         \17528 , \17529 , \17530 , \17531 , \17532 , \17533 , \17534 , \17535 , \17536 , \17537 ,
         \17538 , \17539 , \17540 , \17541 , \17542 , \17543 , \17544 , \17545 , \17546 , \17547 ,
         \17548 , \17549 , \17550 , \17551 , \17552 , \17553 , \17554 , \17555 , \17556 , \17557 ,
         \17558 , \17559 , \17560 , \17561 , \17562 , \17563 , \17564 , \17565 , \17566 , \17567 ,
         \17568 , \17569 , \17570 , \17571 , \17572 , \17573 , \17574 , \17575 , \17576 , \17577 ,
         \17578 , \17579 , \17580 , \17581 , \17582 , \17583 , \17584 , \17585 , \17586 , \17587 ,
         \17588 , \17589 , \17590 , \17591 , \17592 , \17593 , \17594 , \17595 , \17596 , \17597 ,
         \17598 , \17599 , \17600 , \17601 , \17602 , \17603 , \17604 , \17605 , \17606 , \17607 ,
         \17608 , \17609 , \17610 , \17611 , \17612 , \17613 , \17614 , \17615 , \17616 , \17617 ,
         \17618 , \17619 , \17620 , \17621 , \17622 , \17623 , \17624 , \17625 , \17626 , \17627 ,
         \17628 , \17629 , \17630 , \17631 , \17632 , \17633 , \17634 , \17635 , \17636 , \17637 ,
         \17638 , \17639 , \17640 , \17641 , \17642 , \17643 , \17644 , \17645 , \17646 , \17647 ,
         \17648 , \17649 , \17650 , \17651 , \17652 , \17653 , \17654 , \17655 , \17656 , \17657 ,
         \17658 , \17659 , \17660 , \17661 , \17662 , \17663 , \17664 , \17665 , \17666 , \17667 ,
         \17668 , \17669 , \17670 , \17671 , \17672 , \17673 , \17674 , \17675 , \17676 , \17677 ,
         \17678 , \17679 , \17680 , \17681 , \17682 , \17683 , \17684 , \17685 , \17686 , \17687 ,
         \17688 , \17689 , \17690 , \17691 , \17692 , \17693 , \17694 , \17695 , \17696 , \17697 ,
         \17698 , \17699 , \17700 , \17701 , \17702 , \17703 , \17704 , \17705 , \17706 , \17707 ,
         \17708 , \17709 , \17710 , \17711 , \17712 , \17713 , \17714 , \17715 , \17716 , \17717 ,
         \17718 , \17719 , \17720 , \17721 , \17722 , \17723 , \17724 , \17725 , \17726 , \17727 ,
         \17728 , \17729 , \17730 , \17731 , \17732 , \17733 , \17734 , \17735 , \17736 , \17737 ,
         \17738 , \17739 , \17740 , \17741 , \17742 , \17743 , \17744 , \17745 , \17746 , \17747 ,
         \17748 , \17749 , \17750 , \17751 , \17752 , \17753 , \17754 , \17755 , \17756 , \17757 ,
         \17758 , \17759 , \17760 , \17761 , \17762 , \17763 , \17764 , \17765 , \17766 , \17767 ,
         \17768 , \17769 , \17770 , \17771 , \17772 , \17773 , \17774 , \17775 , \17776 , \17777 ,
         \17778 , \17779 , \17780 , \17781 , \17782 , \17783 , \17784 , \17785 , \17786 , \17787 ,
         \17788 , \17789 , \17790 , \17791 , \17792 , \17793 , \17794 , \17795 , \17796 , \17797 ,
         \17798 , \17799 , \17800 , \17801 , \17802 , \17803 , \17804 , \17805 , \17806 , \17807 ,
         \17808 , \17809 , \17810 , \17811 , \17812 , \17813 , \17814 , \17815 , \17816 , \17817 ,
         \17818 , \17819 , \17820 , \17821 , \17822 , \17823 , \17824 , \17825 , \17826 , \17827 ,
         \17828 , \17829 , \17830 , \17831 , \17832 , \17833 , \17834 , \17835 , \17836 , \17837 ,
         \17838 , \17839 , \17840 , \17841 , \17842 , \17843 , \17844 , \17845 , \17846 , \17847 ,
         \17848 , \17849 , \17850 , \17851 , \17852 , \17853 , \17854 , \17855 , \17856 , \17857 ,
         \17858 , \17859 , \17860 , \17861 , \17862 , \17863 , \17864 , \17865 , \17866 , \17867 ,
         \17868 , \17869 , \17870 , \17871 , \17872 , \17873 , \17874 , \17875 , \17876 , \17877 ,
         \17878 , \17879 , \17880 , \17881 , \17882 , \17883 , \17884 , \17885 , \17886 , \17887 ,
         \17888 , \17889 , \17890 , \17891 , \17892 , \17893 , \17894 , \17895 , \17896 , \17897 ,
         \17898 , \17899 , \17900 , \17901 , \17902 , \17903 , \17904 , \17905 , \17906 , \17907 ,
         \17908 , \17909 , \17910 , \17911 , \17912 , \17913 , \17914 , \17915 , \17916 , \17917 ,
         \17918 , \17919 , \17920 , \17921 , \17922 , \17923 , \17924 , \17925 , \17926 , \17927 ,
         \17928 , \17929 , \17930 , \17931 , \17932 , \17933 , \17934 , \17935 , \17936 , \17937 ,
         \17938 , \17939 , \17940 , \17941 , \17942 , \17943 , \17944 , \17945 , \17946 , \17947 ,
         \17948 , \17949 , \17950 , \17951 , \17952 , \17953 , \17954 , \17955 , \17956 , \17957 ,
         \17958 , \17959 , \17960 , \17961 , \17962 , \17963 , \17964 , \17965 , \17966 , \17967 ,
         \17968 , \17969 , \17970 , \17971 , \17972 , \17973 , \17974 , \17975 , \17976 , \17977 ,
         \17978 , \17979 , \17980 , \17981 , \17982 , \17983 , \17984 , \17985 , \17986 , \17987 ,
         \17988 , \17989 , \17990 , \17991 , \17992 , \17993 , \17994 , \17995 , \17996 , \17997 ,
         \17998 , \17999 , \18000 , \18001 , \18002 , \18003 , \18004 , \18005 , \18006 , \18007 ,
         \18008 , \18009 , \18010 , \18011 , \18012 , \18013 , \18014 , \18015 , \18016 , \18017 ,
         \18018 , \18019 , \18020 , \18021 , \18022 , \18023 , \18024 , \18025 , \18026 , \18027 ,
         \18028 , \18029 , \18030 , \18031 , \18032 , \18033 , \18034 , \18035 , \18036 , \18037 ,
         \18038 , \18039 , \18040 , \18041 , \18042 , \18043 , \18044 , \18045 , \18046 , \18047 ,
         \18048 , \18049 , \18050 , \18051 , \18052 , \18053 , \18054 , \18055 , \18056 , \18057 ,
         \18058 , \18059 , \18060 , \18061 , \18062 , \18063 , \18064 , \18065 , \18066 , \18067 ,
         \18068 , \18069 , \18070 , \18071 , \18072 , \18073 , \18074 , \18075 , \18076 , \18077 ,
         \18078 , \18079 , \18080 , \18081 , \18082 , \18083 , \18084 , \18085 , \18086 , \18087 ,
         \18088 , \18089 , \18090 , \18091 , \18092 , \18093 , \18094 , \18095 , \18096 , \18097 ,
         \18098 , \18099 , \18100 , \18101 , \18102 , \18103 , \18104 , \18105 , \18106 , \18107 ,
         \18108 , \18109 , \18110 , \18111 , \18112 , \18113 , \18114 , \18115 , \18116 , \18117 ,
         \18118 , \18119 , \18120 , \18121 , \18122 , \18123 , \18124 , \18125 , \18126 , \18127 ,
         \18128 , \18129 , \18130 , \18131 , \18132 , \18133 , \18134 , \18135 , \18136 , \18137 ,
         \18138 , \18139 , \18140 , \18141 , \18142 , \18143 , \18144 , \18145 , \18146 , \18147 ,
         \18148 , \18149 , \18150 , \18151 , \18152 , \18153 , \18154 , \18155 , \18156 , \18157 ,
         \18158 , \18159 , \18160 , \18161 , \18162 , \18163 , \18164 , \18165 , \18166 , \18167 ,
         \18168 , \18169 , \18170 , \18171 , \18172 , \18173 , \18174 , \18175 , \18176 , \18177 ,
         \18178 , \18179 , \18180 , \18181 , \18182 , \18183 , \18184 , \18185 , \18186 , \18187 ,
         \18188 , \18189 , \18190 , \18191 , \18192 , \18193 , \18194 , \18195 , \18196 , \18197 ,
         \18198 , \18199 , \18200 , \18201 , \18202 , \18203 , \18204 , \18205 , \18206 , \18207 ,
         \18208 , \18209 , \18210 , \18211 , \18212 , \18213 , \18214 , \18215 , \18216 , \18217 ,
         \18218 , \18219 , \18220 , \18221 , \18222 , \18223 , \18224 , \18225 , \18226 , \18227 ,
         \18228 , \18229 , \18230 , \18231 , \18232 , \18233 , \18234 , \18235 , \18236 , \18237 ,
         \18238 , \18239 , \18240 , \18241 , \18242 , \18243 , \18244 , \18245 , \18246 , \18247 ,
         \18248 , \18249 , \18250 , \18251 , \18252 , \18253 , \18254 , \18255 , \18256 , \18257 ,
         \18258 , \18259 , \18260 , \18261 , \18262 , \18263 , \18264 , \18265 , \18266 , \18267 ,
         \18268 , \18269 , \18270 , \18271 , \18272 , \18273 , \18274 , \18275 , \18276 , \18277 ,
         \18278 , \18279 , \18280 , \18281 , \18282 , \18283 , \18284 , \18285 , \18286 , \18287 ,
         \18288 , \18289 , \18290 , \18291 , \18292 , \18293 , \18294 , \18295 , \18296 , \18297 ,
         \18298 , \18299 , \18300 , \18301 , \18302 , \18303 , \18304 , \18305 , \18306 , \18307 ,
         \18308 , \18309 , \18310 , \18311 , \18312 , \18313 , \18314 , \18315 , \18316 , \18317 ,
         \18318 , \18319 , \18320 , \18321 , \18322 , \18323 , \18324 , \18325 , \18326 , \18327 ,
         \18328 , \18329 , \18330 , \18331 , \18332 , \18333 , \18334 , \18335 , \18336 , \18337 ,
         \18338 , \18339 , \18340 , \18341 , \18342 , \18343 , \18344 , \18345 , \18346 , \18347 ,
         \18348 , \18349 , \18350 , \18351 , \18352 , \18353 , \18354 , \18355 , \18356 , \18357 ,
         \18358 , \18359 , \18360 , \18361 , \18362 , \18363 , \18364 , \18365 , \18366 , \18367 ,
         \18368 , \18369 , \18370 , \18371 , \18372 , \18373 , \18374 , \18375 , \18376 , \18377 ,
         \18378 , \18379 , \18380 , \18381 , \18382 , \18383 , \18384 , \18385 , \18386 , \18387 ,
         \18388 , \18389 , \18390 , \18391 , \18392 , \18393 , \18394 , \18395 , \18396 , \18397 ,
         \18398 , \18399 , \18400 , \18401 , \18402 , \18403 , \18404 , \18405 , \18406 , \18407 ,
         \18408 , \18409 , \18410 , \18411 , \18412 , \18413 , \18414 , \18415 , \18416 , \18417 ,
         \18418 , \18419 , \18420 , \18421 , \18422 , \18423 , \18424 , \18425 , \18426 , \18427 ,
         \18428 , \18429 , \18430 , \18431 , \18432 , \18433 , \18434 , \18435 , \18436 , \18437 ,
         \18438 , \18439 , \18440 , \18441 , \18442 , \18443 , \18444 , \18445 , \18446 , \18447 ,
         \18448 , \18449 , \18450 , \18451 , \18452 , \18453 , \18454 , \18455 , \18456 , \18457 ,
         \18458 , \18459 , \18460 , \18461 , \18462 , \18463 , \18464 , \18465 , \18466 , \18467 ,
         \18468 , \18469 , \18470 , \18471 , \18472 , \18473 , \18474 , \18475 , \18476 , \18477 ,
         \18478 , \18479 , \18480 , \18481 , \18482 , \18483 , \18484 , \18485 , \18486 , \18487 ,
         \18488 , \18489 , \18490 , \18491 , \18492 , \18493 , \18494 , \18495 , \18496 , \18497 ,
         \18498 , \18499 , \18500 , \18501 , \18502 , \18503 , \18504 , \18505 , \18506 , \18507 ,
         \18508 , \18509 , \18510 , \18511 , \18512 , \18513 , \18514 , \18515 , \18516 , \18517 ,
         \18518 , \18519 , \18520 , \18521 , \18522 , \18523 , \18524 , \18525 , \18526 , \18527 ,
         \18528 , \18529 , \18530 , \18531 , \18532 , \18533 , \18534 , \18535 , \18536 , \18537 ,
         \18538 , \18539 , \18540 , \18541 , \18542 , \18543 , \18544 , \18545 , \18546 , \18547 ,
         \18548 , \18549 , \18550 , \18551 , \18552 , \18553 , \18554 , \18555 , \18556 , \18557 ,
         \18558 , \18559 , \18560 , \18561 , \18562 , \18563 , \18564 , \18565 , \18566 , \18567 ,
         \18568 , \18569 , \18570 , \18571 , \18572 , \18573 , \18574 , \18575 , \18576 , \18577 ,
         \18578 , \18579 , \18580 , \18581 , \18582 , \18583 , \18584 , \18585 , \18586 , \18587 ,
         \18588 , \18589 , \18590 , \18591 , \18592 , \18593 , \18594 , \18595 , \18596 , \18597 ,
         \18598 , \18599 , \18600 , \18601 , \18602 , \18603 , \18604 , \18605 , \18606 , \18607 ,
         \18608 , \18609 , \18610 , \18611 , \18612 , \18613 , \18614 , \18615 , \18616 , \18617 ,
         \18618 , \18619 , \18620 , \18621 , \18622 , \18623 , \18624 , \18625 , \18626 , \18627 ,
         \18628 , \18629 , \18630 , \18631 , \18632 , \18633 , \18634 , \18635 , \18636 , \18637 ,
         \18638 , \18639 , \18640 , \18641 , \18642 , \18643 , \18644 , \18645 , \18646 , \18647 ,
         \18648 , \18649 , \18650 , \18651 , \18652 , \18653 , \18654 , \18655 , \18656 , \18657 ,
         \18658 , \18659 , \18660 , \18661 , \18662 , \18663 , \18664 , \18665 , \18666 , \18667 ,
         \18668 , \18669 , \18670 , \18671 , \18672 , \18673 , \18674 , \18675 , \18676 , \18677 ,
         \18678 , \18679 , \18680 , \18681 , \18682 , \18683 , \18684 , \18685 , \18686 , \18687 ,
         \18688 , \18689 , \18690 , \18691 , \18692 , \18693 , \18694 , \18695 , \18696 , \18697 ,
         \18698 , \18699 , \18700 , \18701 , \18702 , \18703 , \18704 , \18705 , \18706 , \18707 ,
         \18708 , \18709 , \18710 , \18711 , \18712 , \18713 , \18714 , \18715 , \18716 , \18717 ,
         \18718 , \18719 , \18720 , \18721 , \18722 , \18723 , \18724 , \18725 , \18726 , \18727 ,
         \18728 , \18729 , \18730 , \18731 , \18732 , \18733 , \18734 , \18735 , \18736 , \18737 ,
         \18738 , \18739 , \18740 , \18741 , \18742 , \18743 , \18744 , \18745 , \18746 , \18747 ,
         \18748 , \18749 , \18750 , \18751 , \18752 , \18753 , \18754 , \18755 , \18756 , \18757 ,
         \18758 , \18759 , \18760 , \18761 , \18762 , \18763 , \18764 , \18765 , \18766 , \18767 ,
         \18768 , \18769 , \18770 , \18771 , \18772 , \18773 , \18774 , \18775 , \18776 , \18777 ,
         \18778 , \18779 , \18780 , \18781 , \18782 , \18783 , \18784 , \18785 , \18786 , \18787 ,
         \18788 , \18789 , \18790 , \18791 , \18792 , \18793 , \18794 , \18795 , \18796 , \18797 ,
         \18798 , \18799 , \18800 , \18801 , \18802 , \18803 , \18804 , \18805 , \18806 , \18807 ,
         \18808 , \18809 , \18810 , \18811 , \18812 , \18813 , \18814 , \18815 , \18816 , \18817 ,
         \18818 , \18819 , \18820 , \18821 , \18822 , \18823 , \18824 , \18825 , \18826 , \18827 ,
         \18828 , \18829 , \18830 , \18831 , \18832 , \18833 , \18834 , \18835 , \18836 , \18837 ,
         \18838 , \18839 , \18840 , \18841 , \18842 , \18843 , \18844 , \18845 , \18846 , \18847 ,
         \18848 , \18849 , \18850 , \18851 , \18852 , \18853 , \18854 , \18855 , \18856 , \18857 ,
         \18858 , \18859 , \18860 , \18861 , \18862 , \18863 , \18864 , \18865 , \18866 , \18867 ,
         \18868 , \18869 , \18870 , \18871 , \18872 , \18873 , \18874 , \18875 , \18876 , \18877 ,
         \18878 , \18879 , \18880 , \18881 , \18882 , \18883 , \18884 , \18885 , \18886 , \18887 ,
         \18888 , \18889 , \18890 , \18891 , \18892 , \18893 , \18894 , \18895 , \18896 , \18897 ,
         \18898 , \18899 , \18900 , \18901 , \18902 , \18903 , \18904 , \18905 , \18906 , \18907 ,
         \18908 , \18909 , \18910 , \18911 , \18912 , \18913 , \18914 , \18915 , \18916 , \18917 ,
         \18918 , \18919 , \18920 , \18921 , \18922 , \18923 , \18924 , \18925 , \18926 , \18927 ,
         \18928 , \18929 , \18930 , \18931 , \18932 , \18933 , \18934 , \18935 , \18936 , \18937 ,
         \18938 , \18939 , \18940 , \18941 , \18942 , \18943 , \18944 , \18945 , \18946 , \18947 ,
         \18948 , \18949 , \18950 , \18951 , \18952 , \18953 , \18954 , \18955 , \18956 , \18957 ,
         \18958 , \18959 , \18960 , \18961 , \18962 , \18963 , \18964 , \18965 , \18966 , \18967 ,
         \18968 , \18969 , \18970 , \18971 , \18972 , \18973 , \18974 , \18975 , \18976 , \18977 ,
         \18978 , \18979 , \18980 , \18981 , \18982 , \18983 , \18984 , \18985 , \18986 , \18987 ,
         \18988 , \18989 , \18990 , \18991 , \18992 , \18993 , \18994 , \18995 , \18996 , \18997 ,
         \18998 , \18999 , \19000 , \19001 , \19002 , \19003 , \19004 , \19005 , \19006 , \19007 ,
         \19008 , \19009 , \19010 , \19011 , \19012 , \19013 , \19014 , \19015 , \19016 , \19017 ,
         \19018 , \19019 , \19020 , \19021 , \19022 , \19023 , \19024 , \19025 , \19026 , \19027 ,
         \19028 , \19029 , \19030 , \19031 , \19032 , \19033 , \19034 , \19035 , \19036 , \19037 ,
         \19038 , \19039 , \19040 , \19041 , \19042 , \19043 , \19044 , \19045 , \19046 , \19047 ,
         \19048 , \19049 , \19050 , \19051 , \19052 , \19053 , \19054 , \19055 , \19056 , \19057 ,
         \19058 , \19059 , \19060 , \19061 , \19062 , \19063 , \19064 , \19065 , \19066 , \19067 ,
         \19068 , \19069 , \19070 , \19071 , \19072 , \19073 , \19074 , \19075 , \19076 , \19077 ,
         \19078 , \19079 , \19080 , \19081 , \19082 , \19083 , \19084 , \19085 , \19086 , \19087 ,
         \19088 , \19089 , \19090 , \19091 , \19092 , \19093 , \19094 , \19095 , \19096 , \19097 ,
         \19098 , \19099 , \19100 , \19101 , \19102 , \19103 , \19104 , \19105 , \19106 , \19107 ,
         \19108 , \19109 , \19110 , \19111 , \19112 , \19113 , \19114 , \19115 , \19116 , \19117 ,
         \19118 , \19119 , \19120 , \19121 , \19122 , \19123 , \19124 , \19125 , \19126 , \19127 ,
         \19128 , \19129 , \19130 , \19131 , \19132 , \19133 , \19134 , \19135 , \19136 , \19137 ,
         \19138 , \19139 , \19140 , \19141 , \19142 , \19143 , \19144 , \19145 , \19146 , \19147 ,
         \19148 , \19149 , \19150 , \19151 , \19152 , \19153 , \19154 , \19155 , \19156 , \19157 ,
         \19158 , \19159 , \19160 , \19161 , \19162 , \19163 , \19164 , \19165 , \19166 , \19167 ,
         \19168 , \19169 , \19170 , \19171 , \19172 , \19173 , \19174 , \19175 , \19176 , \19177 ,
         \19178 , \19179 , \19180 , \19181 , \19182 , \19183 , \19184 , \19185 , \19186 , \19187 ,
         \19188 , \19189 , \19190 , \19191 , \19192 , \19193 , \19194 , \19195 , \19196 , \19197 ,
         \19198 , \19199 , \19200 , \19201 , \19202 , \19203 , \19204 , \19205 , \19206 , \19207 ,
         \19208 , \19209 , \19210 , \19211 , \19212 , \19213 , \19214 , \19215 , \19216 , \19217 ,
         \19218 , \19219 , \19220 , \19221 , \19222 , \19223 , \19224 , \19225 , \19226 , \19227 ,
         \19228 , \19229 , \19230 , \19231 , \19232 , \19233 , \19234 , \19235 , \19236 , \19237 ,
         \19238 , \19239 , \19240 , \19241 , \19242 , \19243 , \19244 , \19245 , \19246 , \19247 ,
         \19248 , \19249 , \19250 , \19251 , \19252 , \19253 , \19254 , \19255 , \19256 , \19257 ,
         \19258 , \19259 , \19260 , \19261 , \19262 , \19263 , \19264 , \19265 , \19266 , \19267 ,
         \19268 , \19269 , \19270 , \19271 , \19272 , \19273 , \19274 , \19275 , \19276 , \19277 ,
         \19278 , \19279 , \19280 , \19281 , \19282 , \19283 , \19284 , \19285 , \19286 , \19287 ,
         \19288 , \19289 , \19290 , \19291 , \19292 , \19293 , \19294 , \19295 , \19296 , \19297 ,
         \19298 , \19299 , \19300 , \19301 , \19302 , \19303 , \19304 , \19305 , \19306 , \19307 ,
         \19308 , \19309 , \19310 , \19311 , \19312 , \19313 , \19314 , \19315 , \19316 , \19317 ,
         \19318 , \19319 , \19320 , \19321 , \19322 , \19323 , \19324 , \19325 , \19326 , \19327 ,
         \19328 , \19329 , \19330 , \19331 , \19332 , \19333 , \19334 , \19335 , \19336 , \19337 ,
         \19338 , \19339 , \19340 , \19341 , \19342 , \19343 , \19344 , \19345 , \19346 , \19347 ,
         \19348 , \19349 , \19350 , \19351 , \19352 , \19353 , \19354 , \19355 , \19356 , \19357 ,
         \19358 , \19359 , \19360 , \19361 , \19362 , \19363 , \19364 , \19365 , \19366 , \19367 ,
         \19368 , \19369 , \19370 , \19371 , \19372 , \19373 , \19374 , \19375 , \19376 , \19377 ,
         \19378 , \19379 , \19380 , \19381 , \19382 , \19383 , \19384 , \19385 , \19386 , \19387 ,
         \19388 , \19389 , \19390 , \19391 , \19392 , \19393 , \19394 , \19395 , \19396 , \19397 ,
         \19398 , \19399 , \19400 , \19401 , \19402 , \19403 , \19404 , \19405 , \19406 , \19407 ,
         \19408 , \19409 , \19410 , \19411 , \19412 , \19413 , \19414 , \19415 , \19416 , \19417 ,
         \19418 , \19419 , \19420 , \19421 , \19422 , \19423 , \19424 , \19425 , \19426 , \19427 ,
         \19428 , \19429 , \19430 , \19431 , \19432 , \19433 , \19434 , \19435 , \19436 , \19437 ,
         \19438 , \19439 , \19440 , \19441 , \19442 , \19443 , \19444 , \19445 , \19446 , \19447 ,
         \19448 , \19449 , \19450 , \19451 , \19452 , \19453 , \19454 , \19455 , \19456 , \19457 ,
         \19458 , \19459 , \19460 , \19461 , \19462 , \19463 , \19464 , \19465 , \19466 , \19467 ,
         \19468 , \19469 , \19470 , \19471 , \19472 , \19473 , \19474 , \19475 , \19476 , \19477 ,
         \19478 , \19479 , \19480 , \19481 , \19482 , \19483 , \19484 , \19485 , \19486 , \19487 ,
         \19488 , \19489 , \19490 , \19491 , \19492 , \19493 , \19494 , \19495 , \19496 , \19497 ,
         \19498 , \19499 , \19500 , \19501 , \19502 , \19503 , \19504 , \19505 , \19506 , \19507 ,
         \19508 , \19509 , \19510 , \19511 , \19512 , \19513 , \19514 , \19515 , \19516 , \19517 ,
         \19518 , \19519 , \19520 , \19521 , \19522 , \19523 , \19524 , \19525 , \19526 , \19527 ,
         \19528 , \19529 , \19530 , \19531 , \19532 , \19533 , \19534 , \19535 , \19536 , \19537 ,
         \19538 , \19539 , \19540 , \19541 , \19542 , \19543 , \19544 , \19545 , \19546 , \19547 ,
         \19548 , \19549 , \19550 , \19551 , \19552 , \19553 , \19554 , \19555 , \19556 , \19557 ,
         \19558 , \19559 , \19560 , \19561 , \19562 , \19563 , \19564 , \19565 , \19566 , \19567 ,
         \19568 , \19569 , \19570 , \19571 , \19572 , \19573 , \19574 , \19575 , \19576 , \19577 ,
         \19578 , \19579 , \19580 , \19581 , \19582 , \19583 , \19584 , \19585 , \19586 , \19587 ,
         \19588 , \19589 , \19590 , \19591 , \19592 , \19593 , \19594 , \19595 , \19596 , \19597 ,
         \19598 , \19599 , \19600 , \19601 , \19602 , \19603 , \19604 , \19605 , \19606 , \19607 ,
         \19608 , \19609 , \19610 , \19611 , \19612 , \19613 , \19614 , \19615 , \19616 , \19617 ,
         \19618 , \19619 , \19620 , \19621 , \19622 , \19623 , \19624 , \19625 , \19626 , \19627 ,
         \19628 , \19629 , \19630 , \19631 , \19632 , \19633 , \19634 , \19635 , \19636 , \19637 ,
         \19638 , \19639 , \19640 , \19641 , \19642 , \19643 , \19644 , \19645 , \19646 , \19647 ,
         \19648 , \19649 , \19650 , \19651 , \19652 , \19653 , \19654 , \19655 , \19656 , \19657 ,
         \19658 , \19659 , \19660 , \19661 , \19662 , \19663 , \19664 , \19665 , \19666 , \19667 ,
         \19668 , \19669 , \19670 , \19671 , \19672 , \19673 , \19674 , \19675 , \19676 , \19677 ,
         \19678 , \19679 , \19680 , \19681 , \19682 , \19683 , \19684 , \19685 , \19686 , \19687 ,
         \19688 , \19689 , \19690 , \19691 , \19692 , \19693 , \19694 , \19695 , \19696 , \19697 ,
         \19698 , \19699 , \19700 , \19701 , \19702 , \19703 , \19704 , \19705 , \19706 , \19707 ,
         \19708 , \19709 , \19710 , \19711 , \19712 , \19713 , \19714 , \19715 , \19716 , \19717 ,
         \19718 , \19719 , \19720 , \19721 , \19722 , \19723 , \19724 , \19725 , \19726 , \19727 ,
         \19728 , \19729 , \19730 , \19731 , \19732 , \19733 , \19734 , \19735 , \19736 , \19737 ,
         \19738 , \19739 , \19740 , \19741 , \19742 , \19743 , \19744 , \19745 , \19746 , \19747 ,
         \19748 , \19749 , \19750 , \19751 , \19752 , \19753 , \19754 , \19755 , \19756 , \19757 ,
         \19758 , \19759 , \19760 , \19761 , \19762 , \19763 , \19764 , \19765 , \19766 , \19767 ,
         \19768 , \19769 , \19770 , \19771 , \19772 , \19773 , \19774 , \19775 , \19776 , \19777 ,
         \19778 , \19779 , \19780 , \19781 , \19782 , \19783 , \19784 , \19785 , \19786 , \19787 ,
         \19788 , \19789 , \19790 , \19791 , \19792 , \19793 , \19794 , \19795 , \19796 , \19797 ,
         \19798 , \19799 , \19800 , \19801 , \19802 , \19803 , \19804 , \19805 , \19806 , \19807 ,
         \19808 , \19809 , \19810 , \19811 , \19812 , \19813 , \19814 , \19815 , \19816 , \19817 ,
         \19818 , \19819 , \19820 , \19821 , \19822 , \19823 , \19824 , \19825 , \19826 , \19827 ,
         \19828 , \19829 , \19830 , \19831 , \19832 , \19833 , \19834 , \19835 , \19836 , \19837 ,
         \19838 , \19839 , \19840 , \19841 , \19842 , \19843 , \19844 , \19845 , \19846 , \19847 ,
         \19848 , \19849 , \19850 , \19851 , \19852 , \19853 , \19854 , \19855 , \19856 , \19857 ,
         \19858 , \19859 , \19860 , \19861 , \19862 , \19863 , \19864 , \19865 , \19866 , \19867 ,
         \19868 , \19869 , \19870 , \19871 , \19872 , \19873 , \19874 , \19875 , \19876 , \19877 ,
         \19878 , \19879 , \19880 , \19881 , \19882 , \19883 , \19884 , \19885 , \19886 , \19887 ,
         \19888 , \19889 , \19890 , \19891 , \19892 , \19893 , \19894 , \19895 , \19896 , \19897 ,
         \19898 , \19899 , \19900 , \19901 , \19902 , \19903 , \19904 , \19905 , \19906 , \19907 ,
         \19908 , \19909 , \19910 , \19911 , \19912 , \19913 , \19914 , \19915 , \19916 , \19917 ,
         \19918 , \19919 , \19920 , \19921 , \19922 , \19923 , \19924 , \19925 , \19926 , \19927 ,
         \19928 , \19929 , \19930 , \19931 , \19932 , \19933 , \19934 , \19935 , \19936 , \19937 ,
         \19938 , \19939 , \19940 , \19941 , \19942 , \19943 , \19944 , \19945 , \19946 , \19947 ,
         \19948 , \19949 , \19950 , \19951 , \19952 , \19953 , \19954 , \19955 , \19956 , \19957 ,
         \19958 , \19959 , \19960 , \19961 , \19962 , \19963 , \19964 , \19965 , \19966 , \19967 ,
         \19968 , \19969 , \19970 , \19971 , \19972 , \19973 , \19974 , \19975 , \19976 , \19977 ,
         \19978 , \19979 , \19980 , \19981 , \19982 , \19983 , \19984 , \19985 , \19986 , \19987 ,
         \19988 , \19989 , \19990 , \19991 , \19992 , \19993 , \19994 , \19995 , \19996 , \19997 ,
         \19998 , \19999 , \20000 , \20001 , \20002 , \20003 , \20004 , \20005 , \20006 , \20007 ,
         \20008 , \20009 , \20010 , \20011 , \20012 , \20013 , \20014 , \20015 , \20016 , \20017 ,
         \20018 , \20019 , \20020 , \20021 , \20022 , \20023 , \20024 , \20025 , \20026 , \20027 ,
         \20028 , \20029 , \20030 , \20031 , \20032 , \20033 , \20034 , \20035 , \20036 , \20037 ,
         \20038 , \20039 , \20040 , \20041 , \20042 , \20043 , \20044 , \20045 , \20046 , \20047 ,
         \20048 , \20049 , \20050 , \20051 , \20052 , \20053 , \20054 , \20055 , \20056 , \20057 ,
         \20058 , \20059 , \20060 , \20061 , \20062 , \20063 , \20064 , \20065 , \20066 , \20067 ,
         \20068 , \20069 , \20070 , \20071 , \20072 , \20073 , \20074 , \20075 , \20076 , \20077 ,
         \20078 , \20079 , \20080 , \20081 , \20082 , \20083 , \20084 , \20085 , \20086 , \20087 ,
         \20088 , \20089 , \20090 , \20091 , \20092 , \20093 , \20094 , \20095 , \20096 , \20097 ,
         \20098 , \20099 , \20100 , \20101 , \20102 , \20103 , \20104 , \20105 , \20106 , \20107 ,
         \20108 , \20109 , \20110 , \20111 , \20112 , \20113 , \20114 , \20115 , \20116 , \20117 ,
         \20118 , \20119 , \20120 , \20121 , \20122 , \20123 , \20124 , \20125 , \20126 , \20127 ,
         \20128 , \20129 , \20130 , \20131 , \20132 , \20133 , \20134 , \20135 , \20136 , \20137 ,
         \20138 , \20139 , \20140 , \20141 , \20142 , \20143 , \20144 , \20145 , \20146 , \20147 ,
         \20148 , \20149 , \20150 , \20151 , \20152 , \20153 , \20154 , \20155 , \20156 , \20157 ,
         \20158 , \20159 , \20160 , \20161 , \20162 , \20163 , \20164 , \20165 , \20166 , \20167 ,
         \20168 , \20169 , \20170 , \20171 , \20172 , \20173 , \20174 , \20175 , \20176 , \20177 ,
         \20178 , \20179 , \20180 , \20181 , \20182 , \20183 , \20184 , \20185 , \20186 , \20187 ,
         \20188 , \20189 , \20190 , \20191 , \20192 , \20193 , \20194 , \20195 , \20196 , \20197 ,
         \20198 , \20199 , \20200 , \20201 , \20202 , \20203 , \20204 , \20205 , \20206 , \20207 ,
         \20208 , \20209 , \20210 , \20211 , \20212 , \20213 , \20214 , \20215 , \20216 , \20217 ,
         \20218 , \20219 , \20220 , \20221 , \20222 , \20223 , \20224 , \20225 , \20226 , \20227 ,
         \20228 , \20229 , \20230 , \20231 , \20232 , \20233 , \20234 , \20235 , \20236 , \20237 ,
         \20238 , \20239 , \20240 , \20241 , \20242 , \20243 , \20244 , \20245 , \20246 , \20247 ,
         \20248 , \20249 , \20250 , \20251 , \20252 , \20253 , \20254 , \20255 , \20256 , \20257 ,
         \20258 , \20259 , \20260 , \20261 , \20262 , \20263 , \20264 , \20265 , \20266 , \20267 ,
         \20268 , \20269 , \20270 , \20271 , \20272 , \20273 , \20274 , \20275 , \20276 , \20277 ,
         \20278 , \20279 , \20280 , \20281 , \20282 , \20283 , \20284 , \20285 , \20286 , \20287 ,
         \20288 , \20289 , \20290 , \20291 , \20292 , \20293 , \20294 , \20295 , \20296 , \20297 ,
         \20298 , \20299 , \20300 , \20301 , \20302 , \20303 , \20304 , \20305 , \20306 , \20307 ,
         \20308 , \20309 , \20310 , \20311 , \20312 , \20313 , \20314 , \20315 , \20316 , \20317 ,
         \20318 , \20319 , \20320 , \20321 , \20322 , \20323 , \20324 , \20325 , \20326 , \20327 ,
         \20328 , \20329 , \20330 , \20331 , \20332 , \20333 , \20334 , \20335 , \20336 , \20337 ,
         \20338 , \20339 , \20340 , \20341 , \20342 , \20343 , \20344 , \20345 , \20346 , \20347 ,
         \20348 , \20349 , \20350 , \20351 , \20352 , \20353 , \20354 , \20355 , \20356 , \20357 ,
         \20358 , \20359 , \20360 , \20361 , \20362 , \20363 , \20364 , \20365 , \20366 , \20367 ,
         \20368 , \20369 , \20370 , \20371 , \20372 , \20373 , \20374 , \20375 , \20376 , \20377 ,
         \20378 , \20379 , \20380 , \20381 , \20382 , \20383 , \20384 , \20385 , \20386 , \20387 ,
         \20388 , \20389 , \20390 , \20391 , \20392 , \20393 , \20394 , \20395 , \20396 , \20397 ,
         \20398 , \20399 , \20400 , \20401 , \20402 , \20403 , \20404 , \20405 , \20406 , \20407 ,
         \20408 , \20409 , \20410 , \20411 , \20412 , \20413 , \20414 , \20415 , \20416 , \20417 ,
         \20418 , \20419 , \20420 , \20421 , \20422 , \20423 , \20424 , \20425 , \20426 , \20427 ,
         \20428 , \20429 , \20430 , \20431 , \20432 , \20433 , \20434 , \20435 , \20436 , \20437 ,
         \20438 , \20439 , \20440 , \20441 , \20442 , \20443 , \20444 , \20445 , \20446 , \20447 ,
         \20448 , \20449 , \20450 , \20451 , \20452 , \20453 , \20454 , \20455 , \20456 , \20457 ,
         \20458 , \20459 , \20460 , \20461 , \20462 , \20463 , \20464 , \20465 , \20466 , \20467 ,
         \20468 , \20469 , \20470 , \20471 , \20472 , \20473 , \20474 , \20475 , \20476 , \20477 ,
         \20478 , \20479 , \20480 , \20481 , \20482 , \20483 , \20484 , \20485 , \20486 , \20487 ,
         \20488 , \20489 , \20490 , \20491 , \20492 , \20493 , \20494 , \20495 , \20496 , \20497 ,
         \20498 , \20499 , \20500 , \20501 , \20502 , \20503 , \20504 , \20505 , \20506 , \20507 ,
         \20508 , \20509 , \20510 , \20511 , \20512 , \20513 , \20514 , \20515 , \20516 , \20517 ,
         \20518 , \20519 , \20520 , \20521 , \20522 , \20523 , \20524 , \20525 , \20526 , \20527 ,
         \20528 , \20529 , \20530 , \20531 , \20532 , \20533 , \20534 , \20535 , \20536 , \20537 ,
         \20538 , \20539 , \20540 , \20541 , \20542 , \20543 , \20544 , \20545 , \20546 , \20547 ,
         \20548 , \20549 , \20550 , \20551 , \20552 , \20553 , \20554 , \20555 , \20556 , \20557 ,
         \20558 , \20559 , \20560 , \20561 , \20562 , \20563 , \20564 , \20565 , \20566 , \20567 ,
         \20568 , \20569 , \20570 , \20571 , \20572 , \20573 , \20574 , \20575 , \20576 , \20577 ,
         \20578 , \20579 , \20580 , \20581 , \20582 , \20583 , \20584 , \20585 , \20586 , \20587 ,
         \20588 , \20589 , \20590 , \20591 , \20592 , \20593 , \20594 , \20595 , \20596 , \20597 ,
         \20598 , \20599 , \20600 , \20601 , \20602 , \20603 , \20604 , \20605 , \20606 , \20607 ,
         \20608 , \20609 , \20610 , \20611 , \20612 , \20613 , \20614 , \20615 , \20616 , \20617 ,
         \20618 , \20619 , \20620 , \20621 , \20622 , \20623 , \20624 , \20625 , \20626 , \20627 ,
         \20628 , \20629 , \20630 , \20631 , \20632 , \20633 , \20634 , \20635 , \20636 , \20637 ,
         \20638 , \20639 , \20640 , \20641 , \20642 , \20643 , \20644 , \20645 , \20646 , \20647 ,
         \20648 , \20649 , \20650 , \20651 , \20652 , \20653 , \20654 , \20655 , \20656 , \20657 ,
         \20658 , \20659 , \20660 , \20661 , \20662 , \20663 , \20664 , \20665 , \20666 , \20667 ,
         \20668 , \20669 , \20670 , \20671 , \20672 , \20673 , \20674 , \20675 , \20676 , \20677 ,
         \20678 , \20679 , \20680 , \20681 , \20682 , \20683 , \20684 , \20685 , \20686 , \20687 ,
         \20688 , \20689 , \20690 , \20691 , \20692 , \20693 , \20694 , \20695 , \20696 , \20697 ,
         \20698 , \20699 , \20700 , \20701 , \20702 , \20703 , \20704 , \20705 , \20706 , \20707 ,
         \20708 , \20709 , \20710 , \20711 , \20712 , \20713 , \20714 , \20715 , \20716 , \20717 ,
         \20718 , \20719 , \20720 , \20721 , \20722 , \20723 , \20724 , \20725 , \20726 , \20727 ,
         \20728 , \20729 , \20730 , \20731 , \20732 , \20733 , \20734 , \20735 , \20736 , \20737 ,
         \20738 , \20739 , \20740 , \20741 , \20742 , \20743 , \20744 , \20745 , \20746 , \20747 ,
         \20748 , \20749 , \20750 , \20751 , \20752 , \20753 , \20754 , \20755 , \20756 , \20757 ,
         \20758 , \20759 , \20760 , \20761 , \20762 , \20763 , \20764 , \20765 , \20766 , \20767 ,
         \20768 , \20769 , \20770 , \20771 , \20772 , \20773 , \20774 , \20775 , \20776 , \20777 ,
         \20778 , \20779 , \20780 , \20781 , \20782 , \20783 , \20784 , \20785 , \20786 , \20787 ,
         \20788 , \20789 , \20790 , \20791 , \20792 , \20793 , \20794 , \20795 , \20796 , \20797 ,
         \20798 , \20799 , \20800 , \20801 , \20802 , \20803 , \20804 , \20805 , \20806 , \20807 ,
         \20808 , \20809 , \20810 , \20811 , \20812 , \20813 , \20814 , \20815 , \20816 , \20817 ,
         \20818 , \20819 , \20820 , \20821 , \20822 , \20823 , \20824 , \20825 , \20826 , \20827 ,
         \20828 , \20829 , \20830 , \20831 , \20832 , \20833 , \20834 , \20835 , \20836 , \20837 ,
         \20838 , \20839 , \20840 , \20841 , \20842 , \20843 , \20844 , \20845 , \20846 , \20847 ,
         \20848 , \20849 , \20850 , \20851 , \20852 , \20853 , \20854 , \20855 , \20856 , \20857 ,
         \20858 , \20859 , \20860 , \20861 , \20862 , \20863 , \20864 , \20865 , \20866 , \20867 ,
         \20868 , \20869 , \20870 , \20871 , \20872 , \20873 , \20874 , \20875 , \20876 , \20877 ,
         \20878 , \20879 , \20880 , \20881 , \20882 , \20883 , \20884 , \20885 , \20886 , \20887 ,
         \20888 , \20889 , \20890 , \20891 , \20892 , \20893 , \20894 , \20895 , \20896 , \20897 ,
         \20898 , \20899 , \20900 , \20901 , \20902 , \20903 , \20904 , \20905 , \20906 , \20907 ,
         \20908 , \20909 , \20910 , \20911 , \20912 , \20913 , \20914 , \20915 , \20916 , \20917 ,
         \20918 , \20919 , \20920 , \20921 , \20922 , \20923 , \20924 , \20925 , \20926 , \20927 ,
         \20928 , \20929 , \20930 , \20931 , \20932 , \20933 , \20934 , \20935 , \20936 , \20937 ,
         \20938 , \20939 , \20940 , \20941 , \20942 , \20943 , \20944 , \20945 , \20946 , \20947 ,
         \20948 , \20949 , \20950 , \20951 , \20952 , \20953 , \20954 , \20955 , \20956 , \20957 ,
         \20958 , \20959 , \20960 , \20961 , \20962 , \20963 , \20964 , \20965 , \20966 , \20967 ,
         \20968 , \20969 , \20970 , \20971 , \20972 , \20973 , \20974 , \20975 , \20976 , \20977 ,
         \20978 , \20979 , \20980 , \20981 , \20982 , \20983 , \20984 , \20985 , \20986 , \20987 ,
         \20988 , \20989 , \20990 , \20991 , \20992 , \20993 , \20994 , \20995 , \20996 , \20997 ,
         \20998 , \20999 , \21000 , \21001 , \21002 , \21003 , \21004 , \21005 , \21006 , \21007 ,
         \21008 , \21009 , \21010 , \21011 , \21012 , \21013 , \21014 , \21015 , \21016 , \21017 ,
         \21018 , \21019 , \21020 , \21021 , \21022 , \21023 , \21024 , \21025 , \21026 , \21027 ,
         \21028 , \21029 , \21030 , \21031 , \21032 , \21033 , \21034 , \21035 , \21036 , \21037 ,
         \21038 , \21039 , \21040 , \21041 , \21042 , \21043 , \21044 , \21045 , \21046 , \21047 ,
         \21048 , \21049 , \21050 , \21051 , \21052 , \21053 , \21054 , \21055 , \21056 , \21057 ,
         \21058 , \21059 , \21060 , \21061 , \21062 , \21063 , \21064 , \21065 , \21066 , \21067 ,
         \21068 , \21069 , \21070 , \21071 , \21072 , \21073 , \21074 , \21075 , \21076 , \21077 ,
         \21078 , \21079 , \21080 , \21081 , \21082 , \21083 , \21084 , \21085 , \21086 , \21087 ,
         \21088 , \21089 , \21090 , \21091 , \21092 , \21093 , \21094 , \21095 , \21096 , \21097 ,
         \21098 , \21099 , \21100 , \21101 , \21102 , \21103 , \21104 , \21105 , \21106 , \21107 ,
         \21108 , \21109 , \21110 , \21111 , \21112 , \21113 , \21114 , \21115 , \21116 , \21117 ,
         \21118 , \21119 , \21120 , \21121 , \21122 , \21123 , \21124 , \21125 , \21126 , \21127 ,
         \21128 , \21129 , \21130 , \21131 , \21132 , \21133 , \21134 , \21135 , \21136 , \21137 ,
         \21138 , \21139 , \21140 , \21141 , \21142 , \21143 , \21144 , \21145 , \21146 , \21147 ,
         \21148 , \21149 , \21150 , \21151 , \21152 , \21153 , \21154 , \21155 , \21156 , \21157 ,
         \21158 , \21159 , \21160 , \21161 , \21162 , \21163 , \21164 , \21165 , \21166 , \21167 ,
         \21168 , \21169 , \21170 , \21171 , \21172 , \21173 , \21174 , \21175 , \21176 , \21177 ,
         \21178 , \21179 , \21180 , \21181 , \21182 , \21183 , \21184 , \21185 , \21186 , \21187 ,
         \21188 , \21189 , \21190 , \21191 , \21192 , \21193 , \21194 , \21195 , \21196 , \21197 ,
         \21198 , \21199 , \21200 , \21201 , \21202 , \21203 , \21204 , \21205 , \21206 , \21207 ,
         \21208 , \21209 , \21210 , \21211 , \21212 , \21213 , \21214 , \21215 , \21216 , \21217 ,
         \21218 , \21219 , \21220 , \21221 , \21222 , \21223 , \21224 , \21225 , \21226 , \21227 ,
         \21228 , \21229 , \21230 , \21231 , \21232 , \21233 , \21234 , \21235 , \21236 , \21237 ,
         \21238 , \21239 , \21240 , \21241 , \21242 , \21243 , \21244 , \21245 , \21246 , \21247 ,
         \21248 , \21249 , \21250 , \21251 , \21252 , \21253 , \21254 , \21255 , \21256 , \21257 ,
         \21258 , \21259 , \21260 , \21261 , \21262 , \21263 , \21264 , \21265 , \21266 , \21267 ,
         \21268 , \21269 , \21270 , \21271 , \21272 , \21273 , \21274 , \21275 , \21276 , \21277 ,
         \21278 , \21279 , \21280 , \21281 , \21282 , \21283 , \21284 , \21285 , \21286 , \21287 ,
         \21288 , \21289 , \21290 , \21291 , \21292 , \21293 , \21294 , \21295 , \21296 , \21297 ,
         \21298 , \21299 , \21300 , \21301 , \21302 , \21303 , \21304 , \21305 , \21306 , \21307 ,
         \21308 , \21309 , \21310 , \21311 , \21312 , \21313 , \21314 , \21315 , \21316 , \21317 ,
         \21318 , \21319 , \21320 , \21321 , \21322 , \21323 , \21324 , \21325 , \21326 , \21327 ,
         \21328 , \21329 , \21330 , \21331 , \21332 , \21333 , \21334 , \21335 , \21336 , \21337 ,
         \21338 , \21339 , \21340 , \21341 , \21342 , \21343 , \21344 , \21345 , \21346 , \21347 ,
         \21348 , \21349 , \21350 , \21351 , \21352 , \21353 , \21354 , \21355 , \21356 , \21357 ,
         \21358 , \21359 , \21360 , \21361 , \21362 , \21363 , \21364 , \21365 , \21366 , \21367 ,
         \21368 , \21369 , \21370 , \21371 , \21372 , \21373 , \21374 , \21375 , \21376 , \21377 ,
         \21378 , \21379 , \21380 , \21381 , \21382 , \21383 , \21384 , \21385 , \21386 , \21387 ,
         \21388 , \21389 , \21390 , \21391 , \21392 , \21393 , \21394 , \21395 , \21396 , \21397 ,
         \21398 , \21399 , \21400 , \21401 , \21402 , \21403 , \21404 , \21405 , \21406 , \21407 ,
         \21408 , \21409 , \21410 , \21411 , \21412 , \21413 , \21414 , \21415 , \21416 , \21417 ,
         \21418 , \21419 , \21420 , \21421 , \21422 , \21423 , \21424 , \21425 , \21426 , \21427 ,
         \21428 , \21429 , \21430 , \21431 , \21432 , \21433 , \21434 , \21435 , \21436 , \21437 ,
         \21438 , \21439 , \21440 , \21441 , \21442 , \21443 , \21444 , \21445 , \21446 , \21447 ,
         \21448 , \21449 , \21450 , \21451 , \21452 , \21453 , \21454 , \21455 , \21456 , \21457 ,
         \21458 , \21459 , \21460 , \21461 , \21462 , \21463 , \21464 , \21465 , \21466 , \21467 ,
         \21468 , \21469 , \21470 , \21471 , \21472 , \21473 , \21474 , \21475 , \21476 , \21477 ,
         \21478 , \21479 , \21480 , \21481 , \21482 , \21483 , \21484 , \21485 , \21486 , \21487 ,
         \21488 , \21489 , \21490 , \21491 , \21492 , \21493 , \21494 , \21495 , \21496 , \21497 ,
         \21498 , \21499 , \21500 , \21501 , \21502 , \21503 , \21504 , \21505 , \21506 , \21507 ,
         \21508 , \21509 , \21510 , \21511 , \21512 , \21513 , \21514 , \21515 , \21516 , \21517 ,
         \21518 , \21519 , \21520 , \21521 , \21522 , \21523 , \21524 , \21525 , \21526 , \21527 ,
         \21528 , \21529 , \21530 , \21531 , \21532 , \21533 , \21534 , \21535 , \21536 , \21537 ,
         \21538 , \21539 , \21540 , \21541 , \21542 , \21543 , \21544 , \21545 , \21546 , \21547 ,
         \21548 , \21549 , \21550 , \21551 , \21552 , \21553 , \21554 , \21555 , \21556 , \21557 ,
         \21558 , \21559 , \21560 , \21561 , \21562 , \21563 , \21564 , \21565 , \21566 , \21567 ,
         \21568 , \21569 , \21570 , \21571 , \21572 , \21573 , \21574 , \21575 , \21576 , \21577 ,
         \21578 , \21579 , \21580 , \21581 , \21582 , \21583 , \21584 , \21585 , \21586 , \21587 ,
         \21588 , \21589 , \21590 , \21591 , \21592 , \21593 , \21594 , \21595 , \21596 , \21597 ,
         \21598 , \21599 , \21600 , \21601 , \21602 , \21603 , \21604 , \21605 , \21606 , \21607 ,
         \21608 , \21609 , \21610 , \21611 , \21612 , \21613 , \21614 , \21615 , \21616 , \21617 ,
         \21618 , \21619 , \21620 , \21621 , \21622 , \21623 , \21624 , \21625 , \21626 , \21627 ,
         \21628 , \21629 , \21630 , \21631 , \21632 , \21633 , \21634 , \21635 , \21636 , \21637 ,
         \21638 , \21639 , \21640 , \21641 , \21642 , \21643 , \21644 , \21645 , \21646 , \21647 ,
         \21648 , \21649 , \21650 , \21651 , \21652 , \21653 , \21654 , \21655 , \21656 , \21657 ,
         \21658 , \21659 , \21660 , \21661 , \21662 , \21663 , \21664 , \21665 , \21666 , \21667 ,
         \21668 , \21669 , \21670 , \21671 , \21672 , \21673 , \21674 , \21675 , \21676 , \21677 ,
         \21678 , \21679 , \21680 , \21681 , \21682 , \21683 , \21684 , \21685 , \21686 , \21687 ,
         \21688 , \21689 , \21690 , \21691 , \21692 , \21693 , \21694 , \21695 , \21696 , \21697 ,
         \21698 , \21699 , \21700 , \21701 , \21702 , \21703 , \21704 , \21705 , \21706 , \21707 ,
         \21708 , \21709 , \21710 , \21711 , \21712 , \21713 , \21714 , \21715 , \21716 , \21717 ,
         \21718 , \21719 , \21720 , \21721 , \21722 , \21723 , \21724 , \21725 , \21726 , \21727 ,
         \21728 , \21729 , \21730 , \21731 , \21732 , \21733 , \21734 , \21735 , \21736 , \21737 ,
         \21738 , \21739 , \21740 , \21741 , \21742 , \21743 , \21744 , \21745 , \21746 , \21747 ,
         \21748 , \21749 , \21750 , \21751 , \21752 , \21753 , \21754 , \21755 , \21756 , \21757 ,
         \21758 , \21759 , \21760 , \21761 , \21762 , \21763 , \21764 , \21765 , \21766 , \21767 ,
         \21768 , \21769 , \21770 , \21771 , \21772 , \21773 , \21774 , \21775 , \21776 , \21777 ,
         \21778 , \21779 , \21780 , \21781 , \21782 , \21783 , \21784 , \21785 , \21786 , \21787 ,
         \21788 , \21789 , \21790 , \21791 , \21792 , \21793 , \21794 , \21795 , \21796 , \21797 ,
         \21798 , \21799 , \21800 , \21801 , \21802 , \21803 , \21804 , \21805 , \21806 , \21807 ,
         \21808 , \21809 , \21810 , \21811 , \21812 , \21813 , \21814 , \21815 , \21816 , \21817 ,
         \21818 , \21819 , \21820 , \21821 , \21822 , \21823 , \21824 , \21825 , \21826 , \21827 ,
         \21828 , \21829 , \21830 , \21831 , \21832 , \21833 , \21834 , \21835 , \21836 , \21837 ,
         \21838 , \21839 , \21840 , \21841 , \21842 , \21843 , \21844 , \21845 , \21846 , \21847 ,
         \21848 , \21849 , \21850 , \21851 , \21852 , \21853 , \21854 , \21855 , \21856 , \21857 ,
         \21858 , \21859 , \21860 , \21861 , \21862 , \21863 , \21864 , \21865 , \21866 , \21867 ,
         \21868 , \21869 , \21870 , \21871 , \21872 , \21873 , \21874 , \21875 , \21876 , \21877 ,
         \21878 , \21879 , \21880 , \21881 , \21882 , \21883 , \21884 , \21885 , \21886 , \21887 ,
         \21888 , \21889 , \21890 , \21891 , \21892 , \21893 , \21894 , \21895 , \21896 , \21897 ,
         \21898 , \21899 , \21900 , \21901 , \21902 , \21903 , \21904 , \21905 , \21906 , \21907 ,
         \21908 , \21909 , \21910 , \21911 , \21912 , \21913 , \21914 , \21915 , \21916 , \21917 ,
         \21918 , \21919 , \21920 , \21921 , \21922 , \21923 , \21924 , \21925 , \21926 , \21927 ,
         \21928 , \21929 , \21930 , \21931 , \21932 , \21933 , \21934 , \21935 , \21936 , \21937 ,
         \21938 , \21939 , \21940 , \21941 , \21942 , \21943 , \21944 , \21945 , \21946 , \21947 ,
         \21948 , \21949 , \21950 , \21951 , \21952 , \21953 , \21954 , \21955 , \21956 , \21957 ,
         \21958 , \21959 , \21960 , \21961 , \21962 , \21963 , \21964 , \21965 , \21966 , \21967 ,
         \21968 , \21969 , \21970 , \21971 , \21972 , \21973 , \21974 , \21975 , \21976 , \21977 ,
         \21978 , \21979 , \21980 , \21981 , \21982 , \21983 , \21984 , \21985 , \21986 , \21987 ,
         \21988 , \21989 , \21990 , \21991 , \21992 , \21993 , \21994 , \21995 , \21996 , \21997 ,
         \21998 , \21999 , \22000 , \22001 , \22002 , \22003 , \22004 , \22005 , \22006 , \22007 ,
         \22008 , \22009 , \22010 , \22011 , \22012 , \22013 , \22014 , \22015 , \22016 , \22017 ,
         \22018 , \22019 , \22020 , \22021 , \22022 , \22023 , \22024 , \22025 , \22026 , \22027 ,
         \22028 , \22029 , \22030 , \22031 , \22032 , \22033 , \22034 , \22035 , \22036 , \22037 ,
         \22038 , \22039 , \22040 , \22041 , \22042 , \22043 , \22044 , \22045 , \22046 , \22047 ,
         \22048 , \22049 , \22050 , \22051 , \22052 , \22053 , \22054 , \22055 , \22056 , \22057 ,
         \22058 , \22059 , \22060 , \22061 , \22062 , \22063 , \22064 , \22065 ;
buf \U$labajz2280 ( R_267_b0ecd58, \10828 );
buf \U$labajz2281 ( R_268_b0ece00, \10846 );
buf \U$labajz2282 ( R_269_b0ecea8, \10895 );
buf \U$labajz2283 ( R_26a_b0ecf50, \10928 );
buf \U$labajz2284 ( R_26b_b0ecff8, \10951 );
buf \U$labajz2285 ( R_26c_b0ed0a0, \10959 );
buf \U$labajz2286 ( R_26d_b0ed148, \10993 );
buf \U$labajz2287 ( R_26e_b0ed1f0, \11010 );
buf \U$labajz2288 ( R_26f_b0ed298, \11035 );
buf \U$labajz2289 ( R_270_b0ed340, \11043 );
buf \U$labajz2290 ( R_271_b0ed3e8, \11100 );
buf \U$labajz2291 ( R_272_b0ed490, \11113 );
buf \U$labajz2292 ( R_273_b0ed538, \11129 );
buf \U$labajz2293 ( R_274_b0ed5e0, \11138 );
buf \U$labajz2294 ( R_275_b0ed688, \11171 );
buf \U$labajz2295 ( R_276_b0ed730, \11189 );
buf \U$labajz2296 ( R_277_b0ed7d8, \11208 );
buf \U$labajz2297 ( R_278_b0ed880, \11230 );
buf \U$labajz2298 ( R_279_b0ed928, \11254 );
buf \U$labajz2299 ( R_27a_b0ed9d0, \11266 );
buf \U$labajz2300 ( R_27b_b0eda78, \11296 );
buf \U$labajz2301 ( R_27c_b0edb20, \11308 );
buf \U$labajz2302 ( R_27d_b0edbc8, \11320 );
buf \U$labajz2303 ( R_27e_b0edc70, \11327 );
buf \U$labajz2304 ( R_27f_b0edd18, \11334 );
buf \U$labajz2305 ( R_280_b0eddc0, \11351 );
buf \U$labajz2306 ( R_281_b0ede68, \11363 );
buf \U$labajz2307 ( R_282_b0edf10, \21478 );
buf \U$labajz2308 ( R_283_b0edfb8, \21502 );
buf \U$labajz2309 ( R_284_b0ee060, \21570 );
buf \U$labajz2310 ( R_285_b0ee108, \21602 );
buf \U$labajz2311 ( R_286_b0ee1b0, \21629 );
buf \U$labajz2312 ( R_287_b0ee258, \21646 );
buf \U$labajz2313 ( R_288_b0ee300, \21683 );
buf \U$labajz2314 ( R_289_b0ee3a8, \21697 );
buf \U$labajz2315 ( R_28a_b0ee450, \21720 );
buf \U$labajz2316 ( R_28b_b0ee4f8, \21730 );
buf \U$labajz2317 ( R_28c_b0ee5a0, \21774 );
buf \U$labajz2318 ( R_28d_b0ee648, \21788 );
buf \U$labajz2319 ( R_28e_b0ee6f0, \21815 );
buf \U$labajz2320 ( R_28f_b0ee798, \21831 );
buf \U$labajz2321 ( R_290_b0ee840, \21867 );
buf \U$labajz2322 ( R_291_b0ee8e8, \21876 );
buf \U$labajz2323 ( R_292_b0ee990, \21896 );
buf \U$labajz2324 ( R_293_b0eea38, \21912 );
buf \U$labajz2325 ( R_294_b0eeae0, \21958 );
buf \U$labajz2326 ( R_295_b0eeb88, \21978 );
buf \U$labajz2327 ( R_296_b0eec30, \22001 );
buf \U$labajz2328 ( R_297_b0eecd8, \22015 );
buf \U$labajz2329 ( R_298_b0eed80, \22029 );
buf \U$labajz2330 ( R_299_b0eee28, \22036 );
buf \U$labajz2331 ( R_29a_b0eeed0, \22043 );
buf \U$labajz2332 ( R_29b_b0eef78, \22053 );
buf \U$labajz2333 ( R_29c_b0ef020, \22065 );
not \U$1 ( \671 , RIaa97c98_14);
not \U$2 ( \672 , \671 );
nor \U$3 ( \673 , RIaa9e7f0_243, RIaa9e868_244);
nor \U$4 ( \674 , RIaa9e778_242, RIaa9e9d0_247);
not \U$5 ( \675 , RIaa97d88_16);
nand \U$6 ( \676 , \673 , \674 , \675 );
not \U$7 ( \677 , \676 );
not \U$8 ( \678 , \677 );
not \U$9 ( \679 , \678 );
and \U$10 ( \680 , RIaa97d10_15, RIaa97e00_17);
nand \U$11 ( \681 , RIaa97c20_13, RIaa97c98_14);
nor \U$12 ( \682 , RIaa9e688_240, RIaa9e700_241);
nor \U$13 ( \683 , RIaa9e8e0_245, RIaa9e958_246);
and \U$14 ( \684 , \680 , \681 , \682 , \683 );
nand \U$15 ( \685 , \679 , \684 );
not \U$16 ( \686 , \685 );
not \U$17 ( \687 , \686 );
or \U$18 ( \688 , \672 , \687 );
not \U$19 ( \689 , \678 );
not \U$20 ( \690 , \689 );
not \U$21 ( \691 , \684 );
or \U$22 ( \692 , \690 , \691 );
nand \U$23 ( \693 , \692 , RIaa97c98_14);
nand \U$24 ( \694 , \688 , \693 );
buf \U$25 ( \695 , \694 );
not \U$26 ( \696 , \695 );
not \U$27 ( \697 , \696 );
nor \U$28 ( \698 , RIaa9e8e0_245, RIaa9e958_246);
nor \U$29 ( \699 , RIaa9e688_240, RIaa9e700_241);
and \U$30 ( \700 , \698 , \699 , RIaa97e00_17);
nand \U$31 ( \701 , RIaa97d10_15, RIaa97c20_13, RIaa97c98_14);
and \U$32 ( \702 , \677 , \700 , \701 );
not \U$33 ( \703 , RIaa97d10_15);
and \U$34 ( \704 , \702 , \703 );
not \U$35 ( \705 , \702 );
and \U$36 ( \706 , \705 , RIaa97d10_15);
nor \U$37 ( \707 , \704 , \706 );
buf \U$38 ( \708 , \707 );
not \U$39 ( \709 , \708 );
not \U$40 ( \710 , RIaa97e00_17);
not \U$41 ( \711 , \710 );
not \U$42 ( \712 , \678 );
and \U$43 ( \713 , \682 , \683 );
nand \U$44 ( \714 , \712 , \713 );
not \U$45 ( \715 , \714 );
or \U$46 ( \716 , \711 , \715 );
not \U$47 ( \717 , \702 );
nand \U$48 ( \718 , \716 , \717 );
buf \U$49 ( \719 , \718 );
not \U$50 ( \720 , \719 );
not \U$51 ( \721 , RIaa97c98_14);
not \U$52 ( \722 , \686 );
or \U$53 ( \723 , \721 , \722 );
not \U$54 ( \724 , RIaa97c20_13);
nand \U$55 ( \725 , \723 , \724 );
buf \U$56 ( \726 , \725 );
nand \U$57 ( \727 , \697 , \709 , \720 , \726 );
not \U$58 ( \728 , \727 );
nand \U$59 ( \729 , \728 , RIaa9cf90_191);
not \U$60 ( \730 , \696 );
not \U$61 ( \731 , \726 );
not \U$62 ( \732 , \719 );
not \U$63 ( \733 , \732 );
not \U$64 ( \734 , \707 );
not \U$65 ( \735 , \734 );
and \U$66 ( \736 , \730 , \731 , \733 , \735 );
nand \U$67 ( \737 , \736 , RIaa9d170_195);
nand \U$68 ( \738 , RIaa97d88_16, RIaa9cea0_189);
nand \U$69 ( \739 , \729 , \737 , \738 );
not \U$70 ( \740 , RIaa9d1e8_196);
not \U$71 ( \741 , \734 );
buf \U$72 ( \742 , \694 );
nand \U$73 ( \743 , \741 , \742 , \731 , \720 );
not \U$74 ( \744 , \743 );
not \U$75 ( \745 , \744 );
or \U$76 ( \746 , \740 , \745 );
nor \U$77 ( \747 , \695 , RIaa97d88_16);
buf \U$78 ( \748 , \725 );
not \U$79 ( \749 , \748 );
not \U$80 ( \750 , \734 );
buf \U$81 ( \751 , \718 );
nand \U$82 ( \752 , \747 , \749 , \750 , \751 );
not \U$83 ( \753 , \752 );
nand \U$84 ( \754 , \753 , RIaa9d080_193);
nand \U$85 ( \755 , \746 , \754 );
nor \U$86 ( \756 , \739 , \755 );
not \U$87 ( \757 , RIaa9d0f8_194);
not \U$88 ( \758 , \695 );
not \U$89 ( \759 , \758 );
not \U$90 ( \760 , \726 );
not \U$91 ( \761 , \760 );
buf \U$92 ( \762 , \708 );
not \U$93 ( \763 , \751 );
nand \U$94 ( \764 , \759 , \761 , \762 , \763 );
not \U$95 ( \765 , \764 );
not \U$96 ( \766 , \765 );
or \U$97 ( \767 , \757 , \766 );
buf \U$98 ( \768 , \707 );
not \U$99 ( \769 , \768 );
not \U$100 ( \770 , \769 );
not \U$101 ( \771 , \742 );
not \U$102 ( \772 , \719 );
not \U$103 ( \773 , \772 );
nand \U$104 ( \774 , \770 , \726 , \771 , \773 );
not \U$105 ( \775 , \774 );
nand \U$106 ( \776 , \775 , RIaa9d5a8_204);
nand \U$107 ( \777 , \767 , \776 );
not \U$108 ( \778 , RIaa9d620_205);
not \U$109 ( \779 , \768 );
not \U$110 ( \780 , \779 );
not \U$111 ( \781 , \748 );
not \U$112 ( \782 , \781 );
not \U$113 ( \783 , \742 );
nand \U$114 ( \784 , \780 , \782 , \783 , \763 );
not \U$115 ( \785 , \784 );
not \U$116 ( \786 , \785 );
or \U$117 ( \787 , \778 , \786 );
and \U$118 ( \788 , \726 , \742 , \768 , \751 );
nand \U$119 ( \789 , \788 , RIaa9d2d8_198);
nand \U$120 ( \790 , \787 , \789 );
nor \U$121 ( \791 , \777 , \790 );
not \U$122 ( \792 , RIaa9d008_192);
not \U$123 ( \793 , \742 );
not \U$124 ( \794 , \751 );
nand \U$125 ( \795 , \793 , \741 , \794 , \781 );
not \U$126 ( \796 , \795 );
not \U$127 ( \797 , \796 );
or \U$128 ( \798 , \792 , \797 );
not \U$129 ( \799 , \707 );
nand \U$130 ( \800 , \799 , \718 );
not \U$131 ( \801 , \800 );
not \U$132 ( \802 , \695 );
and \U$133 ( \803 , \801 , \802 , \748 );
nand \U$134 ( \804 , \803 , RIaa9d3c8_200);
nand \U$135 ( \805 , \798 , \804 );
not \U$136 ( \806 , RIaa9d4b8_202);
not \U$137 ( \807 , \751 );
and \U$138 ( \808 , \779 , \731 , \771 , \807 );
not \U$139 ( \809 , \808 );
or \U$140 ( \810 , \806 , \809 );
and \U$141 ( \811 , \801 , \742 , \749 );
nand \U$142 ( \812 , \811 , RIaa9d260_197);
nand \U$143 ( \813 , \810 , \812 );
nor \U$144 ( \814 , \805 , \813 );
not \U$145 ( \815 , RIaa9d350_199);
not \U$146 ( \816 , \719 );
and \U$147 ( \817 , \771 , \816 , \734 , \748 );
not \U$148 ( \818 , \817 );
or \U$149 ( \819 , \815 , \818 );
not \U$150 ( \820 , \800 );
not \U$151 ( \821 , \820 );
nand \U$152 ( \822 , \748 , \695 );
nor \U$153 ( \823 , \821 , \822 );
nand \U$154 ( \824 , \823 , RIaa9cf18_190);
nand \U$155 ( \825 , \819 , \824 );
not \U$156 ( \826 , RIaa9d530_203);
and \U$157 ( \827 , \696 , \820 , \760 );
not \U$158 ( \828 , \827 );
or \U$159 ( \829 , \826 , \828 );
not \U$160 ( \830 , \726 );
and \U$161 ( \831 , \695 , \830 , \769 , \807 );
nand \U$162 ( \832 , \831 , RIaa9d440_201);
nand \U$163 ( \833 , \829 , \832 );
nor \U$164 ( \834 , \825 , \833 );
nand \U$165 ( \835 , \756 , \791 , \814 , \834 );
nand \U$166 ( \836 , RIaa97860_5, RIaa976f8_2, RIaa97770_3, RIaa977e8_4);
not \U$167 ( \837 , RIaa97860_5);
nand \U$168 ( \838 , RIaa97770_3, RIaa977e8_4);
not \U$169 ( \839 , \838 );
nand \U$170 ( \840 , \839 , RIaa976f8_2);
nand \U$171 ( \841 , \837 , \840 );
and \U$172 ( \842 , \836 , \841 );
not \U$173 ( \843 , \842 );
nand \U$174 ( \844 , \835 , \843 );
buf \U$175 ( \845 , \844 );
not \U$176 ( \846 , \845 );
not \U$177 ( \847 , RIaa97770_3);
not \U$178 ( \848 , \847 );
not \U$179 ( \849 , RIaa977e8_4);
not \U$180 ( \850 , \849 );
or \U$181 ( \851 , \848 , \850 );
nand \U$182 ( \852 , \851 , \838 );
not \U$183 ( \853 , \852 );
not \U$184 ( \854 , \853 );
nand \U$185 ( \855 , \728 , RIaa9ba00_145);
nand \U$186 ( \856 , \720 , \742 , \748 , \750 );
not \U$187 ( \857 , \856 );
nand \U$188 ( \858 , \857 , RIaa9b640_137);
nand \U$189 ( \859 , RIaa97d88_16, RIaa9b910_143);
nand \U$190 ( \860 , \855 , \858 , \859 );
not \U$191 ( \861 , RIaa9bd48_152);
not \U$192 ( \862 , \732 );
nand \U$193 ( \863 , \761 , \783 , \762 , \862 );
not \U$194 ( \864 , \863 );
not \U$195 ( \865 , \864 );
or \U$196 ( \866 , \861 , \865 );
and \U$197 ( \867 , \708 , \695 , \748 , \751 );
nand \U$198 ( \868 , \867 , RIaa9ba78_146);
nand \U$199 ( \869 , \866 , \868 );
nor \U$200 ( \870 , \860 , \869 );
not \U$201 ( \871 , RIaa9bb68_148);
not \U$202 ( \872 , \800 );
and \U$203 ( \873 , \872 , \726 , \771 );
not \U$204 ( \874 , \873 );
or \U$205 ( \875 , \871 , \874 );
nand \U$206 ( \876 , \811 , RIaa9b7a8_140);
nand \U$207 ( \877 , \875 , \876 );
not \U$208 ( \878 , RIaa9bdc0_153);
not \U$209 ( \879 , \785 );
or \U$210 ( \880 , \878 , \879 );
and \U$211 ( \881 , \779 , \726 , \816 , \696 );
nand \U$212 ( \882 , \881 , RIaa9baf0_147);
nand \U$213 ( \883 , \880 , \882 );
nor \U$214 ( \884 , \877 , \883 );
not \U$215 ( \885 , RIaa9b730_139);
not \U$216 ( \886 , \744 );
or \U$217 ( \887 , \885 , \886 );
and \U$218 ( \888 , \758 , \830 , \772 , \769 );
nand \U$219 ( \889 , \888 , RIaa9bc58_150);
nand \U$220 ( \890 , \887 , \889 );
not \U$221 ( \891 , RIaa9b6b8_138);
not \U$222 ( \892 , \769 );
not \U$223 ( \893 , \748 );
not \U$224 ( \894 , \802 );
nand \U$225 ( \895 , \892 , \893 , \894 , \773 );
not \U$226 ( \896 , \895 );
not \U$227 ( \897 , \896 );
or \U$228 ( \898 , \891 , \897 );
nand \U$229 ( \899 , \753 , RIaa9b898_142);
nand \U$230 ( \900 , \898 , \899 );
nor \U$231 ( \901 , \890 , \900 );
not \U$232 ( \902 , RIaa9bcd0_151);
and \U$233 ( \903 , \872 , \758 , \830 );
not \U$234 ( \904 , \903 );
or \U$235 ( \905 , \902 , \904 );
nand \U$236 ( \906 , \823 , RIaa9b988_144);
nand \U$237 ( \907 , \905 , \906 );
not \U$238 ( \908 , RIaa9b820_141);
not \U$239 ( \909 , \796 );
or \U$240 ( \910 , \908 , \909 );
and \U$241 ( \911 , \830 , \734 , \732 , \742 );
nand \U$242 ( \912 , \911 , RIaa9bbe0_149);
nand \U$243 ( \913 , \910 , \912 );
nor \U$244 ( \914 , \907 , \913 );
nand \U$245 ( \915 , \870 , \884 , \901 , \914 );
nand \U$246 ( \916 , \854 , \915 );
nand \U$247 ( \917 , \803 , RIaa9b370_131);
nand \U$248 ( \918 , \736 , RIaa9b0a0_125);
nand \U$249 ( \919 , \903 , RIaa9b5c8_136);
nand \U$250 ( \920 , \911 , RIaa9b3e8_132);
nand \U$251 ( \921 , \917 , \918 , \919 , \920 );
nand \U$252 ( \922 , \758 , \893 , \816 , \735 );
not \U$253 ( \923 , \922 );
not \U$254 ( \924 , RIaa9ae48_120);
not \U$255 ( \925 , \924 );
and \U$256 ( \926 , \923 , \925 );
and \U$257 ( \927 , \775 , RIaa9b460_133);
nor \U$258 ( \928 , \926 , \927 );
nand \U$259 ( \929 , \735 , \742 , \893 , \720 );
not \U$260 ( \930 , \929 );
not \U$261 ( \931 , RIaa9b190_127);
not \U$262 ( \932 , \931 );
and \U$263 ( \933 , \930 , \932 );
not \U$264 ( \934 , RIaa9b118_126);
nor \U$265 ( \935 , \934 , \856 );
nor \U$266 ( \936 , \933 , \935 );
nand \U$267 ( \937 , \928 , \936 );
nor \U$268 ( \938 , \921 , \937 );
and \U$269 ( \939 , \735 , \802 , \816 , \726 );
and \U$270 ( \940 , \939 , RIaa9b4d8_134);
and \U$271 ( \941 , \788 , RIaa9b280_129);
nor \U$272 ( \942 , \940 , \941 );
and \U$273 ( \943 , \728 , RIaa9b028_124);
and \U$274 ( \944 , RIaa97d88_16, RIaa9af38_122);
nor \U$275 ( \945 , \943 , \944 );
nand \U$276 ( \946 , \881 , RIaa9b2f8_130);
nand \U$277 ( \947 , \942 , \945 , \946 );
nand \U$278 ( \948 , \753 , RIaa9aec0_121);
nand \U$279 ( \949 , \888 , RIaa9b550_135);
nand \U$280 ( \950 , \823 , RIaa9afb0_123);
nand \U$281 ( \951 , \811 , RIaa9b208_128);
nand \U$282 ( \952 , \948 , \949 , \950 , \951 );
nor \U$283 ( \953 , \947 , \952 );
nand \U$284 ( \954 , \938 , \953 );
not \U$285 ( \955 , RIaa976f8_2);
and \U$286 ( \956 , \838 , \955 );
not \U$287 ( \957 , \838 );
and \U$288 ( \958 , \957 , RIaa976f8_2);
nor \U$289 ( \959 , \956 , \958 );
not \U$290 ( \960 , \959 );
nand \U$291 ( \961 , \954 , \960 );
and \U$292 ( \962 , \916 , \961 );
not \U$293 ( \963 , \962 );
not \U$294 ( \964 , \849 );
nand \U$295 ( \965 , \736 , RIaa9c2e8_164);
nand \U$296 ( \966 , \939 , RIaa9c4c8_168);
not \U$297 ( \967 , \922 );
nand \U$298 ( \968 , \967 , RIaa9c018_158);
nand \U$299 ( \969 , \881 , RIaa9c3d8_166);
and \U$300 ( \970 , \965 , \966 , \968 , \969 );
not \U$301 ( \971 , RIaa9c450_167);
not \U$302 ( \972 , \864 );
or \U$303 ( \973 , \971 , \972 );
nand \U$304 ( \974 , \788 , RIaa9be38_154);
nand \U$305 ( \975 , \973 , \974 );
not \U$306 ( \976 , RIaa9bfa0_157);
not \U$307 ( \977 , \888 );
or \U$308 ( \978 , \976 , \977 );
nand \U$309 ( \979 , \911 , RIaa9beb0_155);
nand \U$310 ( \980 , \978 , \979 );
nor \U$311 ( \981 , \975 , \980 );
nand \U$312 ( \982 , \970 , \981 );
not \U$313 ( \983 , RIaa9c270_163);
not \U$314 ( \984 , \744 );
or \U$315 ( \985 , \983 , \984 );
nand \U$316 ( \986 , \753 , RIaa9c090_159);
nand \U$317 ( \987 , \985 , \986 );
not \U$318 ( \988 , \987 );
and \U$319 ( \989 , RIaa97d88_16, RIaa9c108_160);
not \U$320 ( \990 , \989 );
not \U$321 ( \991 , \727 );
nand \U$322 ( \992 , \991 , RIaa9c180_161);
nand \U$323 ( \993 , \903 , RIaa9bf28_156);
nand \U$324 ( \994 , \990 , \992 , \993 );
not \U$325 ( \995 , \994 );
not \U$326 ( \996 , \764 );
not \U$327 ( \997 , RIaa9c5b8_170);
not \U$328 ( \998 , \997 );
and \U$329 ( \999 , \996 , \998 );
not \U$330 ( \1000 , \822 );
and \U$331 ( \1001 , \1000 , \872 );
and \U$332 ( \1002 , \1001 , RIaa9c1f8_162);
nor \U$333 ( \1003 , \999 , \1002 );
not \U$334 ( \1004 , \803 );
not \U$335 ( \1005 , \1004 );
not \U$336 ( \1006 , RIaa9c360_165);
not \U$337 ( \1007 , \1006 );
and \U$338 ( \1008 , \1005 , \1007 );
not \U$339 ( \1009 , \811 );
not \U$340 ( \1010 , RIaa9c540_169);
nor \U$341 ( \1011 , \1009 , \1010 );
nor \U$342 ( \1012 , \1008 , \1011 );
nand \U$343 ( \1013 , \988 , \995 , \1003 , \1012 );
nor \U$344 ( \1014 , \982 , \1013 );
not \U$345 ( \1015 , \1014 );
or \U$346 ( \1016 , \964 , \1015 );
not \U$347 ( \1017 , RIaa9ce28_188);
not \U$348 ( \1018 , \1017 );
nand \U$349 ( \1019 , \888 , RIaa9c978_178);
nand \U$350 ( \1020 , \803 , RIaa9c9f0_179);
and \U$351 ( \1021 , \872 , \893 , \742 );
nand \U$352 ( \1022 , RIaa9c900_177, \1021 );
nand \U$353 ( \1023 , \911 , RIaa9cdb0_187);
nand \U$354 ( \1024 , \1019 , \1020 , \1022 , \1023 );
not \U$355 ( \1025 , \802 );
not \U$356 ( \1026 , \708 );
nand \U$357 ( \1027 , \1025 , \1026 , \726 , \794 );
not \U$358 ( \1028 , \1027 );
and \U$359 ( \1029 , \1028 , RIaa9c810_175);
and \U$360 ( \1030 , RIaa97d88_16, RIaa9c720_173);
nor \U$361 ( \1031 , \1029 , \1030 );
nand \U$362 ( \1032 , \939 , RIaa9cb58_182);
nand \U$363 ( \1033 , \903 , RIaa9cae0_181);
nand \U$364 ( \1034 , \823 , RIaa9c630_171);
nand \U$365 ( \1035 , \1031 , \1032 , \1033 , \1034 );
nor \U$366 ( \1036 , \1024 , \1035 );
nand \U$367 ( \1037 , \775 , RIaa9ca68_180);
not \U$368 ( \1038 , \929 );
nand \U$369 ( \1039 , \1038 , RIaa9cc48_184);
nand \U$370 ( \1040 , \736 , RIaa9ccc0_185);
nand \U$371 ( \1041 , \857 , RIaa9c888_176);
nand \U$372 ( \1042 , \1037 , \1039 , \1040 , \1041 );
nand \U$373 ( \1043 , \796 , RIaa9c6a8_172);
nand \U$374 ( \1044 , \753 , RIaa9c798_174);
nand \U$375 ( \1045 , \881 , RIaa9cbd0_183);
nand \U$376 ( \1046 , \788 , RIaa9cd38_186);
nand \U$377 ( \1047 , \1043 , \1044 , \1045 , \1046 );
nor \U$378 ( \1048 , \1042 , \1047 );
nand \U$379 ( \1049 , \1036 , \1048 );
not \U$380 ( \1050 , \1049 );
or \U$381 ( \1051 , \1018 , \1050 );
not \U$382 ( \1052 , \980 );
nand \U$383 ( \1053 , \995 , \1003 , \1012 , \1052 );
nor \U$384 ( \1054 , \987 , \975 );
nand \U$385 ( \1055 , \970 , \1054 );
or \U$386 ( \1056 , \1053 , \1055 );
nand \U$387 ( \1057 , \1056 , RIaa977e8_4);
nand \U$388 ( \1058 , \1051 , \1057 );
nand \U$389 ( \1059 , \1016 , \1058 );
not \U$390 ( \1060 , \1059 );
or \U$391 ( \1061 , \963 , \1060 );
not \U$392 ( \1062 , \915 );
nand \U$393 ( \1063 , \1062 , \853 );
not \U$394 ( \1064 , \1063 );
nor \U$395 ( \1065 , \954 , \960 );
not \U$396 ( \1066 , \1065 );
not \U$397 ( \1067 , \1066 );
or \U$398 ( \1068 , \1064 , \1067 );
nand \U$399 ( \1069 , \1068 , \961 );
nand \U$400 ( \1070 , \1061 , \1069 );
not \U$401 ( \1071 , \1070 );
or \U$402 ( \1072 , \846 , \1071 );
buf \U$403 ( \1073 , \835 );
nor \U$404 ( \1074 , \1073 , \843 );
not \U$405 ( \1075 , \1074 );
nand \U$406 ( \1076 , \1072 , \1075 );
not \U$407 ( \1077 , \1076 );
not \U$408 ( \1078 , RIaa9ab78_114);
not \U$409 ( \1079 , \873 );
or \U$410 ( \1080 , \1078 , \1079 );
nand \U$411 ( \1081 , \1021 , RIaa9aa10_111);
nand \U$412 ( \1082 , \1080 , \1081 );
not \U$413 ( \1083 , RIaa9ac68_116);
not \U$414 ( \1084 , \827 );
or \U$415 ( \1085 , \1083 , \1084 );
nand \U$416 ( \1086 , \1001 , RIaa9a7b8_106);
nand \U$417 ( \1087 , \1085 , \1086 );
nor \U$418 ( \1088 , \1082 , \1087 );
not \U$419 ( \1089 , RIaa9a6c8_104);
not \U$420 ( \1090 , \753 );
or \U$421 ( \1091 , \1089 , \1090 );
nand \U$422 ( \1092 , \785 , RIaa9add0_119);
nand \U$423 ( \1093 , \1091 , \1092 );
not \U$424 ( \1094 , \831 );
not \U$425 ( \1095 , RIaa9abf0_115);
or \U$426 ( \1096 , \1094 , \1095 );
not \U$427 ( \1097 , \895 );
nand \U$428 ( \1098 , \1097 , RIaa9a8a8_108);
nand \U$429 ( \1099 , \1096 , \1098 );
nor \U$430 ( \1100 , \1093 , \1099 );
not \U$431 ( \1101 , RIaa9a998_110);
not \U$432 ( \1102 , \744 );
or \U$433 ( \1103 , \1101 , \1102 );
not \U$434 ( \1104 , \764 );
nand \U$435 ( \1105 , \1104 , RIaa9a920_109);
nand \U$436 ( \1106 , \1103 , \1105 );
nand \U$437 ( \1107 , \1028 , RIaa9a830_107);
nand \U$438 ( \1108 , \775 , RIaa9ad58_118);
nand \U$439 ( \1109 , RIaa97d88_16, RIaa9a740_105);
nand \U$440 ( \1110 , \1107 , \1108 , \1109 );
nor \U$441 ( \1111 , \1106 , \1110 );
not \U$442 ( \1112 , RIaa9ab00_113);
not \U$443 ( \1113 , \817 );
or \U$444 ( \1114 , \1112 , \1113 );
nand \U$445 ( \1115 , \867 , RIaa9aa88_112);
nand \U$446 ( \1116 , \1114 , \1115 );
not \U$447 ( \1117 , RIaa9a650_103);
not \U$448 ( \1118 , \796 );
or \U$449 ( \1119 , \1117 , \1118 );
nand \U$450 ( \1120 , \808 , RIaa9ace0_117);
nand \U$451 ( \1121 , \1119 , \1120 );
nor \U$452 ( \1122 , \1116 , \1121 );
nand \U$453 ( \1123 , \1088 , \1100 , \1111 , \1122 );
buf \U$454 ( \1124 , \836 );
not \U$455 ( \1125 , \1124 );
nor \U$456 ( \1126 , \1125 , RIaa978d8_6);
not \U$457 ( \1127 , \1126 );
not \U$458 ( \1128 , \836 );
nand \U$459 ( \1129 , \1128 , RIaa978d8_6);
nand \U$460 ( \1130 , \1127 , \1129 );
nand \U$461 ( \1131 , \1123 , \1130 );
not \U$462 ( \1132 , \1131 );
not \U$463 ( \1133 , \1132 );
not \U$464 ( \1134 , \1130 );
not \U$465 ( \1135 , \1123 );
nand \U$466 ( \1136 , \1134 , \1135 );
buf \U$467 ( \1137 , \1136 );
nand \U$468 ( \1138 , \1133 , \1137 );
not \U$469 ( \1139 , \1138 );
and \U$470 ( \1140 , \1077 , \1139 );
and \U$471 ( \1141 , \1076 , \1138 );
nor \U$472 ( \1142 , \1140 , \1141 );
not \U$473 ( \1143 , \1074 );
nand \U$474 ( \1144 , \1143 , \845 );
not \U$475 ( \1145 , \1144 );
not \U$476 ( \1146 , \1070 );
or \U$477 ( \1147 , \1145 , \1146 );
or \U$478 ( \1148 , \1144 , \1070 );
nand \U$479 ( \1149 , \1147 , \1148 );
not \U$480 ( \1150 , \1149 );
and \U$481 ( \1151 , \1142 , \1150 );
not \U$482 ( \1152 , \1149 );
and \U$483 ( \1153 , \1048 , \1036 );
nor \U$484 ( \1154 , \1153 , RIaa9ce28_188);
not \U$485 ( \1155 , \1154 );
nand \U$486 ( \1156 , \1014 , \849 );
not \U$487 ( \1157 , \1156 );
or \U$488 ( \1158 , \1155 , \1157 );
and \U$489 ( \1159 , \1057 , \916 );
nand \U$490 ( \1160 , \1158 , \1159 );
buf \U$491 ( \1161 , \1063 );
nand \U$492 ( \1162 , \1160 , \1161 );
not \U$493 ( \1163 , \1162 );
buf \U$494 ( \1164 , \954 );
and \U$495 ( \1165 , \1164 , \959 );
not \U$496 ( \1166 , \1164 );
and \U$497 ( \1167 , \1166 , \960 );
nor \U$498 ( \1168 , \1165 , \1167 );
not \U$499 ( \1169 , \1168 );
and \U$500 ( \1170 , \1163 , \1169 );
and \U$501 ( \1171 , \1162 , \1168 );
nor \U$502 ( \1172 , \1170 , \1171 );
not \U$503 ( \1173 , \1172 );
or \U$504 ( \1174 , \1152 , \1173 );
or \U$505 ( \1175 , \1172 , \1149 );
nand \U$506 ( \1176 , \1174 , \1175 );
nor \U$507 ( \1177 , \1151 , \1176 );
not \U$508 ( \1178 , \1150 );
not \U$509 ( \1179 , \1138 );
and \U$510 ( \1180 , \1076 , \1179 );
not \U$511 ( \1181 , \1076 );
and \U$512 ( \1182 , \1181 , \1138 );
nor \U$513 ( \1183 , \1180 , \1182 );
nand \U$514 ( \1184 , \1178 , \1183 );
nand \U$515 ( \1185 , \1177 , \1184 );
buf \U$516 ( \1186 , \1185 );
not \U$517 ( \1187 , \1186 );
not \U$518 ( \1188 , \1187 );
buf \U$519 ( \1189 , \1176 );
not \U$520 ( \1190 , \1189 );
and \U$521 ( \1191 , \1188 , \1190 );
buf \U$522 ( \1192 , \1142 );
buf \U$523 ( \1193 , \1192 );
nor \U$524 ( \1194 , \1191 , \1193 );
and \U$525 ( \1195 , \961 , \844 );
not \U$526 ( \1196 , \1195 );
nor \U$527 ( \1197 , \1196 , \1132 );
not \U$528 ( \1198 , \1197 );
nor \U$529 ( \1199 , \915 , \852 );
nor \U$530 ( \1200 , \1199 , \1065 );
nand \U$531 ( \1201 , \1160 , \1200 );
buf \U$532 ( \1202 , \1201 );
not \U$533 ( \1203 , \1202 );
or \U$534 ( \1204 , \1198 , \1203 );
nand \U$535 ( \1205 , \1137 , \1075 );
not \U$536 ( \1206 , \1132 );
and \U$537 ( \1207 , \1205 , \1206 );
not \U$538 ( \1208 , RIaa9a308_96);
not \U$539 ( \1209 , \765 );
or \U$540 ( \1210 , \1208 , \1209 );
nand \U$541 ( \1211 , \939 , RIaa9a218_94);
nand \U$542 ( \1212 , \1210 , \1211 );
nand \U$543 ( \1213 , \1038 , RIaa9a380_97);
not \U$544 ( \1214 , \1027 );
nand \U$545 ( \1215 , \1214 , RIaa9a038_90);
nand \U$546 ( \1216 , RIaa97d88_16, RIaa99ed0_87);
nand \U$547 ( \1217 , \1213 , \1215 , \1216 );
nor \U$548 ( \1218 , \1212 , \1217 );
not \U$549 ( \1219 , RIaa9a290_95);
not \U$550 ( \1220 , \896 );
or \U$551 ( \1221 , \1219 , \1220 );
nand \U$552 ( \1222 , \864 , RIaa9a0b0_91);
nand \U$553 ( \1223 , \1221 , \1222 );
not \U$554 ( \1224 , RIaa99fc0_89);
not \U$555 ( \1225 , \753 );
or \U$556 ( \1226 , \1224 , \1225 );
nand \U$557 ( \1227 , \867 , RIaa9a470_99);
nand \U$558 ( \1228 , \1226 , \1227 );
nor \U$559 ( \1229 , \1223 , \1228 );
not \U$560 ( \1230 , RIaa99f48_88);
not \U$561 ( \1231 , \1001 );
or \U$562 ( \1232 , \1230 , \1231 );
nand \U$563 ( \1233 , \873 , RIaa9a4e8_100);
nand \U$564 ( \1234 , \1232 , \1233 );
not \U$565 ( \1235 , RIaa9a1a0_93);
not \U$566 ( \1236 , \827 );
or \U$567 ( \1237 , \1235 , \1236 );
nand \U$568 ( \1238 , \1021 , RIaa9a3f8_98);
nand \U$569 ( \1239 , \1237 , \1238 );
nor \U$570 ( \1240 , \1234 , \1239 );
not \U$571 ( \1241 , RIaa99e58_86);
not \U$572 ( \1242 , \796 );
or \U$573 ( \1243 , \1241 , \1242 );
nand \U$574 ( \1244 , \817 , RIaa9a560_101);
nand \U$575 ( \1245 , \1243 , \1244 );
not \U$576 ( \1246 , RIaa9a128_92);
not \U$577 ( \1247 , \808 );
or \U$578 ( \1248 , \1246 , \1247 );
nand \U$579 ( \1249 , \831 , RIaa9a5d8_102);
nand \U$580 ( \1250 , \1248 , \1249 );
nor \U$581 ( \1251 , \1245 , \1250 );
nand \U$582 ( \1252 , \1218 , \1229 , \1240 , \1251 );
not \U$583 ( \1253 , \1252 );
xor \U$584 ( \1254 , \1129 , RIaa97950_7);
not \U$585 ( \1255 , \1254 );
nand \U$586 ( \1256 , \1253 , \1255 );
not \U$587 ( \1257 , \1256 );
nor \U$588 ( \1258 , \1207 , \1257 );
nand \U$589 ( \1259 , \1204 , \1258 );
nand \U$590 ( \1260 , \1252 , \1254 );
not \U$591 ( \1261 , \1260 );
not \U$592 ( \1262 , \1261 );
nand \U$593 ( \1263 , \1259 , \1262 );
not \U$594 ( \1264 , \827 );
not \U$595 ( \1265 , RIaa99b10_79);
or \U$596 ( \1266 , \1264 , \1265 );
not \U$597 ( \1267 , \1001 );
not \U$598 ( \1268 , RIaa999a8_76);
or \U$599 ( \1269 , \1267 , \1268 );
nand \U$600 ( \1270 , \1266 , \1269 );
nand \U$601 ( \1271 , \1214 , RIaa99a20_77);
nand \U$602 ( \1272 , \1021 , RIaa996d8_70);
nand \U$603 ( \1273 , RIaa97d88_16, RIaa99930_75);
nand \U$604 ( \1274 , \1271 , \1272 , \1273 );
nor \U$605 ( \1275 , \1270 , \1274 );
not \U$606 ( \1276 , \895 );
not \U$607 ( \1277 , RIaa99d68_84);
not \U$608 ( \1278 , \1277 );
and \U$609 ( \1279 , \1276 , \1278 );
and \U$610 ( \1280 , \864 , RIaa99b88_80);
nor \U$611 ( \1281 , \1279 , \1280 );
not \U$612 ( \1282 , \1281 );
not \U$613 ( \1283 , RIaa99660_69);
not \U$614 ( \1284 , \744 );
or \U$615 ( \1285 , \1283 , \1284 );
nand \U$616 ( \1286 , \867 , RIaa99cf0_83);
nand \U$617 ( \1287 , \1285 , \1286 );
nor \U$618 ( \1288 , \1282 , \1287 );
nand \U$619 ( \1289 , \785 , RIaa99c00_81);
nand \U$620 ( \1290 , \753 , RIaa998b8_74);
nand \U$621 ( \1291 , RIaa99de0_85, \831 );
nand \U$622 ( \1292 , RIaa99a98_78, \808 );
and \U$623 ( \1293 , \1289 , \1290 , \1291 , \1292 );
not \U$624 ( \1294 , RIaa99c78_82);
not \U$625 ( \1295 , \1104 );
or \U$626 ( \1296 , \1294 , \1295 );
nand \U$627 ( \1297 , \817 , RIaa997c8_72);
nand \U$628 ( \1298 , \1296 , \1297 );
not \U$629 ( \1299 , RIaa99840_73);
not \U$630 ( \1300 , \796 );
or \U$631 ( \1301 , \1299 , \1300 );
nand \U$632 ( \1302 , \873 , RIaa99750_71);
nand \U$633 ( \1303 , \1301 , \1302 );
nor \U$634 ( \1304 , \1298 , \1303 );
nand \U$635 ( \1305 , \1275 , \1288 , \1293 , \1304 );
not \U$636 ( \1306 , \1124 );
and \U$637 ( \1307 , \1306 , RIaa97950_7, RIaa978d8_6);
nor \U$638 ( \1308 , \1307 , RIaa979c8_8);
not \U$639 ( \1309 , \836 );
and \U$640 ( \1310 , \1309 , RIaa979c8_8, RIaa97950_7, RIaa978d8_6);
or \U$641 ( \1311 , \1308 , \1310 );
nand \U$642 ( \1312 , \1305 , \1311 );
not \U$643 ( \1313 , \1312 );
not \U$644 ( \1314 , \1313 );
not \U$645 ( \1315 , \1303 );
buf \U$646 ( \1316 , \827 );
nand \U$647 ( \1317 , \1316 , RIaa99b10_79);
and \U$648 ( \1318 , \1315 , \1281 , \1317 );
not \U$649 ( \1319 , \1001 );
or \U$650 ( \1320 , \1319 , \1268 );
not \U$651 ( \1321 , \1311 );
nand \U$652 ( \1322 , \1320 , \1321 );
nor \U$653 ( \1323 , \1274 , \1322 );
nor \U$654 ( \1324 , \1287 , \1298 );
nand \U$655 ( \1325 , \1318 , \1323 , \1293 , \1324 );
buf \U$656 ( \1326 , \1325 );
nand \U$657 ( \1327 , \1314 , \1326 );
and \U$658 ( \1328 , \1263 , \1327 );
not \U$659 ( \1329 , \1263 );
not \U$660 ( \1330 , \1327 );
and \U$661 ( \1331 , \1329 , \1330 );
nor \U$662 ( \1332 , \1328 , \1331 );
buf \U$663 ( \1333 , \1332 );
not \U$664 ( \1334 , \1333 );
buf \U$665 ( \1335 , \1334 );
not \U$666 ( \1336 , \1332 );
not \U$667 ( \1337 , \1205 );
not \U$668 ( \1338 , \1337 );
nand \U$669 ( \1339 , \1070 , \845 );
not \U$670 ( \1340 , \1339 );
or \U$671 ( \1341 , \1338 , \1340 );
nand \U$672 ( \1342 , \1341 , \1206 );
buf \U$673 ( \1343 , \1252 );
and \U$674 ( \1344 , \1343 , \1255 );
not \U$675 ( \1345 , \1343 );
and \U$676 ( \1346 , \1345 , \1254 );
nor \U$677 ( \1347 , \1344 , \1346 );
not \U$678 ( \1348 , \1347 );
and \U$679 ( \1349 , \1342 , \1348 );
not \U$680 ( \1350 , \1342 );
and \U$681 ( \1351 , \1350 , \1347 );
nor \U$682 ( \1352 , \1349 , \1351 );
and \U$683 ( \1353 , \1336 , \1352 );
not \U$684 ( \1354 , \1336 );
not \U$685 ( \1355 , \1352 );
and \U$686 ( \1356 , \1354 , \1355 );
nor \U$687 ( \1357 , \1353 , \1356 );
not \U$688 ( \1358 , \1183 );
not \U$689 ( \1359 , \1352 );
not \U$690 ( \1360 , \1359 );
or \U$691 ( \1361 , \1358 , \1360 );
nand \U$692 ( \1362 , \1352 , \1142 );
nand \U$693 ( \1363 , \1361 , \1362 );
nand \U$694 ( \1364 , \1357 , \1363 );
nor \U$695 ( \1365 , \1335 , \1364 );
not \U$696 ( \1366 , \1365 );
not \U$697 ( \1367 , \1366 );
not \U$698 ( \1368 , \1367 );
buf \U$699 ( \1369 , \782 );
not \U$700 ( \1370 , \1369 );
not \U$701 ( \1371 , \862 );
buf \U$702 ( \1372 , \714 );
not \U$703 ( \1373 , \1372 );
nand \U$704 ( \1374 , \1371 , \1373 );
nor \U$705 ( \1375 , \780 , \1374 );
buf \U$706 ( \1376 , \759 );
and \U$707 ( \1377 , \1375 , \1376 );
not \U$708 ( \1378 , \1377 );
or \U$709 ( \1379 , \1370 , \1378 );
buf \U$710 ( \1380 , \1374 );
not \U$711 ( \1381 , \1376 );
or \U$712 ( \1382 , \1380 , \1381 , \780 );
not \U$713 ( \1383 , \1369 );
nand \U$714 ( \1384 , \1382 , \1383 );
nand \U$715 ( \1385 , \1379 , \1384 );
buf \U$716 ( \1386 , \1385 );
not \U$717 ( \1387 , \1386 );
buf \U$718 ( \1388 , \1376 );
not \U$719 ( \1389 , \1388 );
buf \U$720 ( \1390 , \1375 );
not \U$721 ( \1391 , \1390 );
or \U$722 ( \1392 , \1389 , \1391 );
or \U$723 ( \1393 , \1388 , \1390 );
nand \U$724 ( \1394 , \1392 , \1393 );
not \U$725 ( \1395 , \1394 );
buf \U$726 ( \1396 , \1395 );
not \U$727 ( \1397 , \1396 );
not \U$728 ( \1398 , \780 );
and \U$729 ( \1399 , \1398 , \1373 );
not \U$730 ( \1400 , \1398 );
and \U$731 ( \1401 , \1400 , \1380 );
nor \U$732 ( \1402 , \1399 , \1401 );
not \U$733 ( \1403 , \1402 );
buf \U$734 ( \1404 , \821 );
nand \U$735 ( \1405 , \1403 , \1404 );
not \U$736 ( \1406 , \1373 );
nand \U$737 ( \1407 , \1406 , \1371 );
buf \U$738 ( \1408 , \717 );
nand \U$739 ( \1409 , \1407 , \1408 );
and \U$740 ( \1410 , \1405 , \1409 );
buf \U$741 ( \1411 , \1410 );
and \U$742 ( \1412 , \1387 , \1397 , \1411 );
buf \U$743 ( \1413 , \1412 );
not \U$744 ( \1414 , \1413 );
not \U$745 ( \1415 , \1414 );
not \U$746 ( \1416 , RIaa9f6f0_275);
not \U$747 ( \1417 , \1416 );
and \U$748 ( \1418 , \1415 , \1417 );
not \U$749 ( \1419 , \1395 );
buf \U$750 ( \1420 , \1419 );
not \U$751 ( \1421 , \1404 );
nor \U$752 ( \1422 , \1421 , \1402 );
buf \U$753 ( \1423 , \1422 );
not \U$754 ( \1424 , \1409 );
and \U$755 ( \1425 , \1423 , \1424 );
nand \U$756 ( \1426 , \1387 , \1420 , \1425 );
not \U$757 ( \1427 , RIaa9f768_276);
nor \U$758 ( \1428 , \1426 , \1427 );
nor \U$759 ( \1429 , \1418 , \1428 );
not \U$760 ( \1430 , \1385 );
not \U$761 ( \1431 , \1430 );
not \U$762 ( \1432 , \1431 );
and \U$763 ( \1433 , \1422 , \1409 );
and \U$764 ( \1434 , \1432 , \1397 , \1433 );
not \U$765 ( \1435 , \1434 );
not \U$766 ( \1436 , \1435 );
buf \U$767 ( \1437 , \1436 );
and \U$768 ( \1438 , \1437 , RIaa9f3a8_268);
nand \U$769 ( \1439 , \1410 , \1395 );
not \U$770 ( \1440 , \1430 );
nor \U$771 ( \1441 , \1439 , \1440 );
not \U$772 ( \1442 , \1441 );
not \U$773 ( \1443 , \1442 );
not \U$774 ( \1444 , \1443 );
not \U$775 ( \1445 , RIaa9f600_273);
or \U$776 ( \1446 , \1444 , \1445 );
nor \U$777 ( \1447 , \1432 , \1439 );
not \U$778 ( \1448 , \1447 );
not \U$779 ( \1449 , \1448 );
nand \U$780 ( \1450 , \1449 , RIaa9f2b8_266);
nand \U$781 ( \1451 , \1446 , \1450 );
nor \U$782 ( \1452 , \1438 , \1451 );
nand \U$783 ( \1453 , \1429 , \1452 );
not \U$784 ( \1454 , \1387 );
buf \U$785 ( \1455 , \1405 );
and \U$786 ( \1456 , \1455 , \1424 );
nand \U$787 ( \1457 , \1454 , \1420 , \1456 );
not \U$788 ( \1458 , \1457 );
and \U$789 ( \1459 , \1458 , RIaa9f330_267);
nand \U$790 ( \1460 , \1411 , \1420 , \1431 );
not \U$791 ( \1461 , \1460 );
not \U$792 ( \1462 , \1461 );
not \U$793 ( \1463 , \1462 );
and \U$794 ( \1464 , \1463 , RIaa9f420_269);
nor \U$795 ( \1465 , \1459 , \1464 );
not \U$796 ( \1466 , \1395 );
nor \U$797 ( \1467 , \1466 , \1409 );
nor \U$798 ( \1468 , \1385 , \1423 );
nand \U$799 ( \1469 , \1467 , \1468 );
not \U$800 ( \1470 , \1469 );
and \U$801 ( \1471 , \1470 , RIaa9f9c0_281);
buf \U$802 ( \1472 , \1455 );
and \U$803 ( \1473 , \1386 , \1396 , \1472 , \1424 );
buf \U$804 ( \1474 , \1473 );
and \U$805 ( \1475 , \1474 , RIaa9f948_280);
nor \U$806 ( \1476 , \1471 , \1475 );
nand \U$807 ( \1477 , \1465 , \1476 );
nor \U$808 ( \1478 , \1453 , \1477 );
and \U$809 ( \1479 , \1456 , \1419 , \1430 );
buf \U$810 ( \1480 , \1479 );
and \U$811 ( \1481 , \1480 , RIaa9f678_274);
and \U$812 ( \1482 , \1396 , \1430 , \1433 );
buf \U$813 ( \1483 , \1482 );
not \U$814 ( \1484 , \1483 );
not \U$815 ( \1485 , RIaa9f8d0_279);
or \U$816 ( \1486 , \1484 , \1485 );
not \U$817 ( \1487 , \1369 );
not \U$818 ( \1488 , \1377 );
or \U$819 ( \1489 , \1487 , \1488 );
not \U$820 ( \1490 , RIaa97d88_16);
nand \U$821 ( \1491 , \1489 , \1490 );
and \U$822 ( \1492 , \1491 , RIaa9f588_272);
not \U$823 ( \1493 , RIaa9f240_265);
buf \U$824 ( \1494 , \753 );
not \U$825 ( \1495 , \1494 );
nor \U$826 ( \1496 , \1493 , \1495 );
nor \U$827 ( \1497 , \1492 , \1496 );
nand \U$828 ( \1498 , \1486 , \1497 );
nor \U$829 ( \1499 , \1481 , \1498 );
not \U$830 ( \1500 , \1396 );
and \U$831 ( \1501 , \1500 , \1440 , \1433 );
buf \U$832 ( \1502 , \1501 );
and \U$833 ( \1503 , \1502 , RIaa9f510_271);
not \U$834 ( \1504 , \1467 );
not \U$835 ( \1505 , \1504 );
nor \U$836 ( \1506 , \1472 , \1440 );
nand \U$837 ( \1507 , \1505 , \1506 );
not \U$838 ( \1508 , \1507 );
and \U$839 ( \1509 , RIaa9f7e0_277, \1508 );
nor \U$840 ( \1510 , \1503 , \1509 );
and \U$841 ( \1511 , \1431 , \1396 , \1423 , \1424 );
buf \U$842 ( \1512 , \1511 );
and \U$843 ( \1513 , \1512 , RIaa9f858_278);
nand \U$844 ( \1514 , \1396 , \1433 );
or \U$845 ( \1515 , \1514 , \1387 );
not \U$846 ( \1516 , \1515 );
and \U$847 ( \1517 , \1516 , RIaa9f498_270);
nor \U$848 ( \1518 , \1513 , \1517 );
and \U$849 ( \1519 , \1499 , \1510 , \1518 );
and \U$850 ( \1520 , \1478 , \1519 );
not \U$851 ( \1521 , \1520 );
not \U$852 ( \1522 , \1521 );
not \U$853 ( \1523 , \1522 );
or \U$854 ( \1524 , \1368 , \1523 );
and \U$855 ( \1525 , \1458 , RIaa9eca0_253);
and \U$856 ( \1526 , \1463 , RIaa9ee08_256);
nor \U$857 ( \1527 , \1525 , \1526 );
and \U$858 ( \1528 , \1413 , RIaa9eef8_258);
and \U$859 ( \1529 , RIaa9ed90_255, \1516 );
not \U$860 ( \1530 , \1482 );
not \U$861 ( \1531 , \1530 );
and \U$862 ( \1532 , \1531 , RIaa9f1c8_264);
nor \U$863 ( \1533 , \1528 , \1529 , \1532 );
and \U$864 ( \1534 , \1470 , RIaa9efe8_260);
and \U$865 ( \1535 , \1474 , RIaa9ef70_259);
nor \U$866 ( \1536 , \1534 , \1535 );
nand \U$867 ( \1537 , \1527 , \1533 , \1536 );
not \U$868 ( \1538 , \1537 );
and \U$869 ( \1539 , \1437 , RIaa9ed18_254);
not \U$870 ( \1540 , RIaa9eb38_250);
not \U$871 ( \1541 , \1442 );
not \U$872 ( \1542 , \1541 );
or \U$873 ( \1543 , \1540 , \1542 );
and \U$874 ( \1544 , \1491 , RIaa9ebb0_251);
not \U$875 ( \1545 , RIaa9ea48_248);
nor \U$876 ( \1546 , \1545 , \1495 );
nor \U$877 ( \1547 , \1544 , \1546 );
nand \U$878 ( \1548 , \1543 , \1547 );
nor \U$879 ( \1549 , \1539 , \1548 );
and \U$880 ( \1550 , \1420 , \1432 , \1425 );
buf \U$881 ( \1551 , \1550 );
and \U$882 ( \1552 , \1551 , RIaa9f0d8_262);
and \U$883 ( \1553 , \1480 , RIaa9ee80_257);
nor \U$884 ( \1554 , \1552 , \1553 );
and \U$885 ( \1555 , \1502 , RIaa9eac0_249);
not \U$886 ( \1556 , RIaa9f150_263);
not \U$887 ( \1557 , \1504 );
and \U$888 ( \1558 , \1440 , \1423 );
nand \U$889 ( \1559 , \1557 , \1558 );
not \U$890 ( \1560 , \1559 );
not \U$891 ( \1561 , \1560 );
nor \U$892 ( \1562 , \1556 , \1561 );
nor \U$893 ( \1563 , \1555 , \1562 );
not \U$894 ( \1564 , \1507 );
not \U$895 ( \1565 , \1564 );
not \U$896 ( \1566 , \1565 );
and \U$897 ( \1567 , \1566 , RIaa9f060_261);
and \U$898 ( \1568 , \1449 , RIaa9ec28_252);
nor \U$899 ( \1569 , \1567 , \1568 );
and \U$900 ( \1570 , \1549 , \1554 , \1563 , \1569 );
nand \U$901 ( \1571 , \1538 , \1570 );
not \U$902 ( \1572 , \1571 );
not \U$903 ( \1573 , \1572 );
not \U$904 ( \1574 , \1363 );
not \U$905 ( \1575 , \1333 );
nand \U$906 ( \1576 , \1574 , \1575 );
not \U$907 ( \1577 , \1576 );
not \U$908 ( \1578 , \1577 );
not \U$909 ( \1579 , \1578 );
and \U$910 ( \1580 , \1573 , \1579 );
not \U$911 ( \1581 , \1573 );
nor \U$912 ( \1582 , \1334 , \1363 );
buf \U$913 ( \1583 , \1582 );
buf \U$914 ( \1584 , \1583 );
and \U$915 ( \1585 , \1581 , \1584 );
nor \U$916 ( \1586 , \1580 , \1585 );
nand \U$917 ( \1587 , \1524 , \1586 );
not \U$918 ( \1588 , \1575 );
nor \U$919 ( \1589 , \1364 , \1588 );
not \U$920 ( \1590 , \1589 );
not \U$921 ( \1591 , \1590 );
not \U$922 ( \1592 , \1591 );
nor \U$923 ( \1593 , \1592 , \1522 );
nor \U$924 ( \1594 , \1587 , \1593 );
xor \U$925 ( \1595 , \1194 , \1594 );
not \U$926 ( \1596 , \1595 );
not \U$927 ( \1597 , RIaa97b30_11);
not \U$928 ( \1598 , \1597 );
nand \U$929 ( \1599 , \1310 , RIaa97ba8_12);
not \U$930 ( \1600 , \1599 );
or \U$931 ( \1601 , \1598 , \1600 );
not \U$932 ( \1602 , \1599 );
nand \U$933 ( \1603 , \1602 , RIaa97b30_11);
nand \U$934 ( \1604 , \1601 , \1603 );
not \U$935 ( \1605 , \1604 );
not \U$936 ( \1606 , \1605 );
not \U$937 ( \1607 , RIaa9de18_222);
buf \U$938 ( \1608 , \1214 );
not \U$939 ( \1609 , \1608 );
or \U$940 ( \1610 , \1607 , \1609 );
nand \U$941 ( \1611 , RIaa97d88_16, RIaa9db48_216);
nand \U$942 ( \1612 , \1610 , \1611 );
buf \U$943 ( \1613 , \1021 );
not \U$944 ( \1614 , \1613 );
not \U$945 ( \1615 , RIaa9d968_212);
nor \U$946 ( \1616 , \1614 , \1615 );
nor \U$947 ( \1617 , \1612 , \1616 );
not \U$948 ( \1618 , \1264 );
not \U$949 ( \1619 , RIaa9dbc0_217);
not \U$950 ( \1620 , \1619 );
and \U$951 ( \1621 , \1618 , \1620 );
not \U$952 ( \1622 , \1319 );
and \U$953 ( \1623 , \1622 , RIaa9dda0_221);
nor \U$954 ( \1624 , \1621 , \1623 );
nand \U$955 ( \1625 , \1617 , \1624 );
buf \U$956 ( \1626 , \785 );
nand \U$957 ( \1627 , \1626 , RIaa9dd28_220);
nand \U$958 ( \1628 , \1494 , RIaa9dad0_215);
buf \U$959 ( \1629 , \831 );
nand \U$960 ( \1630 , \1629 , RIaa9d800_209);
buf \U$961 ( \1631 , \808 );
nand \U$962 ( \1632 , \1631 , RIaa9dc38_218);
nand \U$963 ( \1633 , \1627 , \1628 , \1630 , \1632 );
nor \U$964 ( \1634 , \1625 , \1633 );
buf \U$965 ( \1635 , \1104 );
nand \U$966 ( \1636 , \1635 , RIaa9d710_207);
buf \U$967 ( \1637 , \864 );
nand \U$968 ( \1638 , \1637 , RIaa9dcb0_219);
buf \U$969 ( \1639 , \895 );
not \U$970 ( \1640 , \1639 );
nand \U$971 ( \1641 , \1640 , RIaa9d788_208);
buf \U$972 ( \1642 , \867 );
nand \U$973 ( \1643 , \1642 , RIaa9d698_206);
nand \U$974 ( \1644 , \1636 , \1638 , \1641 , \1643 );
buf \U$975 ( \1645 , \796 );
nand \U$976 ( \1646 , \1645 , RIaa9da58_214);
buf \U$977 ( \1647 , \744 );
nand \U$978 ( \1648 , \1647 , RIaa9d9e0_213);
buf \U$979 ( \1649 , \873 );
nand \U$980 ( \1650 , \1649 , RIaa9d878_210);
buf \U$981 ( \1651 , \817 );
nand \U$982 ( \1652 , \1651 , RIaa9d8f0_211);
nand \U$983 ( \1653 , \1646 , \1648 , \1650 , \1652 );
nor \U$984 ( \1654 , \1644 , \1653 );
nand \U$985 ( \1655 , \1634 , \1654 );
not \U$986 ( \1656 , \1655 );
not \U$987 ( \1657 , \1656 );
or \U$988 ( \1658 , \1606 , \1657 );
nand \U$989 ( \1659 , \1629 , RIaa994f8_66);
nand \U$990 ( \1660 , \1608 , RIaa99048_56);
nand \U$991 ( \1661 , RIaa97d88_16, RIaa98f58_54);
nand \U$992 ( \1662 , \1659 , \1660 , \1661 );
not \U$993 ( \1663 , RIaa99570_67);
not \U$994 ( \1664 , \1647 );
or \U$995 ( \1665 , \1663 , \1664 );
nand \U$996 ( \1666 , \1635 , RIaa990c0_57);
nand \U$997 ( \1667 , \1665 , \1666 );
nor \U$998 ( \1668 , \1662 , \1667 );
not \U$999 ( \1669 , RIaa99138_58);
not \U$1000 ( \1670 , \1639 );
not \U$1001 ( \1671 , \1670 );
or \U$1002 ( \1672 , \1669 , \1671 );
nand \U$1003 ( \1673 , \1637 , RIaa99390_63);
nand \U$1004 ( \1674 , \1672 , \1673 );
not \U$1005 ( \1675 , RIaa98ee0_53);
not \U$1006 ( \1676 , \1494 );
or \U$1007 ( \1677 , \1675 , \1676 );
nand \U$1008 ( \1678 , \1642 , RIaa99480_65);
nand \U$1009 ( \1679 , \1677 , \1678 );
nor \U$1010 ( \1680 , \1674 , \1679 );
not \U$1011 ( \1681 , RIaa98fd0_55);
not \U$1012 ( \1682 , \1319 );
not \U$1013 ( \1683 , \1682 );
or \U$1014 ( \1684 , \1681 , \1683 );
nand \U$1015 ( \1685 , \1613 , RIaa995e8_68);
nand \U$1016 ( \1686 , \1684 , \1685 );
not \U$1017 ( \1687 , RIaa99318_62);
not \U$1018 ( \1688 , \1316 );
or \U$1019 ( \1689 , \1687 , \1688 );
nand \U$1020 ( \1690 , \1649 , RIaa991b0_59);
nand \U$1021 ( \1691 , \1689 , \1690 );
nor \U$1022 ( \1692 , \1686 , \1691 );
not \U$1023 ( \1693 , RIaa99408_64);
not \U$1024 ( \1694 , \1626 );
or \U$1025 ( \1695 , \1693 , \1694 );
nand \U$1026 ( \1696 , \1631 , RIaa992a0_61);
nand \U$1027 ( \1697 , \1695 , \1696 );
not \U$1028 ( \1698 , RIaa98e68_52);
not \U$1029 ( \1699 , \1645 );
or \U$1030 ( \1700 , \1698 , \1699 );
nand \U$1031 ( \1701 , \1651 , RIaa99228_60);
nand \U$1032 ( \1702 , \1700 , \1701 );
nor \U$1033 ( \1703 , \1697 , \1702 );
nand \U$1034 ( \1704 , \1668 , \1680 , \1692 , \1703 );
not \U$1035 ( \1705 , \1704 );
nor \U$1036 ( \1706 , \1310 , RIaa97ba8_12);
not \U$1037 ( \1707 , \1706 );
nand \U$1038 ( \1708 , \1707 , \1599 );
buf \U$1039 ( \1709 , \1708 );
not \U$1040 ( \1710 , \1709 );
nand \U$1041 ( \1711 , \1705 , \1710 );
nand \U$1042 ( \1712 , \1658 , \1711 );
not \U$1043 ( \1713 , \1712 );
and \U$1044 ( \1714 , \1131 , \1195 , \1260 , \1312 );
nand \U$1045 ( \1715 , \1704 , \1709 );
nand \U$1046 ( \1716 , \1202 , \1714 , \1715 );
and \U$1047 ( \1717 , \1326 , \1261 );
nor \U$1048 ( \1718 , \1717 , \1313 );
not \U$1049 ( \1719 , \1074 );
not \U$1050 ( \1720 , \1131 );
or \U$1051 ( \1721 , \1719 , \1720 );
and \U$1052 ( \1722 , \1136 , \1256 , \1325 );
nand \U$1053 ( \1723 , \1721 , \1722 );
nand \U$1054 ( \1724 , \1718 , \1723 , \1715 );
nand \U$1055 ( \1725 , \1713 , \1716 , \1724 );
nand \U$1056 ( \1726 , \1655 , \1604 );
buf \U$1057 ( \1727 , \1726 );
nand \U$1058 ( \1728 , \1725 , \1727 );
not \U$1059 ( \1729 , RIaa9e160_229);
not \U$1060 ( \1730 , \1608 );
or \U$1061 ( \1731 , \1729 , \1730 );
nand \U$1062 ( \1732 , RIaa97d88_16, RIaa9df80_225);
nand \U$1063 ( \1733 , \1731 , \1732 );
not \U$1064 ( \1734 , RIaa9e3b8_234);
not \U$1065 ( \1735 , \1649 );
nor \U$1066 ( \1736 , \1734 , \1735 );
nor \U$1067 ( \1737 , \1733 , \1736 );
and \U$1068 ( \1738 , \1645 , RIaa9de90_223);
and \U$1069 ( \1739 , \1629 , RIaa9e610_239);
nor \U$1070 ( \1740 , \1738 , \1739 );
nand \U$1071 ( \1741 , \1737 , \1740 );
not \U$1072 ( \1742 , RIaa9e2c8_232);
not \U$1073 ( \1743 , \1642 );
nor \U$1074 ( \1744 , \1742 , \1743 );
not \U$1075 ( \1745 , \1640 );
not \U$1076 ( \1746 , RIaa9e598_238);
nor \U$1077 ( \1747 , \1745 , \1746 );
nor \U$1078 ( \1748 , \1744 , \1747 );
and \U$1079 ( \1749 , \1637 , RIaa9e1d8_230);
not \U$1080 ( \1750 , RIaa9df08_224);
nor \U$1081 ( \1751 , \1495 , \1750 );
nor \U$1082 ( \1752 , \1749 , \1751 );
nand \U$1083 ( \1753 , \1748 , \1752 );
nor \U$1084 ( \1754 , \1741 , \1753 );
buf \U$1085 ( \1755 , \1647 );
nand \U$1086 ( \1756 , \1755 , RIaa9e520_237);
nand \U$1087 ( \1757 , RIaa9e340_233, \1635 );
nand \U$1088 ( \1758 , \1626 , RIaa9e250_231);
nand \U$1089 ( \1759 , \1651 , RIaa9e430_235);
nand \U$1090 ( \1760 , \1756 , \1757 , \1758 , \1759 );
nand \U$1091 ( \1761 , \1622 , RIaa9e0e8_228);
nand \U$1092 ( \1762 , \1316 , RIaa9dff8_226);
nand \U$1093 ( \1763 , \1613 , RIaa9e4a8_236);
nand \U$1094 ( \1764 , \1631 , RIaa9e070_227);
nand \U$1095 ( \1765 , \1761 , \1762 , \1763 , \1764 );
nor \U$1096 ( \1766 , \1760 , \1765 );
nand \U$1097 ( \1767 , \1754 , \1766 );
buf \U$1098 ( \1768 , \1767 );
not \U$1099 ( \1769 , RIaa97ab8_10);
and \U$1100 ( \1770 , \1603 , \1769 );
not \U$1101 ( \1771 , \1603 );
and \U$1102 ( \1772 , \1771 , RIaa97ab8_10);
nor \U$1103 ( \1773 , \1770 , \1772 );
not \U$1104 ( \1774 , \1773 );
and \U$1105 ( \1775 , \1768 , \1774 );
not \U$1106 ( \1776 , \1768 );
and \U$1107 ( \1777 , \1776 , \1773 );
nor \U$1108 ( \1778 , \1775 , \1777 );
and \U$1109 ( \1779 , \1728 , \1778 );
not \U$1110 ( \1780 , \1728 );
not \U$1111 ( \1781 , \1778 );
and \U$1112 ( \1782 , \1780 , \1781 );
nor \U$1113 ( \1783 , \1779 , \1782 );
not \U$1114 ( \1784 , \1783 );
buf \U$1115 ( \1785 , \1711 );
nand \U$1116 ( \1786 , \1716 , \1724 , \1785 );
not \U$1117 ( \1787 , \1786 );
not \U$1118 ( \1788 , \1605 );
not \U$1119 ( \1789 , \1656 );
or \U$1120 ( \1790 , \1788 , \1789 );
nand \U$1121 ( \1791 , \1790 , \1727 );
not \U$1122 ( \1792 , \1791 );
and \U$1123 ( \1793 , \1787 , \1792 );
and \U$1124 ( \1794 , \1786 , \1791 );
nor \U$1125 ( \1795 , \1793 , \1794 );
not \U$1126 ( \1796 , \1795 );
not \U$1127 ( \1797 , \1796 );
and \U$1128 ( \1798 , \1784 , \1797 );
and \U$1129 ( \1799 , \1796 , \1783 );
nor \U$1130 ( \1800 , \1798 , \1799 );
not \U$1131 ( \1801 , \1800 );
not \U$1132 ( \1802 , \1783 );
nand \U$1133 ( \1803 , \1767 , \1774 );
and \U$1134 ( \1804 , \1726 , \1715 , \1803 );
not \U$1135 ( \1805 , \1804 );
not \U$1136 ( \1806 , \1714 );
not \U$1137 ( \1807 , \1201 );
or \U$1138 ( \1808 , \1806 , \1807 );
nand \U$1139 ( \1809 , \1723 , \1718 );
nand \U$1140 ( \1810 , \1808 , \1809 );
not \U$1141 ( \1811 , \1810 );
or \U$1142 ( \1812 , \1805 , \1811 );
nand \U$1143 ( \1813 , \1726 , \1803 );
not \U$1144 ( \1814 , \1813 );
and \U$1145 ( \1815 , \1814 , \1712 );
nor \U$1146 ( \1816 , \1768 , \1774 );
nor \U$1147 ( \1817 , \1815 , \1816 );
nand \U$1148 ( \1818 , \1812 , \1817 );
not \U$1149 ( \1819 , \1818 );
not \U$1150 ( \1820 , \1603 );
and \U$1151 ( \1821 , \1820 , RIaa97ab8_10);
nor \U$1152 ( \1822 , \1821 , RIaa97a40_9);
and \U$1153 ( \1823 , RIaa97a40_9, RIaa97ab8_10, RIaa97b30_11, RIaa97ba8_12);
and \U$1154 ( \1824 , \1310 , \1823 );
nor \U$1155 ( \1825 , \1822 , \1824 );
buf \U$1156 ( \1826 , \1825 );
not \U$1157 ( \1827 , \1826 );
not \U$1158 ( \1828 , \1745 );
not \U$1159 ( \1829 , RIaa98b20_45);
not \U$1160 ( \1830 , \1829 );
and \U$1161 ( \1831 , \1828 , \1830 );
buf \U$1162 ( \1832 , \1637 );
and \U$1163 ( \1833 , \1832 , RIaa989b8_42);
nor \U$1164 ( \1834 , \1831 , \1833 );
not \U$1165 ( \1835 , RIaa98c88_48);
nor \U$1166 ( \1836 , \1835 , \1743 );
not \U$1167 ( \1837 , RIaa98a30_43);
not \U$1168 ( \1838 , \1626 );
nor \U$1169 ( \1839 , \1837 , \1838 );
nor \U$1170 ( \1840 , \1836 , \1839 );
nand \U$1171 ( \1841 , \1834 , \1840 );
not \U$1172 ( \1842 , \1635 );
not \U$1173 ( \1843 , \1842 );
nand \U$1174 ( \1844 , \1843 , RIaa98aa8_44);
nand \U$1175 ( \1845 , \1755 , RIaa98df0_51);
buf \U$1176 ( \1846 , \1631 );
nand \U$1177 ( \1847 , \1846 , RIaa98940_41);
nand \U$1178 ( \1848 , \1651 , RIaa98c10_47);
nand \U$1179 ( \1849 , \1844 , \1845 , \1847 , \1848 );
nor \U$1180 ( \1850 , \1841 , \1849 );
not \U$1181 ( \1851 , RIaa98670_35);
not \U$1182 ( \1852 , \1645 );
nor \U$1183 ( \1853 , \1851 , \1852 );
not \U$1184 ( \1854 , RIaa98850_39);
not \U$1185 ( \1855 , \1608 );
or \U$1186 ( \1856 , \1854 , \1855 );
nand \U$1187 ( \1857 , RIaa97d88_16, RIaa98760_37);
nand \U$1188 ( \1858 , \1856 , \1857 );
nor \U$1189 ( \1859 , \1853 , \1858 );
and \U$1190 ( \1860 , \1494 , RIaa986e8_36);
buf \U$1191 ( \1861 , \1629 );
and \U$1192 ( \1862 , \1861 , RIaa98d00_49);
nor \U$1193 ( \1863 , \1860 , \1862 );
nand \U$1194 ( \1864 , \1859 , \1863 );
not \U$1195 ( \1865 , RIaa98b98_46);
nor \U$1196 ( \1866 , \1865 , \1735 );
not \U$1197 ( \1867 , RIaa987d8_38);
not \U$1198 ( \1868 , \1682 );
nor \U$1199 ( \1869 , \1867 , \1868 );
nor \U$1200 ( \1870 , \1866 , \1869 );
buf \U$1201 ( \1871 , \1264 );
not \U$1202 ( \1872 , \1871 );
and \U$1203 ( \1873 , \1872 , RIaa988c8_40);
buf \U$1204 ( \1874 , \1613 );
and \U$1205 ( \1875 , \1874 , RIaa98d78_50);
nor \U$1206 ( \1876 , \1873 , \1875 );
nand \U$1207 ( \1877 , \1870 , \1876 );
nor \U$1208 ( \1878 , \1864 , \1877 );
nand \U$1209 ( \1879 , \1850 , \1878 );
not \U$1210 ( \1880 , \1879 );
not \U$1211 ( \1881 , \1880 );
or \U$1212 ( \1882 , \1827 , \1881 );
or \U$1213 ( \1883 , \1880 , \1826 );
nand \U$1214 ( \1884 , \1882 , \1883 );
and \U$1215 ( \1885 , \1819 , \1884 );
not \U$1216 ( \1886 , \1819 );
not \U$1217 ( \1887 , \1884 );
and \U$1218 ( \1888 , \1886 , \1887 );
nor \U$1219 ( \1889 , \1885 , \1888 );
nor \U$1220 ( \1890 , \1802 , \1889 );
not \U$1221 ( \1891 , \1890 );
not \U$1222 ( \1892 , \1783 );
nand \U$1223 ( \1893 , \1892 , \1889 );
nand \U$1224 ( \1894 , \1891 , \1893 );
nor \U$1225 ( \1895 , \1801 , \1894 );
not \U$1226 ( \1896 , \1889 );
buf \U$1227 ( \1897 , \1896 );
not \U$1228 ( \1898 , \1897 );
and \U$1229 ( \1899 , \1895 , \1898 );
buf \U$1230 ( \1900 , \1899 );
not \U$1231 ( \1901 , \1900 );
and \U$1232 ( \1902 , \1437 , RIaaa1ce8_356);
and \U$1233 ( \1903 , \1480 , RIaaa1e50_359);
nor \U$1234 ( \1904 , \1902 , \1903 );
nand \U$1235 ( \1905 , \1550 , RIaaa2030_363);
and \U$1236 ( \1906 , \1470 , RIaaa1fb8_362);
and \U$1237 ( \1907 , \1474 , RIaaa1f40_361);
nor \U$1238 ( \1908 , \1906 , \1907 );
nand \U$1239 ( \1909 , \1904 , \1905 , \1908 );
and \U$1240 ( \1910 , \1458 , RIaaa1c70_355);
and \U$1241 ( \1911 , \1463 , RIaaa1d60_357);
nor \U$1242 ( \1912 , \1910 , \1911 );
nand \U$1243 ( \1913 , \1413 , RIaaa1ec8_360);
and \U$1244 ( \1914 , \1541 , RIaaa1b80_353);
and \U$1245 ( \1915 , \1449 , RIaaa1bf8_354);
nor \U$1246 ( \1916 , \1914 , \1915 );
and \U$1247 ( \1917 , \1913 , \1916 );
nand \U$1248 ( \1918 , \1912 , \1917 );
nor \U$1249 ( \1919 , \1909 , \1918 );
buf \U$1250 ( \1920 , \1508 );
and \U$1251 ( \1921 , \1920 , RIaaa20a8_364);
and \U$1252 ( \1922 , \1502 , RIaaa1a90_351);
nor \U$1253 ( \1923 , \1921 , \1922 );
and \U$1254 ( \1924 , \1512 , RIaaa2120_365);
and \U$1255 ( \1925 , \1516 , RIaaa1dd8_358);
nor \U$1256 ( \1926 , \1924 , \1925 );
not \U$1257 ( \1927 , \1530 );
and \U$1258 ( \1928 , \1927 , RIaaa2198_366);
not \U$1259 ( \1929 , RIaaa1b08_352);
not \U$1260 ( \1930 , \1491 );
or \U$1261 ( \1931 , \1929 , \1930 );
nand \U$1262 ( \1932 , \1494 , RIaaa1a18_350);
nand \U$1263 ( \1933 , \1931 , \1932 );
nor \U$1264 ( \1934 , \1928 , \1933 );
and \U$1265 ( \1935 , \1923 , \1926 , \1934 );
nand \U$1266 ( \1936 , \1919 , \1935 );
buf \U$1267 ( \1937 , \1936 );
buf \U$1268 ( \1938 , \1937 );
or \U$1269 ( \1939 , \1901 , \1938 );
not \U$1270 ( \1940 , \1896 );
not \U$1271 ( \1941 , \1940 );
nand \U$1272 ( \1942 , \1941 , \1801 );
buf \U$1273 ( \1943 , \1942 );
not \U$1274 ( \1944 , \1943 );
not \U$1275 ( \1945 , \1561 );
not \U$1276 ( \1946 , RIaaa1130_331);
not \U$1277 ( \1947 , \1946 );
and \U$1278 ( \1948 , \1945 , \1947 );
and \U$1279 ( \1949 , \1502 , RIaaa0f50_327);
nor \U$1280 ( \1950 , \1948 , \1949 );
not \U$1281 ( \1951 , \1435 );
and \U$1282 ( \1952 , \1951 , RIaaa0a28_316);
and \U$1283 ( \1953 , \1411 , \1420 , \1387 );
and \U$1284 ( \1954 , \1953 , RIaaa0b90_319);
nor \U$1285 ( \1955 , \1952 , \1954 );
and \U$1286 ( \1956 , \1480 , RIaaa0b18_318);
not \U$1287 ( \1957 , RIaaa1040_329);
not \U$1288 ( \1958 , \1443 );
or \U$1289 ( \1959 , \1957 , \1958 );
not \U$1290 ( \1960 , \1448 );
nand \U$1291 ( \1961 , \1960 , RIaaa0c80_321);
nand \U$1292 ( \1962 , \1959 , \1961 );
nor \U$1293 ( \1963 , \1956 , \1962 );
nand \U$1294 ( \1964 , \1551 , RIaaa0cf8_322);
nand \U$1295 ( \1965 , \1950 , \1955 , \1963 , \1964 );
and \U$1296 ( \1966 , \1458 , RIaaa0c08_320);
and \U$1297 ( \1967 , \1463 , RIaaa0ed8_326);
nor \U$1298 ( \1968 , \1966 , \1967 );
nand \U$1299 ( \1969 , \1508 , RIaaa0d70_323);
and \U$1300 ( \1970 , \1516 , RIaaa0aa0_317);
not \U$1301 ( \1971 , RIaaa0fc8_328);
not \U$1302 ( \1972 , \1491 );
or \U$1303 ( \1973 , \1971 , \1972 );
not \U$1304 ( \1974 , RIaaa11a8_332);
nor \U$1305 ( \1975 , \1974 , \1495 );
not \U$1306 ( \1976 , \1975 );
nand \U$1307 ( \1977 , \1973 , \1976 );
nor \U$1308 ( \1978 , \1970 , \1977 );
nand \U$1309 ( \1979 , \1483 , RIaaa10b8_330);
and \U$1310 ( \1980 , \1969 , \1978 , \1979 );
and \U$1311 ( \1981 , \1470 , RIaaa0e60_325);
and \U$1312 ( \1982 , \1474 , RIaaa0de8_324);
nor \U$1313 ( \1983 , \1981 , \1982 );
nand \U$1314 ( \1984 , \1968 , \1980 , \1983 );
nor \U$1315 ( \1985 , \1965 , \1984 );
buf \U$1316 ( \1986 , \1985 );
not \U$1317 ( \1987 , \1986 );
not \U$1318 ( \1988 , \1987 );
not \U$1319 ( \1989 , \1988 );
and \U$1320 ( \1990 , \1944 , \1989 );
buf \U$1321 ( \1991 , \1889 );
and \U$1322 ( \1992 , \1801 , \1991 );
buf \U$1323 ( \1993 , \1992 );
not \U$1324 ( \1994 , \1985 );
not \U$1325 ( \1995 , \1994 );
not \U$1326 ( \1996 , \1995 );
not \U$1327 ( \1997 , \1996 );
and \U$1328 ( \1998 , \1993 , \1997 );
nor \U$1329 ( \1999 , \1990 , \1998 );
nand \U$1330 ( \2000 , \1939 , \1999 );
not \U$1331 ( \2001 , \1938 );
and \U$1332 ( \2002 , \1895 , \1897 );
not \U$1333 ( \2003 , \2002 );
nor \U$1334 ( \2004 , \2001 , \2003 );
nor \U$1335 ( \2005 , \2000 , \2004 );
not \U$1336 ( \2006 , \2005 );
and \U$1337 ( \2007 , \1596 , \2006 );
and \U$1338 ( \2008 , \1595 , \2005 );
nor \U$1339 ( \2009 , \2007 , \2008 );
not \U$1340 ( \2010 , \2009 );
not \U$1341 ( \2011 , \2010 );
and \U$1342 ( \2012 , \1824 , RIaa97680_1);
not \U$1343 ( \2013 , \2012 );
not \U$1344 ( \2014 , \1755 );
not \U$1345 ( \2015 , \2014 );
not \U$1346 ( \2016 , RIaa98508_32);
not \U$1347 ( \2017 , \2016 );
and \U$1348 ( \2018 , \2015 , \2017 );
not \U$1349 ( \2019 , RIaa98328_28);
buf \U$1350 ( \2020 , \1842 );
nor \U$1351 ( \2021 , \2019 , \2020 );
nor \U$1352 ( \2022 , \2018 , \2021 );
buf \U$1353 ( \2023 , \1626 );
and \U$1354 ( \2024 , \2023 , RIaa98238_26);
not \U$1355 ( \2025 , RIaa98418_30);
not \U$1356 ( \2026 , \1651 );
nor \U$1357 ( \2027 , \2025 , \2026 );
nor \U$1358 ( \2028 , \2024 , \2027 );
nand \U$1359 ( \2029 , \2022 , \2028 );
not \U$1360 ( \2030 , \1495 );
not \U$1361 ( \2031 , RIaa97e78_18);
not \U$1362 ( \2032 , \2031 );
and \U$1363 ( \2033 , \2030 , \2032 );
and \U$1364 ( \2034 , \1832 , RIaa981c0_25);
nor \U$1365 ( \2035 , \2033 , \2034 );
not \U$1366 ( \2036 , \1861 );
not \U$1367 ( \2037 , \2036 );
not \U$1368 ( \2038 , RIaa985f8_34);
not \U$1369 ( \2039 , \2038 );
and \U$1370 ( \2040 , \2037 , \2039 );
and \U$1371 ( \2041 , \1642 , RIaa982b0_27);
nor \U$1372 ( \2042 , \2040 , \2041 );
nand \U$1373 ( \2043 , \2035 , \2042 );
nor \U$1374 ( \2044 , \2029 , \2043 );
not \U$1375 ( \2045 , RIaa98580_33);
not \U$1376 ( \2046 , \1640 );
nor \U$1377 ( \2047 , \2045 , \2046 );
not \U$1378 ( \2048 , RIaa97ef0_19);
nor \U$1379 ( \2049 , \2048 , \1852 );
nor \U$1380 ( \2050 , \2047 , \2049 );
not \U$1381 ( \2051 , RIaa98058_22);
not \U$1382 ( \2052 , \1846 );
nor \U$1383 ( \2053 , \2051 , \2052 );
not \U$1384 ( \2054 , RIaa98148_24);
not \U$1385 ( \2055 , \1608 );
or \U$1386 ( \2056 , \2054 , \2055 );
nand \U$1387 ( \2057 , RIaa97d88_16, RIaa97f68_20);
nand \U$1388 ( \2058 , \2056 , \2057 );
nor \U$1389 ( \2059 , \2053 , \2058 );
nand \U$1390 ( \2060 , \2050 , \2059 );
buf \U$1391 ( \2061 , \1316 );
nand \U$1392 ( \2062 , \2061 , RIaa97fe0_21);
buf \U$1393 ( \2063 , \1735 );
not \U$1394 ( \2064 , \2063 );
nand \U$1395 ( \2065 , \2064 , RIaa983a0_29);
buf \U$1396 ( \2066 , \1682 );
nand \U$1397 ( \2067 , \2066 , RIaa980d0_23);
not \U$1398 ( \2068 , \1874 );
not \U$1399 ( \2069 , \2068 );
nand \U$1400 ( \2070 , \2069 , RIaa98490_31);
nand \U$1401 ( \2071 , \2062 , \2065 , \2067 , \2070 );
nor \U$1402 ( \2072 , \2060 , \2071 );
and \U$1403 ( \2073 , \2044 , \2072 );
not \U$1404 ( \2074 , \2073 );
not \U$1405 ( \2075 , \2074 );
xnor \U$1406 ( \2076 , \1824 , RIaa97680_1);
not \U$1407 ( \2077 , \2076 );
and \U$1408 ( \2078 , \2075 , \2077 );
not \U$1409 ( \2079 , \1826 );
nand \U$1410 ( \2080 , \2079 , \1879 );
not \U$1411 ( \2081 , \2080 );
not \U$1412 ( \2082 , \1818 );
or \U$1413 ( \2083 , \2081 , \2082 );
nand \U$1414 ( \2084 , \1880 , \1826 );
nand \U$1415 ( \2085 , \2083 , \2084 );
not \U$1416 ( \2086 , \2076 );
not \U$1417 ( \2087 , \2073 );
or \U$1418 ( \2088 , \2086 , \2087 );
or \U$1419 ( \2089 , \2073 , \2076 );
nand \U$1420 ( \2090 , \2088 , \2089 );
and \U$1421 ( \2091 , \2085 , \2090 );
nor \U$1422 ( \2092 , \2078 , \2091 );
xor \U$1423 ( \2093 , \2013 , \2092 );
not \U$1424 ( \2094 , \2085 );
nand \U$1425 ( \2095 , \2094 , \2090 );
not \U$1426 ( \2096 , \2090 );
nand \U$1427 ( \2097 , \2096 , \2085 );
nand \U$1428 ( \2098 , \2095 , \2097 );
xnor \U$1429 ( \2099 , \2093 , \2098 );
xnor \U$1430 ( \2100 , \2098 , \1991 );
nand \U$1431 ( \2101 , \2099 , \2100 );
not \U$1432 ( \2102 , \2101 );
buf \U$1433 ( \2103 , \2102 );
not \U$1434 ( \2104 , \2103 );
not \U$1435 ( \2105 , \2092 );
nor \U$1436 ( \2106 , \2105 , \2012 );
not \U$1437 ( \2107 , \2106 );
nand \U$1438 ( \2108 , \2105 , \2012 );
nand \U$1439 ( \2109 , \2107 , \2108 );
buf \U$1440 ( \2110 , \2109 );
not \U$1441 ( \2111 , \2110 );
buf \U$1442 ( \2112 , \1564 );
nand \U$1443 ( \2113 , \2112 , RIaaa2cd8_390);
and \U$1444 ( \2114 , \1516 , RIaaa2af8_386);
not \U$1445 ( \2115 , RIaaa3110_399);
not \U$1446 ( \2116 , \1491 );
or \U$1447 ( \2117 , \2115 , \2116 );
nand \U$1448 ( \2118 , \1494 , RIaaa3188_400);
nand \U$1449 ( \2119 , \2117 , \2118 );
nor \U$1450 ( \2120 , \2114 , \2119 );
nand \U$1451 ( \2121 , \1531 , RIaaa2f30_395);
and \U$1452 ( \2122 , \2113 , \2120 , \2121 );
and \U$1453 ( \2123 , \1458 , RIaaa2c60_389);
and \U$1454 ( \2124 , \1463 , RIaaa2eb8_394);
nor \U$1455 ( \2125 , \2123 , \2124 );
and \U$1456 ( \2126 , \1470 , RIaaa2dc8_392);
and \U$1457 ( \2127 , \1474 , RIaaa2e40_393);
nor \U$1458 ( \2128 , \2126 , \2127 );
nand \U$1459 ( \2129 , \2122 , \2125 , \2128 );
not \U$1460 ( \2130 , \1561 );
not \U$1461 ( \2131 , RIaaa2fa8_396);
not \U$1462 ( \2132 , \2131 );
and \U$1463 ( \2133 , \2130 , \2132 );
buf \U$1464 ( \2134 , \1502 );
and \U$1465 ( \2135 , \2134 , RIaaa3020_397);
nor \U$1466 ( \2136 , \2133 , \2135 );
and \U$1467 ( \2137 , \1413 , RIaaa2a08_384);
not \U$1468 ( \2138 , \1443 );
not \U$1469 ( \2139 , RIaaa3098_398);
or \U$1470 ( \2140 , \2138 , \2139 );
not \U$1471 ( \2141 , \1448 );
nand \U$1472 ( \2142 , \2141 , RIaaa2be8_388);
nand \U$1473 ( \2143 , \2140 , \2142 );
nor \U$1474 ( \2144 , \2137 , \2143 );
and \U$1475 ( \2145 , \1951 , RIaaa2b70_387);
and \U$1476 ( \2146 , \1480 , RIaaa2a80_385);
nor \U$1477 ( \2147 , \2145 , \2146 );
nand \U$1478 ( \2148 , \1551 , RIaaa2d50_391);
nand \U$1479 ( \2149 , \2136 , \2144 , \2147 , \2148 );
nor \U$1480 ( \2150 , \2129 , \2149 );
buf \U$1481 ( \2151 , \2150 );
not \U$1482 ( \2152 , \2151 );
not \U$1483 ( \2153 , \2152 );
buf \U$1484 ( \2154 , \2153 );
and \U$1485 ( \2155 , \2111 , \2154 );
not \U$1486 ( \2156 , \2111 );
and \U$1487 ( \2157 , \2156 , \2152 );
or \U$1488 ( \2158 , \2155 , \2157 );
nor \U$1489 ( \2159 , \2104 , \2158 );
buf \U$1490 ( \2160 , \2109 );
buf \U$1491 ( \2161 , \2160 );
not \U$1492 ( \2162 , \2161 );
not \U$1493 ( \2163 , \2100 );
buf \U$1494 ( \2164 , \2163 );
nand \U$1495 ( \2165 , \2162 , \2164 );
nand \U$1496 ( \2166 , \1502 , RIaaa1298_334);
nand \U$1497 ( \2167 , \1413 , RIaaa16d0_343);
nand \U$1498 ( \2168 , \1512 , RIaaa1928_348);
nand \U$1499 ( \2169 , \2166 , \2167 , \2168 );
nand \U$1500 ( \2170 , \1480 , RIaaa1658_342);
nand \U$1501 ( \2171 , \1550 , RIaaa1838_346);
nand \U$1502 ( \2172 , \1951 , RIaaa14f0_339);
not \U$1503 ( \2173 , \1442 );
buf \U$1504 ( \2174 , \2173 );
and \U$1505 ( \2175 , \2174 , RIaaa1388_336);
and \U$1506 ( \2176 , \1449 , RIaaa1400_337);
nor \U$1507 ( \2177 , \2175 , \2176 );
nand \U$1508 ( \2178 , \2170 , \2171 , \2172 , \2177 );
nor \U$1509 ( \2179 , \2169 , \2178 );
not \U$1510 ( \2180 , \1530 );
not \U$1511 ( \2181 , RIaaa19a0_349);
not \U$1512 ( \2182 , \2181 );
and \U$1513 ( \2183 , \2180 , \2182 );
and \U$1514 ( \2184 , \1474 , RIaaa1748_344);
nor \U$1515 ( \2185 , \2183 , \2184 );
and \U$1516 ( \2186 , \1516 , RIaaa15e0_341);
not \U$1517 ( \2187 , RIaaa1310_335);
not \U$1518 ( \2188 , \1491 );
or \U$1519 ( \2189 , \2187 , \2188 );
not \U$1520 ( \2190 , RIaaa1220_333);
nor \U$1521 ( \2191 , \2190 , \1495 );
not \U$1522 ( \2192 , \2191 );
nand \U$1523 ( \2193 , \2189 , \2192 );
nor \U$1524 ( \2194 , \2186 , \2193 );
nand \U$1525 ( \2195 , \2185 , \2194 );
not \U$1526 ( \2196 , RIaaa1478_338);
not \U$1527 ( \2197 , \1458 );
or \U$1528 ( \2198 , \2196 , \2197 );
not \U$1529 ( \2199 , \1460 );
nand \U$1530 ( \2200 , \2199 , RIaaa1568_340);
nand \U$1531 ( \2201 , \2198 , \2200 );
not \U$1532 ( \2202 , RIaaa17c0_345);
not \U$1533 ( \2203 , \1470 );
or \U$1534 ( \2204 , \2202 , \2203 );
nand \U$1535 ( \2205 , \1508 , RIaaa18b0_347);
nand \U$1536 ( \2206 , \2204 , \2205 );
nor \U$1537 ( \2207 , \2195 , \2201 , \2206 );
nand \U$1538 ( \2208 , \2179 , \2207 );
not \U$1539 ( \2209 , \2208 );
buf \U$1540 ( \2210 , \2209 );
or \U$1541 ( \2211 , \2165 , \2210 );
nand \U$1542 ( \2212 , \2163 , \2161 );
not \U$1543 ( \2213 , \2212 );
buf \U$1544 ( \2214 , \2210 );
nand \U$1545 ( \2215 , \2213 , \2214 );
nand \U$1546 ( \2216 , \2211 , \2215 );
nor \U$1547 ( \2217 , \2159 , \2216 );
buf \U$1548 ( \2218 , \2217 );
not \U$1549 ( \2219 , \2218 );
not \U$1550 ( \2220 , \2219 );
or \U$1551 ( \2221 , \2011 , \2220 );
not \U$1552 ( \2222 , \2218 );
not \U$1553 ( \2223 , \2009 );
or \U$1554 ( \2224 , \2222 , \2223 );
not \U$1555 ( \2225 , \2210 );
not \U$1556 ( \2226 , \2225 );
not \U$1557 ( \2227 , \2002 );
or \U$1558 ( \2228 , \2226 , \2227 );
and \U$1559 ( \2229 , \1900 , \2214 );
not \U$1560 ( \2230 , \1937 );
not \U$1561 ( \2231 , \2230 );
not \U$1562 ( \2232 , \1992 );
or \U$1563 ( \2233 , \2231 , \2232 );
not \U$1564 ( \2234 , \1800 );
and \U$1565 ( \2235 , \2234 , \1897 );
nand \U$1566 ( \2236 , \2235 , \1938 );
nand \U$1567 ( \2237 , \2233 , \2236 );
nor \U$1568 ( \2238 , \2229 , \2237 );
nand \U$1569 ( \2239 , \2228 , \2238 );
not \U$1570 ( \2240 , \2239 );
not \U$1571 ( \2241 , \1590 );
and \U$1572 ( \2242 , \1480 , RIaa9ff60_293);
not \U$1573 ( \2243 , RIaa9fba0_285);
not \U$1574 ( \2244 , \1502 );
or \U$1575 ( \2245 , \2243 , \2244 );
nand \U$1576 ( \2246 , \1512 , RIaa9fa38_282);
nand \U$1577 ( \2247 , \2245 , \2246 );
nor \U$1578 ( \2248 , \2242 , \2247 );
and \U$1579 ( \2249 , \1437 , RIaaa0050_295);
and \U$1580 ( \2250 , \1413 , RIaa9ffd8_294);
nor \U$1581 ( \2251 , \2249 , \2250 );
and \U$1582 ( \2252 , \1551 , RIaa9fe70_291);
and \U$1583 ( \2253 , RIaa9fc90_287, \1541 );
and \U$1584 ( \2254 , \1449 , RIaaa01b8_298);
nor \U$1585 ( \2255 , \2252 , \2253 , \2254 );
and \U$1586 ( \2256 , \2248 , \2251 , \2255 );
and \U$1587 ( \2257 , \1458 , RIaaa0140_297);
and \U$1588 ( \2258 , \1463 , RIaa9fdf8_290);
nor \U$1589 ( \2259 , \2257 , \2258 );
and \U$1590 ( \2260 , \1531 , RIaa9fab0_283);
not \U$1591 ( \2261 , RIaa9fc18_286);
not \U$1592 ( \2262 , \1491 );
or \U$1593 ( \2263 , \2261 , \2262 );
nand \U$1594 ( \2264 , \1494 , RIaa9fb28_284);
nand \U$1595 ( \2265 , \2263 , \2264 );
nor \U$1596 ( \2266 , \2260 , \2265 );
not \U$1597 ( \2267 , \2266 );
not \U$1598 ( \2268 , RIaa9fd08_288);
not \U$1599 ( \2269 , \1474 );
or \U$1600 ( \2270 , \2268 , \2269 );
nand \U$1601 ( \2271 , \1516 , RIaaa00c8_296);
nand \U$1602 ( \2272 , \2270 , \2271 );
nor \U$1603 ( \2273 , \2267 , \2272 );
and \U$1604 ( \2274 , \1920 , RIaa9fee8_292);
and \U$1605 ( \2275 , \1470 , RIaa9fd80_289);
nor \U$1606 ( \2276 , \2274 , \2275 );
and \U$1607 ( \2277 , \2259 , \2273 , \2276 );
nand \U$1608 ( \2278 , \2256 , \2277 );
not \U$1609 ( \2279 , \2278 );
buf \U$1610 ( \2280 , \2279 );
not \U$1611 ( \2281 , \2280 );
nand \U$1612 ( \2282 , \2241 , \2281 );
not \U$1613 ( \2283 , \2282 );
not \U$1614 ( \2284 , \2280 );
nor \U$1615 ( \2285 , \1575 , \1364 );
not \U$1616 ( \2286 , \2285 );
or \U$1617 ( \2287 , \2284 , \2286 );
buf \U$1618 ( \2288 , \1520 );
and \U$1619 ( \2289 , \2288 , \1583 );
not \U$1620 ( \2290 , \2288 );
not \U$1621 ( \2291 , \1576 );
and \U$1622 ( \2292 , \2290 , \2291 );
nor \U$1623 ( \2293 , \2289 , \2292 );
nand \U$1624 ( \2294 , \2287 , \2293 );
nor \U$1625 ( \2295 , \2283 , \2294 );
not \U$1626 ( \2296 , \1795 );
nand \U$1627 ( \2297 , \1711 , \1715 );
xor \U$1628 ( \2298 , \2297 , \1810 );
not \U$1629 ( \2299 , \2298 );
and \U$1630 ( \2300 , \2296 , \2299 );
and \U$1631 ( \2301 , \1795 , \2298 );
nor \U$1632 ( \2302 , \2300 , \2301 );
not \U$1633 ( \2303 , \1332 );
not \U$1634 ( \2304 , \2298 );
and \U$1635 ( \2305 , \2303 , \2304 );
and \U$1636 ( \2306 , \1332 , \2298 );
nor \U$1637 ( \2307 , \2305 , \2306 );
nand \U$1638 ( \2308 , \2302 , \2307 );
not \U$1639 ( \2309 , \2308 );
buf \U$1640 ( \2310 , \1795 );
nand \U$1641 ( \2311 , \2309 , \2310 );
not \U$1642 ( \2312 , \2311 );
nand \U$1643 ( \2313 , \2312 , \1987 );
not \U$1644 ( \2314 , \2313 );
not \U$1645 ( \2315 , \1995 );
buf \U$1646 ( \2316 , \2308 );
buf \U$1647 ( \2317 , \2310 );
nor \U$1648 ( \2318 , \2316 , \2317 );
not \U$1649 ( \2319 , \2318 );
or \U$1650 ( \2320 , \2315 , \2319 );
not \U$1651 ( \2321 , RIaaa05f0_307);
not \U$1652 ( \2322 , \1413 );
or \U$1653 ( \2323 , \2321 , \2322 );
and \U$1654 ( \2324 , \1512 , RIaaa0938_314);
and \U$1655 ( \2325 , \2134 , RIaaa0758_310);
nor \U$1656 ( \2326 , \2324 , \2325 );
nand \U$1657 ( \2327 , \2323 , \2326 );
and \U$1658 ( \2328 , \1437 , RIaaa0488_304);
and \U$1659 ( \2329 , \1480 , RIaaa0578_306);
nor \U$1660 ( \2330 , \2328 , \2329 );
and \U$1661 ( \2331 , \1551 , RIaaa0230_299);
not \U$1662 ( \2332 , RIaaa06e0_309);
not \U$1663 ( \2333 , \1960 );
or \U$1664 ( \2334 , \2332 , \2333 );
nand \U$1665 ( \2335 , \1443 , RIaaa0848_312);
nand \U$1666 ( \2336 , \2334 , \2335 );
nor \U$1667 ( \2337 , \2331 , \2336 );
nand \U$1668 ( \2338 , \2330 , \2337 );
nor \U$1669 ( \2339 , \2327 , \2338 );
and \U$1670 ( \2340 , \1470 , RIaaa0398_302);
and \U$1671 ( \2341 , \1474 , RIaaa0320_301);
nor \U$1672 ( \2342 , \2340 , \2341 );
nand \U$1673 ( \2343 , \1458 , RIaaa0668_308);
buf \U$1674 ( \2344 , \1461 );
nand \U$1675 ( \2345 , \2344 , RIaaa0410_303);
nand \U$1676 ( \2346 , \2342 , \2343 , \2345 );
and \U$1677 ( \2347 , \2112 , RIaaa02a8_300);
and \U$1678 ( \2348 , \1531 , RIaaa08c0_313);
nor \U$1679 ( \2349 , \2347 , \2348 );
and \U$1680 ( \2350 , \1516 , RIaaa0500_305);
not \U$1681 ( \2351 , RIaaa07d0_311);
not \U$1682 ( \2352 , \1491 );
or \U$1683 ( \2353 , \2351 , \2352 );
nand \U$1684 ( \2354 , \1494 , RIaaa09b0_315);
nand \U$1685 ( \2355 , \2353 , \2354 );
nor \U$1686 ( \2356 , \2350 , \2355 );
nand \U$1687 ( \2357 , \2349 , \2356 );
nor \U$1688 ( \2358 , \2346 , \2357 );
nand \U$1689 ( \2359 , \2339 , \2358 );
not \U$1690 ( \2360 , \2359 );
not \U$1691 ( \2361 , \2310 );
or \U$1692 ( \2362 , \2360 , \2361 );
buf \U$1693 ( \2363 , \2359 );
or \U$1694 ( \2364 , \2317 , \2363 );
nand \U$1695 ( \2365 , \2362 , \2364 );
not \U$1696 ( \2366 , \2307 );
buf \U$1697 ( \2367 , \2366 );
nand \U$1698 ( \2368 , \2365 , \2367 );
nand \U$1699 ( \2369 , \2320 , \2368 );
nor \U$1700 ( \2370 , \2314 , \2369 );
and \U$1701 ( \2371 , \2295 , \2370 );
not \U$1702 ( \2372 , \2295 );
not \U$1703 ( \2373 , \2370 );
and \U$1704 ( \2374 , \2372 , \2373 );
nor \U$1705 ( \2375 , \2371 , \2374 );
not \U$1706 ( \2376 , \2375 );
or \U$1707 ( \2377 , \2240 , \2376 );
not \U$1708 ( \2378 , \2282 );
or \U$1709 ( \2379 , \2294 , \2378 );
not \U$1710 ( \2380 , \2313 );
or \U$1711 ( \2381 , \2369 , \2380 );
nand \U$1712 ( \2382 , \2379 , \2381 );
nand \U$1713 ( \2383 , \2377 , \2382 );
buf \U$1714 ( \2384 , \2383 );
nand \U$1715 ( \2385 , \2224 , \2384 );
nand \U$1716 ( \2386 , \2221 , \2385 );
not \U$1717 ( \2387 , \2386 );
nor \U$1718 ( \2388 , \2316 , \2317 );
not \U$1719 ( \2389 , \2388 );
not \U$1720 ( \2390 , \2389 );
not \U$1721 ( \2391 , \2279 );
buf \U$1722 ( \2392 , \2391 );
not \U$1723 ( \2393 , \2392 );
and \U$1724 ( \2394 , \2390 , \2393 );
nand \U$1725 ( \2395 , \2366 , \2310 );
buf \U$1726 ( \2396 , \2395 );
or \U$1727 ( \2397 , \2396 , \1522 );
not \U$1728 ( \2398 , \2310 );
nand \U$1729 ( \2399 , \2398 , \2366 );
buf \U$1730 ( \2400 , \2399 );
not \U$1731 ( \2401 , \1522 );
or \U$1732 ( \2402 , \2400 , \2401 );
nand \U$1733 ( \2403 , \2397 , \2402 );
nor \U$1734 ( \2404 , \2394 , \2403 );
buf \U$1735 ( \2405 , \2311 );
not \U$1736 ( \2406 , \2405 );
nand \U$1737 ( \2407 , \2406 , \2392 );
nand \U$1738 ( \2408 , \2404 , \2407 );
not \U$1739 ( \2409 , \2408 );
buf \U$1740 ( \2410 , \1996 );
nand \U$1741 ( \2411 , \2002 , \2410 );
not \U$1742 ( \2412 , \2411 );
not \U$1743 ( \2413 , \1900 );
not \U$1744 ( \2414 , \1997 );
or \U$1745 ( \2415 , \2413 , \2414 );
not \U$1746 ( \2416 , \2363 );
and \U$1747 ( \2417 , \1993 , \2416 );
nor \U$1748 ( \2418 , \1942 , \2416 );
nor \U$1749 ( \2419 , \2417 , \2418 );
nand \U$1750 ( \2420 , \2415 , \2419 );
nor \U$1751 ( \2421 , \2412 , \2420 );
not \U$1752 ( \2422 , \2421 );
or \U$1753 ( \2423 , \2409 , \2422 );
not \U$1754 ( \2424 , \2411 );
not \U$1755 ( \2425 , \2420 );
not \U$1756 ( \2426 , \2425 );
or \U$1757 ( \2427 , \2424 , \2426 );
not \U$1758 ( \2428 , \2408 );
nand \U$1759 ( \2429 , \2427 , \2428 );
nand \U$1760 ( \2430 , \2423 , \2429 );
buf \U$1761 ( \2431 , \2430 );
buf \U$1762 ( \2432 , \2160 );
not \U$1763 ( \2433 , \2432 );
not \U$1764 ( \2434 , \2433 );
nand \U$1765 ( \2435 , \2434 , \2103 );
nor \U$1766 ( \2436 , \2435 , \2225 );
not \U$1767 ( \2437 , \2436 );
not \U$1768 ( \2438 , \2165 );
and \U$1769 ( \2439 , \2438 , \1938 );
nor \U$1770 ( \2440 , \2212 , \1938 );
nor \U$1771 ( \2441 , \2439 , \2440 );
not \U$1772 ( \2442 , \2101 );
and \U$1773 ( \2443 , \2442 , \2433 );
nand \U$1774 ( \2444 , \2443 , \2225 );
nand \U$1775 ( \2445 , \2437 , \2441 , \2444 );
xor \U$1776 ( \2446 , \2431 , \2445 );
buf \U$1777 ( \2447 , \2108 );
not \U$1778 ( \2448 , \2447 );
nand \U$1779 ( \2449 , \1413 , RIaaa24e0_373);
nand \U$1780 ( \2450 , \1436 , RIaaa2558_374);
and \U$1781 ( \2451 , \2449 , \2450 );
not \U$1782 ( \2452 , \1561 );
not \U$1783 ( \2453 , RIaaa2738_378);
not \U$1784 ( \2454 , \2453 );
and \U$1785 ( \2455 , \2452 , \2454 );
and \U$1786 ( \2456 , \2134 , RIaaa2828_380);
nor \U$1787 ( \2457 , \2455 , \2456 );
and \U$1788 ( \2458 , \1551 , RIaaa2300_369);
not \U$1789 ( \2459 , RIaaa26c0_377);
not \U$1790 ( \2460 , \1960 );
or \U$1791 ( \2461 , \2459 , \2460 );
nand \U$1792 ( \2462 , \2174 , RIaaa2918_382);
nand \U$1793 ( \2463 , \2461 , \2462 );
nor \U$1794 ( \2464 , \2458 , \2463 );
nand \U$1795 ( \2465 , \1480 , RIaaa2468_372);
nand \U$1796 ( \2466 , \2451 , \2457 , \2464 , \2465 );
and \U$1797 ( \2467 , \1920 , RIaaa2378_370);
and \U$1798 ( \2468 , \1474 , RIaaa2288_368);
nor \U$1799 ( \2469 , \2467 , \2468 );
and \U$1800 ( \2470 , \1458 , RIaaa2648_376);
and \U$1801 ( \2471 , \2344 , RIaaa23f0_371);
nor \U$1802 ( \2472 , \2470 , \2471 );
and \U$1803 ( \2473 , \1470 , RIaaa2210_367);
and \U$1804 ( \2474 , \1516 , RIaaa25d0_375);
nor \U$1805 ( \2475 , \2473 , \2474 );
and \U$1806 ( \2476 , \1927 , RIaaa27b0_379);
not \U$1807 ( \2477 , RIaaa28a0_381);
not \U$1808 ( \2478 , \1491 );
or \U$1809 ( \2479 , \2477 , \2478 );
nand \U$1810 ( \2480 , \1494 , RIaaa2990_383);
nand \U$1811 ( \2481 , \2479 , \2480 );
nor \U$1812 ( \2482 , \2476 , \2481 );
nand \U$1813 ( \2483 , \2469 , \2472 , \2475 , \2482 );
nor \U$1814 ( \2484 , \2466 , \2483 );
not \U$1815 ( \2485 , \2484 );
buf \U$1816 ( \2486 , \2485 );
nand \U$1817 ( \2487 , \2448 , \2486 );
not \U$1818 ( \2488 , \2487 );
not \U$1819 ( \2489 , \2405 );
not \U$1820 ( \2490 , \2416 );
and \U$1821 ( \2491 , \2489 , \2490 );
not \U$1822 ( \2492 , \2416 );
not \U$1823 ( \2493 , \2390 );
or \U$1824 ( \2494 , \2492 , \2493 );
not \U$1825 ( \2495 , \2399 );
and \U$1826 ( \2496 , \2280 , \2495 );
not \U$1827 ( \2497 , \2280 );
not \U$1828 ( \2498 , \2396 );
and \U$1829 ( \2499 , \2497 , \2498 );
nor \U$1830 ( \2500 , \2496 , \2499 );
nand \U$1831 ( \2501 , \2494 , \2500 );
nor \U$1832 ( \2502 , \2491 , \2501 );
not \U$1833 ( \2503 , \2502 );
or \U$1834 ( \2504 , \2488 , \2503 );
not \U$1835 ( \2505 , \1573 );
not \U$1836 ( \2506 , \1186 );
nand \U$1837 ( \2507 , \2506 , \1193 );
not \U$1838 ( \2508 , \2507 );
buf \U$1839 ( \2509 , \2508 );
not \U$1840 ( \2510 , \2509 );
or \U$1841 ( \2511 , \2505 , \2510 );
not \U$1842 ( \2512 , \1185 );
buf \U$1843 ( \2513 , \1183 );
nand \U$1844 ( \2514 , \2512 , \2513 );
not \U$1845 ( \2515 , \2514 );
buf \U$1846 ( \2516 , \2515 );
not \U$1847 ( \2517 , \1573 );
and \U$1848 ( \2518 , \2516 , \2517 );
not \U$1849 ( \2519 , \1142 );
nand \U$1850 ( \2520 , \2519 , \1189 );
not \U$1851 ( \2521 , \2520 );
nor \U$1852 ( \2522 , \2518 , \2521 );
nand \U$1853 ( \2523 , \2511 , \2522 );
nand \U$1854 ( \2524 , \2504 , \2523 );
not \U$1855 ( \2525 , \2524 );
nand \U$1856 ( \2526 , \2446 , \2525 );
and \U$1857 ( \2527 , \2387 , \2526 );
nor \U$1858 ( \2528 , \2446 , \2525 );
nor \U$1859 ( \2529 , \2527 , \2528 );
not \U$1860 ( \2530 , \2529 );
buf \U$1861 ( \2531 , \1364 );
not \U$1862 ( \2532 , \2531 );
buf \U$1863 ( \2533 , \1582 );
not \U$1864 ( \2534 , \2533 );
not \U$1865 ( \2535 , \2534 );
or \U$1866 ( \2536 , \2532 , \2535 );
buf \U$1867 ( \2537 , \1363 );
not \U$1868 ( \2538 , \1335 );
and \U$1869 ( \2539 , \2537 , \2538 , \1573 );
and \U$1870 ( \2540 , \1335 , \2517 );
nor \U$1871 ( \2541 , \2539 , \2540 );
nand \U$1872 ( \2542 , \2536 , \2541 );
not \U$1873 ( \2543 , \2542 );
buf \U$1874 ( \2544 , \2005 );
and \U$1875 ( \2545 , \1194 , \1594 );
or \U$1876 ( \2546 , \2544 , \2545 );
or \U$1877 ( \2547 , \1594 , \1194 );
nand \U$1878 ( \2548 , \2546 , \2547 );
not \U$1879 ( \2549 , \2548 );
or \U$1880 ( \2550 , \2543 , \2549 );
not \U$1881 ( \2551 , \2154 );
nand \U$1882 ( \2552 , \2448 , \2551 );
nand \U$1883 ( \2553 , \2550 , \2552 );
not \U$1884 ( \2554 , \2553 );
not \U$1885 ( \2555 , \2416 );
not \U$1886 ( \2556 , \1901 );
not \U$1887 ( \2557 , \2556 );
or \U$1888 ( \2558 , \2555 , \2557 );
and \U$1889 ( \2559 , \1993 , \2393 );
nor \U$1890 ( \2560 , \1943 , \2393 );
nor \U$1891 ( \2561 , \2559 , \2560 );
nand \U$1892 ( \2562 , \2558 , \2561 );
buf \U$1893 ( \2563 , \2002 );
not \U$1894 ( \2564 , \2563 );
nor \U$1895 ( \2565 , \2564 , \2416 );
nor \U$1896 ( \2566 , \2562 , \2565 );
not \U$1897 ( \2567 , \2566 );
not \U$1898 ( \2568 , \2537 );
not \U$1899 ( \2569 , \2531 );
or \U$1900 ( \2570 , \2568 , \2569 );
nand \U$1901 ( \2571 , \2570 , \2538 );
nor \U$1902 ( \2572 , \2316 , \2317 );
not \U$1903 ( \2573 , \2572 );
not \U$1904 ( \2574 , \2573 );
and \U$1905 ( \2575 , \2574 , \1522 );
not \U$1906 ( \2576 , \1572 );
and \U$1907 ( \2577 , \2576 , \2396 );
not \U$1908 ( \2578 , \2576 );
and \U$1909 ( \2579 , \2578 , \2400 );
nor \U$1910 ( \2580 , \2577 , \2579 );
nor \U$1911 ( \2581 , \2575 , \2580 );
not \U$1912 ( \2582 , \2311 );
buf \U$1913 ( \2583 , \2582 );
nand \U$1914 ( \2584 , \2583 , \2401 );
nand \U$1915 ( \2585 , \2581 , \2584 );
xor \U$1916 ( \2586 , \2571 , \2585 );
not \U$1917 ( \2587 , \2586 );
and \U$1918 ( \2588 , \2567 , \2587 );
and \U$1919 ( \2589 , \2586 , \2566 );
nor \U$1920 ( \2590 , \2588 , \2589 );
and \U$1921 ( \2591 , \2443 , \1938 );
nor \U$1922 ( \2592 , \2435 , \1938 );
nor \U$1923 ( \2593 , \2591 , \2592 );
and \U$1924 ( \2594 , \2410 , \2438 );
not \U$1925 ( \2595 , \2410 );
not \U$1926 ( \2596 , \2212 );
and \U$1927 ( \2597 , \2595 , \2596 );
nor \U$1928 ( \2598 , \2594 , \2597 );
nand \U$1929 ( \2599 , \2593 , \2598 );
not \U$1930 ( \2600 , \2225 );
not \U$1931 ( \2601 , \2448 );
or \U$1932 ( \2602 , \2600 , \2601 );
nand \U$1933 ( \2603 , \2602 , \2542 );
or \U$1934 ( \2604 , \2599 , \2603 );
nand \U$1935 ( \2605 , \2599 , \2603 );
nand \U$1936 ( \2606 , \2604 , \2605 );
xor \U$1937 ( \2607 , \2590 , \2606 );
not \U$1938 ( \2608 , \2421 );
not \U$1939 ( \2609 , \2428 );
and \U$1940 ( \2610 , \2608 , \2609 );
and \U$1941 ( \2611 , \2445 , \2431 );
nor \U$1942 ( \2612 , \2610 , \2611 );
xor \U$1943 ( \2613 , \2607 , \2612 );
not \U$1944 ( \2614 , \2613 );
or \U$1945 ( \2615 , \2554 , \2614 );
or \U$1946 ( \2616 , \2613 , \2553 );
nand \U$1947 ( \2617 , \2615 , \2616 );
not \U$1948 ( \2618 , \2617 );
or \U$1949 ( \2619 , \2530 , \2618 );
or \U$1950 ( \2620 , \2529 , \2617 );
nand \U$1951 ( \2621 , \2619 , \2620 );
and \U$1952 ( \2622 , \2542 , \2552 );
xor \U$1953 ( \2623 , \2548 , \2622 );
not \U$1954 ( \2624 , \2623 );
xor \U$1955 ( \2625 , \2524 , \2430 );
xor \U$1956 ( \2626 , \2625 , \2445 );
and \U$1957 ( \2627 , \2626 , \2386 );
not \U$1958 ( \2628 , \2626 );
and \U$1959 ( \2629 , \2628 , \2387 );
nor \U$1960 ( \2630 , \2627 , \2629 );
not \U$1961 ( \2631 , \2630 );
or \U$1962 ( \2632 , \2624 , \2631 );
or \U$1963 ( \2633 , \2623 , \2630 );
nand \U$1964 ( \2634 , \2632 , \2633 );
not \U$1965 ( \2635 , \2523 );
not \U$1966 ( \2636 , \2635 );
not \U$1967 ( \2637 , \2154 );
nand \U$1968 ( \2638 , \2637 , \2438 );
not \U$1969 ( \2639 , \2486 );
buf \U$1970 ( \2640 , \2160 );
and \U$1971 ( \2641 , \2639 , \2640 );
not \U$1972 ( \2642 , \2639 );
and \U$1973 ( \2643 , \2642 , \2111 );
or \U$1974 ( \2644 , \2641 , \2643 );
nand \U$1975 ( \2645 , \2103 , \2644 );
nand \U$1976 ( \2646 , \2596 , \2154 );
nand \U$1977 ( \2647 , \2638 , \2645 , \2646 );
not \U$1978 ( \2648 , \2647 );
or \U$1979 ( \2649 , \2636 , \2648 );
and \U$1980 ( \2650 , \1458 , RIaaa3f20_429);
and \U$1981 ( \2651 , \2344 , RIaaa3f98_430);
nor \U$1982 ( \2652 , \2650 , \2651 );
not \U$1983 ( \2653 , RIaaa3cc8_424);
not \U$1984 ( \2654 , \1474 );
or \U$1985 ( \2655 , \2653 , \2654 );
nand \U$1986 ( \2656 , \1531 , RIaaa3c50_423);
nand \U$1987 ( \2657 , \2655 , \2656 );
not \U$1988 ( \2658 , RIaaa4010_431);
not \U$1989 ( \2659 , \1516 );
or \U$1990 ( \2660 , \2658 , \2659 );
and \U$1991 ( \2661 , \1491 , RIaaa4100_433);
nand \U$1992 ( \2662 , \1494 , RIaaa3db8_426);
not \U$1993 ( \2663 , \2662 );
nor \U$1994 ( \2664 , \2661 , \2663 );
nand \U$1995 ( \2665 , \2660 , \2664 );
nor \U$1996 ( \2666 , \2657 , \2665 );
and \U$1997 ( \2667 , \1566 , RIaaa3b60_421);
and \U$1998 ( \2668 , \1470 , RIaaa3d40_425);
nor \U$1999 ( \2669 , \2667 , \2668 );
and \U$2000 ( \2670 , \2652 , \2666 , \2669 );
and \U$2001 ( \2671 , \1551 , RIaaa3ae8_420);
and \U$2002 ( \2672 , \1413 , RIaaa3a70_419);
nor \U$2003 ( \2673 , \2671 , \2672 );
and \U$2004 ( \2674 , \1480 , RIaaa39f8_418);
and \U$2005 ( \2675 , \2174 , RIaaa4178_434);
and \U$2006 ( \2676 , \1960 , RIaaa3e30_427);
nor \U$2007 ( \2677 , \2674 , \2675 , \2676 );
nand \U$2008 ( \2678 , \2673 , \2677 );
not \U$2009 ( \2679 , \1561 );
not \U$2010 ( \2680 , RIaaa3bd8_422);
not \U$2011 ( \2681 , \2680 );
and \U$2012 ( \2682 , \2679 , \2681 );
and \U$2013 ( \2683 , \1502 , RIaaa4088_432);
nor \U$2014 ( \2684 , \2682 , \2683 );
nand \U$2015 ( \2685 , \1951 , RIaaa3ea8_428);
nand \U$2016 ( \2686 , \2684 , \2685 );
nor \U$2017 ( \2687 , \2678 , \2686 );
nand \U$2018 ( \2688 , \2670 , \2687 );
buf \U$2019 ( \2689 , \2688 );
not \U$2020 ( \2690 , \2689 );
not \U$2021 ( \2691 , \2690 );
and \U$2022 ( \2692 , \2448 , \2691 );
not \U$2023 ( \2693 , \2692 );
nand \U$2024 ( \2694 , \2649 , \2693 );
and \U$2025 ( \2695 , \2502 , \2523 );
not \U$2026 ( \2696 , \2502 );
and \U$2027 ( \2697 , \2696 , \2635 );
nor \U$2028 ( \2698 , \2695 , \2697 );
nand \U$2029 ( \2699 , \2698 , \2487 );
nand \U$2030 ( \2700 , \2694 , \2699 );
not \U$2031 ( \2701 , \2700 );
xor \U$2032 ( \2702 , \2217 , \2383 );
xnor \U$2033 ( \2703 , \2702 , \2009 );
not \U$2034 ( \2704 , \2703 );
or \U$2035 ( \2705 , \2701 , \2704 );
not \U$2036 ( \2706 , \2694 );
not \U$2037 ( \2707 , \2699 );
nand \U$2038 ( \2708 , \2706 , \2707 );
nand \U$2039 ( \2709 , \2705 , \2708 );
nand \U$2040 ( \2710 , \2634 , \2709 );
not \U$2041 ( \2711 , \2623 );
nand \U$2042 ( \2712 , \2711 , \2630 );
nand \U$2043 ( \2713 , \2710 , \2712 );
nand \U$2044 ( \2714 , \2621 , \2713 );
not \U$2045 ( \2715 , \2709 );
not \U$2046 ( \2716 , \2634 );
not \U$2047 ( \2717 , \2716 );
or \U$2048 ( \2718 , \2715 , \2717 );
not \U$2049 ( \2719 , \2709 );
nand \U$2050 ( \2720 , \2719 , \2634 );
nand \U$2051 ( \2721 , \2718 , \2720 );
buf \U$2052 ( \2722 , \1062 );
xor \U$2053 ( \2723 , \852 , \2722 );
not \U$2054 ( \2724 , \1059 );
xnor \U$2055 ( \2725 , \2723 , \2724 );
not \U$2056 ( \2726 , \2725 );
not \U$2057 ( \2727 , \849 );
buf \U$2058 ( \2728 , \1014 );
not \U$2059 ( \2729 , \2728 );
or \U$2060 ( \2730 , \2727 , \2729 );
buf \U$2061 ( \2731 , \1057 );
nand \U$2062 ( \2732 , \2730 , \2731 );
buf \U$2063 ( \2733 , \1154 );
not \U$2064 ( \2734 , \2733 );
and \U$2065 ( \2735 , \2732 , \2734 );
not \U$2066 ( \2736 , \2732 );
and \U$2067 ( \2737 , \2736 , \2733 );
nor \U$2068 ( \2738 , \2735 , \2737 );
not \U$2069 ( \2739 , \2738 );
or \U$2070 ( \2740 , \2726 , \2739 );
or \U$2071 ( \2741 , \2725 , \2738 );
nand \U$2072 ( \2742 , \2740 , \2741 );
not \U$2073 ( \2743 , \1172 );
not \U$2074 ( \2744 , \2725 );
and \U$2075 ( \2745 , \2743 , \2744 );
not \U$2076 ( \2746 , \2743 );
and \U$2077 ( \2747 , \2746 , \2725 );
nor \U$2078 ( \2748 , \2745 , \2747 );
nand \U$2079 ( \2749 , \2742 , \2748 );
buf \U$2080 ( \2750 , \2749 );
buf \U$2081 ( \2751 , \2750 );
not \U$2082 ( \2752 , \2751 );
buf \U$2083 ( \2753 , \1172 );
nor \U$2084 ( \2754 , \2742 , \2753 );
not \U$2085 ( \2755 , \2754 );
not \U$2086 ( \2756 , \2755 );
or \U$2087 ( \2757 , \2752 , \2756 );
buf \U$2088 ( \2758 , \2753 );
not \U$2089 ( \2759 , \2758 );
not \U$2090 ( \2760 , \2759 );
not \U$2091 ( \2761 , \2576 );
and \U$2092 ( \2762 , \2760 , \2761 );
not \U$2093 ( \2763 , \2725 );
not \U$2094 ( \2764 , \2738 );
or \U$2095 ( \2765 , \2763 , \2764 );
not \U$2096 ( \2766 , \2744 );
not \U$2097 ( \2767 , \2738 );
not \U$2098 ( \2768 , \2767 );
or \U$2099 ( \2769 , \2766 , \2768 );
nand \U$2100 ( \2770 , \2765 , \2769 );
buf \U$2101 ( \2771 , \2770 );
buf \U$2102 ( \2772 , \2771 );
nor \U$2103 ( \2773 , \1572 , \2758 );
and \U$2104 ( \2774 , \2772 , \2773 );
nor \U$2105 ( \2775 , \2762 , \2774 );
nand \U$2106 ( \2776 , \2757 , \2775 );
not \U$2107 ( \2777 , \2776 );
not \U$2108 ( \2778 , \1938 );
not \U$2109 ( \2779 , \2583 );
or \U$2110 ( \2780 , \2778 , \2779 );
and \U$2111 ( \2781 , \2390 , \2001 );
and \U$2112 ( \2782 , \1996 , \2396 );
not \U$2113 ( \2783 , \1996 );
and \U$2114 ( \2784 , \2783 , \2400 );
nor \U$2115 ( \2785 , \2782 , \2784 );
nor \U$2116 ( \2786 , \2781 , \2785 );
nand \U$2117 ( \2787 , \2780 , \2786 );
xor \U$2118 ( \2788 , \2777 , \2787 );
not \U$2119 ( \2789 , \2551 );
not \U$2120 ( \2790 , \2563 );
or \U$2121 ( \2791 , \2789 , \2790 );
and \U$2122 ( \2792 , \2556 , \2154 );
and \U$2123 ( \2793 , \1993 , \2214 );
and \U$2124 ( \2794 , \2235 , \2225 );
nor \U$2125 ( \2795 , \2792 , \2793 , \2794 );
nand \U$2126 ( \2796 , \2791 , \2795 );
and \U$2127 ( \2797 , \2788 , \2796 );
and \U$2128 ( \2798 , \2777 , \2787 );
or \U$2129 ( \2799 , \2797 , \2798 );
not \U$2130 ( \2800 , \2799 );
buf \U$2131 ( \2801 , \1366 );
not \U$2132 ( \2802 , \2801 );
and \U$2133 ( \2803 , \2802 , \2416 );
buf \U$2134 ( \2804 , \2291 );
not \U$2135 ( \2805 , \2804 );
not \U$2136 ( \2806 , \2391 );
or \U$2137 ( \2807 , \2805 , \2806 );
not \U$2138 ( \2808 , \1584 );
or \U$2139 ( \2809 , \2808 , \2392 );
nand \U$2140 ( \2810 , \2807 , \2809 );
nor \U$2141 ( \2811 , \2803 , \2810 );
buf \U$2142 ( \2812 , \1591 );
not \U$2143 ( \2813 , \2416 );
nand \U$2144 ( \2814 , \2812 , \2813 );
nand \U$2145 ( \2815 , \2811 , \2814 );
not \U$2146 ( \2816 , \2815 );
nand \U$2147 ( \2817 , \2750 , \2771 );
and \U$2148 ( \2818 , \2817 , \2759 );
not \U$2149 ( \2819 , \2401 );
not \U$2150 ( \2820 , \2509 );
or \U$2151 ( \2821 , \2819 , \2820 );
not \U$2152 ( \2822 , \2514 );
buf \U$2153 ( \2823 , \2822 );
and \U$2154 ( \2824 , \2823 , \1522 );
not \U$2155 ( \2825 , \1571 );
not \U$2156 ( \2826 , \1142 );
not \U$2157 ( \2827 , \1189 );
nor \U$2158 ( \2828 , \2826 , \2827 );
not \U$2159 ( \2829 , \2828 );
not \U$2160 ( \2830 , \2829 );
not \U$2161 ( \2831 , \2830 );
or \U$2162 ( \2832 , \2825 , \2831 );
not \U$2163 ( \2833 , \2521 );
or \U$2164 ( \2834 , \2833 , \2576 );
nand \U$2165 ( \2835 , \2832 , \2834 );
nor \U$2166 ( \2836 , \2824 , \2835 );
nand \U$2167 ( \2837 , \2821 , \2836 );
xnor \U$2168 ( \2838 , \2818 , \2837 );
not \U$2169 ( \2839 , \2838 );
or \U$2170 ( \2840 , \2816 , \2839 );
not \U$2171 ( \2841 , \2818 );
nand \U$2172 ( \2842 , \2841 , \2837 );
nand \U$2173 ( \2843 , \2840 , \2842 );
and \U$2174 ( \2844 , \2375 , \2239 );
not \U$2175 ( \2845 , \2375 );
not \U$2176 ( \2846 , \2239 );
and \U$2177 ( \2847 , \2845 , \2846 );
nor \U$2178 ( \2848 , \2844 , \2847 );
xor \U$2179 ( \2849 , \2843 , \2848 );
not \U$2180 ( \2850 , \2849 );
nor \U$2181 ( \2851 , \2800 , \2850 );
and \U$2182 ( \2852 , \2843 , \2848 );
nor \U$2183 ( \2853 , \2851 , \2852 );
not \U$2184 ( \2854 , \2703 );
not \U$2185 ( \2855 , \2699 );
not \U$2186 ( \2856 , \2706 );
or \U$2187 ( \2857 , \2855 , \2856 );
nand \U$2188 ( \2858 , \2694 , \2707 );
nand \U$2189 ( \2859 , \2857 , \2858 );
not \U$2190 ( \2860 , \2859 );
and \U$2191 ( \2861 , \2854 , \2860 );
and \U$2192 ( \2862 , \2703 , \2859 );
nor \U$2193 ( \2863 , \2861 , \2862 );
xor \U$2194 ( \2864 , \2853 , \2863 );
not \U$2195 ( \2865 , \2799 );
not \U$2196 ( \2866 , \2849 );
not \U$2197 ( \2867 , \2866 );
or \U$2198 ( \2868 , \2865 , \2867 );
or \U$2199 ( \2869 , \2850 , \2799 );
nand \U$2200 ( \2870 , \2868 , \2869 );
and \U$2201 ( \2871 , \1951 , RIaaa32f0_403);
and \U$2202 ( \2872 , \1413 , RIaaa3890_415);
nor \U$2203 ( \2873 , \2871 , \2872 );
and \U$2204 ( \2874 , RIaaa34d0_407, \1502 );
and \U$2205 ( \2875 , \1512 , RIaaa3638_410);
not \U$2206 ( \2876 , RIaaa3728_412);
nor \U$2207 ( \2877 , \2876 , \1426 );
nor \U$2208 ( \2878 , \2874 , \2875 , \2877 );
and \U$2209 ( \2879 , \1541 , RIaaa35c0_409);
not \U$2210 ( \2880 , \1419 );
and \U$2211 ( \2881 , \1440 , \2880 , \1410 );
and \U$2212 ( \2882 , \2881 , RIaaa3278_402);
nor \U$2213 ( \2883 , \2879 , \2882 );
nand \U$2214 ( \2884 , \1480 , RIaaa3818_414);
and \U$2215 ( \2885 , \2883 , \2884 );
nand \U$2216 ( \2886 , \2873 , \2878 , \2885 );
and \U$2217 ( \2887 , \2199 , RIaaa33e0_405);
and \U$2218 ( \2888 , \1458 , RIaaa3368_404);
nor \U$2219 ( \2889 , \2887 , \2888 );
and \U$2220 ( \2890 , \1566 , RIaaa37a0_413);
and \U$2221 ( \2891 , \1470 , RIaaa3980_417);
nor \U$2222 ( \2892 , \2890 , \2891 );
and \U$2223 ( \2893 , \1474 , RIaaa3908_416);
not \U$2224 ( \2894 , RIaaa36b0_411);
nor \U$2225 ( \2895 , \2894 , \1530 );
nor \U$2226 ( \2896 , \2893 , \2895 );
and \U$2227 ( \2897 , \1516 , RIaaa3458_406);
not \U$2228 ( \2898 , RIaaa3548_408);
not \U$2229 ( \2899 , \1491 );
or \U$2230 ( \2900 , \2898 , \2899 );
nand \U$2231 ( \2901 , \1494 , RIaaa3200_401);
nand \U$2232 ( \2902 , \2900 , \2901 );
nor \U$2233 ( \2903 , \2897 , \2902 );
nand \U$2234 ( \2904 , \2889 , \2892 , \2896 , \2903 );
nor \U$2235 ( \2905 , \2886 , \2904 );
buf \U$2236 ( \2906 , \2905 );
buf \U$2237 ( \2907 , \2906 );
not \U$2238 ( \2908 , \2907 );
and \U$2239 ( \2909 , \2448 , \2908 );
not \U$2240 ( \2910 , \2909 );
not \U$2241 ( \2911 , \2690 );
not \U$2242 ( \2912 , \2432 );
or \U$2243 ( \2913 , \2911 , \2912 );
not \U$2244 ( \2914 , \2688 );
not \U$2245 ( \2915 , \2914 );
not \U$2246 ( \2916 , \2915 );
or \U$2247 ( \2917 , \2432 , \2916 );
nand \U$2248 ( \2918 , \2913 , \2917 );
not \U$2249 ( \2919 , \2918 );
buf \U$2250 ( \2920 , \2442 );
not \U$2251 ( \2921 , \2920 );
or \U$2252 ( \2922 , \2919 , \2921 );
nand \U$2253 ( \2923 , \2644 , \2164 );
nand \U$2254 ( \2924 , \2922 , \2923 );
not \U$2255 ( \2925 , \2924 );
or \U$2256 ( \2926 , \2910 , \2925 );
not \U$2257 ( \2927 , \2924 );
not \U$2258 ( \2928 , \2927 );
not \U$2259 ( \2929 , \2909 );
not \U$2260 ( \2930 , \2929 );
or \U$2261 ( \2931 , \2928 , \2930 );
or \U$2262 ( \2932 , \2808 , \2813 );
nand \U$2263 ( \2933 , \2813 , \1579 );
nand \U$2264 ( \2934 , \2932 , \2933 );
not \U$2265 ( \2935 , \2934 );
not \U$2266 ( \2936 , \2410 );
nand \U$2267 ( \2937 , \2936 , \2802 );
nand \U$2268 ( \2938 , \2812 , \2410 );
nand \U$2269 ( \2939 , \2935 , \2937 , \2938 );
not \U$2270 ( \2940 , \2939 );
not \U$2271 ( \2941 , \2777 );
not \U$2272 ( \2942 , \2392 );
buf \U$2273 ( \2943 , \2507 );
not \U$2274 ( \2944 , \2943 );
not \U$2275 ( \2945 , \2944 );
or \U$2276 ( \2946 , \2942 , \2945 );
not \U$2277 ( \2947 , \2391 );
and \U$2278 ( \2948 , \2823 , \2947 );
buf \U$2279 ( \2949 , \2520 );
or \U$2280 ( \2950 , \2949 , \1521 );
not \U$2281 ( \2951 , \2829 );
nand \U$2282 ( \2952 , \2951 , \1521 );
nand \U$2283 ( \2953 , \2950 , \2952 );
nor \U$2284 ( \2954 , \2948 , \2953 );
nand \U$2285 ( \2955 , \2946 , \2954 );
not \U$2286 ( \2956 , \2955 );
or \U$2287 ( \2957 , \2941 , \2956 );
or \U$2288 ( \2958 , \2777 , \2955 );
nand \U$2289 ( \2959 , \2957 , \2958 );
not \U$2290 ( \2960 , \2959 );
or \U$2291 ( \2961 , \2940 , \2960 );
nand \U$2292 ( \2962 , \2776 , \2955 );
nand \U$2293 ( \2963 , \2961 , \2962 );
nand \U$2294 ( \2964 , \2931 , \2963 );
nand \U$2295 ( \2965 , \2926 , \2964 );
not \U$2296 ( \2966 , \2523 );
not \U$2297 ( \2967 , \2692 );
and \U$2298 ( \2968 , \2966 , \2967 );
and \U$2299 ( \2969 , \2523 , \2692 );
nor \U$2300 ( \2970 , \2968 , \2969 );
xnor \U$2301 ( \2971 , \2647 , \2970 );
or \U$2302 ( \2972 , \2965 , \2971 );
and \U$2303 ( \2973 , \2870 , \2972 );
and \U$2304 ( \2974 , \2965 , \2971 );
nor \U$2305 ( \2975 , \2973 , \2974 );
and \U$2306 ( \2976 , \2864 , \2975 );
and \U$2307 ( \2977 , \2853 , \2863 );
or \U$2308 ( \2978 , \2976 , \2977 );
nand \U$2309 ( \2979 , \2721 , \2978 );
nand \U$2310 ( \2980 , \2714 , \2979 );
not \U$2311 ( \2981 , \2154 );
not \U$2312 ( \2982 , \1992 );
or \U$2313 ( \2983 , \2981 , \2982 );
not \U$2314 ( \2984 , \1942 );
not \U$2315 ( \2985 , \2151 );
and \U$2316 ( \2986 , \2984 , \2985 );
not \U$2317 ( \2987 , \2486 );
not \U$2318 ( \2988 , \1897 );
or \U$2319 ( \2989 , \2987 , \2988 );
not \U$2320 ( \2990 , \2486 );
not \U$2321 ( \2991 , \2990 );
or \U$2322 ( \2992 , \2991 , \1897 );
nand \U$2323 ( \2993 , \2989 , \2992 );
buf \U$2324 ( \2994 , \1895 );
and \U$2325 ( \2995 , \2993 , \2994 );
nor \U$2326 ( \2996 , \2986 , \2995 );
nand \U$2327 ( \2997 , \2983 , \2996 );
not \U$2328 ( \2998 , \2997 );
not \U$2329 ( \2999 , \2210 );
not \U$2330 ( \3000 , \2574 );
or \U$2331 ( \3001 , \2999 , \3000 );
not \U$2332 ( \3002 , \2498 );
not \U$2333 ( \3003 , \3002 );
and \U$2334 ( \3004 , \1938 , \3003 );
not \U$2335 ( \3005 , \1938 );
and \U$2336 ( \3006 , \3005 , \2495 );
nor \U$2337 ( \3007 , \3004 , \3006 );
nand \U$2338 ( \3008 , \3001 , \3007 );
not \U$2339 ( \3009 , \2583 );
nor \U$2340 ( \3010 , \3009 , \2214 );
nor \U$2341 ( \3011 , \3008 , \3010 );
not \U$2342 ( \3012 , \3011 );
not \U$2343 ( \3013 , \3012 );
or \U$2344 ( \3014 , \2998 , \3013 );
not \U$2345 ( \3015 , \2997 );
not \U$2346 ( \3016 , \3015 );
not \U$2347 ( \3017 , \3011 );
or \U$2348 ( \3018 , \3016 , \3017 );
not \U$2349 ( \3019 , \2768 );
not \U$2350 ( \3020 , \3019 );
not \U$2351 ( \3021 , \3020 );
not \U$2352 ( \3022 , \1522 );
not \U$2353 ( \3023 , \2753 );
not \U$2354 ( \3024 , \3023 );
nor \U$2355 ( \3025 , \2749 , \3024 );
buf \U$2356 ( \3026 , \3025 );
not \U$2357 ( \3027 , \3026 );
or \U$2358 ( \3028 , \3022 , \3027 );
nor \U$2359 ( \3029 , \2770 , \3023 );
not \U$2360 ( \3030 , \3029 );
not \U$2361 ( \3031 , \3030 );
and \U$2362 ( \3032 , \3031 , \2576 );
not \U$2363 ( \3033 , \2755 );
and \U$2364 ( \3034 , \3033 , \1572 );
nor \U$2365 ( \3035 , \3032 , \3034 );
nand \U$2366 ( \3036 , \3028 , \3035 );
nor \U$2367 ( \3037 , \2749 , \2759 );
buf \U$2368 ( \3038 , \3037 );
and \U$2369 ( \3039 , \3038 , \1521 );
nor \U$2370 ( \3040 , \3036 , \3039 );
nand \U$2371 ( \3041 , \3021 , \3040 );
nand \U$2372 ( \3042 , \3018 , \3041 );
nand \U$2373 ( \3043 , \3014 , \3042 );
xor \U$2374 ( \3044 , \2838 , \2815 );
xor \U$2375 ( \3045 , \3043 , \3044 );
xor \U$2376 ( \3046 , \2777 , \2787 );
xor \U$2377 ( \3047 , \3046 , \2796 );
xor \U$2378 ( \3048 , \3045 , \3047 );
not \U$2379 ( \3049 , \2508 );
not \U$2380 ( \3050 , \3049 );
not \U$2381 ( \3051 , \2416 );
and \U$2382 ( \3052 , \3050 , \3051 );
not \U$2383 ( \3053 , \2363 );
not \U$2384 ( \3054 , \3053 );
not \U$2385 ( \3055 , \2515 );
or \U$2386 ( \3056 , \3054 , \3055 );
and \U$2387 ( \3057 , \2279 , \2521 );
not \U$2388 ( \3058 , \2279 );
and \U$2389 ( \3059 , \3058 , \2951 );
nor \U$2390 ( \3060 , \3057 , \3059 );
nand \U$2391 ( \3061 , \3056 , \3060 );
nor \U$2392 ( \3062 , \3052 , \3061 );
not \U$2393 ( \3063 , \3062 );
not \U$2394 ( \3064 , RIaa9ce28_188);
not \U$2395 ( \3065 , \1049 );
not \U$2396 ( \3066 , \3065 );
or \U$2397 ( \3067 , \3064 , \3066 );
nand \U$2398 ( \3068 , \3067 , \2734 );
not \U$2399 ( \3069 , \3068 );
nand \U$2400 ( \3070 , \3069 , \2767 );
not \U$2401 ( \3071 , \3070 );
not \U$2402 ( \3072 , \3071 );
not \U$2403 ( \3073 , \1572 );
or \U$2404 ( \3074 , \3072 , \3073 );
nand \U$2405 ( \3075 , \2767 , \3068 );
not \U$2406 ( \3076 , \3075 );
not \U$2407 ( \3077 , \3076 );
nand \U$2408 ( \3078 , \3074 , \3077 );
not \U$2409 ( \3079 , \2391 );
not \U$2410 ( \3080 , \3038 );
or \U$2411 ( \3081 , \3079 , \3080 );
and \U$2412 ( \3082 , \3026 , \2280 );
or \U$2413 ( \3083 , \2755 , \1521 );
nand \U$2414 ( \3084 , \3031 , \1521 );
nand \U$2415 ( \3085 , \3083 , \3084 );
nor \U$2416 ( \3086 , \3082 , \3085 );
nand \U$2417 ( \3087 , \3081 , \3086 );
and \U$2418 ( \3088 , \3078 , \3087 );
nand \U$2419 ( \3089 , \3063 , \3088 );
not \U$2420 ( \3090 , \3089 );
not \U$2421 ( \3091 , \2001 );
not \U$2422 ( \3092 , \1366 );
not \U$2423 ( \3093 , \3092 );
or \U$2424 ( \3094 , \3091 , \3093 );
and \U$2425 ( \3095 , \1988 , \1584 );
not \U$2426 ( \3096 , \1988 );
and \U$2427 ( \3097 , \3096 , \1579 );
nor \U$2428 ( \3098 , \3095 , \3097 );
nand \U$2429 ( \3099 , \3094 , \3098 );
buf \U$2430 ( \3100 , \1590 );
nor \U$2431 ( \3101 , \3100 , \2001 );
nor \U$2432 ( \3102 , \3099 , \3101 );
not \U$2433 ( \3103 , \3102 );
or \U$2434 ( \3104 , \3090 , \3103 );
not \U$2435 ( \3105 , \3078 );
not \U$2436 ( \3106 , \3087 );
or \U$2437 ( \3107 , \3105 , \3106 );
nand \U$2438 ( \3108 , \3107 , \3062 );
nand \U$2439 ( \3109 , \3104 , \3108 );
not \U$2440 ( \3110 , \2907 );
not \U$2441 ( \3111 , \2640 );
or \U$2442 ( \3112 , \3110 , \3111 );
not \U$2443 ( \3113 , \2908 );
or \U$2444 ( \3114 , \3113 , \2161 );
nand \U$2445 ( \3115 , \3112 , \3114 );
not \U$2446 ( \3116 , \3115 );
not \U$2447 ( \3117 , \2103 );
or \U$2448 ( \3118 , \3116 , \3117 );
nand \U$2449 ( \3119 , \2918 , \2164 );
nand \U$2450 ( \3120 , \3118 , \3119 );
and \U$2451 ( \3121 , \1458 , RIaaa4448_440);
and \U$2452 ( \3122 , \2344 , RIaaa4538_442);
nor \U$2453 ( \3123 , \3121 , \3122 );
and \U$2454 ( \3124 , \1502 , RIaaa4268_436);
not \U$2455 ( \3125 , \1960 );
not \U$2456 ( \3126 , RIaaa43d0_439);
or \U$2457 ( \3127 , \3125 , \3126 );
and \U$2458 ( \3128 , \1491 , RIaaa42e0_437);
nand \U$2459 ( \3129 , \1494 , RIaaa41f0_435);
not \U$2460 ( \3130 , \3129 );
nor \U$2461 ( \3131 , \3128 , \3130 );
nand \U$2462 ( \3132 , \3127 , \3131 );
nor \U$2463 ( \3133 , \3124 , \3132 );
nand \U$2464 ( \3134 , \3123 , \3133 );
nand \U$2465 ( \3135 , \1480 , RIaaa4628_444);
nand \U$2466 ( \3136 , \1550 , RIaaa4808_448);
not \U$2467 ( \3137 , \1515 );
not \U$2468 ( \3138 , RIaaa45b0_443);
not \U$2469 ( \3139 , \3138 );
and \U$2470 ( \3140 , \3137 , \3139 );
and \U$2471 ( \3141 , \1474 , RIaaa4718_446);
nor \U$2472 ( \3142 , \3140 , \3141 );
nand \U$2473 ( \3143 , \1951 , RIaaa44c0_441);
nand \U$2474 ( \3144 , \3135 , \3136 , \3142 , \3143 );
nor \U$2475 ( \3145 , \3134 , \3144 );
and \U$2476 ( \3146 , \1512 , RIaaa48f8_450);
and \U$2477 ( \3147 , \1541 , RIaaa4358_438);
and \U$2478 ( \3148 , \1483 , RIaaa4970_451);
nor \U$2479 ( \3149 , \3146 , \3147 , \3148 );
and \U$2480 ( \3150 , \2112 , RIaaa4880_449);
and \U$2481 ( \3151 , \1470 , RIaaa4790_447);
nor \U$2482 ( \3152 , \3150 , \3151 );
nand \U$2483 ( \3153 , \1413 , RIaaa46a0_445);
and \U$2484 ( \3154 , \3149 , \3152 , \3153 );
nand \U$2485 ( \3155 , \3145 , \3154 );
buf \U$2486 ( \3156 , \3155 );
buf \U$2487 ( \3157 , \3156 );
and \U$2488 ( \3158 , \2448 , \3157 );
nand \U$2489 ( \3159 , \3120 , \3158 );
not \U$2490 ( \3160 , \3159 );
nor \U$2491 ( \3161 , \3120 , \3158 );
nor \U$2492 ( \3162 , \3160 , \3161 );
and \U$2493 ( \3163 , \3109 , \3162 );
not \U$2494 ( \3164 , \3109 );
and \U$2495 ( \3165 , \3164 , \3161 );
nor \U$2496 ( \3166 , \3163 , \3165 );
not \U$2497 ( \3167 , RIaaa6248_504);
not \U$2498 ( \3168 , \1502 );
or \U$2499 ( \3169 , \3167 , \3168 );
nand \U$2500 ( \3170 , \1512 , RIaaa66f8_514);
nand \U$2501 ( \3171 , \3169 , \3170 );
and \U$2502 ( \3172 , \1480 , RIaaa6860_517);
nor \U$2503 ( \3173 , \3171 , \3172 );
not \U$2504 ( \3174 , RIaaa67e8_516);
not \U$2505 ( \3175 , \1953 );
nor \U$2506 ( \3176 , \3174 , \3175 );
not \U$2507 ( \3177 , RIaaa6680_513);
nor \U$2508 ( \3178 , \3177 , \1426 );
nor \U$2509 ( \3179 , \3176 , \3178 );
and \U$2510 ( \3180 , \1951 , RIaaa64a0_509);
and \U$2511 ( \3181 , RIaaa6338_506, \1541 );
and \U$2512 ( \3182 , \2881 , RIaaa63b0_507);
nor \U$2513 ( \3183 , \3180 , \3181 , \3182 );
and \U$2514 ( \3184 , \3173 , \3179 , \3183 );
not \U$2515 ( \3185 , RIaaa6950_519);
nor \U$2516 ( \3186 , \3185 , \1469 );
not \U$2517 ( \3187 , \3186 );
not \U$2518 ( \3188 , RIaaa6608_512);
nor \U$2519 ( \3189 , \1565 , \3188 );
not \U$2520 ( \3190 , \3189 );
nand \U$2521 ( \3191 , \2199 , RIaaa6590_511);
nand \U$2522 ( \3192 , \1458 , RIaaa6428_508);
nand \U$2523 ( \3193 , \3187 , \3190 , \3191 , \3192 );
not \U$2524 ( \3194 , \1530 );
not \U$2525 ( \3195 , RIaaa6770_515);
not \U$2526 ( \3196 , \3195 );
and \U$2527 ( \3197 , \3194 , \3196 );
and \U$2528 ( \3198 , \1474 , RIaaa68d8_518);
nor \U$2529 ( \3199 , \3197 , \3198 );
and \U$2530 ( \3200 , \1516 , RIaaa6518_510);
not \U$2531 ( \3201 , RIaaa62c0_505);
not \U$2532 ( \3202 , \1491 );
or \U$2533 ( \3203 , \3201 , \3202 );
nand \U$2534 ( \3204 , \1494 , RIaaa61d0_503);
nand \U$2535 ( \3205 , \3203 , \3204 );
nor \U$2536 ( \3206 , \3200 , \3205 );
nand \U$2537 ( \3207 , \3199 , \3206 );
nor \U$2538 ( \3208 , \3193 , \3207 );
nand \U$2539 ( \3209 , \3184 , \3208 );
not \U$2540 ( \3210 , \3209 );
buf \U$2541 ( \3211 , \3210 );
not \U$2542 ( \3212 , \3211 );
nand \U$2543 ( \3213 , \2448 , \3212 );
not \U$2544 ( \3214 , \3213 );
not \U$2545 ( \3215 , \3156 );
not \U$2546 ( \3216 , \3215 );
not \U$2547 ( \3217 , \2161 );
or \U$2548 ( \3218 , \3216 , \3217 );
not \U$2549 ( \3219 , \2640 );
nand \U$2550 ( \3220 , \3219 , \3156 );
nand \U$2551 ( \3221 , \3218 , \3220 );
not \U$2552 ( \3222 , \3221 );
not \U$2553 ( \3223 , \2103 );
or \U$2554 ( \3224 , \3222 , \3223 );
nand \U$2555 ( \3225 , \3115 , \2164 );
nand \U$2556 ( \3226 , \3224 , \3225 );
nand \U$2557 ( \3227 , \3214 , \3226 );
not \U$2558 ( \3228 , \3227 );
not \U$2559 ( \3229 , \2210 );
not \U$2560 ( \3230 , \3092 );
or \U$2561 ( \3231 , \3229 , \3230 );
not \U$2562 ( \3232 , \1583 );
not \U$2563 ( \3233 , \3232 );
and \U$2564 ( \3234 , \2230 , \3233 );
not \U$2565 ( \3235 , \2230 );
and \U$2566 ( \3236 , \3235 , \1579 );
nor \U$2567 ( \3237 , \3234 , \3236 );
nand \U$2568 ( \3238 , \3231 , \3237 );
not \U$2569 ( \3239 , \2241 );
nor \U$2570 ( \3240 , \3239 , \2210 );
nor \U$2571 ( \3241 , \3238 , \3240 );
not \U$2572 ( \3242 , \3241 );
not \U$2573 ( \3243 , \2363 );
not \U$2574 ( \3244 , \3038 );
or \U$2575 ( \3245 , \3243 , \3244 );
and \U$2576 ( \3246 , \3026 , \3053 );
not \U$2577 ( \3247 , \2770 );
nand \U$2578 ( \3248 , \3247 , \2758 );
or \U$2579 ( \3249 , \2279 , \3248 );
not \U$2580 ( \3250 , \2755 );
nand \U$2581 ( \3251 , \2279 , \3250 );
nand \U$2582 ( \3252 , \3249 , \3251 );
nor \U$2583 ( \3253 , \3246 , \3252 );
nand \U$2584 ( \3254 , \3245 , \3253 );
not \U$2585 ( \3255 , \3071 );
not \U$2586 ( \3256 , \2288 );
or \U$2587 ( \3257 , \3255 , \3256 );
and \U$2588 ( \3258 , \2768 , \3068 );
buf \U$2589 ( \3259 , \3258 );
and \U$2590 ( \3260 , \3259 , \1571 );
nor \U$2591 ( \3261 , \3077 , \1571 );
nor \U$2592 ( \3262 , \3260 , \3261 );
nand \U$2593 ( \3263 , \3257 , \3262 );
and \U$2594 ( \3264 , \3254 , \3263 );
not \U$2595 ( \3265 , \1988 );
nand \U$2596 ( \3266 , \3265 , \2944 );
and \U$2597 ( \3267 , \2823 , \1988 );
or \U$2598 ( \3268 , \2949 , \2363 );
not \U$2599 ( \3269 , \2359 );
not \U$2600 ( \3270 , \3269 );
nand \U$2601 ( \3271 , \3270 , \2951 );
nand \U$2602 ( \3272 , \3268 , \3271 );
nor \U$2603 ( \3273 , \3267 , \3272 );
nand \U$2604 ( \3274 , \3266 , \3273 );
xor \U$2605 ( \3275 , \3264 , \3274 );
and \U$2606 ( \3276 , \3242 , \3275 );
and \U$2607 ( \3277 , \3264 , \3274 );
nor \U$2608 ( \3278 , \3276 , \3277 );
not \U$2609 ( \3279 , \3278 );
or \U$2610 ( \3280 , \3228 , \3279 );
not \U$2611 ( \3281 , \3226 );
nand \U$2612 ( \3282 , \3281 , \3213 );
nand \U$2613 ( \3283 , \3280 , \3282 );
nand \U$2614 ( \3284 , \3166 , \3283 );
not \U$2615 ( \3285 , \3284 );
xor \U$2616 ( \3286 , \3062 , \3088 );
xor \U$2617 ( \3287 , \3286 , \3102 );
not \U$2618 ( \3288 , \3287 );
xor \U$2619 ( \3289 , \3078 , \3087 );
not \U$2620 ( \3290 , \3289 );
not \U$2621 ( \3291 , \2639 );
not \U$2622 ( \3292 , \2572 );
or \U$2623 ( \3293 , \3291 , \3292 );
not \U$2624 ( \3294 , \2151 );
not \U$2625 ( \3295 , \2396 );
and \U$2626 ( \3296 , \3294 , \3295 );
not \U$2627 ( \3297 , \3294 );
and \U$2628 ( \3298 , \3297 , \2495 );
nor \U$2629 ( \3299 , \3296 , \3298 );
nand \U$2630 ( \3300 , \3293 , \3299 );
not \U$2631 ( \3301 , \2486 );
nor \U$2632 ( \3302 , \2405 , \3301 );
nor \U$2633 ( \3303 , \3300 , \3302 );
not \U$2634 ( \3304 , \3303 );
or \U$2635 ( \3305 , \3290 , \3304 );
or \U$2636 ( \3306 , \3289 , \3303 );
nand \U$2637 ( \3307 , \3305 , \3306 );
not \U$2638 ( \3308 , \3307 );
and \U$2639 ( \3309 , \1900 , \2907 );
not \U$2640 ( \3310 , \2235 );
not \U$2641 ( \3311 , \2915 );
or \U$2642 ( \3312 , \3310 , \3311 );
not \U$2643 ( \3313 , \2691 );
nand \U$2644 ( \3314 , \3313 , \1993 );
nand \U$2645 ( \3315 , \3312 , \3314 );
nor \U$2646 ( \3316 , \3309 , \3315 );
not \U$2647 ( \3317 , \2907 );
nand \U$2648 ( \3318 , \3317 , \2563 );
nand \U$2649 ( \3319 , \3316 , \3318 );
not \U$2650 ( \3320 , \3319 );
or \U$2651 ( \3321 , \3308 , \3320 );
not \U$2652 ( \3322 , \3303 );
nand \U$2653 ( \3323 , \3322 , \3289 );
nand \U$2654 ( \3324 , \3321 , \3323 );
not \U$2655 ( \3325 , \3324 );
or \U$2656 ( \3326 , \3288 , \3325 );
or \U$2657 ( \3327 , \3287 , \3324 );
and \U$2658 ( \3328 , \2574 , \2153 );
or \U$2659 ( \3329 , \2396 , \2210 );
or \U$2660 ( \3330 , \2400 , \2225 );
nand \U$2661 ( \3331 , \3329 , \3330 );
nor \U$2662 ( \3332 , \3328 , \3331 );
nand \U$2663 ( \3333 , \2406 , \2551 );
nand \U$2664 ( \3334 , \3332 , \3333 );
and \U$2665 ( \3335 , \1900 , \2690 );
and \U$2666 ( \3336 , \2486 , \2235 );
not \U$2667 ( \3337 , \2486 );
and \U$2668 ( \3338 , \3337 , \1992 );
or \U$2669 ( \3339 , \3336 , \3338 );
nor \U$2670 ( \3340 , \3335 , \3339 );
not \U$2671 ( \3341 , \2003 );
nand \U$2672 ( \3342 , \3341 , \2691 );
nand \U$2673 ( \3343 , \3340 , \3342 );
xor \U$2674 ( \3344 , \3334 , \3343 );
not \U$2675 ( \3345 , \3040 );
nand \U$2676 ( \3346 , \3345 , \3020 );
nand \U$2677 ( \3347 , \3346 , \3041 );
xor \U$2678 ( \3348 , \3344 , \3347 );
nand \U$2679 ( \3349 , \3327 , \3348 );
nand \U$2680 ( \3350 , \3326 , \3349 );
not \U$2681 ( \3351 , \3350 );
or \U$2682 ( \3352 , \3285 , \3351 );
not \U$2683 ( \3353 , \3283 );
not \U$2684 ( \3354 , \3166 );
nand \U$2685 ( \3355 , \3353 , \3354 );
nand \U$2686 ( \3356 , \3352 , \3355 );
xor \U$2687 ( \3357 , \3048 , \3356 );
or \U$2688 ( \3358 , \3161 , \3109 );
nand \U$2689 ( \3359 , \3358 , \3159 );
xor \U$2690 ( \3360 , \2909 , \2924 );
xor \U$2691 ( \3361 , \3360 , \2963 );
xor \U$2692 ( \3362 , \3359 , \3361 );
not \U$2693 ( \3363 , \2939 );
not \U$2694 ( \3364 , \3363 );
not \U$2695 ( \3365 , \2959 );
and \U$2696 ( \3366 , \3364 , \3365 );
and \U$2697 ( \3367 , \2959 , \3363 );
nor \U$2698 ( \3368 , \3366 , \3367 );
not \U$2699 ( \3369 , \3368 );
not \U$2700 ( \3370 , \3369 );
not \U$2701 ( \3371 , \3012 );
and \U$2702 ( \3372 , \3041 , \2997 );
not \U$2703 ( \3373 , \3041 );
and \U$2704 ( \3374 , \3373 , \3015 );
nor \U$2705 ( \3375 , \3372 , \3374 );
not \U$2706 ( \3376 , \3375 );
or \U$2707 ( \3377 , \3371 , \3376 );
or \U$2708 ( \3378 , \3375 , \3012 );
nand \U$2709 ( \3379 , \3377 , \3378 );
not \U$2710 ( \3380 , \3379 );
not \U$2711 ( \3381 , \3380 );
or \U$2712 ( \3382 , \3370 , \3381 );
not \U$2713 ( \3383 , \3379 );
not \U$2714 ( \3384 , \3368 );
or \U$2715 ( \3385 , \3383 , \3384 );
xor \U$2716 ( \3386 , \3334 , \3343 );
and \U$2717 ( \3387 , \3386 , \3347 );
and \U$2718 ( \3388 , \3334 , \3343 );
or \U$2719 ( \3389 , \3387 , \3388 );
nand \U$2720 ( \3390 , \3385 , \3389 );
nand \U$2721 ( \3391 , \3382 , \3390 );
xor \U$2722 ( \3392 , \3362 , \3391 );
and \U$2723 ( \3393 , \3357 , \3392 );
and \U$2724 ( \3394 , \3048 , \3356 );
or \U$2725 ( \3395 , \3393 , \3394 );
not \U$2726 ( \3396 , \3395 );
not \U$2727 ( \3397 , \2870 );
not \U$2728 ( \3398 , \2971 );
not \U$2729 ( \3399 , \2965 );
or \U$2730 ( \3400 , \3398 , \3399 );
or \U$2731 ( \3401 , \2965 , \2971 );
nand \U$2732 ( \3402 , \3400 , \3401 );
not \U$2733 ( \3403 , \3402 );
and \U$2734 ( \3404 , \3397 , \3403 );
and \U$2735 ( \3405 , \2870 , \3402 );
nor \U$2736 ( \3406 , \3404 , \3405 );
not \U$2737 ( \3407 , \3406 );
xor \U$2738 ( \3408 , \3043 , \3044 );
and \U$2739 ( \3409 , \3408 , \3047 );
and \U$2740 ( \3410 , \3043 , \3044 );
or \U$2741 ( \3411 , \3409 , \3410 );
xor \U$2742 ( \3412 , \3359 , \3361 );
and \U$2743 ( \3413 , \3412 , \3391 );
and \U$2744 ( \3414 , \3359 , \3361 );
or \U$2745 ( \3415 , \3413 , \3414 );
xor \U$2746 ( \3416 , \3411 , \3415 );
not \U$2747 ( \3417 , \3416 );
or \U$2748 ( \3418 , \3407 , \3417 );
or \U$2749 ( \3419 , \3416 , \3406 );
nand \U$2750 ( \3420 , \3418 , \3419 );
not \U$2751 ( \3421 , \3420 );
nand \U$2752 ( \3422 , \3396 , \3421 );
xor \U$2753 ( \3423 , \2853 , \2863 );
xor \U$2754 ( \3424 , \3423 , \2975 );
not \U$2755 ( \3425 , \3406 );
and \U$2756 ( \3426 , \3416 , \3425 );
and \U$2757 ( \3427 , \3411 , \3415 );
nor \U$2758 ( \3428 , \3426 , \3427 );
nand \U$2759 ( \3429 , \3424 , \3428 );
nand \U$2760 ( \3430 , \3422 , \3429 );
nor \U$2761 ( \3431 , \2980 , \3430 );
buf \U$2762 ( \3432 , \3431 );
not \U$2763 ( \3433 , \2393 );
not \U$2764 ( \3434 , \2556 );
or \U$2765 ( \3435 , \3433 , \3434 );
not \U$2766 ( \3436 , \1943 );
not \U$2767 ( \3437 , \1522 );
and \U$2768 ( \3438 , \3436 , \3437 );
not \U$2769 ( \3439 , \1993 );
nor \U$2770 ( \3440 , \3439 , \2401 );
nor \U$2771 ( \3441 , \3438 , \3440 );
nand \U$2772 ( \3442 , \3435 , \3441 );
and \U$2773 ( \3443 , \2563 , \2392 );
nor \U$2774 ( \3444 , \3442 , \3443 );
xor \U$2775 ( \3445 , \3444 , \2605 );
or \U$2776 ( \3446 , \2562 , \2565 );
and \U$2777 ( \3447 , \3446 , \2586 );
and \U$2778 ( \3448 , \2571 , \2585 );
nor \U$2779 ( \3449 , \3447 , \3448 );
xnor \U$2780 ( \3450 , \3445 , \3449 );
not \U$2781 ( \3451 , \3450 );
not \U$2782 ( \3452 , \1573 );
not \U$2783 ( \3453 , \2583 );
or \U$2784 ( \3454 , \3452 , \3453 );
and \U$2785 ( \3455 , \2574 , \2517 );
not \U$2786 ( \3456 , \1938 );
not \U$2787 ( \3457 , \2448 );
or \U$2788 ( \3458 , \3456 , \3457 );
nand \U$2789 ( \3459 , \3458 , \2400 );
nor \U$2790 ( \3460 , \3455 , \3459 );
nand \U$2791 ( \3461 , \3454 , \3460 );
not \U$2792 ( \3462 , \2435 );
not \U$2793 ( \3463 , \3462 );
or \U$2794 ( \3464 , \3463 , \2410 );
buf \U$2795 ( \3465 , \2443 );
nand \U$2796 ( \3466 , \3465 , \2410 );
and \U$2797 ( \3467 , \2438 , \2813 );
not \U$2798 ( \3468 , \2596 );
nor \U$2799 ( \3469 , \3468 , \2813 );
nor \U$2800 ( \3470 , \3467 , \3469 );
nand \U$2801 ( \3471 , \3464 , \3466 , \3470 );
xor \U$2802 ( \3472 , \3461 , \3471 );
nand \U$2803 ( \3473 , \3451 , \3472 );
not \U$2804 ( \3474 , \3472 );
not \U$2805 ( \3475 , \3474 );
not \U$2806 ( \3476 , \3450 );
or \U$2807 ( \3477 , \3475 , \3476 );
xor \U$2808 ( \3478 , \2590 , \2606 );
and \U$2809 ( \3479 , \3478 , \2612 );
and \U$2810 ( \3480 , \2590 , \2606 );
or \U$2811 ( \3481 , \3479 , \3480 );
not \U$2812 ( \3482 , \3481 );
nand \U$2813 ( \3483 , \3477 , \3482 );
and \U$2814 ( \3484 , \3473 , \3483 );
not \U$2815 ( \3485 , \3484 );
nand \U$2816 ( \3486 , \3471 , \3461 );
not \U$2817 ( \3487 , \3449 );
not \U$2818 ( \3488 , \3444 );
and \U$2819 ( \3489 , \3487 , \3488 );
and \U$2820 ( \3490 , \3449 , \3444 );
nor \U$2821 ( \3491 , \3489 , \3490 );
not \U$2822 ( \3492 , \3491 );
not \U$2823 ( \3493 , \2605 );
and \U$2824 ( \3494 , \3492 , \3493 );
not \U$2825 ( \3495 , \3444 );
nor \U$2826 ( \3496 , \3495 , \3449 );
nor \U$2827 ( \3497 , \3494 , \3496 );
xor \U$2828 ( \3498 , \3486 , \3497 );
not \U$2829 ( \3499 , \2410 );
not \U$2830 ( \3500 , \2448 );
or \U$2831 ( \3501 , \3499 , \3500 );
nand \U$2832 ( \3502 , \3501 , \3444 );
not \U$2833 ( \3503 , \2367 );
not \U$2834 ( \3504 , \3503 );
not \U$2835 ( \3505 , \2316 );
or \U$2836 ( \3506 , \3504 , \3505 );
not \U$2837 ( \3507 , \2317 );
nand \U$2838 ( \3508 , \3506 , \3507 );
not \U$2839 ( \3509 , \2994 );
not \U$2840 ( \3510 , \3509 );
buf \U$2841 ( \3511 , \2234 );
not \U$2842 ( \3512 , \3511 );
not \U$2843 ( \3513 , \1991 );
buf \U$2844 ( \3514 , \3513 );
not \U$2845 ( \3515 , \3514 );
and \U$2846 ( \3516 , \3515 , \2517 );
not \U$2847 ( \3517 , \3515 );
and \U$2848 ( \3518 , \3517 , \1573 );
nor \U$2849 ( \3519 , \3516 , \3518 );
nor \U$2850 ( \3520 , \3512 , \3519 );
or \U$2851 ( \3521 , \3510 , \3520 );
xnor \U$2852 ( \3522 , \2401 , \3515 );
nand \U$2853 ( \3523 , \3512 , \3522 );
nand \U$2854 ( \3524 , \3521 , \3523 );
not \U$2855 ( \3525 , \3524 );
xor \U$2856 ( \3526 , \3508 , \3525 );
or \U$2857 ( \3527 , \3463 , \2813 );
nand \U$2858 ( \3528 , \3465 , \2813 );
and \U$2859 ( \3529 , \2438 , \2392 );
nor \U$2860 ( \3530 , \3468 , \2392 );
nor \U$2861 ( \3531 , \3529 , \3530 );
nand \U$2862 ( \3532 , \3527 , \3528 , \3531 );
xor \U$2863 ( \3533 , \3526 , \3532 );
xor \U$2864 ( \3534 , \3502 , \3533 );
xnor \U$2865 ( \3535 , \3498 , \3534 );
not \U$2866 ( \3536 , \3535 );
or \U$2867 ( \3537 , \3485 , \3536 );
xor \U$2868 ( \3538 , \3472 , \3481 );
xnor \U$2869 ( \3539 , \3538 , \3451 );
not \U$2870 ( \3540 , \3539 );
not \U$2871 ( \3541 , \2529 );
not \U$2872 ( \3542 , \3541 );
not \U$2873 ( \3543 , \2617 );
or \U$2874 ( \3544 , \3542 , \3543 );
not \U$2875 ( \3545 , \2553 );
nand \U$2876 ( \3546 , \3545 , \2613 );
nand \U$2877 ( \3547 , \3544 , \3546 );
nand \U$2878 ( \3548 , \3540 , \3547 );
nand \U$2879 ( \3549 , \3537 , \3548 );
xor \U$2880 ( \3550 , \3497 , \3486 );
not \U$2881 ( \3551 , \3534 );
and \U$2882 ( \3552 , \3550 , \3551 );
and \U$2883 ( \3553 , \3497 , \3486 );
or \U$2884 ( \3554 , \3552 , \3553 );
xor \U$2885 ( \3555 , \3508 , \3525 );
and \U$2886 ( \3556 , \3555 , \3532 );
and \U$2887 ( \3557 , \3508 , \3525 );
or \U$2888 ( \3558 , \3556 , \3557 );
not \U$2889 ( \3559 , \3558 );
and \U$2890 ( \3560 , \2393 , \3462 );
not \U$2891 ( \3561 , \2393 );
and \U$2892 ( \3562 , \3561 , \3465 );
nor \U$2893 ( \3563 , \3560 , \3562 );
and \U$2894 ( \3564 , \2438 , \2401 );
nor \U$2895 ( \3565 , \3468 , \2401 );
nor \U$2896 ( \3566 , \3564 , \3565 );
and \U$2897 ( \3567 , \3563 , \3566 );
not \U$2898 ( \3568 , \1573 );
not \U$2899 ( \3569 , \2563 );
or \U$2900 ( \3570 , \3568 , \3569 );
and \U$2901 ( \3571 , \2556 , \2517 );
nor \U$2902 ( \3572 , \3571 , \1993 );
nand \U$2903 ( \3573 , \3570 , \3572 );
and \U$2904 ( \3574 , \2448 , \2813 );
nor \U$2905 ( \3575 , \3573 , \3574 );
xor \U$2906 ( \3576 , \3567 , \3575 );
xor \U$2907 ( \3577 , \3559 , \3576 );
nand \U$2908 ( \3578 , \3533 , \3502 );
xor \U$2909 ( \3579 , \3577 , \3578 );
and \U$2910 ( \3580 , \3554 , \3579 );
nor \U$2911 ( \3581 , \3549 , \3580 );
xor \U$2912 ( \3582 , \3559 , \3576 );
and \U$2913 ( \3583 , \3582 , \3578 );
and \U$2914 ( \3584 , \3559 , \3576 );
or \U$2915 ( \3585 , \3583 , \3584 );
buf \U$2916 ( \3586 , \1892 );
not \U$2917 ( \3587 , \3586 );
not \U$2918 ( \3588 , \3507 );
or \U$2919 ( \3589 , \3587 , \3588 );
nand \U$2920 ( \3590 , \3589 , \1898 );
not \U$2921 ( \3591 , \3590 );
not \U$2922 ( \3592 , \3591 );
nand \U$2923 ( \3593 , \2448 , \2392 );
nand \U$2924 ( \3594 , \3592 , \3593 );
or \U$2925 ( \3595 , \2433 , \2517 );
or \U$2926 ( \3596 , \2434 , \1573 );
nand \U$2927 ( \3597 , \3595 , \3596 , \2164 );
not \U$2928 ( \3598 , \3597 );
not \U$2929 ( \3599 , \2920 );
not \U$2930 ( \3600 , \3599 );
or \U$2931 ( \3601 , \3598 , \3600 );
and \U$2932 ( \3602 , \2401 , \2434 );
not \U$2933 ( \3603 , \2401 );
and \U$2934 ( \3604 , \3603 , \2433 );
nor \U$2935 ( \3605 , \3602 , \3604 );
or \U$2936 ( \3606 , \3605 , \2164 );
nand \U$2937 ( \3607 , \3601 , \3606 );
xnor \U$2938 ( \3608 , \3594 , \3607 );
not \U$2939 ( \3609 , \3608 );
not \U$2940 ( \3610 , \3573 );
and \U$2941 ( \3611 , \3609 , \3610 );
and \U$2942 ( \3612 , \3608 , \3573 );
nor \U$2943 ( \3613 , \3611 , \3612 );
not \U$2944 ( \3614 , \3567 );
and \U$2945 ( \3615 , \3575 , \3614 );
nor \U$2946 ( \3616 , \3615 , \3574 );
xnor \U$2947 ( \3617 , \3613 , \3616 );
nand \U$2948 ( \3618 , \3585 , \3617 );
and \U$2949 ( \3619 , \3432 , \3581 , \3618 );
not \U$2950 ( \3620 , \3283 );
not \U$2951 ( \3621 , \3354 );
or \U$2952 ( \3622 , \3620 , \3621 );
or \U$2953 ( \3623 , \3283 , \3354 );
nand \U$2954 ( \3624 , \3622 , \3623 );
not \U$2955 ( \3625 , \3624 );
not \U$2956 ( \3626 , \3350 );
and \U$2957 ( \3627 , \3625 , \3626 );
and \U$2958 ( \3628 , \3624 , \3350 );
nor \U$2959 ( \3629 , \3627 , \3628 );
not \U$2960 ( \3630 , \3629 );
not \U$2961 ( \3631 , \3368 );
not \U$2962 ( \3632 , \3380 );
or \U$2963 ( \3633 , \3631 , \3632 );
nand \U$2964 ( \3634 , \3369 , \3379 );
nand \U$2965 ( \3635 , \3633 , \3634 );
buf \U$2966 ( \3636 , \3389 );
xor \U$2967 ( \3637 , \3635 , \3636 );
not \U$2968 ( \3638 , \3637 );
not \U$2969 ( \3639 , RIaaa57f8_482);
not \U$2970 ( \3640 , \1512 );
or \U$2971 ( \3641 , \3639 , \3640 );
not \U$2972 ( \3642 , \1502 );
not \U$2973 ( \3643 , RIaaa54b0_475);
or \U$2974 ( \3644 , \3642 , \3643 );
nand \U$2975 ( \3645 , \3641 , \3644 );
and \U$2976 ( \3646 , RIaaa5618_478, \1480 );
nor \U$2977 ( \3647 , \3645 , \3646 );
nand \U$2978 ( \3648 , \1436 , RIaaa52d0_471);
and \U$2979 ( \3649 , \1541 , RIaaa5528_476);
and \U$2980 ( \3650 , \1449 , RIaaa5258_470);
nor \U$2981 ( \3651 , \3649 , \3650 );
and \U$2982 ( \3652 , \3648 , \3651 );
and \U$2983 ( \3653 , \1551 , RIaaa5708_480);
and \U$2984 ( \3654 , \1413 , RIaaa5690_479);
nor \U$2985 ( \3655 , \3653 , \3654 );
nand \U$2986 ( \3656 , \3647 , \3652 , \3655 );
and \U$2987 ( \3657 , \1458 , RIaaa5348_472);
and \U$2988 ( \3658 , \2344 , RIaaa53c0_473);
nor \U$2989 ( \3659 , \3657 , \3658 );
and \U$2990 ( \3660 , \1470 , RIaaa58e8_484);
and \U$2991 ( \3661 , \1474 , RIaaa5960_485);
nor \U$2992 ( \3662 , \3660 , \3661 );
and \U$2993 ( \3663 , \2112 , RIaaa5780_481);
and \U$2994 ( \3664 , \1516 , RIaaa5438_474);
nor \U$2995 ( \3665 , \3663 , \3664 );
and \U$2996 ( \3666 , \1531 , RIaaa5870_483);
not \U$2997 ( \3667 , RIaaa55a0_477);
not \U$2998 ( \3668 , \1491 );
or \U$2999 ( \3669 , \3667 , \3668 );
not \U$3000 ( \3670 , RIaaa51e0_469);
nor \U$3001 ( \3671 , \3670 , \1495 );
not \U$3002 ( \3672 , \3671 );
nand \U$3003 ( \3673 , \3669 , \3672 );
nor \U$3004 ( \3674 , \3666 , \3673 );
nand \U$3005 ( \3675 , \3659 , \3662 , \3665 , \3674 );
nor \U$3006 ( \3676 , \3656 , \3675 );
buf \U$3007 ( \3677 , \3676 );
buf \U$3008 ( \3678 , \3677 );
not \U$3009 ( \3679 , \3678 );
and \U$3010 ( \3680 , \2448 , \3679 );
not \U$3011 ( \3681 , \3211 );
not \U$3012 ( \3682 , \2161 );
or \U$3013 ( \3683 , \3681 , \3682 );
not \U$3014 ( \3684 , \3212 );
or \U$3015 ( \3685 , \2161 , \3684 );
nand \U$3016 ( \3686 , \3683 , \3685 );
not \U$3017 ( \3687 , \3686 );
not \U$3018 ( \3688 , \2103 );
or \U$3019 ( \3689 , \3687 , \3688 );
nand \U$3020 ( \3690 , \3221 , \2164 );
nand \U$3021 ( \3691 , \3689 , \3690 );
xor \U$3022 ( \3692 , \3680 , \3691 );
and \U$3023 ( \3693 , \2515 , \2230 );
not \U$3024 ( \3694 , \2951 );
not \U$3025 ( \3695 , \1987 );
or \U$3026 ( \3696 , \3694 , \3695 );
or \U$3027 ( \3697 , \2520 , \1996 );
nand \U$3028 ( \3698 , \3696 , \3697 );
nor \U$3029 ( \3699 , \3693 , \3698 );
nand \U$3030 ( \3700 , \2508 , \1937 );
nand \U$3031 ( \3701 , \3699 , \3700 );
and \U$3032 ( \3702 , \3259 , \1521 );
nor \U$3033 ( \3703 , \1521 , \3077 );
nor \U$3034 ( \3704 , \3702 , \3703 );
nand \U$3035 ( \3705 , \3071 , \2279 );
nand \U$3036 ( \3706 , \3704 , \3705 );
not \U$3037 ( \3707 , \3706 );
nand \U$3038 ( \3708 , \3038 , \1996 );
not \U$3039 ( \3709 , \3708 );
not \U$3040 ( \3710 , \1986 );
not \U$3041 ( \3711 , \3026 );
or \U$3042 ( \3712 , \3710 , \3711 );
and \U$3043 ( \3713 , \3029 , \2359 );
nor \U$3044 ( \3714 , \2755 , \2359 );
nor \U$3045 ( \3715 , \3713 , \3714 );
nand \U$3046 ( \3716 , \3712 , \3715 );
nor \U$3047 ( \3717 , \3709 , \3716 );
nor \U$3048 ( \3718 , \3707 , \3717 );
xor \U$3049 ( \3719 , \3701 , \3718 );
not \U$3050 ( \3720 , \2152 );
not \U$3051 ( \3721 , \1591 );
or \U$3052 ( \3722 , \3720 , \3721 );
not \U$3053 ( \3723 , \2801 );
and \U$3054 ( \3724 , \3723 , \2154 );
or \U$3055 ( \3725 , \3232 , \2225 );
nand \U$3056 ( \3726 , \2291 , \2225 );
nand \U$3057 ( \3727 , \3725 , \3726 );
nor \U$3058 ( \3728 , \3724 , \3727 );
nand \U$3059 ( \3729 , \3722 , \3728 );
and \U$3060 ( \3730 , \3719 , \3729 );
and \U$3061 ( \3731 , \3701 , \3718 );
or \U$3062 ( \3732 , \3730 , \3731 );
and \U$3063 ( \3733 , \3692 , \3732 );
and \U$3064 ( \3734 , \3680 , \3691 );
nor \U$3065 ( \3735 , \3733 , \3734 );
xnor \U$3066 ( \3736 , \3226 , \3213 );
not \U$3067 ( \3737 , \3736 );
not \U$3068 ( \3738 , \3278 );
and \U$3069 ( \3739 , \3737 , \3738 );
and \U$3070 ( \3740 , \3278 , \3736 );
nor \U$3071 ( \3741 , \3739 , \3740 );
xor \U$3072 ( \3742 , \3735 , \3741 );
not \U$3073 ( \3743 , \3319 );
not \U$3074 ( \3744 , \3743 );
not \U$3075 ( \3745 , \3307 );
and \U$3076 ( \3746 , \3744 , \3745 );
and \U$3077 ( \3747 , \3307 , \3743 );
nor \U$3078 ( \3748 , \3746 , \3747 );
not \U$3079 ( \3749 , \3275 );
not \U$3080 ( \3750 , \3241 );
and \U$3081 ( \3751 , \3749 , \3750 );
and \U$3082 ( \3752 , \3275 , \3241 );
nor \U$3083 ( \3753 , \3751 , \3752 );
nand \U$3084 ( \3754 , \3748 , \3753 );
not \U$3085 ( \3755 , \2907 );
not \U$3086 ( \3756 , \1993 );
or \U$3087 ( \3757 , \3755 , \3756 );
not \U$3088 ( \3758 , \1943 );
not \U$3089 ( \3759 , \2907 );
and \U$3090 ( \3760 , \3758 , \3759 );
and \U$3091 ( \3761 , \3157 , \1897 );
not \U$3092 ( \3762 , \3157 );
and \U$3093 ( \3763 , \3762 , \1898 );
nor \U$3094 ( \3764 , \3761 , \3763 );
not \U$3095 ( \3765 , \3764 );
and \U$3096 ( \3766 , \3510 , \3765 );
nor \U$3097 ( \3767 , \3760 , \3766 );
nand \U$3098 ( \3768 , \3757 , \3767 );
not \U$3099 ( \3769 , \3768 );
xnor \U$3100 ( \3770 , \3254 , \3263 );
not \U$3101 ( \3771 , \3770 );
not \U$3102 ( \3772 , \2915 );
not \U$3103 ( \3773 , \2406 );
or \U$3104 ( \3774 , \3772 , \3773 );
not \U$3105 ( \3775 , \2389 );
not \U$3106 ( \3776 , \2689 );
and \U$3107 ( \3777 , \3775 , \3776 );
and \U$3108 ( \3778 , \2486 , \2396 );
not \U$3109 ( \3779 , \2486 );
and \U$3110 ( \3780 , \3779 , \2399 );
nor \U$3111 ( \3781 , \3778 , \3780 );
nor \U$3112 ( \3782 , \3777 , \3781 );
nand \U$3113 ( \3783 , \3774 , \3782 );
not \U$3114 ( \3784 , \3783 );
or \U$3115 ( \3785 , \3771 , \3784 );
or \U$3116 ( \3786 , \3770 , \3783 );
nand \U$3117 ( \3787 , \3785 , \3786 );
not \U$3118 ( \3788 , \3787 );
or \U$3119 ( \3789 , \3769 , \3788 );
not \U$3120 ( \3790 , \3770 );
nand \U$3121 ( \3791 , \3790 , \3783 );
nand \U$3122 ( \3792 , \3789 , \3791 );
and \U$3123 ( \3793 , \3754 , \3792 );
nor \U$3124 ( \3794 , \3748 , \3753 );
nor \U$3125 ( \3795 , \3793 , \3794 );
and \U$3126 ( \3796 , \3742 , \3795 );
and \U$3127 ( \3797 , \3735 , \3741 );
or \U$3128 ( \3798 , \3796 , \3797 );
not \U$3129 ( \3799 , \3798 );
or \U$3130 ( \3800 , \3638 , \3799 );
or \U$3131 ( \3801 , \3798 , \3637 );
nand \U$3132 ( \3802 , \3800 , \3801 );
not \U$3133 ( \3803 , \3802 );
or \U$3134 ( \3804 , \3630 , \3803 );
or \U$3135 ( \3805 , \3629 , \3802 );
nand \U$3136 ( \3806 , \3804 , \3805 );
xor \U$3137 ( \3807 , \3287 , \3324 );
xnor \U$3138 ( \3808 , \3807 , \3348 );
not \U$3139 ( \3809 , \3732 );
and \U$3140 ( \3810 , \3692 , \3809 );
not \U$3141 ( \3811 , \3692 );
and \U$3142 ( \3812 , \3811 , \3732 );
nor \U$3143 ( \3813 , \3810 , \3812 );
not \U$3144 ( \3814 , \2486 );
not \U$3145 ( \3815 , \3100 );
not \U$3146 ( \3816 , \3815 );
or \U$3147 ( \3817 , \3814 , \3816 );
and \U$3148 ( \3818 , \2802 , \2639 );
or \U$3149 ( \3819 , \2534 , \2152 );
not \U$3150 ( \3820 , \1578 );
nand \U$3151 ( \3821 , \3820 , \3294 );
nand \U$3152 ( \3822 , \3819 , \3821 );
nor \U$3153 ( \3823 , \3818 , \3822 );
nand \U$3154 ( \3824 , \3817 , \3823 );
not \U$3155 ( \3825 , \3824 );
not \U$3156 ( \3826 , \2210 );
not \U$3157 ( \3827 , \2515 );
or \U$3158 ( \3828 , \3826 , \3827 );
and \U$3159 ( \3829 , \1937 , \2830 );
not \U$3160 ( \3830 , \1937 );
and \U$3161 ( \3831 , \3830 , \2521 );
nor \U$3162 ( \3832 , \3829 , \3831 );
nand \U$3163 ( \3833 , \3828 , \3832 );
nor \U$3164 ( \3834 , \2943 , \2210 );
nor \U$3165 ( \3835 , \3833 , \3834 );
not \U$3166 ( \3836 , \3835 );
not \U$3167 ( \3837 , \1937 );
not \U$3168 ( \3838 , \3038 );
or \U$3169 ( \3839 , \3837 , \3838 );
and \U$3170 ( \3840 , \3026 , \2230 );
or \U$3171 ( \3841 , \1995 , \3248 );
nand \U$3172 ( \3842 , \2754 , \1986 );
nand \U$3173 ( \3843 , \3841 , \3842 );
nor \U$3174 ( \3844 , \3840 , \3843 );
nand \U$3175 ( \3845 , \3839 , \3844 );
not \U$3176 ( \3846 , \3269 );
not \U$3177 ( \3847 , \3071 );
or \U$3178 ( \3848 , \3846 , \3847 );
and \U$3179 ( \3849 , \3259 , \2278 );
nor \U$3180 ( \3850 , \3075 , \2278 );
nor \U$3181 ( \3851 , \3849 , \3850 );
nand \U$3182 ( \3852 , \3848 , \3851 );
and \U$3183 ( \3853 , \3845 , \3852 );
not \U$3184 ( \3854 , \3853 );
or \U$3185 ( \3855 , \3836 , \3854 );
or \U$3186 ( \3856 , \3853 , \3835 );
nand \U$3187 ( \3857 , \3855 , \3856 );
not \U$3188 ( \3858 , \3857 );
or \U$3189 ( \3859 , \3825 , \3858 );
not \U$3190 ( \3860 , \3835 );
nand \U$3191 ( \3861 , \3860 , \3853 );
nand \U$3192 ( \3862 , \3859 , \3861 );
buf \U$3193 ( \3863 , \3862 );
not \U$3194 ( \3864 , \3678 );
not \U$3195 ( \3865 , \2110 );
or \U$3196 ( \3866 , \3864 , \3865 );
or \U$3197 ( \3867 , \3678 , \2110 );
nand \U$3198 ( \3868 , \3866 , \3867 );
not \U$3199 ( \3869 , \3868 );
not \U$3200 ( \3870 , \2442 );
or \U$3201 ( \3871 , \3869 , \3870 );
nand \U$3202 ( \3872 , \3686 , \2164 );
nand \U$3203 ( \3873 , \3871 , \3872 );
not \U$3204 ( \3874 , \3873 );
not \U$3205 ( \3875 , RIaaa4e98_462);
not \U$3206 ( \3876 , \1480 );
or \U$3207 ( \3877 , \3875 , \3876 );
not \U$3208 ( \3878 , \1561 );
not \U$3209 ( \3879 , RIaaa49e8_452);
not \U$3210 ( \3880 , \3879 );
and \U$3211 ( \3881 , \3878 , \3880 );
and \U$3212 ( \3882 , \1502 , RIaaa4b50_455);
nor \U$3213 ( \3883 , \3881 , \3882 );
nand \U$3214 ( \3884 , \3877 , \3883 );
nand \U$3215 ( \3885 , \1413 , RIaaa4e20_461);
nand \U$3216 ( \3886 , \1550 , RIaaa50f0_467);
nand \U$3217 ( \3887 , \1436 , RIaaa4f88_464);
and \U$3218 ( \3888 , \1449 , RIaaa5000_465);
and \U$3219 ( \3889 , RIaaa4c40_457, \1541 );
nor \U$3220 ( \3890 , \3888 , \3889 );
nand \U$3221 ( \3891 , \3885 , \3886 , \3887 , \3890 );
nor \U$3222 ( \3892 , \3884 , \3891 );
and \U$3223 ( \3893 , RIaaa4cb8_458, \1470 );
not \U$3224 ( \3894 , RIaaa4a60_453);
nor \U$3225 ( \3895 , \3894 , \1530 );
nor \U$3226 ( \3896 , \3893 , \3895 );
and \U$3227 ( \3897 , \1516 , RIaaa4f10_463);
not \U$3228 ( \3898 , RIaaa4bc8_456);
not \U$3229 ( \3899 , \1491 );
or \U$3230 ( \3900 , \3898 , \3899 );
nand \U$3231 ( \3901 , \1494 , RIaaa4ad8_454);
nand \U$3232 ( \3902 , \3900 , \3901 );
nor \U$3233 ( \3903 , \3897 , \3902 );
nand \U$3234 ( \3904 , \3896 , \3903 );
and \U$3235 ( \3905 , \1508 , RIaaa5168_468);
and \U$3236 ( \3906 , \1474 , RIaaa4d30_459);
nor \U$3237 ( \3907 , \3905 , \3906 );
nand \U$3238 ( \3908 , \2199 , RIaaa4da8_460);
nand \U$3239 ( \3909 , \1458 , RIaaa5078_466);
nand \U$3240 ( \3910 , \3907 , \3908 , \3909 );
nor \U$3241 ( \3911 , \3904 , \3910 );
nand \U$3242 ( \3912 , \3892 , \3911 );
not \U$3243 ( \3913 , \3912 );
buf \U$3244 ( \3914 , \3913 );
not \U$3245 ( \3915 , \3914 );
nand \U$3246 ( \3916 , \2448 , \3915 );
not \U$3247 ( \3917 , \3916 );
and \U$3248 ( \3918 , \3874 , \3917 );
and \U$3249 ( \3919 , \3873 , \3916 );
nor \U$3250 ( \3920 , \3918 , \3919 );
not \U$3251 ( \3921 , \3920 );
and \U$3252 ( \3922 , \3863 , \3921 );
not \U$3253 ( \3923 , \3873 );
nor \U$3254 ( \3924 , \3923 , \3916 );
nor \U$3255 ( \3925 , \3922 , \3924 );
xor \U$3256 ( \3926 , \3813 , \3925 );
not \U$3257 ( \3927 , \3787 );
not \U$3258 ( \3928 , \3768 );
not \U$3259 ( \3929 , \3928 );
and \U$3260 ( \3930 , \3927 , \3929 );
and \U$3261 ( \3931 , \3787 , \3928 );
nor \U$3262 ( \3932 , \3930 , \3931 );
xor \U$3263 ( \3933 , \3701 , \3718 );
xor \U$3264 ( \3934 , \3933 , \3729 );
not \U$3265 ( \3935 , \3934 );
nand \U$3266 ( \3936 , \3932 , \3935 );
not \U$3267 ( \3937 , \3212 );
not \U$3268 ( \3938 , \3341 );
or \U$3269 ( \3939 , \3937 , \3938 );
not \U$3270 ( \3940 , \3764 );
not \U$3271 ( \3941 , \3512 );
and \U$3272 ( \3942 , \3940 , \3941 );
and \U$3273 ( \3943 , \1900 , \3684 );
nor \U$3274 ( \3944 , \3942 , \3943 );
nand \U$3275 ( \3945 , \3939 , \3944 );
not \U$3276 ( \3946 , \3945 );
not \U$3277 ( \3947 , \2405 );
not \U$3278 ( \3948 , \2907 );
and \U$3279 ( \3949 , \3947 , \3948 );
not \U$3280 ( \3950 , \2907 );
not \U$3281 ( \3951 , \2572 );
or \U$3282 ( \3952 , \3950 , \3951 );
and \U$3283 ( \3953 , \2916 , \2495 );
not \U$3284 ( \3954 , \2916 );
and \U$3285 ( \3955 , \3954 , \2498 );
nor \U$3286 ( \3956 , \3953 , \3955 );
nand \U$3287 ( \3957 , \3952 , \3956 );
nor \U$3288 ( \3958 , \3949 , \3957 );
not \U$3289 ( \3959 , \3958 );
not \U$3290 ( \3960 , \3706 );
not \U$3291 ( \3961 , \3708 );
nor \U$3292 ( \3962 , \3961 , \3716 );
not \U$3293 ( \3963 , \3962 );
or \U$3294 ( \3964 , \3960 , \3963 );
not \U$3295 ( \3965 , \3706 );
not \U$3296 ( \3966 , \3716 );
nand \U$3297 ( \3967 , \3966 , \3708 );
nand \U$3298 ( \3968 , \3965 , \3967 );
nand \U$3299 ( \3969 , \3964 , \3968 );
not \U$3300 ( \3970 , \3969 );
or \U$3301 ( \3971 , \3959 , \3970 );
or \U$3302 ( \3972 , \3969 , \3958 );
nand \U$3303 ( \3973 , \3971 , \3972 );
not \U$3304 ( \3974 , \3973 );
or \U$3305 ( \3975 , \3946 , \3974 );
not \U$3306 ( \3976 , \3958 );
nand \U$3307 ( \3977 , \3976 , \3969 );
nand \U$3308 ( \3978 , \3975 , \3977 );
buf \U$3309 ( \3979 , \3978 );
and \U$3310 ( \3980 , \3936 , \3979 );
nor \U$3311 ( \3981 , \3932 , \3935 );
nor \U$3312 ( \3982 , \3980 , \3981 );
and \U$3313 ( \3983 , \3926 , \3982 );
and \U$3314 ( \3984 , \3813 , \3925 );
or \U$3315 ( \3985 , \3983 , \3984 );
xor \U$3316 ( \3986 , \3808 , \3985 );
xor \U$3317 ( \3987 , \3735 , \3741 );
xor \U$3318 ( \3988 , \3987 , \3795 );
and \U$3319 ( \3989 , \3986 , \3988 );
and \U$3320 ( \3990 , \3808 , \3985 );
or \U$3321 ( \3991 , \3989 , \3990 );
nand \U$3322 ( \3992 , \3806 , \3991 );
xor \U$3323 ( \3993 , \3048 , \3356 );
xor \U$3324 ( \3994 , \3993 , \3392 );
not \U$3325 ( \3995 , \3994 );
not \U$3326 ( \3996 , \3629 );
not \U$3327 ( \3997 , \3996 );
not \U$3328 ( \3998 , \3802 );
or \U$3329 ( \3999 , \3997 , \3998 );
not \U$3330 ( \4000 , \3637 );
nand \U$3331 ( \4001 , \4000 , \3798 );
nand \U$3332 ( \4002 , \3999 , \4001 );
nand \U$3333 ( \4003 , \3995 , \4002 );
nand \U$3334 ( \4004 , \3992 , \4003 );
not \U$3335 ( \4005 , \4004 );
xor \U$3336 ( \4006 , \3808 , \3985 );
xor \U$3337 ( \4007 , \4006 , \3988 );
xor \U$3338 ( \4008 , \3813 , \3925 );
xor \U$3339 ( \4009 , \4008 , \3982 );
not \U$3340 ( \4010 , \4009 );
not \U$3341 ( \4011 , \3753 );
not \U$3342 ( \4012 , \3792 );
or \U$3343 ( \4013 , \4011 , \4012 );
or \U$3344 ( \4014 , \3753 , \3792 );
nand \U$3345 ( \4015 , \4013 , \4014 );
not \U$3346 ( \4016 , \3748 );
xnor \U$3347 ( \4017 , \4015 , \4016 );
not \U$3348 ( \4018 , \4017 );
not \U$3349 ( \4019 , \3945 );
not \U$3350 ( \4020 , \3973 );
not \U$3351 ( \4021 , \4020 );
or \U$3352 ( \4022 , \4019 , \4021 );
not \U$3353 ( \4023 , \3945 );
nand \U$3354 ( \4024 , \4023 , \3973 );
nand \U$3355 ( \4025 , \4022 , \4024 );
not \U$3356 ( \4026 , \4025 );
not \U$3357 ( \4027 , \3857 );
and \U$3358 ( \4028 , \3824 , \4027 );
not \U$3359 ( \4029 , \3824 );
and \U$3360 ( \4030 , \4029 , \3857 );
or \U$3361 ( \4031 , \4028 , \4030 );
not \U$3362 ( \4032 , \4031 );
or \U$3363 ( \4033 , \4026 , \4032 );
or \U$3364 ( \4034 , \4025 , \4031 );
not \U$3365 ( \4035 , \2994 );
not \U$3366 ( \4036 , \3677 );
nor \U$3367 ( \4037 , \1897 , \4036 );
not \U$3368 ( \4038 , \4037 );
or \U$3369 ( \4039 , \4035 , \4038 );
nor \U$3370 ( \4040 , \1898 , \3678 );
and \U$3371 ( \4041 , \2994 , \4040 );
buf \U$3372 ( \4042 , \3209 );
nor \U$3373 ( \4043 , \3513 , \4042 );
not \U$3374 ( \4044 , \4043 );
not \U$3375 ( \4045 , \2234 );
or \U$3376 ( \4046 , \4044 , \4045 );
nor \U$3377 ( \4047 , \1940 , \3210 );
nand \U$3378 ( \4048 , \2234 , \4047 );
nand \U$3379 ( \4049 , \4046 , \4048 );
nor \U$3380 ( \4050 , \4041 , \4049 );
nand \U$3381 ( \4051 , \4039 , \4050 );
not \U$3382 ( \4052 , \2406 );
not \U$3383 ( \4053 , \3156 );
or \U$3384 ( \4054 , \4052 , \4053 );
not \U$3385 ( \4055 , \3157 );
and \U$3386 ( \4056 , \2390 , \4055 );
nand \U$3387 ( \4057 , \2366 , \2310 );
not \U$3388 ( \4058 , \4057 );
not \U$3389 ( \4059 , \4058 );
not \U$3390 ( \4060 , \2906 );
not \U$3391 ( \4061 , \4060 );
or \U$3392 ( \4062 , \4059 , \4061 );
or \U$3393 ( \4063 , \2400 , \2908 );
nand \U$3394 ( \4064 , \4062 , \4063 );
nor \U$3395 ( \4065 , \4056 , \4064 );
nand \U$3396 ( \4066 , \4054 , \4065 );
xor \U$3397 ( \4067 , \4051 , \4066 );
not \U$3398 ( \4068 , \3852 );
not \U$3399 ( \4069 , \4068 );
buf \U$3400 ( \4070 , \3845 );
not \U$3401 ( \4071 , \4070 );
or \U$3402 ( \4072 , \4069 , \4071 );
or \U$3403 ( \4073 , \4070 , \4068 );
nand \U$3404 ( \4074 , \4072 , \4073 );
and \U$3405 ( \4075 , \4067 , \4074 );
and \U$3406 ( \4076 , \4051 , \4066 );
or \U$3407 ( \4077 , \4075 , \4076 );
buf \U$3408 ( \4078 , \4077 );
nand \U$3409 ( \4079 , \4034 , \4078 );
nand \U$3410 ( \4080 , \4033 , \4079 );
not \U$3411 ( \4081 , \3862 );
not \U$3412 ( \4082 , \3920 );
and \U$3413 ( \4083 , \4081 , \4082 );
and \U$3414 ( \4084 , \3920 , \3862 );
nor \U$3415 ( \4085 , \4083 , \4084 );
not \U$3416 ( \4086 , \4085 );
nand \U$3417 ( \4087 , \4080 , \4086 );
not \U$3418 ( \4088 , \2153 );
not \U$3419 ( \4089 , \2515 );
or \U$3420 ( \4090 , \4088 , \4089 );
and \U$3421 ( \4091 , \2210 , \2521 );
not \U$3422 ( \4092 , \2210 );
and \U$3423 ( \4093 , \4092 , \2951 );
nor \U$3424 ( \4094 , \4091 , \4093 );
nand \U$3425 ( \4095 , \4090 , \4094 );
nor \U$3426 ( \4096 , \2943 , \2153 );
nor \U$3427 ( \4097 , \4095 , \4096 );
not \U$3428 ( \4098 , \4097 );
not \U$3429 ( \4099 , \2225 );
not \U$3430 ( \4100 , \3038 );
or \U$3431 ( \4101 , \4099 , \4100 );
and \U$3432 ( \4102 , \3026 , \2210 );
and \U$3433 ( \4103 , \1936 , \3031 );
not \U$3434 ( \4104 , \1936 );
and \U$3435 ( \4105 , \4104 , \3250 );
or \U$3436 ( \4106 , \4103 , \4105 );
nor \U$3437 ( \4107 , \4102 , \4106 );
nand \U$3438 ( \4108 , \4101 , \4107 );
not \U$3439 ( \4109 , \1988 );
not \U$3440 ( \4110 , \3071 );
or \U$3441 ( \4111 , \4109 , \4110 );
and \U$3442 ( \4112 , \3259 , \2363 );
nor \U$3443 ( \4113 , \3077 , \2363 );
nor \U$3444 ( \4114 , \4112 , \4113 );
nand \U$3445 ( \4115 , \4111 , \4114 );
nand \U$3446 ( \4116 , \4108 , \4115 );
not \U$3447 ( \4117 , \4116 );
or \U$3448 ( \4118 , \4098 , \4117 );
nand \U$3449 ( \4119 , \3723 , \2916 );
nand \U$3450 ( \4120 , \3815 , \2915 );
and \U$3451 ( \4121 , \3301 , \1584 );
not \U$3452 ( \4122 , \3301 );
and \U$3453 ( \4123 , \4122 , \1579 );
nor \U$3454 ( \4124 , \4121 , \4123 );
nand \U$3455 ( \4125 , \4119 , \4120 , \4124 );
nand \U$3456 ( \4126 , \4118 , \4125 );
or \U$3457 ( \4127 , \4116 , \4097 );
nand \U$3458 ( \4128 , \4126 , \4127 );
not \U$3459 ( \4129 , \3914 );
not \U$3460 ( \4130 , \2160 );
or \U$3461 ( \4131 , \4129 , \4130 );
or \U$3462 ( \4132 , \2640 , \3914 );
nand \U$3463 ( \4133 , \4131 , \4132 );
nand \U$3464 ( \4134 , \4133 , \2102 );
nand \U$3465 ( \4135 , \3868 , \2163 );
nand \U$3466 ( \4136 , \4134 , \4135 );
not \U$3467 ( \4137 , \4136 );
not \U$3468 ( \4138 , RIaaa5e10_495);
not \U$3469 ( \4139 , \1501 );
or \U$3470 ( \4140 , \4138 , \4139 );
nand \U$3471 ( \4141 , \1511 , RIaaa5ca8_492);
nand \U$3472 ( \4142 , \4140 , \4141 );
not \U$3473 ( \4143 , \1479 );
not \U$3474 ( \4144 , RIaaa59d8_486);
nor \U$3475 ( \4145 , \4143 , \4144 );
nor \U$3476 ( \4146 , \4142 , \4145 );
not \U$3477 ( \4147 , \1426 );
not \U$3478 ( \4148 , RIaaa60e0_501);
not \U$3479 ( \4149 , \4148 );
and \U$3480 ( \4150 , \4147 , \4149 );
nor \U$3481 ( \4151 , \1386 , \1396 );
nand \U$3482 ( \4152 , \4151 , \1433 );
not \U$3483 ( \4153 , RIaaa5b40_489);
nor \U$3484 ( \4154 , \4152 , \4153 );
nor \U$3485 ( \4155 , \4150 , \4154 );
and \U$3486 ( \4156 , \1953 , RIaaa5a50_487);
not \U$3487 ( \4157 , RIaaa5f00_497);
not \U$3488 ( \4158 , \1443 );
or \U$3489 ( \4159 , \4157 , \4158 );
nand \U$3490 ( \4160 , \2881 , RIaaa5bb8_490);
nand \U$3491 ( \4161 , \4159 , \4160 );
nor \U$3492 ( \4162 , \4156 , \4161 );
and \U$3493 ( \4163 , \4146 , \4155 , \4162 );
nand \U$3494 ( \4164 , \1564 , RIaaa6158_502);
nand \U$3495 ( \4165 , \1470 , RIaaa5f78_498);
nand \U$3496 ( \4166 , \1431 , \1396 , \1433 );
not \U$3497 ( \4167 , \4166 );
and \U$3498 ( \4168 , \4167 , RIaaa5ac8_488);
not \U$3499 ( \4169 , RIaaa5e88_496);
not \U$3500 ( \4170 , \1491 );
or \U$3501 ( \4171 , \4169 , \4170 );
nand \U$3502 ( \4172 , \1494 , RIaaa5d98_494);
nand \U$3503 ( \4173 , \4171 , \4172 );
nor \U$3504 ( \4174 , \4168 , \4173 );
nand \U$3505 ( \4175 , \4164 , \4165 , \4174 );
and \U$3506 ( \4176 , \1440 , \1472 );
nand \U$3507 ( \4177 , \1557 , \4176 );
not \U$3508 ( \4178 , \4177 );
not \U$3509 ( \4179 , RIaaa5ff0_499);
not \U$3510 ( \4180 , \4179 );
and \U$3511 ( \4181 , \4178 , \4180 );
and \U$3512 ( \4182 , \1482 , RIaaa5d20_493);
nor \U$3513 ( \4183 , \4181 , \4182 );
nand \U$3514 ( \4184 , \1461 , RIaaa6068_500);
not \U$3515 ( \4185 , \1396 );
and \U$3516 ( \4186 , \1386 , \4185 , \1456 );
nand \U$3517 ( \4187 , \4186 , RIaaa5c30_491);
nand \U$3518 ( \4188 , \4183 , \4184 , \4187 );
nor \U$3519 ( \4189 , \4175 , \4188 );
nand \U$3520 ( \4190 , \4163 , \4189 );
buf \U$3521 ( \4191 , \4190 );
buf \U$3522 ( \4192 , \4191 );
not \U$3523 ( \4193 , \4192 );
buf \U$3524 ( \4194 , \4193 );
not \U$3525 ( \4195 , \4194 );
nand \U$3526 ( \4196 , \2448 , \4195 );
not \U$3527 ( \4197 , \4196 );
and \U$3528 ( \4198 , \4137 , \4197 );
and \U$3529 ( \4199 , \4136 , \4196 );
nor \U$3530 ( \4200 , \4198 , \4199 );
not \U$3531 ( \4201 , \4200 );
and \U$3532 ( \4202 , \4128 , \4201 );
and \U$3533 ( \4203 , \4134 , \4135 );
nor \U$3534 ( \4204 , \4203 , \4196 );
nor \U$3535 ( \4205 , \4202 , \4204 );
buf \U$3536 ( \4206 , \4205 );
and \U$3537 ( \4207 , \4087 , \4206 );
nor \U$3538 ( \4208 , \4080 , \4086 );
nor \U$3539 ( \4209 , \4207 , \4208 );
not \U$3540 ( \4210 , \4209 );
or \U$3541 ( \4211 , \4018 , \4210 );
and \U$3542 ( \4212 , \4087 , \4206 );
nor \U$3543 ( \4213 , \4212 , \4208 );
or \U$3544 ( \4214 , \4213 , \4017 );
nand \U$3545 ( \4215 , \4211 , \4214 );
not \U$3546 ( \4216 , \4215 );
or \U$3547 ( \4217 , \4010 , \4216 );
not \U$3548 ( \4218 , \4213 );
nand \U$3549 ( \4219 , \4218 , \4017 );
nand \U$3550 ( \4220 , \4217 , \4219 );
nand \U$3551 ( \4221 , \4007 , \4220 );
not \U$3552 ( \4222 , \4221 );
not \U$3553 ( \4223 , \4222 );
not \U$3554 ( \4224 , \4009 );
not \U$3555 ( \4225 , \4224 );
not \U$3556 ( \4226 , \4215 );
or \U$3557 ( \4227 , \4225 , \4226 );
or \U$3558 ( \4228 , \4224 , \4215 );
nand \U$3559 ( \4229 , \4227 , \4228 );
not \U$3560 ( \4230 , \4080 );
not \U$3561 ( \4231 , \4205 );
not \U$3562 ( \4232 , \4085 );
not \U$3563 ( \4233 , \4232 );
or \U$3564 ( \4234 , \4231 , \4233 );
not \U$3565 ( \4235 , \4085 );
or \U$3566 ( \4236 , \4235 , \4205 );
nand \U$3567 ( \4237 , \4234 , \4236 );
not \U$3568 ( \4238 , \4237 );
or \U$3569 ( \4239 , \4230 , \4238 );
buf \U$3570 ( \4240 , \4080 );
or \U$3571 ( \4241 , \4237 , \4240 );
nand \U$3572 ( \4242 , \4239 , \4241 );
not \U$3573 ( \4243 , \4242 );
not \U$3574 ( \4244 , \4128 );
not \U$3575 ( \4245 , \4200 );
or \U$3576 ( \4246 , \4244 , \4245 );
or \U$3577 ( \4247 , \4128 , \4200 );
nand \U$3578 ( \4248 , \4246 , \4247 );
not \U$3579 ( \4249 , \4248 );
not \U$3580 ( \4250 , \2486 );
and \U$3581 ( \4251 , \1187 , \1193 );
not \U$3582 ( \4252 , \4251 );
or \U$3583 ( \4253 , \4250 , \4252 );
not \U$3584 ( \4254 , \2485 );
and \U$3585 ( \4255 , \2822 , \4254 );
and \U$3586 ( \4256 , \2150 , \2520 );
not \U$3587 ( \4257 , \2150 );
not \U$3588 ( \4258 , \1183 );
nand \U$3589 ( \4259 , \4258 , \1189 );
and \U$3590 ( \4260 , \4257 , \4259 );
nor \U$3591 ( \4261 , \4256 , \4260 );
nor \U$3592 ( \4262 , \4255 , \4261 );
nand \U$3593 ( \4263 , \4253 , \4262 );
not \U$3594 ( \4264 , \4263 );
not \U$3595 ( \4265 , \4264 );
not \U$3596 ( \4266 , \1590 );
not \U$3597 ( \4267 , \2907 );
and \U$3598 ( \4268 , \4266 , \4267 );
not \U$3599 ( \4269 , \2907 );
not \U$3600 ( \4270 , \2285 );
or \U$3601 ( \4271 , \4269 , \4270 );
and \U$3602 ( \4272 , \2914 , \1582 );
not \U$3603 ( \4273 , \2914 );
not \U$3604 ( \4274 , \1363 );
nand \U$3605 ( \4275 , \4274 , \1575 );
not \U$3606 ( \4276 , \4275 );
and \U$3607 ( \4277 , \4273 , \4276 );
nor \U$3608 ( \4278 , \4272 , \4277 );
nand \U$3609 ( \4279 , \4271 , \4278 );
nor \U$3610 ( \4280 , \4268 , \4279 );
not \U$3611 ( \4281 , \4280 );
or \U$3612 ( \4282 , \4265 , \4281 );
not \U$3613 ( \4283 , \2152 );
not \U$3614 ( \4284 , \3038 );
or \U$3615 ( \4285 , \4283 , \4284 );
nor \U$3616 ( \4286 , \2749 , \2758 );
and \U$3617 ( \4287 , \4286 , \2151 );
or \U$3618 ( \4288 , \3248 , \2209 );
nand \U$3619 ( \4289 , \2754 , \2209 );
nand \U$3620 ( \4290 , \4288 , \4289 );
nor \U$3621 ( \4291 , \4287 , \4290 );
nand \U$3622 ( \4292 , \4285 , \4291 );
not \U$3623 ( \4293 , \1936 );
not \U$3624 ( \4294 , \3071 );
or \U$3625 ( \4295 , \4293 , \4294 );
not \U$3626 ( \4296 , \3068 );
not \U$3627 ( \4297 , \1994 );
or \U$3628 ( \4298 , \4296 , \4297 );
nand \U$3629 ( \4299 , \4298 , \3020 );
nand \U$3630 ( \4300 , \4295 , \4299 );
not \U$3631 ( \4301 , \1985 );
nand \U$3632 ( \4302 , \4301 , \3019 );
and \U$3633 ( \4303 , \4302 , \3068 );
nor \U$3634 ( \4304 , \4303 , \3071 );
nor \U$3635 ( \4305 , \4300 , \4304 );
and \U$3636 ( \4306 , \4292 , \4305 );
nand \U$3637 ( \4307 , \4282 , \4306 );
not \U$3638 ( \4308 , \4307 );
not \U$3639 ( \4309 , \2447 );
nand \U$3640 ( \4310 , \1470 , RIaaa6d10_527);
and \U$3641 ( \4311 , \4167 , RIaaa6a40_521);
not \U$3642 ( \4312 , RIaaa7058_534);
not \U$3643 ( \4313 , \1491 );
or \U$3644 ( \4314 , \4312 , \4313 );
nand \U$3645 ( \4315 , \1494 , RIaaa7148_536);
nand \U$3646 ( \4316 , \4314 , \4315 );
nor \U$3647 ( \4317 , \4311 , \4316 );
nand \U$3648 ( \4318 , \1564 , RIaaa6e00_529);
and \U$3649 ( \4319 , \4310 , \4317 , \4318 );
and \U$3650 ( \4320 , \4186 , RIaaa6ba8_524);
and \U$3651 ( \4321 , \1461 , RIaaa6e78_530);
nor \U$3652 ( \4322 , \4320 , \4321 );
not \U$3653 ( \4323 , \4177 );
not \U$3654 ( \4324 , RIaaa6c98_526);
not \U$3655 ( \4325 , \4324 );
and \U$3656 ( \4326 , \4323 , \4325 );
and \U$3657 ( \4327 , \1927 , RIaaa6f68_532);
nor \U$3658 ( \4328 , \4326 , \4327 );
nand \U$3659 ( \4329 , \4319 , \4322 , \4328 );
not \U$3660 ( \4330 , RIaaa6ab8_522);
not \U$3661 ( \4331 , \1953 );
or \U$3662 ( \4332 , \4330 , \4331 );
not \U$3663 ( \4333 , \2173 );
not \U$3664 ( \4334 , RIaaa70d0_535);
nor \U$3665 ( \4335 , \4333 , \4334 );
not \U$3666 ( \4336 , \2881 );
not \U$3667 ( \4337 , RIaaa6c20_525);
nor \U$3668 ( \4338 , \4336 , \4337 );
nor \U$3669 ( \4339 , \4335 , \4338 );
nand \U$3670 ( \4340 , \4332 , \4339 );
not \U$3671 ( \4341 , RIaaa69c8_520);
not \U$3672 ( \4342 , \1434 );
or \U$3673 ( \4343 , \4341 , \4342 );
nand \U$3674 ( \4344 , \1550 , RIaaa6d88_528);
nand \U$3675 ( \4345 , \4343 , \4344 );
nor \U$3676 ( \4346 , \4340 , \4345 );
not \U$3677 ( \4347 , RIaaa6fe0_533);
not \U$3678 ( \4348 , \1502 );
or \U$3679 ( \4349 , \4347 , \4348 );
nand \U$3680 ( \4350 , \1512 , RIaaa6ef0_531);
nand \U$3681 ( \4351 , \4349 , \4350 );
not \U$3682 ( \4352 , RIaaa6b30_523);
nor \U$3683 ( \4353 , \4352 , \4143 );
nor \U$3684 ( \4354 , \4351 , \4353 );
nand \U$3685 ( \4355 , \4346 , \4354 );
nor \U$3686 ( \4356 , \4329 , \4355 );
buf \U$3687 ( \4357 , \4356 );
buf \U$3688 ( \4358 , \4357 );
buf \U$3689 ( \4359 , \4358 );
not \U$3690 ( \4360 , \4359 );
and \U$3691 ( \4361 , \4309 , \4360 );
not \U$3692 ( \4362 , \4264 );
not \U$3693 ( \4363 , \4280 );
and \U$3694 ( \4364 , \4362 , \4363 );
nor \U$3695 ( \4365 , \4361 , \4364 );
not \U$3696 ( \4366 , \4365 );
or \U$3697 ( \4367 , \4308 , \4366 );
not \U$3698 ( \4368 , \2442 );
not \U$3699 ( \4369 , \4194 );
not \U$3700 ( \4370 , \2110 );
or \U$3701 ( \4371 , \4369 , \4370 );
not \U$3702 ( \4372 , \4191 );
buf \U$3703 ( \4373 , \4372 );
or \U$3704 ( \4374 , \2110 , \4373 );
nand \U$3705 ( \4375 , \4371 , \4374 );
not \U$3706 ( \4376 , \4375 );
or \U$3707 ( \4377 , \4368 , \4376 );
nand \U$3708 ( \4378 , \4133 , \2164 );
nand \U$3709 ( \4379 , \4377 , \4378 );
nand \U$3710 ( \4380 , \4367 , \4379 );
nand \U$3711 ( \4381 , \4249 , \4380 );
not \U$3712 ( \4382 , \4097 );
not \U$3713 ( \4383 , \4116 );
or \U$3714 ( \4384 , \4382 , \4383 );
nand \U$3715 ( \4385 , \4384 , \4127 );
not \U$3716 ( \4386 , \4125 );
xor \U$3717 ( \4387 , \4385 , \4386 );
not \U$3718 ( \4388 , \3212 );
not \U$3719 ( \4389 , \2582 );
or \U$3720 ( \4390 , \4388 , \4389 );
and \U$3721 ( \4391 , \3211 , \2572 );
not \U$3722 ( \4392 , \2310 );
nand \U$3723 ( \4393 , \4392 , \2366 );
or \U$3724 ( \4394 , \4393 , \3156 );
nand \U$3725 ( \4395 , \4058 , \3156 );
nand \U$3726 ( \4396 , \4394 , \4395 );
nor \U$3727 ( \4397 , \4391 , \4396 );
nand \U$3728 ( \4398 , \4390 , \4397 );
not \U$3729 ( \4399 , \4398 );
not \U$3730 ( \4400 , \1942 );
not \U$3731 ( \4401 , \3678 );
and \U$3732 ( \4402 , \4400 , \4401 );
not \U$3733 ( \4403 , \3913 );
not \U$3734 ( \4404 , \4403 );
not \U$3735 ( \4405 , \1896 );
or \U$3736 ( \4406 , \4404 , \4405 );
or \U$3737 ( \4407 , \4403 , \3513 );
nand \U$3738 ( \4408 , \4406 , \4407 );
and \U$3739 ( \4409 , \2994 , \4408 );
nor \U$3740 ( \4410 , \4402 , \4409 );
not \U$3741 ( \4411 , \3679 );
nand \U$3742 ( \4412 , \4411 , \1992 );
nand \U$3743 ( \4413 , \4410 , \4412 );
not \U$3744 ( \4414 , \4413 );
or \U$3745 ( \4415 , \4399 , \4414 );
xor \U$3746 ( \4416 , \4108 , \4115 );
not \U$3747 ( \4417 , \4416 );
nand \U$3748 ( \4418 , \4415 , \4417 );
or \U$3749 ( \4419 , \4413 , \4398 );
nand \U$3750 ( \4420 , \4418 , \4419 );
not \U$3751 ( \4421 , \4420 );
or \U$3752 ( \4422 , \4387 , \4421 );
xor \U$3753 ( \4423 , \4051 , \4066 );
xor \U$3754 ( \4424 , \4423 , \4074 );
nand \U$3755 ( \4425 , \4422 , \4424 );
nand \U$3756 ( \4426 , \4387 , \4421 );
nand \U$3757 ( \4427 , \4425 , \4426 );
and \U$3758 ( \4428 , \4381 , \4427 );
not \U$3759 ( \4429 , \4248 );
nor \U$3760 ( \4430 , \4429 , \4380 );
nor \U$3761 ( \4431 , \4428 , \4430 );
not \U$3762 ( \4432 , \4431 );
xor \U$3763 ( \4433 , \3934 , \3978 );
xnor \U$3764 ( \4434 , \4433 , \3932 );
not \U$3765 ( \4435 , \4434 );
or \U$3766 ( \4436 , \4432 , \4435 );
or \U$3767 ( \4437 , \4431 , \4434 );
nand \U$3768 ( \4438 , \4436 , \4437 );
not \U$3769 ( \4439 , \4438 );
or \U$3770 ( \4440 , \4243 , \4439 );
not \U$3771 ( \4441 , \4434 );
nand \U$3772 ( \4442 , \4441 , \4431 );
nand \U$3773 ( \4443 , \4440 , \4442 );
nand \U$3774 ( \4444 , \4229 , \4443 );
and \U$3775 ( \4445 , \4005 , \4223 , \4444 );
not \U$3776 ( \4446 , \4445 );
xor \U$3777 ( \4447 , \4248 , \4380 );
xnor \U$3778 ( \4448 , \4447 , \4427 );
not \U$3779 ( \4449 , \4448 );
xor \U$3780 ( \4450 , \4077 , \4031 );
xnor \U$3781 ( \4451 , \4450 , \4025 );
not \U$3782 ( \4452 , \4451 );
not \U$3783 ( \4453 , \2447 );
and \U$3784 ( \4454 , \1951 , RIaaa8408_576);
not \U$3785 ( \4455 , RIaaa87c8_584);
nor \U$3786 ( \4456 , \4455 , \1426 );
nor \U$3787 ( \4457 , \4454 , \4456 );
and \U$3788 ( \4458 , \2199 , RIaaa84f8_578);
not \U$3789 ( \4459 , RIaaa8390_575);
not \U$3790 ( \4460 , \2881 );
or \U$3791 ( \4461 , \4459 , \4460 );
nand \U$3792 ( \4462 , \1541 , RIaaa8318_574);
nand \U$3793 ( \4463 , \4461 , \4462 );
nor \U$3794 ( \4464 , \4458 , \4463 );
and \U$3795 ( \4465 , \4457 , \4464 );
nand \U$3796 ( \4466 , \1413 , RIaaa8660_581);
nand \U$3797 ( \4467 , RIaaa8228_572, \1502 );
nand \U$3798 ( \4468 , \1512 , RIaaa88b8_586);
and \U$3799 ( \4469 , \4466 , \4467 , \4468 );
not \U$3800 ( \4470 , \1530 );
not \U$3801 ( \4471 , RIaaa8930_587);
not \U$3802 ( \4472 , \4471 );
and \U$3803 ( \4473 , \4470 , \4472 );
and \U$3804 ( \4474 , \1470 , RIaaa8750_583);
nor \U$3805 ( \4475 , \4473 , \4474 );
nand \U$3806 ( \4476 , \1458 , RIaaa8480_577);
and \U$3807 ( \4477 , \1508 , RIaaa8840_585);
buf \U$3808 ( \4478 , \1473 );
and \U$3809 ( \4479 , \4478 , RIaaa86d8_582);
nor \U$3810 ( \4480 , \4477 , \4479 );
and \U$3811 ( \4481 , \4475 , \4476 , \4480 );
and \U$3812 ( \4482 , \1480 , RIaaa85e8_580);
not \U$3813 ( \4483 , RIaaa8570_579);
not \U$3814 ( \4484 , \4167 );
or \U$3815 ( \4485 , \4483 , \4484 );
and \U$3816 ( \4486 , \1491 , RIaaa82a0_573);
not \U$3817 ( \4487 , RIaaa81b0_571);
nor \U$3818 ( \4488 , \4487 , \1495 );
nor \U$3819 ( \4489 , \4486 , \4488 );
nand \U$3820 ( \4490 , \4485 , \4489 );
nor \U$3821 ( \4491 , \4482 , \4490 );
nand \U$3822 ( \4492 , \4465 , \4469 , \4481 , \4491 );
buf \U$3823 ( \4493 , \4492 );
not \U$3824 ( \4494 , \4493 );
not \U$3825 ( \4495 , \4494 );
and \U$3826 ( \4496 , \4453 , \4495 );
not \U$3827 ( \4497 , \2907 );
nand \U$3828 ( \4498 , \4497 , \2508 );
and \U$3829 ( \4499 , \2822 , \2907 );
not \U$3830 ( \4500 , \2830 );
not \U$3831 ( \4501 , \2915 );
or \U$3832 ( \4502 , \4500 , \4501 );
or \U$3833 ( \4503 , \2833 , \2689 );
nand \U$3834 ( \4504 , \4502 , \4503 );
nor \U$3835 ( \4505 , \4499 , \4504 );
nand \U$3836 ( \4506 , \4498 , \4505 );
not \U$3837 ( \4507 , \2210 );
not \U$3838 ( \4508 , \3071 );
or \U$3839 ( \4509 , \4507 , \4508 );
and \U$3840 ( \4510 , \3259 , \1937 );
nor \U$3841 ( \4511 , \3077 , \1937 );
nor \U$3842 ( \4512 , \4510 , \4511 );
nand \U$3843 ( \4513 , \4509 , \4512 );
and \U$3844 ( \4514 , \4506 , \4513 );
nor \U$3845 ( \4515 , \4496 , \4514 );
not \U$3846 ( \4516 , \4513 );
nand \U$3847 ( \4517 , \4516 , \4505 , \4498 );
not \U$3848 ( \4518 , \3301 );
not \U$3849 ( \4519 , \3026 );
or \U$3850 ( \4520 , \4518 , \4519 );
buf \U$3851 ( \4521 , \3029 );
and \U$3852 ( \4522 , \2152 , \4521 );
not \U$3853 ( \4523 , \2152 );
and \U$3854 ( \4524 , \4523 , \3033 );
nor \U$3855 ( \4525 , \4522 , \4524 );
nand \U$3856 ( \4526 , \4520 , \4525 );
not \U$3857 ( \4527 , \4526 );
nand \U$3858 ( \4528 , \3038 , \2991 );
nand \U$3859 ( \4529 , \4527 , \4528 );
nand \U$3860 ( \4530 , \4517 , \4529 );
nand \U$3861 ( \4531 , \4515 , \4530 );
not \U$3862 ( \4532 , \3175 );
not \U$3863 ( \4533 , RIaaa7670_547);
not \U$3864 ( \4534 , \4533 );
and \U$3865 ( \4535 , \4532 , \4534 );
and \U$3866 ( \4536 , \1502 , RIaaa7238_538);
nor \U$3867 ( \4537 , \4535 , \4536 );
and \U$3868 ( \4538 , \1436 , RIaaa7490_543);
not \U$3869 ( \4539 , RIaaa75f8_546);
nor \U$3870 ( \4540 , \4539 , \4143 );
nor \U$3871 ( \4541 , \4538 , \4540 );
not \U$3872 ( \4542 , \1559 );
not \U$3873 ( \4543 , RIaaa78c8_552);
not \U$3874 ( \4544 , \4543 );
and \U$3875 ( \4545 , \4542 , \4544 );
not \U$3876 ( \4546 , RIaaa7328_540);
not \U$3877 ( \4547 , \2173 );
or \U$3878 ( \4548 , \4546 , \4547 );
nand \U$3879 ( \4549 , \2881 , RIaaa73a0_541);
nand \U$3880 ( \4550 , \4548 , \4549 );
nor \U$3881 ( \4551 , \4545 , \4550 );
nand \U$3882 ( \4552 , \1550 , RIaaa77d8_550);
nand \U$3883 ( \4553 , \4537 , \4541 , \4551 , \4552 );
nand \U$3884 ( \4554 , \1564 , RIaaa7850_551);
nand \U$3885 ( \4555 , \4478 , RIaaa76e8_548);
and \U$3886 ( \4556 , \4167 , RIaaa7580_545);
not \U$3887 ( \4557 , RIaaa72b0_539);
not \U$3888 ( \4558 , \1491 );
or \U$3889 ( \4559 , \4557 , \4558 );
nand \U$3890 ( \4560 , \1494 , RIaaa71c0_537);
nand \U$3891 ( \4561 , \4559 , \4560 );
nor \U$3892 ( \4562 , \4556 , \4561 );
nand \U$3893 ( \4563 , \4554 , \4555 , \4562 );
not \U$3894 ( \4564 , \4563 );
not \U$3895 ( \4565 , \1460 );
not \U$3896 ( \4566 , RIaaa7508_544);
not \U$3897 ( \4567 , \4566 );
and \U$3898 ( \4568 , \4565 , \4567 );
and \U$3899 ( \4569 , \4186 , RIaaa7418_542);
nor \U$3900 ( \4570 , \4568 , \4569 );
and \U$3901 ( \4571 , \1927 , RIaaa7940_553);
and \U$3902 ( \4572 , \1470 , RIaaa7760_549);
nor \U$3903 ( \4573 , \4571 , \4572 );
nand \U$3904 ( \4574 , \4564 , \4570 , \4573 );
nor \U$3905 ( \4575 , \4553 , \4574 );
buf \U$3906 ( \4576 , \4575 );
not \U$3907 ( \4577 , \4576 );
not \U$3908 ( \4578 , \2432 );
or \U$3909 ( \4579 , \4577 , \4578 );
or \U$3910 ( \4580 , \2432 , \4576 );
nand \U$3911 ( \4581 , \4579 , \4580 );
not \U$3912 ( \4582 , \4581 );
not \U$3913 ( \4583 , \2920 );
or \U$3914 ( \4584 , \4582 , \4583 );
not \U$3915 ( \4585 , \4359 );
not \U$3916 ( \4586 , \2110 );
or \U$3917 ( \4587 , \4585 , \4586 );
or \U$3918 ( \4588 , \2110 , \4359 );
nand \U$3919 ( \4589 , \4587 , \4588 );
nand \U$3920 ( \4590 , \4589 , \2164 );
nand \U$3921 ( \4591 , \4584 , \4590 );
nand \U$3922 ( \4592 , \4531 , \4591 );
not \U$3923 ( \4593 , \4592 );
not \U$3924 ( \4594 , \4593 );
xor \U$3925 ( \4595 , \4263 , \4306 );
xnor \U$3926 ( \4596 , \4595 , \4363 );
not \U$3927 ( \4597 , \4596 );
not \U$3928 ( \4598 , \4597 );
not \U$3929 ( \4599 , \4372 );
not \U$3930 ( \4600 , \1940 );
or \U$3931 ( \4601 , \4599 , \4600 );
or \U$3932 ( \4602 , \1991 , \4372 );
nand \U$3933 ( \4603 , \4601 , \4602 );
not \U$3934 ( \4604 , \4603 );
not \U$3935 ( \4605 , \1895 );
or \U$3936 ( \4606 , \4604 , \4605 );
nand \U$3937 ( \4607 , \2234 , \4408 );
nand \U$3938 ( \4608 , \4606 , \4607 );
not \U$3939 ( \4609 , \3678 );
not \U$3940 ( \4610 , \2318 );
or \U$3941 ( \4611 , \4609 , \4610 );
not \U$3942 ( \4612 , \4393 );
and \U$3943 ( \4613 , \3211 , \4612 );
not \U$3944 ( \4614 , \3211 );
and \U$3945 ( \4615 , \4614 , \4058 );
nor \U$3946 ( \4616 , \4613 , \4615 );
nand \U$3947 ( \4617 , \4611 , \4616 );
not \U$3948 ( \4618 , \4617 );
nand \U$3949 ( \4619 , \2312 , \3679 );
nand \U$3950 ( \4620 , \4618 , \4619 );
xor \U$3951 ( \4621 , \4608 , \4620 );
not \U$3952 ( \4622 , \4305 );
not \U$3953 ( \4623 , \4622 );
not \U$3954 ( \4624 , \4292 );
or \U$3955 ( \4625 , \4623 , \4624 );
or \U$3956 ( \4626 , \4292 , \4622 );
nand \U$3957 ( \4627 , \4625 , \4626 );
and \U$3958 ( \4628 , \4621 , \4627 );
and \U$3959 ( \4629 , \4608 , \4620 );
or \U$3960 ( \4630 , \4628 , \4629 );
not \U$3961 ( \4631 , \4630 );
not \U$3962 ( \4632 , \4631 );
or \U$3963 ( \4633 , \4598 , \4632 );
nand \U$3964 ( \4634 , \4596 , \4630 );
nand \U$3965 ( \4635 , \4633 , \4634 );
not \U$3966 ( \4636 , \4635 );
or \U$3967 ( \4637 , \4594 , \4636 );
not \U$3968 ( \4638 , \4631 );
nand \U$3969 ( \4639 , \4638 , \4597 );
nand \U$3970 ( \4640 , \4637 , \4639 );
not \U$3971 ( \4641 , \4640 );
not \U$3972 ( \4642 , \4379 );
nand \U$3973 ( \4643 , \4365 , \4307 );
not \U$3974 ( \4644 , \4643 );
not \U$3975 ( \4645 , \4644 );
or \U$3976 ( \4646 , \4642 , \4645 );
or \U$3977 ( \4647 , \4644 , \4379 );
nand \U$3978 ( \4648 , \4646 , \4647 );
not \U$3979 ( \4649 , \4648 );
and \U$3980 ( \4650 , \2823 , \2690 );
or \U$3981 ( \4651 , \2949 , \2486 );
nand \U$3982 ( \4652 , \2951 , \2486 );
nand \U$3983 ( \4653 , \4651 , \4652 );
nor \U$3984 ( \4654 , \4650 , \4653 );
nand \U$3985 ( \4655 , \2944 , \2915 );
nand \U$3986 ( \4656 , \4654 , \4655 );
not \U$3987 ( \4657 , \4656 );
not \U$3988 ( \4658 , \2285 );
not \U$3989 ( \4659 , \4658 );
not \U$3990 ( \4660 , \3156 );
and \U$3991 ( \4661 , \4659 , \4660 );
and \U$3992 ( \4662 , \2907 , \3232 );
not \U$3993 ( \4663 , \2907 );
not \U$3994 ( \4664 , \2291 );
and \U$3995 ( \4665 , \4663 , \4664 );
nor \U$3996 ( \4666 , \4662 , \4665 );
nor \U$3997 ( \4667 , \4661 , \4666 );
nand \U$3998 ( \4668 , \2241 , \3157 );
nand \U$3999 ( \4669 , \4667 , \4668 );
not \U$4000 ( \4670 , \4669 );
or \U$4001 ( \4671 , \4657 , \4670 );
not \U$4002 ( \4672 , \4576 );
nand \U$4003 ( \4673 , \2448 , \4672 );
nand \U$4004 ( \4674 , \4671 , \4673 );
nand \U$4005 ( \4675 , \2442 , \4589 );
nand \U$4006 ( \4676 , \4375 , \2164 );
and \U$4007 ( \4677 , \4675 , \4676 );
not \U$4008 ( \4678 , \4677 );
and \U$4009 ( \4679 , \4674 , \4678 );
not \U$4010 ( \4680 , \4673 );
and \U$4011 ( \4681 , \4669 , \4656 , \4680 );
nor \U$4012 ( \4682 , \4679 , \4681 );
not \U$4013 ( \4683 , \4682 );
and \U$4014 ( \4684 , \4649 , \4683 );
and \U$4015 ( \4685 , \4648 , \4682 );
nor \U$4016 ( \4686 , \4684 , \4685 );
not \U$4017 ( \4687 , \4686 );
not \U$4018 ( \4688 , \4687 );
or \U$4019 ( \4689 , \4641 , \4688 );
not \U$4020 ( \4690 , \4682 );
nand \U$4021 ( \4691 , \4690 , \4648 );
nand \U$4022 ( \4692 , \4689 , \4691 );
not \U$4023 ( \4693 , \4692 );
or \U$4024 ( \4694 , \4452 , \4693 );
or \U$4025 ( \4695 , \4692 , \4451 );
nand \U$4026 ( \4696 , \4694 , \4695 );
not \U$4027 ( \4697 , \4696 );
or \U$4028 ( \4698 , \4449 , \4697 );
or \U$4029 ( \4699 , \4448 , \4696 );
nand \U$4030 ( \4700 , \4698 , \4699 );
xor \U$4031 ( \4701 , \4420 , \4424 );
xor \U$4032 ( \4702 , \4701 , \4387 );
xor \U$4033 ( \4703 , \4674 , \4677 );
not \U$4034 ( \4704 , \4703 );
xor \U$4035 ( \4705 , \4413 , \4398 );
xor \U$4036 ( \4706 , \4705 , \4416 );
not \U$4037 ( \4707 , \4706 );
or \U$4038 ( \4708 , \4704 , \4707 );
or \U$4039 ( \4709 , \4706 , \4703 );
nand \U$4040 ( \4710 , \4708 , \4709 );
not \U$4041 ( \4711 , \4710 );
and \U$4042 ( \4712 , \4635 , \4593 );
not \U$4043 ( \4713 , \4635 );
and \U$4044 ( \4714 , \4713 , \4592 );
nor \U$4045 ( \4715 , \4712 , \4714 );
not \U$4046 ( \4716 , \4715 );
or \U$4047 ( \4717 , \4711 , \4716 );
not \U$4048 ( \4718 , \4703 );
nand \U$4049 ( \4719 , \4718 , \4706 );
nand \U$4050 ( \4720 , \4717 , \4719 );
not \U$4051 ( \4721 , \4720 );
xor \U$4052 ( \4722 , \4702 , \4721 );
not \U$4053 ( \4723 , \4640 );
not \U$4054 ( \4724 , \4686 );
and \U$4055 ( \4725 , \4723 , \4724 );
and \U$4056 ( \4726 , \4640 , \4686 );
nor \U$4057 ( \4727 , \4725 , \4726 );
and \U$4058 ( \4728 , \4722 , \4727 );
and \U$4059 ( \4729 , \4702 , \4721 );
or \U$4060 ( \4730 , \4728 , \4729 );
nand \U$4061 ( \4731 , \4700 , \4730 );
not \U$4062 ( \4732 , \4242 );
not \U$4063 ( \4733 , \4438 );
not \U$4064 ( \4734 , \4733 );
or \U$4065 ( \4735 , \4732 , \4734 );
not \U$4066 ( \4736 , \4242 );
nand \U$4067 ( \4737 , \4736 , \4438 );
nand \U$4068 ( \4738 , \4735 , \4737 );
not \U$4069 ( \4739 , \4696 );
not \U$4070 ( \4740 , \4448 );
not \U$4071 ( \4741 , \4740 );
or \U$4072 ( \4742 , \4739 , \4741 );
not \U$4073 ( \4743 , \4692 );
nand \U$4074 ( \4744 , \4743 , \4451 );
nand \U$4075 ( \4745 , \4742 , \4744 );
nand \U$4076 ( \4746 , \4738 , \4745 );
nand \U$4077 ( \4747 , \4731 , \4746 );
not \U$4078 ( \4748 , \4747 );
not \U$4079 ( \4749 , \3678 );
not \U$4080 ( \4750 , \3092 );
or \U$4081 ( \4751 , \4749 , \4750 );
and \U$4082 ( \4752 , \3684 , \1584 );
not \U$4083 ( \4753 , \3684 );
and \U$4084 ( \4754 , \4753 , \2804 );
nor \U$4085 ( \4755 , \4752 , \4754 );
nand \U$4086 ( \4756 , \4751 , \4755 );
nor \U$4087 ( \4757 , \3239 , \3678 );
nor \U$4088 ( \4758 , \4756 , \4757 );
not \U$4089 ( \4759 , \4758 );
not \U$4090 ( \4760 , \1559 );
not \U$4091 ( \4761 , RIaaa7d00_561);
not \U$4092 ( \4762 , \4761 );
and \U$4093 ( \4763 , \4760 , \4762 );
not \U$4094 ( \4764 , RIaaa7f58_566);
nor \U$4095 ( \4765 , \4177 , \4764 );
nor \U$4096 ( \4766 , \4763 , \4765 );
not \U$4097 ( \4767 , RIaaa7fd0_567);
not \U$4098 ( \4768 , \4767 );
not \U$4099 ( \4769 , \1469 );
and \U$4100 ( \4770 , \4768 , \4769 );
and \U$4101 ( \4771 , \1960 , RIaaa7b98_558);
nor \U$4102 ( \4772 , \4770 , \4771 );
not \U$4103 ( \4773 , \4166 );
not \U$4104 ( \4774 , RIaaa7b20_557);
not \U$4105 ( \4775 , \4774 );
and \U$4106 ( \4776 , \4773 , \4775 );
and \U$4107 ( \4777 , \1541 , RIaaa7df0_563);
nor \U$4108 ( \4778 , \4776 , \4777 );
and \U$4109 ( \4779 , \1482 , RIaaa7c88_560);
not \U$4110 ( \4780 , RIaaa7e68_564);
not \U$4111 ( \4781 , \1491 );
or \U$4112 ( \4782 , \4780 , \4781 );
nand \U$4113 ( \4783 , \1494 , RIaaa7ee0_565);
nand \U$4114 ( \4784 , \4782 , \4783 );
nor \U$4115 ( \4785 , \4779 , \4784 );
and \U$4116 ( \4786 , \4766 , \4772 , \4778 , \4785 );
not \U$4117 ( \4787 , RIaaa7d78_562);
not \U$4118 ( \4788 , \1502 );
or \U$4119 ( \4789 , \4787 , \4788 );
nand \U$4120 ( \4790 , \1461 , RIaaa8048_568);
nand \U$4121 ( \4791 , \4789 , \4790 );
not \U$4122 ( \4792 , RIaaa7c10_559);
not \U$4123 ( \4793 , \4186 );
or \U$4124 ( \4794 , \4792 , \4793 );
nand \U$4125 ( \4795 , \1564 , RIaaa8138_570);
nand \U$4126 ( \4796 , \4794 , \4795 );
nor \U$4127 ( \4797 , \4791 , \4796 );
not \U$4128 ( \4798 , \1426 );
not \U$4129 ( \4799 , RIaaa80c0_569);
not \U$4130 ( \4800 , \4799 );
and \U$4131 ( \4801 , \4798 , \4800 );
not \U$4132 ( \4802 , RIaaa7aa8_556);
nor \U$4133 ( \4803 , \4152 , \4802 );
nor \U$4134 ( \4804 , \4801 , \4803 );
and \U$4135 ( \4805 , \1413 , RIaaa7a30_555);
and \U$4136 ( \4806 , \1479 , RIaaa79b8_554);
nor \U$4137 ( \4807 , \4805 , \4806 );
nand \U$4138 ( \4808 , \4786 , \4797 , \4804 , \4807 );
not \U$4139 ( \4809 , \4808 );
buf \U$4140 ( \4810 , \4809 );
nand \U$4141 ( \4811 , \1897 , \4810 );
and \U$4142 ( \4812 , \4811 , \2098 );
buf \U$4143 ( \4813 , \4808 );
not \U$4144 ( \4814 , \4813 );
nor \U$4145 ( \4815 , \3514 , \4814 );
nor \U$4146 ( \4816 , \4812 , \4815 );
and \U$4147 ( \4817 , \2432 , \4816 );
and \U$4148 ( \4818 , \2516 , \3215 );
or \U$4149 ( \4819 , \2908 , \2949 );
nand \U$4150 ( \4820 , \2908 , \2830 );
nand \U$4151 ( \4821 , \4819 , \4820 );
nor \U$4152 ( \4822 , \4818 , \4821 );
nand \U$4153 ( \4823 , \2508 , \3157 );
nand \U$4154 ( \4824 , \4822 , \4823 );
xor \U$4155 ( \4825 , \4817 , \4824 );
and \U$4156 ( \4826 , \4759 , \4825 );
and \U$4157 ( \4827 , \4817 , \4824 );
nor \U$4158 ( \4828 , \4826 , \4827 );
buf \U$4159 ( \4829 , \4506 );
not \U$4160 ( \4830 , \4829 );
not \U$4161 ( \4831 , \4513 );
not \U$4162 ( \4832 , \4528 );
nor \U$4163 ( \4833 , \4832 , \4526 );
not \U$4164 ( \4834 , \4833 );
or \U$4165 ( \4835 , \4831 , \4834 );
or \U$4166 ( \4836 , \4833 , \4513 );
nand \U$4167 ( \4837 , \4835 , \4836 );
not \U$4168 ( \4838 , \4837 );
or \U$4169 ( \4839 , \4830 , \4838 );
or \U$4170 ( \4840 , \4837 , \4829 );
nand \U$4171 ( \4841 , \4839 , \4840 );
nor \U$4172 ( \4842 , \4828 , \4841 );
not \U$4173 ( \4843 , \4842 );
nand \U$4174 ( \4844 , \4828 , \4841 );
nand \U$4175 ( \4845 , \4843 , \4844 );
not \U$4176 ( \4846 , \4672 );
not \U$4177 ( \4847 , \3341 );
or \U$4178 ( \4848 , \4846 , \4847 );
and \U$4179 ( \4849 , \1900 , \4576 );
not \U$4180 ( \4850 , \4358 );
not \U$4181 ( \4851 , \3514 );
not \U$4182 ( \4852 , \4851 );
or \U$4183 ( \4853 , \4850 , \4852 );
not \U$4184 ( \4854 , \4358 );
nand \U$4185 ( \4855 , \1897 , \4854 );
nand \U$4186 ( \4856 , \4853 , \4855 );
not \U$4187 ( \4857 , \4856 );
nor \U$4188 ( \4858 , \4857 , \3512 );
nor \U$4189 ( \4859 , \4849 , \4858 );
nand \U$4190 ( \4860 , \4848 , \4859 );
not \U$4191 ( \4861 , \4860 );
not \U$4192 ( \4862 , \2151 );
not \U$4193 ( \4863 , \3071 );
nor \U$4194 ( \4864 , \4862 , \4863 );
and \U$4195 ( \4865 , \2209 , \3076 );
not \U$4196 ( \4866 , \2209 );
and \U$4197 ( \4867 , \4866 , \3258 );
or \U$4198 ( \4868 , \4865 , \4867 );
nor \U$4199 ( \4869 , \4864 , \4868 );
and \U$4200 ( \4870 , \3026 , \2914 );
not \U$4201 ( \4871 , \2754 );
buf \U$4202 ( \4872 , \2484 );
not \U$4203 ( \4873 , \4872 );
or \U$4204 ( \4874 , \4871 , \4873 );
or \U$4205 ( \4875 , \4254 , \3248 );
nand \U$4206 ( \4876 , \4874 , \4875 );
nor \U$4207 ( \4877 , \4870 , \4876 );
nand \U$4208 ( \4878 , \3038 , \2689 );
and \U$4209 ( \4879 , \4877 , \4878 );
xor \U$4210 ( \4880 , \4869 , \4879 );
not \U$4211 ( \4881 , \2311 );
not \U$4212 ( \4882 , \4373 );
and \U$4213 ( \4883 , \4881 , \4882 );
not \U$4214 ( \4884 , \4372 );
not \U$4215 ( \4885 , \2318 );
or \U$4216 ( \4886 , \4884 , \4885 );
and \U$4217 ( \4887 , \4403 , \4058 );
not \U$4218 ( \4888 , \4403 );
and \U$4219 ( \4889 , \4888 , \4612 );
nor \U$4220 ( \4890 , \4887 , \4889 );
nand \U$4221 ( \4891 , \4886 , \4890 );
nor \U$4222 ( \4892 , \4883 , \4891 );
xnor \U$4223 ( \4893 , \4880 , \4892 );
not \U$4224 ( \4894 , \4893 );
or \U$4225 ( \4895 , \4861 , \4894 );
not \U$4226 ( \4896 , \4892 );
not \U$4227 ( \4897 , \4879 );
and \U$4228 ( \4898 , \4897 , \4869 );
not \U$4229 ( \4899 , \4897 );
not \U$4230 ( \4900 , \4869 );
and \U$4231 ( \4901 , \4899 , \4900 );
or \U$4232 ( \4902 , \4898 , \4901 );
nand \U$4233 ( \4903 , \4896 , \4902 );
nand \U$4234 ( \4904 , \4895 , \4903 );
and \U$4235 ( \4905 , \4845 , \4904 );
not \U$4236 ( \4906 , \4845 );
not \U$4237 ( \4907 , \4904 );
and \U$4238 ( \4908 , \4906 , \4907 );
nor \U$4239 ( \4909 , \4905 , \4908 );
not \U$4240 ( \4910 , \4576 );
not \U$4241 ( \4911 , \1993 );
or \U$4242 ( \4912 , \4910 , \4911 );
not \U$4243 ( \4913 , \1943 );
not \U$4244 ( \4914 , \4576 );
and \U$4245 ( \4915 , \4913 , \4914 );
not \U$4246 ( \4916 , \4494 );
not \U$4247 ( \4917 , \3515 );
or \U$4248 ( \4918 , \4916 , \4917 );
nand \U$4249 ( \4919 , \1897 , \4493 );
nand \U$4250 ( \4920 , \4918 , \4919 );
and \U$4251 ( \4921 , \3510 , \4920 );
nor \U$4252 ( \4922 , \4915 , \4921 );
nand \U$4253 ( \4923 , \4912 , \4922 );
not \U$4254 ( \4924 , \4923 );
and \U$4255 ( \4925 , \3259 , \3294 );
nor \U$4256 ( \4926 , \3077 , \3294 );
nor \U$4257 ( \4927 , \4925 , \4926 );
nand \U$4258 ( \4928 , \3071 , \2990 );
nand \U$4259 ( \4929 , \4927 , \4928 );
not \U$4260 ( \4930 , \4814 );
and \U$4261 ( \4931 , \2163 , \4930 );
xor \U$4262 ( \4932 , \4929 , \4931 );
not \U$4263 ( \4933 , \2908 );
not \U$4264 ( \4934 , \3038 );
or \U$4265 ( \4935 , \4933 , \4934 );
and \U$4266 ( \4936 , \3026 , \2907 );
and \U$4267 ( \4937 , \2689 , \4521 );
not \U$4268 ( \4938 , \2689 );
and \U$4269 ( \4939 , \4938 , \3033 );
or \U$4270 ( \4940 , \4937 , \4939 );
nor \U$4271 ( \4941 , \4936 , \4940 );
nand \U$4272 ( \4942 , \4935 , \4941 );
xor \U$4273 ( \4943 , \4932 , \4942 );
not \U$4274 ( \4944 , \4943 );
and \U$4275 ( \4945 , \2574 , \4359 );
or \U$4276 ( \4946 , \3002 , \4194 );
or \U$4277 ( \4947 , \4195 , \2400 );
nand \U$4278 ( \4948 , \4946 , \4947 );
nor \U$4279 ( \4949 , \4945 , \4948 );
not \U$4280 ( \4950 , \4359 );
nand \U$4281 ( \4951 , \4950 , \2583 );
and \U$4282 ( \4952 , \4949 , \4951 );
nand \U$4283 ( \4953 , \4944 , \4952 );
not \U$4284 ( \4954 , \4953 );
or \U$4285 ( \4955 , \4924 , \4954 );
not \U$4286 ( \4956 , \4952 );
nand \U$4287 ( \4957 , \4956 , \4943 );
nand \U$4288 ( \4958 , \4955 , \4957 );
not \U$4289 ( \4959 , \4958 );
xor \U$4290 ( \4960 , \4825 , \4758 );
not \U$4291 ( \4961 , \4960 );
and \U$4292 ( \4962 , \4893 , \4860 );
not \U$4293 ( \4963 , \4893 );
not \U$4294 ( \4964 , \4860 );
and \U$4295 ( \4965 , \4963 , \4964 );
nor \U$4296 ( \4966 , \4962 , \4965 );
not \U$4297 ( \4967 , \4966 );
or \U$4298 ( \4968 , \4961 , \4967 );
or \U$4299 ( \4969 , \4966 , \4960 );
nand \U$4300 ( \4970 , \4968 , \4969 );
not \U$4301 ( \4971 , \4970 );
or \U$4302 ( \4972 , \4959 , \4971 );
not \U$4303 ( \4973 , \4960 );
nand \U$4304 ( \4974 , \4973 , \4966 );
nand \U$4305 ( \4975 , \4972 , \4974 );
not \U$4306 ( \4976 , \4975 );
xor \U$4307 ( \4977 , \4909 , \4976 );
not \U$4308 ( \4978 , \2920 );
not \U$4309 ( \4979 , \2161 );
not \U$4310 ( \4980 , \4494 );
and \U$4311 ( \4981 , \4979 , \4980 );
and \U$4312 ( \4982 , \2432 , \4494 );
nor \U$4313 ( \4983 , \4981 , \4982 );
not \U$4314 ( \4984 , \4983 );
not \U$4315 ( \4985 , \4984 );
or \U$4316 ( \4986 , \4978 , \4985 );
nand \U$4317 ( \4987 , \4581 , \2164 );
nand \U$4318 ( \4988 , \4986 , \4987 );
and \U$4319 ( \4989 , \3510 , \4856 );
and \U$4320 ( \4990 , \3511 , \4603 );
nor \U$4321 ( \4991 , \4989 , \4990 );
not \U$4322 ( \4992 , \4991 );
not \U$4323 ( \4993 , \3915 );
not \U$4324 ( \4994 , \2406 );
or \U$4325 ( \4995 , \4993 , \4994 );
and \U$4326 ( \4996 , \2390 , \3914 );
or \U$4327 ( \4997 , \2399 , \3679 );
nand \U$4328 ( \4998 , \4058 , \4036 );
nand \U$4329 ( \4999 , \4997 , \4998 );
nor \U$4330 ( \5000 , \4996 , \4999 );
nand \U$4331 ( \5001 , \4995 , \5000 );
not \U$4332 ( \5002 , \5001 );
or \U$4333 ( \5003 , \4992 , \5002 );
or \U$4334 ( \5004 , \5001 , \4991 );
nand \U$4335 ( \5005 , \5003 , \5004 );
not \U$4336 ( \5006 , \5005 );
and \U$4337 ( \5007 , \4988 , \5006 );
not \U$4338 ( \5008 , \4988 );
and \U$4339 ( \5009 , \5008 , \5005 );
nor \U$4340 ( \5010 , \5007 , \5009 );
not \U$4341 ( \5011 , \5010 );
nand \U$4342 ( \5012 , \4897 , \4900 );
not \U$4343 ( \5013 , \5012 );
nand \U$4344 ( \5014 , \2802 , \3684 );
nand \U$4345 ( \5015 , \2241 , \3212 );
and \U$4346 ( \5016 , \1579 , \3157 );
and \U$4347 ( \5017 , \3233 , \4055 );
nor \U$4348 ( \5018 , \5016 , \5017 );
nand \U$4349 ( \5019 , \5014 , \5015 , \5018 );
nand \U$4350 ( \5020 , \5013 , \5019 );
not \U$4351 ( \5021 , \5019 );
buf \U$4352 ( \5022 , \5012 );
nand \U$4353 ( \5023 , \5021 , \5022 );
and \U$4354 ( \5024 , \5020 , \5023 );
not \U$4355 ( \5025 , \4810 );
and \U$4356 ( \5026 , \2448 , \5025 );
nor \U$4357 ( \5027 , \5024 , \5026 );
not \U$4358 ( \5028 , \5027 );
nand \U$4359 ( \5029 , \5011 , \5028 );
nand \U$4360 ( \5030 , \5010 , \5027 );
nand \U$4361 ( \5031 , \5029 , \5030 );
not \U$4362 ( \5032 , \5025 );
not \U$4363 ( \5033 , \2443 );
or \U$4364 ( \5034 , \5032 , \5033 );
not \U$4365 ( \5035 , \4983 );
not \U$4366 ( \5036 , \2164 );
not \U$4367 ( \5037 , \5036 );
and \U$4368 ( \5038 , \5035 , \5037 );
and \U$4369 ( \5039 , \3462 , \4810 );
nor \U$4370 ( \5040 , \5038 , \5039 );
nand \U$4371 ( \5041 , \5034 , \5040 );
not \U$4372 ( \5042 , \5041 );
xor \U$4373 ( \5043 , \4929 , \4931 );
and \U$4374 ( \5044 , \5043 , \4942 );
and \U$4375 ( \5045 , \4929 , \4931 );
or \U$4376 ( \5046 , \5044 , \5045 );
not \U$4377 ( \5047 , \5046 );
not \U$4378 ( \5048 , \3914 );
not \U$4379 ( \5049 , \1365 );
or \U$4380 ( \5050 , \5048 , \5049 );
and \U$4381 ( \5051 , \3677 , \2533 );
not \U$4382 ( \5052 , \3677 );
and \U$4383 ( \5053 , \5052 , \2291 );
nor \U$4384 ( \5054 , \5051 , \5053 );
nand \U$4385 ( \5055 , \5050 , \5054 );
not \U$4386 ( \5056 , \5055 );
nand \U$4387 ( \5057 , \1591 , \3915 );
nand \U$4388 ( \5058 , \5056 , \5057 );
not \U$4389 ( \5059 , \5058 );
not \U$4390 ( \5060 , \3155 );
not \U$4391 ( \5061 , \5060 );
not \U$4392 ( \5062 , \4286 );
or \U$4393 ( \5063 , \5061 , \5062 );
and \U$4394 ( \5064 , \2905 , \2754 );
not \U$4395 ( \5065 , \2905 );
and \U$4396 ( \5066 , \5065 , \3029 );
nor \U$4397 ( \5067 , \5064 , \5066 );
nand \U$4398 ( \5068 , \5063 , \5067 );
and \U$4399 ( \5069 , \3037 , \3155 );
or \U$4400 ( \5070 , \5068 , \5069 );
not \U$4401 ( \5071 , \3077 );
not \U$4402 ( \5072 , \2485 );
and \U$4403 ( \5073 , \5071 , \5072 );
not \U$4404 ( \5074 , \4872 );
and \U$4405 ( \5075 , \3259 , \5074 );
nor \U$4406 ( \5076 , \5073 , \5075 );
nand \U$4407 ( \5077 , \3071 , \2914 );
nand \U$4408 ( \5078 , \5076 , \5077 );
and \U$4409 ( \5079 , \5070 , \5078 );
not \U$4410 ( \5080 , \5079 );
not \U$4411 ( \5081 , \3211 );
not \U$4412 ( \5082 , \2822 );
or \U$4413 ( \5083 , \5081 , \5082 );
and \U$4414 ( \5084 , \3156 , \2830 );
not \U$4415 ( \5085 , \3156 );
and \U$4416 ( \5086 , \5085 , \2521 );
nor \U$4417 ( \5087 , \5084 , \5086 );
nand \U$4418 ( \5088 , \5083 , \5087 );
not \U$4419 ( \5089 , \3211 );
and \U$4420 ( \5090 , \4251 , \5089 );
nor \U$4421 ( \5091 , \5088 , \5090 );
not \U$4422 ( \5092 , \5091 );
or \U$4423 ( \5093 , \5080 , \5092 );
not \U$4424 ( \5094 , \5078 );
not \U$4425 ( \5095 , \5070 );
or \U$4426 ( \5096 , \5094 , \5095 );
or \U$4427 ( \5097 , \5088 , \5090 );
nand \U$4428 ( \5098 , \5096 , \5097 );
nand \U$4429 ( \5099 , \5093 , \5098 );
not \U$4430 ( \5100 , \5099 );
or \U$4431 ( \5101 , \5059 , \5100 );
or \U$4432 ( \5102 , \5090 , \5088 );
buf \U$4433 ( \5103 , \5070 );
nand \U$4434 ( \5104 , \5102 , \5103 , \5078 );
nand \U$4435 ( \5105 , \5101 , \5104 );
not \U$4436 ( \5106 , \5105 );
not \U$4437 ( \5107 , \5106 );
or \U$4438 ( \5108 , \5047 , \5107 );
not \U$4439 ( \5109 , \5046 );
nand \U$4440 ( \5110 , \5105 , \5109 );
nand \U$4441 ( \5111 , \5108 , \5110 );
not \U$4442 ( \5112 , \5111 );
or \U$4443 ( \5113 , \5042 , \5112 );
not \U$4444 ( \5114 , \5106 );
nand \U$4445 ( \5115 , \5114 , \5046 );
nand \U$4446 ( \5116 , \5113 , \5115 );
and \U$4447 ( \5117 , \5031 , \5116 );
not \U$4448 ( \5118 , \5031 );
not \U$4449 ( \5119 , \5116 );
and \U$4450 ( \5120 , \5118 , \5119 );
nor \U$4451 ( \5121 , \5117 , \5120 );
xor \U$4452 ( \5122 , \4977 , \5121 );
and \U$4453 ( \5123 , \5111 , \5041 );
not \U$4454 ( \5124 , \5111 );
not \U$4455 ( \5125 , \5041 );
and \U$4456 ( \5126 , \5124 , \5125 );
nor \U$4457 ( \5127 , \5123 , \5126 );
xor \U$4458 ( \5128 , \5099 , \5058 );
not \U$4459 ( \5129 , \5128 );
nand \U$4460 ( \5130 , \1367 , \4373 );
and \U$4461 ( \5131 , \3914 , \1584 );
not \U$4462 ( \5132 , \3914 );
and \U$4463 ( \5133 , \5132 , \1579 );
nor \U$4464 ( \5134 , \5131 , \5133 );
nand \U$4465 ( \5135 , \5130 , \5134 );
nor \U$4466 ( \5136 , \1592 , \4194 );
nor \U$4467 ( \5137 , \5135 , \5136 );
not \U$4468 ( \5138 , \5137 );
not \U$4469 ( \5139 , \5138 );
not \U$4470 ( \5140 , \2317 );
nor \U$4471 ( \5141 , \5140 , \3586 );
not \U$4472 ( \5142 , \5141 );
not \U$4473 ( \5143 , \4813 );
buf \U$4474 ( \5144 , \5143 );
not \U$4475 ( \5145 , \5144 );
and \U$4476 ( \5146 , \5142 , \5145 );
nor \U$4477 ( \5147 , \5146 , \3590 );
not \U$4478 ( \5148 , \5147 );
not \U$4479 ( \5149 , \3678 );
nand \U$4480 ( \5150 , \5149 , \2508 );
not \U$4481 ( \5151 , \5150 );
not \U$4482 ( \5152 , \3678 );
not \U$4483 ( \5153 , \2515 );
or \U$4484 ( \5154 , \5152 , \5153 );
and \U$4485 ( \5155 , \3211 , \2521 );
not \U$4486 ( \5156 , \3211 );
and \U$4487 ( \5157 , \5156 , \2951 );
nor \U$4488 ( \5158 , \5155 , \5157 );
nand \U$4489 ( \5159 , \5154 , \5158 );
nor \U$4490 ( \5160 , \5151 , \5159 );
not \U$4491 ( \5161 , \5160 );
or \U$4492 ( \5162 , \5148 , \5161 );
not \U$4493 ( \5163 , \5150 );
or \U$4494 ( \5164 , \5159 , \5163 );
not \U$4495 ( \5165 , \5147 );
nand \U$4496 ( \5166 , \5164 , \5165 );
nand \U$4497 ( \5167 , \5162 , \5166 );
not \U$4498 ( \5168 , \5167 );
or \U$4499 ( \5169 , \5139 , \5168 );
or \U$4500 ( \5170 , \5159 , \5163 );
nand \U$4501 ( \5171 , \5170 , \5147 );
nand \U$4502 ( \5172 , \5169 , \5171 );
not \U$4503 ( \5173 , \5172 );
or \U$4504 ( \5174 , \5129 , \5173 );
or \U$4505 ( \5175 , \5172 , \5128 );
not \U$4506 ( \5176 , \5078 );
not \U$4507 ( \5177 , \5176 );
not \U$4508 ( \5178 , \5103 );
or \U$4509 ( \5179 , \5177 , \5178 );
or \U$4510 ( \5180 , \5176 , \5103 );
nand \U$4511 ( \5181 , \5179 , \5180 );
and \U$4512 ( \5182 , \2572 , \4576 );
not \U$4513 ( \5183 , \4359 );
or \U$4514 ( \5184 , \5183 , \2400 );
not \U$4515 ( \5185 , \4358 );
nand \U$4516 ( \5186 , \2498 , \5185 );
nand \U$4517 ( \5187 , \5184 , \5186 );
nor \U$4518 ( \5188 , \5182 , \5187 );
not \U$4519 ( \5189 , \4576 );
nand \U$4520 ( \5190 , \5189 , \2583 );
nand \U$4521 ( \5191 , \5188 , \5190 );
xor \U$4522 ( \5192 , \5181 , \5191 );
not \U$4523 ( \5193 , \5025 );
and \U$4524 ( \5194 , \5193 , \1900 );
not \U$4525 ( \5195 , \4920 );
nor \U$4526 ( \5196 , \5195 , \3512 );
nor \U$4527 ( \5197 , \5194 , \5196 );
nand \U$4528 ( \5198 , \3341 , \5025 );
nand \U$4529 ( \5199 , \5197 , \5198 );
and \U$4530 ( \5200 , \5192 , \5199 );
and \U$4531 ( \5201 , \5181 , \5191 );
nor \U$4532 ( \5202 , \5200 , \5201 );
not \U$4533 ( \5203 , \5202 );
nand \U$4534 ( \5204 , \5175 , \5203 );
nand \U$4535 ( \5205 , \5174 , \5204 );
xor \U$4536 ( \5206 , \5127 , \5205 );
buf \U$4537 ( \5207 , \5206 );
not \U$4538 ( \5208 , \4970 );
not \U$4539 ( \5209 , \4958 );
not \U$4540 ( \5210 , \5209 );
and \U$4541 ( \5211 , \5208 , \5210 );
and \U$4542 ( \5212 , \5209 , \4970 );
nor \U$4543 ( \5213 , \5211 , \5212 );
not \U$4544 ( \5214 , \5213 );
and \U$4545 ( \5215 , \5207 , \5214 );
and \U$4546 ( \5216 , \5127 , \5205 );
nor \U$4547 ( \5217 , \5215 , \5216 );
nand \U$4548 ( \5218 , \5122 , \5217 );
not \U$4549 ( \5219 , \5218 );
xor \U$4550 ( \5220 , \5128 , \5172 );
xor \U$4551 ( \5221 , \5220 , \5202 );
xor \U$4552 ( \5222 , \4923 , \4952 );
xnor \U$4553 ( \5223 , \5222 , \4943 );
not \U$4554 ( \5224 , \5223 );
nand \U$4555 ( \5225 , \5221 , \5224 );
and \U$4556 ( \5226 , \3915 , \2508 );
not \U$4557 ( \5227 , \3914 );
not \U$4558 ( \5228 , \2515 );
or \U$4559 ( \5229 , \5227 , \5228 );
and \U$4560 ( \5230 , \2521 , \3678 );
nor \U$4561 ( \5231 , \4259 , \3678 );
nor \U$4562 ( \5232 , \5230 , \5231 );
nand \U$4563 ( \5233 , \5229 , \5232 );
nor \U$4564 ( \5234 , \5226 , \5233 );
not \U$4565 ( \5235 , \5234 );
and \U$4566 ( \5236 , \3026 , \3678 );
not \U$4567 ( \5237 , \4042 );
or \U$4568 ( \5238 , \3248 , \5237 );
nand \U$4569 ( \5239 , \3250 , \5237 );
nand \U$4570 ( \5240 , \5238 , \5239 );
nor \U$4571 ( \5241 , \5236 , \5240 );
nand \U$4572 ( \5242 , \3038 , \3679 );
nand \U$4573 ( \5243 , \5241 , \5242 );
not \U$4574 ( \5244 , \3215 );
not \U$4575 ( \5245 , \3071 );
or \U$4576 ( \5246 , \5244 , \5245 );
not \U$4577 ( \5247 , \3077 );
not \U$4578 ( \5248 , \2906 );
not \U$4579 ( \5249 , \5248 );
and \U$4580 ( \5250 , \5247 , \5249 );
and \U$4581 ( \5251 , \3259 , \4060 );
nor \U$4582 ( \5252 , \5250 , \5251 );
nand \U$4583 ( \5253 , \5246 , \5252 );
and \U$4584 ( \5254 , \5243 , \5253 );
not \U$4585 ( \5255 , \5254 );
or \U$4586 ( \5256 , \5235 , \5255 );
or \U$4587 ( \5257 , \5254 , \5234 );
nand \U$4588 ( \5258 , \5256 , \5257 );
not \U$4589 ( \5259 , \5258 );
not \U$4590 ( \5260 , \4359 );
not \U$4591 ( \5261 , \2802 );
or \U$4592 ( \5262 , \5260 , \5261 );
and \U$4593 ( \5263 , \4194 , \2533 );
not \U$4594 ( \5264 , \4194 );
and \U$4595 ( \5265 , \5264 , \1579 );
nor \U$4596 ( \5266 , \5263 , \5265 );
nand \U$4597 ( \5267 , \5262 , \5266 );
not \U$4598 ( \5268 , \3815 );
nor \U$4599 ( \5269 , \5268 , \4359 );
nor \U$4600 ( \5270 , \5267 , \5269 );
not \U$4601 ( \5271 , \5270 );
not \U$4602 ( \5272 , \5271 );
or \U$4603 ( \5273 , \5259 , \5272 );
not \U$4604 ( \5274 , \5234 );
nand \U$4605 ( \5275 , \5274 , \5254 );
nand \U$4606 ( \5276 , \5273 , \5275 );
not \U$4607 ( \5277 , \5276 );
xor \U$4608 ( \5278 , \5137 , \5167 );
and \U$4609 ( \5279 , \3511 , \5025 );
not \U$4610 ( \5280 , \5279 );
and \U$4611 ( \5281 , \3259 , \2688 );
nor \U$4612 ( \5282 , \2688 , \3075 );
nor \U$4613 ( \5283 , \5281 , \5282 );
nand \U$4614 ( \5284 , \3071 , \2906 );
and \U$4615 ( \5285 , \5283 , \5284 );
not \U$4616 ( \5286 , \5285 );
not \U$4617 ( \5287 , \3212 );
not \U$4618 ( \5288 , \3038 );
or \U$4619 ( \5289 , \5287 , \5288 );
and \U$4620 ( \5290 , \3026 , \3211 );
and \U$4621 ( \5291 , \3156 , \3029 );
not \U$4622 ( \5292 , \3156 );
and \U$4623 ( \5293 , \5292 , \3033 );
or \U$4624 ( \5294 , \5291 , \5293 );
nor \U$4625 ( \5295 , \5290 , \5294 );
nand \U$4626 ( \5296 , \5289 , \5295 );
not \U$4627 ( \5297 , \5296 );
or \U$4628 ( \5298 , \5286 , \5297 );
or \U$4629 ( \5299 , \5296 , \5285 );
nand \U$4630 ( \5300 , \5298 , \5299 );
not \U$4631 ( \5301 , \5300 );
or \U$4632 ( \5302 , \5280 , \5301 );
not \U$4633 ( \5303 , \5285 );
nand \U$4634 ( \5304 , \5303 , \5296 );
nand \U$4635 ( \5305 , \5302 , \5304 );
xnor \U$4636 ( \5306 , \5278 , \5305 );
not \U$4637 ( \5307 , \5306 );
or \U$4638 ( \5308 , \5277 , \5307 );
xor \U$4639 ( \5309 , \5167 , \5138 );
nand \U$4640 ( \5310 , \5309 , \5305 );
nand \U$4641 ( \5311 , \5308 , \5310 );
buf \U$4642 ( \5312 , \5311 );
and \U$4643 ( \5313 , \5225 , \5312 );
nor \U$4644 ( \5314 , \5221 , \5224 );
nor \U$4645 ( \5315 , \5313 , \5314 );
not \U$4646 ( \5316 , \5315 );
not \U$4647 ( \5317 , \5213 );
not \U$4648 ( \5318 , \5206 );
or \U$4649 ( \5319 , \5317 , \5318 );
or \U$4650 ( \5320 , \5206 , \5213 );
nand \U$4651 ( \5321 , \5319 , \5320 );
nand \U$4652 ( \5322 , \5316 , \5321 );
xor \U$4653 ( \5323 , \5223 , \5311 );
xnor \U$4654 ( \5324 , \5323 , \5221 );
buf \U$4655 ( \5325 , \5306 );
and \U$4656 ( \5326 , \5325 , \5276 );
not \U$4657 ( \5327 , \5325 );
not \U$4658 ( \5328 , \5276 );
and \U$4659 ( \5329 , \5327 , \5328 );
nor \U$4660 ( \5330 , \5326 , \5329 );
not \U$4661 ( \5331 , \5330 );
xor \U$4662 ( \5332 , \5192 , \5199 );
not \U$4663 ( \5333 , \5332 );
xor \U$4664 ( \5334 , \5285 , \5279 );
xnor \U$4665 ( \5335 , \5334 , \5296 );
not \U$4666 ( \5336 , \2583 );
not \U$4667 ( \5337 , \5336 );
not \U$4668 ( \5338 , \4494 );
and \U$4669 ( \5339 , \5337 , \5338 );
not \U$4670 ( \5340 , \4494 );
not \U$4671 ( \5341 , \2574 );
or \U$4672 ( \5342 , \5340 , \5341 );
and \U$4673 ( \5343 , \4672 , \3295 );
not \U$4674 ( \5344 , \4672 );
and \U$4675 ( \5345 , \5344 , \2495 );
nor \U$4676 ( \5346 , \5343 , \5345 );
nand \U$4677 ( \5347 , \5342 , \5346 );
nor \U$4678 ( \5348 , \5339 , \5347 );
not \U$4679 ( \5349 , \5348 );
not \U$4680 ( \5350 , \4193 );
not \U$4681 ( \5351 , \5350 );
not \U$4682 ( \5352 , \4251 );
or \U$4683 ( \5353 , \5351 , \5352 );
and \U$4684 ( \5354 , \2822 , \4193 );
and \U$4685 ( \5355 , \3913 , \2520 );
not \U$4686 ( \5356 , \3913 );
and \U$4687 ( \5357 , \5356 , \4259 );
nor \U$4688 ( \5358 , \5355 , \5357 );
nor \U$4689 ( \5359 , \5354 , \5358 );
nand \U$4690 ( \5360 , \5353 , \5359 );
not \U$4691 ( \5361 , \5360 );
not \U$4692 ( \5362 , \4810 );
buf \U$4693 ( \5363 , \2298 );
not \U$4694 ( \5364 , \5363 );
or \U$4695 ( \5365 , \5362 , \5364 );
nand \U$4696 ( \5366 , \5365 , \2538 );
not \U$4697 ( \5367 , \5363 );
nand \U$4698 ( \5368 , \5367 , \4813 );
nand \U$4699 ( \5369 , \3507 , \5366 , \5368 );
nand \U$4700 ( \5370 , \5361 , \5369 );
not \U$4701 ( \5371 , \5370 );
xor \U$4702 ( \5372 , \5253 , \5243 );
not \U$4703 ( \5373 , \5372 );
or \U$4704 ( \5374 , \5371 , \5373 );
not \U$4705 ( \5375 , \5369 );
nand \U$4706 ( \5376 , \5375 , \5360 );
nand \U$4707 ( \5377 , \5374 , \5376 );
xor \U$4708 ( \5378 , \5349 , \5377 );
nand \U$4709 ( \5379 , \5335 , \5378 );
not \U$4710 ( \5380 , \5379 );
and \U$4711 ( \5381 , \5349 , \5377 );
nor \U$4712 ( \5382 , \5380 , \5381 );
not \U$4713 ( \5383 , \5382 );
or \U$4714 ( \5384 , \5333 , \5383 );
not \U$4715 ( \5385 , \5381 );
not \U$4716 ( \5386 , \5385 );
not \U$4717 ( \5387 , \5379 );
or \U$4718 ( \5388 , \5386 , \5387 );
not \U$4719 ( \5389 , \5332 );
nand \U$4720 ( \5390 , \5388 , \5389 );
nand \U$4721 ( \5391 , \5384 , \5390 );
not \U$4722 ( \5392 , \5391 );
or \U$4723 ( \5393 , \5331 , \5392 );
not \U$4724 ( \5394 , \5385 );
not \U$4725 ( \5395 , \5379 );
or \U$4726 ( \5396 , \5394 , \5395 );
nand \U$4727 ( \5397 , \5396 , \5332 );
nand \U$4728 ( \5398 , \5393 , \5397 );
nand \U$4729 ( \5399 , \5324 , \5398 );
nand \U$4730 ( \5400 , \5322 , \5399 );
not \U$4731 ( \5401 , \5321 );
buf \U$4732 ( \5402 , \5315 );
nand \U$4733 ( \5403 , \5401 , \5402 );
nand \U$4734 ( \5404 , \5400 , \5403 );
not \U$4735 ( \5405 , \5404 );
not \U$4736 ( \5406 , \5405 );
or \U$4737 ( \5407 , \5219 , \5406 );
not \U$4738 ( \5408 , \5030 );
not \U$4739 ( \5409 , \5116 );
or \U$4740 ( \5410 , \5408 , \5409 );
nand \U$4741 ( \5411 , \5410 , \5029 );
not \U$4742 ( \5412 , \5020 );
xor \U$4743 ( \5413 , \4669 , \4656 );
not \U$4744 ( \5414 , \5413 );
or \U$4745 ( \5415 , \5412 , \5414 );
or \U$4746 ( \5416 , \5413 , \5020 );
nand \U$4747 ( \5417 , \5415 , \5416 );
not \U$4748 ( \5418 , \4988 );
not \U$4749 ( \5419 , \5005 );
or \U$4750 ( \5420 , \5418 , \5419 );
not \U$4751 ( \5421 , \4991 );
nand \U$4752 ( \5422 , \5421 , \5001 );
nand \U$4753 ( \5423 , \5420 , \5422 );
xor \U$4754 ( \5424 , \5417 , \5423 );
xor \U$4755 ( \5425 , \5411 , \5424 );
xor \U$4756 ( \5426 , \4608 , \4620 );
xor \U$4757 ( \5427 , \5426 , \4627 );
nor \U$4758 ( \5428 , \4531 , \4591 );
not \U$4759 ( \5429 , \5428 );
nand \U$4760 ( \5430 , \5429 , \4592 );
xor \U$4761 ( \5431 , \5427 , \5430 );
not \U$4762 ( \5432 , \4904 );
not \U$4763 ( \5433 , \4844 );
or \U$4764 ( \5434 , \5432 , \5433 );
not \U$4765 ( \5435 , \4842 );
nand \U$4766 ( \5436 , \5434 , \5435 );
xor \U$4767 ( \5437 , \5431 , \5436 );
xor \U$4768 ( \5438 , \5425 , \5437 );
xor \U$4769 ( \5439 , \4909 , \4976 );
and \U$4770 ( \5440 , \5439 , \5121 );
and \U$4771 ( \5441 , \4909 , \4976 );
or \U$4772 ( \5442 , \5440 , \5441 );
nor \U$4773 ( \5443 , \5438 , \5442 );
nor \U$4774 ( \5444 , \5122 , \5217 );
nor \U$4775 ( \5445 , \5443 , \5444 );
nand \U$4776 ( \5446 , \5407 , \5445 );
xor \U$4777 ( \5447 , \4702 , \4721 );
xor \U$4778 ( \5448 , \5447 , \4727 );
not \U$4779 ( \5449 , \5423 );
not \U$4780 ( \5450 , \5417 );
or \U$4781 ( \5451 , \5449 , \5450 );
not \U$4782 ( \5452 , \5020 );
nand \U$4783 ( \5453 , \5452 , \5413 );
nand \U$4784 ( \5454 , \5451 , \5453 );
not \U$4785 ( \5455 , \5427 );
not \U$4786 ( \5456 , \5455 );
not \U$4787 ( \5457 , \5430 );
or \U$4788 ( \5458 , \5456 , \5457 );
nand \U$4789 ( \5459 , \5458 , \5436 );
not \U$4790 ( \5460 , \5428 );
nand \U$4791 ( \5461 , \5460 , \4592 , \5427 );
nand \U$4792 ( \5462 , \5459 , \5461 );
xor \U$4793 ( \5463 , \5454 , \5462 );
xor \U$4794 ( \5464 , \4715 , \4710 );
and \U$4795 ( \5465 , \5463 , \5464 );
and \U$4796 ( \5466 , \5454 , \5462 );
or \U$4797 ( \5467 , \5465 , \5466 );
not \U$4798 ( \5468 , \5467 );
nand \U$4799 ( \5469 , \5448 , \5468 );
xor \U$4800 ( \5470 , \5454 , \5462 );
xor \U$4801 ( \5471 , \5470 , \5464 );
not \U$4802 ( \5472 , \5471 );
not \U$4803 ( \5473 , \5437 );
and \U$4804 ( \5474 , \5425 , \5473 );
and \U$4805 ( \5475 , \5411 , \5424 );
nor \U$4806 ( \5476 , \5474 , \5475 );
nand \U$4807 ( \5477 , \5472 , \5476 );
nand \U$4808 ( \5478 , \5469 , \5477 );
not \U$4809 ( \5479 , \5478 );
nand \U$4810 ( \5480 , \5438 , \5442 );
buf \U$4811 ( \5481 , \5480 );
nand \U$4812 ( \5482 , \4748 , \5446 , \5479 , \5481 );
not \U$4813 ( \5483 , \5398 );
not \U$4814 ( \5484 , \5324 );
nand \U$4815 ( \5485 , \5483 , \5484 );
and \U$4816 ( \5486 , \5485 , \5403 );
not \U$4817 ( \5487 , \5330 );
and \U$4818 ( \5488 , \5391 , \5487 );
not \U$4819 ( \5489 , \5391 );
and \U$4820 ( \5490 , \5489 , \5330 );
nor \U$4821 ( \5491 , \5488 , \5490 );
xor \U$4822 ( \5492 , \5348 , \5335 );
xnor \U$4823 ( \5493 , \5492 , \5377 );
not \U$4824 ( \5494 , \5258 );
not \U$4825 ( \5495 , \5270 );
and \U$4826 ( \5496 , \5494 , \5495 );
and \U$4827 ( \5497 , \5270 , \5258 );
nor \U$4828 ( \5498 , \5496 , \5497 );
not \U$4829 ( \5499 , \5498 );
not \U$4830 ( \5500 , \5144 );
not \U$4831 ( \5501 , \5500 );
not \U$4832 ( \5502 , \2582 );
or \U$4833 ( \5503 , \5501 , \5502 );
buf \U$4834 ( \5504 , \2318 );
and \U$4835 ( \5505 , \5504 , \5144 );
or \U$4836 ( \5506 , \2396 , \4494 );
or \U$4837 ( \5507 , \4393 , \4493 );
nand \U$4838 ( \5508 , \5506 , \5507 );
nor \U$4839 ( \5509 , \5505 , \5508 );
nand \U$4840 ( \5510 , \5503 , \5509 );
not \U$4841 ( \5511 , \5510 );
buf \U$4842 ( \5512 , \5511 );
not \U$4843 ( \5513 , \5512 );
not \U$4844 ( \5514 , \5513 );
buf \U$4845 ( \5515 , \2285 );
and \U$4846 ( \5516 , \5515 , \4576 );
not \U$4847 ( \5517 , \1583 );
not \U$4848 ( \5518 , \4358 );
or \U$4849 ( \5519 , \5517 , \5518 );
nand \U$4850 ( \5520 , \4854 , \4276 );
nand \U$4851 ( \5521 , \5519 , \5520 );
nor \U$4852 ( \5522 , \5516 , \5521 );
nand \U$4853 ( \5523 , \2241 , \4672 );
nand \U$4854 ( \5524 , \5522 , \5523 );
not \U$4855 ( \5525 , \5524 );
not \U$4856 ( \5526 , \5525 );
not \U$4857 ( \5527 , \5526 );
or \U$4858 ( \5528 , \5514 , \5527 );
not \U$4859 ( \5529 , \3071 );
nor \U$4860 ( \5530 , \5529 , \5089 );
not \U$4861 ( \5531 , \3076 );
not \U$4862 ( \5532 , \5060 );
or \U$4863 ( \5533 , \5531 , \5532 );
not \U$4864 ( \5534 , \3259 );
or \U$4865 ( \5535 , \5534 , \3215 );
nand \U$4866 ( \5536 , \5533 , \5535 );
nor \U$4867 ( \5537 , \5530 , \5536 );
nand \U$4868 ( \5538 , \2367 , \5500 );
xor \U$4869 ( \5539 , \5537 , \5538 );
not \U$4870 ( \5540 , \3914 );
not \U$4871 ( \5541 , \3026 );
or \U$4872 ( \5542 , \5540 , \5541 );
and \U$4873 ( \5543 , \3677 , \3250 );
not \U$4874 ( \5544 , \3677 );
and \U$4875 ( \5545 , \5544 , \3031 );
nor \U$4876 ( \5546 , \5543 , \5545 );
nand \U$4877 ( \5547 , \5542 , \5546 );
and \U$4878 ( \5548 , \3038 , \3915 );
nor \U$4879 ( \5549 , \5547 , \5548 );
and \U$4880 ( \5550 , \5539 , \5549 );
and \U$4881 ( \5551 , \5537 , \5538 );
or \U$4882 ( \5552 , \5550 , \5551 );
not \U$4883 ( \5553 , \5552 );
nand \U$4884 ( \5554 , \5525 , \5512 );
nand \U$4885 ( \5555 , \5553 , \5554 );
nand \U$4886 ( \5556 , \5528 , \5555 );
not \U$4887 ( \5557 , \5556 );
and \U$4888 ( \5558 , \5499 , \5557 );
and \U$4889 ( \5559 , \5498 , \5556 );
nor \U$4890 ( \5560 , \5558 , \5559 );
not \U$4891 ( \5561 , \5560 );
and \U$4892 ( \5562 , \5493 , \5561 );
not \U$4893 ( \5563 , \5556 );
nor \U$4894 ( \5564 , \5563 , \5498 );
nor \U$4895 ( \5565 , \5562 , \5564 );
nand \U$4896 ( \5566 , \5491 , \5565 );
not \U$4897 ( \5567 , \5566 );
nor \U$4898 ( \5568 , \5560 , \5493 );
not \U$4899 ( \5569 , \5568 );
nand \U$4900 ( \5570 , \5560 , \5493 );
xor \U$4901 ( \5571 , \5524 , \5511 );
xnor \U$4902 ( \5572 , \5571 , \5552 );
not \U$4903 ( \5573 , \5572 );
not \U$4904 ( \5574 , \5369 );
not \U$4905 ( \5575 , \5360 );
or \U$4906 ( \5576 , \5574 , \5575 );
or \U$4907 ( \5577 , \5360 , \5369 );
nand \U$4908 ( \5578 , \5576 , \5577 );
xor \U$4909 ( \5579 , \5372 , \5578 );
not \U$4910 ( \5580 , \4808 );
not \U$4911 ( \5581 , \2513 );
or \U$4912 ( \5582 , \5580 , \5581 );
not \U$4913 ( \5583 , \1334 );
nand \U$4914 ( \5584 , \5582 , \5583 );
not \U$4915 ( \5585 , \5584 );
not \U$4916 ( \5586 , \4808 );
and \U$4917 ( \5587 , \1192 , \5586 );
not \U$4918 ( \5588 , \1355 );
nor \U$4919 ( \5589 , \5587 , \5588 );
not \U$4920 ( \5590 , \5589 );
and \U$4921 ( \5591 , \3258 , \3209 );
nor \U$4922 ( \5592 , \3075 , \3209 );
nor \U$4923 ( \5593 , \5591 , \5592 );
nand \U$4924 ( \5594 , \3071 , \3676 );
nand \U$4925 ( \5595 , \5593 , \5594 );
nand \U$4926 ( \5596 , \5585 , \5590 , \5595 );
buf \U$4927 ( \5597 , \5596 );
not \U$4928 ( \5598 , \5597 );
not \U$4929 ( \5599 , \5183 );
not \U$4930 ( \5600 , \2508 );
or \U$4931 ( \5601 , \5599 , \5600 );
and \U$4932 ( \5602 , \2822 , \4358 );
not \U$4933 ( \5603 , \4192 );
not \U$4934 ( \5604 , \2951 );
or \U$4935 ( \5605 , \5603 , \5604 );
not \U$4936 ( \5606 , \4372 );
or \U$4937 ( \5607 , \2833 , \5606 );
nand \U$4938 ( \5608 , \5605 , \5607 );
nor \U$4939 ( \5609 , \5602 , \5608 );
nand \U$4940 ( \5610 , \5601 , \5609 );
not \U$4941 ( \5611 , \5610 );
not \U$4942 ( \5612 , \5611 );
or \U$4943 ( \5613 , \5598 , \5612 );
not \U$4944 ( \5614 , \3092 );
not \U$4945 ( \5615 , \4494 );
or \U$4946 ( \5616 , \5614 , \5615 );
and \U$4947 ( \5617 , \4576 , \2533 );
not \U$4948 ( \5618 , \4576 );
and \U$4949 ( \5619 , \5618 , \2291 );
nor \U$4950 ( \5620 , \5617 , \5619 );
nand \U$4951 ( \5621 , \5616 , \5620 );
nor \U$4952 ( \5622 , \3239 , \4494 );
nor \U$4953 ( \5623 , \5621 , \5622 );
not \U$4954 ( \5624 , \5623 );
nand \U$4955 ( \5625 , \5613 , \5624 );
not \U$4956 ( \5626 , \5597 );
nand \U$4957 ( \5627 , \5626 , \5610 );
nand \U$4958 ( \5628 , \5625 , \5627 );
or \U$4959 ( \5629 , \5579 , \5628 );
and \U$4960 ( \5630 , \5573 , \5629 );
and \U$4961 ( \5631 , \5628 , \5579 );
nor \U$4962 ( \5632 , \5630 , \5631 );
nand \U$4963 ( \5633 , \5569 , \5570 , \5632 );
not \U$4964 ( \5634 , \5633 );
nor \U$4965 ( \5635 , \5589 , \5584 );
nor \U$4966 ( \5636 , \5635 , \5595 );
not \U$4967 ( \5637 , \5636 );
nand \U$4968 ( \5638 , \5637 , \5596 );
not \U$4969 ( \5639 , \4193 );
not \U$4970 ( \5640 , \3026 );
or \U$4971 ( \5641 , \5639 , \5640 );
and \U$4972 ( \5642 , \3913 , \3033 );
not \U$4973 ( \5643 , \3913 );
and \U$4974 ( \5644 , \5643 , \3031 );
nor \U$4975 ( \5645 , \5642 , \5644 );
nand \U$4976 ( \5646 , \5641 , \5645 );
and \U$4977 ( \5647 , \3038 , \4192 );
nor \U$4978 ( \5648 , \5646 , \5647 );
xor \U$4979 ( \5649 , \5638 , \5648 );
not \U$4980 ( \5650 , \4576 );
not \U$4981 ( \5651 , \2515 );
or \U$4982 ( \5652 , \5650 , \5651 );
and \U$4983 ( \5653 , \4358 , \2521 );
not \U$4984 ( \5654 , \4358 );
and \U$4985 ( \5655 , \5654 , \2830 );
nor \U$4986 ( \5656 , \5653 , \5655 );
nand \U$4987 ( \5657 , \5652 , \5656 );
nor \U$4988 ( \5658 , \2943 , \4576 );
nor \U$4989 ( \5659 , \5657 , \5658 );
and \U$4990 ( \5660 , \5649 , \5659 );
and \U$4991 ( \5661 , \5638 , \5648 );
or \U$4992 ( \5662 , \5660 , \5661 );
xor \U$4993 ( \5663 , \5537 , \5538 );
xor \U$4994 ( \5664 , \5663 , \5549 );
xor \U$4995 ( \5665 , \5662 , \5664 );
xor \U$4996 ( \5666 , \5596 , \5610 );
xnor \U$4997 ( \5667 , \5666 , \5623 );
xor \U$4998 ( \5668 , \5665 , \5667 );
xor \U$4999 ( \5669 , \5638 , \5648 );
xor \U$5000 ( \5670 , \5669 , \5659 );
not \U$5001 ( \5671 , \5670 );
nor \U$5002 ( \5672 , \2537 , \5143 );
not \U$5003 ( \5673 , \3913 );
not \U$5004 ( \5674 , \3071 );
or \U$5005 ( \5675 , \5673 , \5674 );
and \U$5006 ( \5676 , \3676 , \3076 );
not \U$5007 ( \5677 , \3676 );
and \U$5008 ( \5678 , \5677 , \3258 );
nor \U$5009 ( \5679 , \5676 , \5678 );
nand \U$5010 ( \5680 , \5675 , \5679 );
nand \U$5011 ( \5681 , \5672 , \5680 );
not \U$5012 ( \5682 , \5681 );
not \U$5013 ( \5683 , \4358 );
not \U$5014 ( \5684 , \3026 );
or \U$5015 ( \5685 , \5683 , \5684 );
and \U$5016 ( \5686 , \4372 , \3250 );
not \U$5017 ( \5687 , \4372 );
and \U$5018 ( \5688 , \5687 , \4521 );
nor \U$5019 ( \5689 , \5686 , \5688 );
nand \U$5020 ( \5690 , \5685 , \5689 );
and \U$5021 ( \5691 , \3038 , \5185 );
nor \U$5022 ( \5692 , \5690 , \5691 );
not \U$5023 ( \5693 , \5692 );
or \U$5024 ( \5694 , \5682 , \5693 );
nor \U$5025 ( \5695 , \5672 , \5680 );
not \U$5026 ( \5696 , \5695 );
nand \U$5027 ( \5697 , \5694 , \5696 );
not \U$5028 ( \5698 , \1590 );
and \U$5029 ( \5699 , \5698 , \5500 );
not \U$5030 ( \5700 , \4810 );
not \U$5031 ( \5701 , \1365 );
or \U$5032 ( \5702 , \5700 , \5701 );
and \U$5033 ( \5703 , \4494 , \2533 );
not \U$5034 ( \5704 , \4494 );
and \U$5035 ( \5705 , \5704 , \1577 );
nor \U$5036 ( \5706 , \5703 , \5705 );
nand \U$5037 ( \5707 , \5702 , \5706 );
nor \U$5038 ( \5708 , \5699 , \5707 );
nand \U$5039 ( \5709 , \5697 , \5708 );
and \U$5040 ( \5710 , \5671 , \5709 );
nor \U$5041 ( \5711 , \5708 , \5697 );
nor \U$5042 ( \5712 , \5710 , \5711 );
nand \U$5043 ( \5713 , \5668 , \5712 );
not \U$5044 ( \5714 , \5713 );
not \U$5045 ( \5715 , \4493 );
not \U$5046 ( \5716 , \2508 );
or \U$5047 ( \5717 , \5715 , \5716 );
and \U$5048 ( \5718 , \2822 , \4494 );
and \U$5049 ( \5719 , \4575 , \2520 );
not \U$5050 ( \5720 , \4575 );
and \U$5051 ( \5721 , \5720 , \4259 );
nor \U$5052 ( \5722 , \5719 , \5721 );
nor \U$5053 ( \5723 , \5718 , \5722 );
nand \U$5054 ( \5724 , \5717 , \5723 );
not \U$5055 ( \5725 , \3912 );
not \U$5056 ( \5726 , \3075 );
and \U$5057 ( \5727 , \5725 , \5726 );
and \U$5058 ( \5728 , \3258 , \4403 );
nor \U$5059 ( \5729 , \5727 , \5728 );
nand \U$5060 ( \5730 , \3071 , \4372 );
nand \U$5061 ( \5731 , \5729 , \5730 );
not \U$5062 ( \5732 , \4808 );
not \U$5063 ( \5733 , \2758 );
not \U$5064 ( \5734 , \5733 );
or \U$5065 ( \5735 , \5732 , \5734 );
not \U$5066 ( \5736 , \4808 );
not \U$5067 ( \5737 , \5736 );
not \U$5068 ( \5738 , \2758 );
or \U$5069 ( \5739 , \5737 , \5738 );
not \U$5070 ( \5740 , \1150 );
nand \U$5071 ( \5741 , \5739 , \5740 );
nand \U$5072 ( \5742 , \5735 , \5741 );
nor \U$5073 ( \5743 , \1193 , \5742 );
and \U$5074 ( \5744 , \5731 , \5743 );
nand \U$5075 ( \5745 , \5724 , \5744 );
not \U$5076 ( \5746 , \5745 );
not \U$5077 ( \5747 , \5695 );
nand \U$5078 ( \5748 , \5747 , \5681 );
not \U$5079 ( \5749 , \5748 );
and \U$5080 ( \5750 , \5692 , \5749 );
not \U$5081 ( \5751 , \5692 );
and \U$5082 ( \5752 , \5751 , \5748 );
nor \U$5083 ( \5753 , \5750 , \5752 );
not \U$5084 ( \5754 , \5753 );
or \U$5085 ( \5755 , \5746 , \5754 );
nor \U$5086 ( \5756 , \5724 , \5744 );
not \U$5087 ( \5757 , \5756 );
nand \U$5088 ( \5758 , \5755 , \5757 );
not \U$5089 ( \5759 , \5758 );
not \U$5090 ( \5760 , \5711 );
nand \U$5091 ( \5761 , \5760 , \5709 );
and \U$5092 ( \5762 , \5761 , \5671 );
not \U$5093 ( \5763 , \5761 );
and \U$5094 ( \5764 , \5763 , \5670 );
nor \U$5095 ( \5765 , \5762 , \5764 );
not \U$5096 ( \5766 , \5765 );
or \U$5097 ( \5767 , \5759 , \5766 );
not \U$5098 ( \5768 , \2833 );
not \U$5099 ( \5769 , \4493 );
and \U$5100 ( \5770 , \5768 , \5769 );
buf \U$5101 ( \5771 , \2830 );
and \U$5102 ( \5772 , \5771 , \4493 );
nor \U$5103 ( \5773 , \5770 , \5772 );
not \U$5104 ( \5774 , \4814 );
not \U$5105 ( \5775 , \2513 );
or \U$5106 ( \5776 , \5774 , \5775 );
or \U$5107 ( \5777 , \2513 , \4814 );
nand \U$5108 ( \5778 , \5776 , \5777 );
nand \U$5109 ( \5779 , \5778 , \1187 );
nand \U$5110 ( \5780 , \5773 , \5779 );
not \U$5111 ( \5781 , \5780 );
not \U$5112 ( \5782 , \5781 );
xor \U$5113 ( \5783 , \5731 , \5743 );
and \U$5114 ( \5784 , \4357 , \5733 );
not \U$5115 ( \5785 , \4357 );
and \U$5116 ( \5786 , \5785 , \2758 );
nor \U$5117 ( \5787 , \5784 , \5786 );
and \U$5118 ( \5788 , \2751 , \5787 );
not \U$5119 ( \5789 , \4575 );
not \U$5120 ( \5790 , \3024 );
or \U$5121 ( \5791 , \5789 , \5790 );
or \U$5122 ( \5792 , \2758 , \4575 );
nand \U$5123 ( \5793 , \5791 , \5792 );
and \U$5124 ( \5794 , \2771 , \5793 );
nor \U$5125 ( \5795 , \5788 , \5794 );
nand \U$5126 ( \5796 , \5795 , \2817 );
not \U$5127 ( \5797 , \5796 );
and \U$5128 ( \5798 , \5783 , \5797 );
not \U$5129 ( \5799 , \5783 );
and \U$5130 ( \5800 , \5799 , \5796 );
nor \U$5131 ( \5801 , \5798 , \5800 );
not \U$5132 ( \5802 , \5801 );
or \U$5133 ( \5803 , \5782 , \5802 );
not \U$5134 ( \5804 , \5783 );
nand \U$5135 ( \5805 , \5804 , \5796 );
nand \U$5136 ( \5806 , \5803 , \5805 );
not \U$5137 ( \5807 , \5806 );
not \U$5138 ( \5808 , \5756 );
nand \U$5139 ( \5809 , \5808 , \5745 );
not \U$5140 ( \5810 , \5753 );
and \U$5141 ( \5811 , \5809 , \5810 );
not \U$5142 ( \5812 , \5809 );
and \U$5143 ( \5813 , \5812 , \5753 );
nor \U$5144 ( \5814 , \5811 , \5813 );
not \U$5145 ( \5815 , \5814 );
or \U$5146 ( \5816 , \5807 , \5815 );
and \U$5147 ( \5817 , \3258 , \4190 );
nor \U$5148 ( \5818 , \4190 , \3075 );
nor \U$5149 ( \5819 , \5817 , \5818 );
nand \U$5150 ( \5820 , \3071 , \4356 );
nand \U$5151 ( \5821 , \5819 , \5820 );
not \U$5152 ( \5822 , \5821 );
not \U$5153 ( \5823 , \4809 );
nand \U$5154 ( \5824 , \5823 , \1189 );
nand \U$5155 ( \5825 , \5822 , \5824 );
not \U$5156 ( \5826 , \5825 );
not \U$5157 ( \5827 , \5821 );
nor \U$5158 ( \5828 , \5827 , \5824 );
nor \U$5159 ( \5829 , \5826 , \5828 );
not \U$5160 ( \5830 , \5829 );
nand \U$5161 ( \5831 , \2750 , \5793 );
and \U$5162 ( \5832 , \4492 , \2758 );
not \U$5163 ( \5833 , \4492 );
and \U$5164 ( \5834 , \5833 , \5733 );
nor \U$5165 ( \5835 , \5832 , \5834 );
nand \U$5166 ( \5836 , \2771 , \5835 );
and \U$5167 ( \5837 , \2817 , \5831 , \5836 );
not \U$5168 ( \5838 , \5837 );
or \U$5169 ( \5839 , \5830 , \5838 );
or \U$5170 ( \5840 , \5829 , \5837 );
nand \U$5171 ( \5841 , \5839 , \5840 );
nand \U$5172 ( \5842 , \2766 , \3020 );
nand \U$5173 ( \5843 , \5842 , \4808 );
not \U$5174 ( \5844 , \2766 );
nand \U$5175 ( \5845 , \5844 , \3019 );
nand \U$5176 ( \5846 , \5843 , \5845 , \5733 );
not \U$5177 ( \5847 , \5846 );
not \U$5178 ( \5848 , \3071 );
nor \U$5179 ( \5849 , \4553 , \4574 );
not \U$5180 ( \5850 , \5849 );
not \U$5181 ( \5851 , \3019 );
or \U$5182 ( \5852 , \5850 , \5851 );
or \U$5183 ( \5853 , \3019 , \5849 );
nand \U$5184 ( \5854 , \5852 , \5853 );
not \U$5185 ( \5855 , \5854 );
or \U$5186 ( \5856 , \5848 , \5855 );
not \U$5187 ( \5857 , \4356 );
and \U$5188 ( \5858 , \3258 , \5857 );
nor \U$5189 ( \5859 , \3075 , \5857 );
nor \U$5190 ( \5860 , \5858 , \5859 );
nand \U$5191 ( \5861 , \5856 , \5860 );
nand \U$5192 ( \5862 , \5847 , \5861 );
nor \U$5193 ( \5863 , \5841 , \5862 );
not \U$5194 ( \5864 , \5825 );
not \U$5195 ( \5865 , \5837 );
or \U$5196 ( \5866 , \5864 , \5865 );
not \U$5197 ( \5867 , \5828 );
nand \U$5198 ( \5868 , \5866 , \5867 );
nor \U$5199 ( \5869 , \5863 , \5868 );
not \U$5200 ( \5870 , \5869 );
nand \U$5201 ( \5871 , \5841 , \5862 );
and \U$5202 ( \5872 , \3038 , \5025 );
xnor \U$5203 ( \5873 , \5861 , \5846 );
and \U$5204 ( \5874 , \2772 , \4930 );
nand \U$5205 ( \5875 , \5854 , \3068 );
and \U$5206 ( \5876 , \5875 , \4863 );
and \U$5207 ( \5877 , \4809 , \3020 );
nor \U$5208 ( \5878 , \5876 , \5877 );
or \U$5209 ( \5879 , \5875 , \5143 );
nand \U$5210 ( \5880 , \5879 , \4493 );
nand \U$5211 ( \5881 , \5878 , \5880 );
nor \U$5212 ( \5882 , \5874 , \5881 );
and \U$5213 ( \5883 , \5873 , \5882 );
nor \U$5214 ( \5884 , \5872 , \5883 );
nand \U$5215 ( \5885 , \3026 , \4810 );
and \U$5216 ( \5886 , \4493 , \3031 );
not \U$5217 ( \5887 , \4493 );
and \U$5218 ( \5888 , \5887 , \3250 );
nor \U$5219 ( \5889 , \5886 , \5888 );
nand \U$5220 ( \5890 , \5884 , \5885 , \5889 );
or \U$5221 ( \5891 , \5873 , \5882 );
nand \U$5222 ( \5892 , \5871 , \5890 , \5891 );
not \U$5223 ( \5893 , \5892 );
or \U$5224 ( \5894 , \5870 , \5893 );
xor \U$5225 ( \5895 , \5780 , \5801 );
nand \U$5226 ( \5896 , \5894 , \5895 );
not \U$5227 ( \5897 , \5863 );
not \U$5228 ( \5898 , \5897 );
not \U$5229 ( \5899 , \5892 );
or \U$5230 ( \5900 , \5898 , \5899 );
nand \U$5231 ( \5901 , \5900 , \5868 );
nand \U$5232 ( \5902 , \5896 , \5901 );
nand \U$5233 ( \5903 , \5816 , \5902 );
not \U$5234 ( \5904 , \5814 );
not \U$5235 ( \5905 , \5806 );
nand \U$5236 ( \5906 , \5904 , \5905 );
nand \U$5237 ( \5907 , \5903 , \5906 );
nand \U$5238 ( \5908 , \5767 , \5907 );
not \U$5239 ( \5909 , \5765 );
not \U$5240 ( \5910 , \5758 );
nand \U$5241 ( \5911 , \5909 , \5910 );
nand \U$5242 ( \5912 , \5908 , \5911 );
not \U$5243 ( \5913 , \5912 );
or \U$5244 ( \5914 , \5714 , \5913 );
not \U$5245 ( \5915 , \5668 );
not \U$5246 ( \5916 , \5712 );
nand \U$5247 ( \5917 , \5915 , \5916 );
nand \U$5248 ( \5918 , \5914 , \5917 );
not \U$5249 ( \5919 , \5918 );
xor \U$5250 ( \5920 , \5662 , \5664 );
and \U$5251 ( \5921 , \5920 , \5667 );
and \U$5252 ( \5922 , \5662 , \5664 );
or \U$5253 ( \5923 , \5921 , \5922 );
not \U$5254 ( \5924 , \5923 );
not \U$5255 ( \5925 , \5572 );
xor \U$5256 ( \5926 , \5628 , \5579 );
not \U$5257 ( \5927 , \5926 );
or \U$5258 ( \5928 , \5925 , \5927 );
or \U$5259 ( \5929 , \5926 , \5572 );
nand \U$5260 ( \5930 , \5928 , \5929 );
not \U$5261 ( \5931 , \5930 );
or \U$5262 ( \5932 , \5924 , \5931 );
or \U$5263 ( \5933 , \5930 , \5923 );
nand \U$5264 ( \5934 , \5932 , \5933 );
not \U$5265 ( \5935 , \5934 );
or \U$5266 ( \5936 , \5919 , \5935 );
not \U$5267 ( \5937 , \5923 );
nand \U$5268 ( \5938 , \5937 , \5930 );
nand \U$5269 ( \5939 , \5936 , \5938 );
not \U$5270 ( \5940 , \5939 );
or \U$5271 ( \5941 , \5634 , \5940 );
not \U$5272 ( \5942 , \5568 );
nand \U$5273 ( \5943 , \5942 , \5570 );
not \U$5274 ( \5944 , \5632 );
nand \U$5275 ( \5945 , \5943 , \5944 );
nand \U$5276 ( \5946 , \5941 , \5945 );
not \U$5277 ( \5947 , \5946 );
or \U$5278 ( \5948 , \5567 , \5947 );
not \U$5279 ( \5949 , \5491 );
not \U$5280 ( \5950 , \5565 );
nand \U$5281 ( \5951 , \5949 , \5950 );
nand \U$5282 ( \5952 , \5948 , \5951 );
nand \U$5283 ( \5953 , \5486 , \5952 , \5218 );
not \U$5284 ( \5954 , \5953 );
not \U$5285 ( \5955 , \5480 );
nor \U$5286 ( \5956 , \5955 , \5478 );
nand \U$5287 ( \5957 , \5954 , \5956 , \4748 );
not \U$5288 ( \5958 , \4747 );
not \U$5289 ( \5959 , \5448 );
nand \U$5290 ( \5960 , \5959 , \5467 );
not \U$5291 ( \5961 , \5476 );
nand \U$5292 ( \5962 , \5961 , \5471 );
and \U$5293 ( \5963 , \5960 , \5962 );
nor \U$5294 ( \5964 , \5959 , \5467 );
nor \U$5295 ( \5965 , \5963 , \5964 );
and \U$5296 ( \5966 , \5958 , \5965 );
nor \U$5297 ( \5967 , \4730 , \4700 );
not \U$5298 ( \5968 , \5967 );
not \U$5299 ( \5969 , \4746 );
or \U$5300 ( \5970 , \5968 , \5969 );
not \U$5301 ( \5971 , \4738 );
not \U$5302 ( \5972 , \4745 );
nand \U$5303 ( \5973 , \5971 , \5972 );
nand \U$5304 ( \5974 , \5970 , \5973 );
nor \U$5305 ( \5975 , \5966 , \5974 );
nand \U$5306 ( \5976 , \5482 , \5957 , \5975 );
not \U$5307 ( \5977 , \5976 );
or \U$5308 ( \5978 , \4446 , \5977 );
nor \U$5309 ( \5979 , \4229 , \4443 );
nand \U$5310 ( \5980 , \4221 , \5979 );
not \U$5311 ( \5981 , \5980 );
nor \U$5312 ( \5982 , \4007 , \4220 );
nor \U$5313 ( \5983 , \3806 , \3991 );
nor \U$5314 ( \5984 , \5982 , \5983 );
not \U$5315 ( \5985 , \5984 );
or \U$5316 ( \5986 , \5981 , \5985 );
nand \U$5317 ( \5987 , \5986 , \4005 );
not \U$5318 ( \5988 , \4002 );
buf \U$5319 ( \5989 , \3994 );
nand \U$5320 ( \5990 , \5988 , \5989 );
nand \U$5321 ( \5991 , \5987 , \5990 );
not \U$5322 ( \5992 , \5991 );
nand \U$5323 ( \5993 , \5978 , \5992 );
nand \U$5324 ( \5994 , \3619 , \5993 );
not \U$5325 ( \5995 , \3581 );
not \U$5326 ( \5996 , \2714 );
not \U$5327 ( \5997 , \3424 );
not \U$5328 ( \5998 , \3428 );
nand \U$5329 ( \5999 , \5997 , \5998 );
nand \U$5330 ( \6000 , \3420 , \3395 );
nand \U$5331 ( \6001 , \5999 , \6000 );
nand \U$5332 ( \6002 , \6001 , \3429 );
not \U$5333 ( \6003 , \2720 );
not \U$5334 ( \6004 , \2634 );
nand \U$5335 ( \6005 , \6004 , \2709 );
not \U$5336 ( \6006 , \6005 );
or \U$5337 ( \6007 , \6003 , \6006 );
nand \U$5338 ( \6008 , \6007 , \2978 );
not \U$5339 ( \6009 , \6008 );
or \U$5340 ( \6010 , \6002 , \6009 );
not \U$5341 ( \6011 , \2721 );
not \U$5342 ( \6012 , \2978 );
nand \U$5343 ( \6013 , \6011 , \6012 );
nand \U$5344 ( \6014 , \6010 , \6013 );
not \U$5345 ( \6015 , \6014 );
or \U$5346 ( \6016 , \5996 , \6015 );
not \U$5347 ( \6017 , \2621 );
nand \U$5348 ( \6018 , \6017 , \2710 , \2712 );
nand \U$5349 ( \6019 , \6016 , \6018 );
not \U$5350 ( \6020 , \6019 );
or \U$5351 ( \6021 , \5995 , \6020 );
and \U$5352 ( \6022 , \3484 , \3535 );
not \U$5353 ( \6023 , \3547 );
nand \U$5354 ( \6024 , \6023 , \3539 );
or \U$5355 ( \6025 , \6022 , \6024 );
or \U$5356 ( \6026 , \3535 , \3484 );
nand \U$5357 ( \6027 , \6025 , \6026 );
not \U$5358 ( \6028 , \3580 );
and \U$5359 ( \6029 , \6027 , \6028 );
or \U$5360 ( \6030 , \3554 , \3579 );
not \U$5361 ( \6031 , \6030 );
nor \U$5362 ( \6032 , \6029 , \6031 );
nand \U$5363 ( \6033 , \6021 , \6032 );
and \U$5364 ( \6034 , \6033 , \3618 );
nor \U$5365 ( \6035 , \3585 , \3617 );
nor \U$5366 ( \6036 , \6034 , \6035 );
and \U$5367 ( \6037 , \5994 , \6036 );
and \U$5368 ( \6038 , \3465 , \1573 );
or \U$5369 ( \6039 , \3463 , \1573 );
nand \U$5370 ( \6040 , \6039 , \3468 );
nor \U$5371 ( \6041 , \6038 , \6040 );
nand \U$5372 ( \6042 , \2448 , \2401 );
nand \U$5373 ( \6043 , \6041 , \6042 );
or \U$5374 ( \6044 , \2920 , \2164 );
and \U$5375 ( \6045 , \2448 , \1573 );
nor \U$5376 ( \6046 , \6045 , \2433 );
nand \U$5377 ( \6047 , \6044 , \6046 );
or \U$5378 ( \6048 , \6047 , \6042 );
nand \U$5379 ( \6049 , \6043 , \6048 );
and \U$5380 ( \6050 , \3607 , \3593 );
nor \U$5381 ( \6051 , \6050 , \3591 );
xor \U$5382 ( \6052 , \6049 , \6051 );
and \U$5383 ( \6053 , \3567 , \3575 );
nor \U$5384 ( \6054 , \6053 , \3608 );
nor \U$5385 ( \6055 , \6052 , \6054 );
nor \U$5386 ( \6056 , \6037 , \6055 );
not \U$5387 ( \6057 , \6042 );
not \U$5388 ( \6058 , \6047 );
or \U$5389 ( \6059 , \6057 , \6058 );
nand \U$5390 ( \6060 , \6059 , \6048 );
not \U$5391 ( \6061 , \6060 );
and \U$5392 ( \6062 , \6049 , \6051 );
not \U$5393 ( \6063 , \6041 );
and \U$5394 ( \6064 , \6063 , \6042 );
nor \U$5395 ( \6065 , \6062 , \6064 );
not \U$5396 ( \6066 , \6065 );
or \U$5397 ( \6067 , \6061 , \6066 );
or \U$5398 ( \6068 , \6065 , \6060 );
nand \U$5399 ( \6069 , \6067 , \6068 );
nand \U$5400 ( \6070 , \6052 , \6054 );
buf \U$5401 ( \6071 , \1704 );
nor \U$5402 ( \6072 , \849 , RIaaa89a8_588);
and \U$5403 ( \6073 , RIaa97770_3, \6072 );
and \U$5404 ( \6074 , \6073 , RIaa976f8_2);
nand \U$5405 ( \6075 , \6074 , RIaa97860_5);
not \U$5406 ( \6076 , \6075 );
nand \U$5407 ( \6077 , \6076 , RIaa978d8_6);
not \U$5408 ( \6078 , \6077 );
nand \U$5409 ( \6079 , \6078 , RIaa97950_7);
not \U$5410 ( \6080 , \6079 );
nand \U$5411 ( \6081 , \6080 , RIaa979c8_8);
not \U$5412 ( \6082 , \6081 );
not \U$5413 ( \6083 , RIaa97ba8_12);
and \U$5414 ( \6084 , \6082 , \6083 );
and \U$5415 ( \6085 , \6081 , RIaa97ba8_12);
nor \U$5416 ( \6086 , \6084 , \6085 );
and \U$5417 ( \6087 , \6071 , \6086 );
or \U$5418 ( \6088 , \6074 , RIaa97860_5);
nand \U$5419 ( \6089 , \6088 , \6075 );
and \U$5420 ( \6090 , \1073 , \6089 );
not \U$5421 ( \6091 , RIaa978d8_6);
not \U$5422 ( \6092 , \6075 );
or \U$5423 ( \6093 , \6091 , \6092 );
or \U$5424 ( \6094 , \6075 , RIaa978d8_6);
nand \U$5425 ( \6095 , \6093 , \6094 );
or \U$5426 ( \6096 , \1135 , \6095 );
not \U$5427 ( \6097 , \6077 );
not \U$5428 ( \6098 , RIaa97950_7);
and \U$5429 ( \6099 , \6097 , \6098 );
and \U$5430 ( \6100 , \6077 , RIaa97950_7);
nor \U$5431 ( \6101 , \6099 , \6100 );
and \U$5432 ( \6102 , \1343 , \6101 );
buf \U$5433 ( \6103 , \1305 );
not \U$5434 ( \6104 , \6079 );
not \U$5435 ( \6105 , RIaa979c8_8);
and \U$5436 ( \6106 , \6104 , \6105 );
and \U$5437 ( \6107 , \6079 , RIaa979c8_8);
nor \U$5438 ( \6108 , \6106 , \6107 );
and \U$5439 ( \6109 , \6103 , \6108 );
nor \U$5440 ( \6110 , \6102 , \6109 );
nand \U$5441 ( \6111 , \6096 , \6110 );
nor \U$5442 ( \6112 , \6090 , \6111 );
buf \U$5443 ( \6113 , \2728 );
and \U$5444 ( \6114 , \849 , RIaaa89a8_588);
nor \U$5445 ( \6115 , \6114 , \6072 );
or \U$5446 ( \6116 , \6113 , \6115 );
xor \U$5447 ( \6117 , RIaa97770_3, \6072 );
buf \U$5448 ( \6118 , \2722 );
or \U$5449 ( \6119 , \6117 , \6118 );
buf \U$5450 ( \6120 , \1164 );
or \U$5451 ( \6121 , \6073 , RIaa976f8_2);
not \U$5452 ( \6122 , \6074 );
nand \U$5453 ( \6123 , \6121 , \6122 );
nand \U$5454 ( \6124 , \6120 , \6123 );
nand \U$5455 ( \6125 , \6116 , \6119 , \6124 );
and \U$5456 ( \6126 , \6113 , \6115 );
nor \U$5457 ( \6127 , \6126 , \2734 );
or \U$5458 ( \6128 , \6125 , \6127 );
or \U$5459 ( \6129 , \6123 , \6120 );
nand \U$5460 ( \6130 , \6124 , \6118 , \6117 );
nand \U$5461 ( \6131 , \6128 , \6129 , \6130 );
and \U$5462 ( \6132 , \6112 , \6131 );
or \U$5463 ( \6133 , \6111 , \1073 , \6089 );
and \U$5464 ( \6134 , \6110 , \1135 , \6095 );
or \U$5465 ( \6135 , \6109 , \1343 , \6101 );
or \U$5466 ( \6136 , \6103 , \6108 );
nand \U$5467 ( \6137 , \6135 , \6136 );
nor \U$5468 ( \6138 , \6134 , \6137 );
nand \U$5469 ( \6139 , \6133 , \6138 );
nor \U$5470 ( \6140 , \6132 , \6139 );
nor \U$5471 ( \6141 , \6087 , \6140 );
nor \U$5472 ( \6142 , \6071 , \6086 );
or \U$5473 ( \6143 , \6141 , \6142 );
not \U$5474 ( \6144 , RIaa97ba8_12);
nor \U$5475 ( \6145 , \6144 , \6081 );
xor \U$5476 ( \6146 , RIaa97b30_11, \6145 );
or \U$5477 ( \6147 , \6146 , \1656 );
not \U$5478 ( \6148 , \1768 );
not \U$5479 ( \6149 , \6148 );
and \U$5480 ( \6150 , RIaa97b30_11, \6145 );
and \U$5481 ( \6151 , \6150 , RIaa97ab8_10);
not \U$5482 ( \6152 , \6150 );
and \U$5483 ( \6153 , \6152 , \1769 );
nor \U$5484 ( \6154 , \6151 , \6153 );
not \U$5485 ( \6155 , \6154 );
and \U$5486 ( \6156 , \6149 , \6155 );
and \U$5487 ( \6157 , \6150 , RIaa97ab8_10);
nor \U$5488 ( \6158 , \6157 , RIaa97a40_9);
not \U$5489 ( \6159 , \1823 );
nor \U$5490 ( \6160 , \6159 , \6081 );
nor \U$5491 ( \6161 , \6158 , \6160 );
nor \U$5492 ( \6162 , \1880 , \6161 );
nor \U$5493 ( \6163 , \6156 , \6162 );
nand \U$5494 ( \6164 , \6143 , \6147 , \6163 );
nand \U$5495 ( \6165 , \6163 , \1656 , \6146 );
not \U$5496 ( \6166 , \6162 );
and \U$5497 ( \6167 , \6166 , \6148 , \6154 );
and \U$5498 ( \6168 , \1880 , \6161 );
nor \U$5499 ( \6169 , \6167 , \6168 );
and \U$5500 ( \6170 , \6164 , \6165 , \6169 );
not \U$5501 ( \6171 , RIaa97d10_15);
nand \U$5502 ( \6172 , \6171 , RIaa97c20_13, RIaa97c98_14, RIaa97e00_17);
not \U$5503 ( \6173 , \6172 );
not \U$5504 ( \6174 , \997 );
and \U$5505 ( \6175 , \6173 , \6174 );
nand \U$5506 ( \6176 , \671 , \703 , \710 , RIaa97c20_13);
not \U$5507 ( \6177 , \6176 );
and \U$5508 ( \6178 , \6177 , RIaa9c450_167);
nor \U$5509 ( \6179 , \6175 , \6178 );
not \U$5510 ( \6180 , RIaa97c98_14);
not \U$5511 ( \6181 , RIaa97e00_17);
nand \U$5512 ( \6182 , \6180 , \6181 , RIaa97c20_13, RIaa97d10_15);
not \U$5513 ( \6183 , \6182 );
and \U$5514 ( \6184 , \6183 , RIaa9c360_165);
not \U$5515 ( \6185 , RIaa9c270_163);
not \U$5516 ( \6186 , RIaa97c20_13);
not \U$5517 ( \6187 , RIaa97d10_15);
nand \U$5518 ( \6188 , \6186 , \6187 , RIaa97c98_14, RIaa97e00_17);
nor \U$5519 ( \6189 , \6185 , \6188 );
nor \U$5520 ( \6190 , \6184 , \6189 );
nand \U$5521 ( \6191 , \6179 , \6190 );
not \U$5522 ( \6192 , RIaa97c98_14);
not \U$5523 ( \6193 , RIaa97d10_15);
nand \U$5524 ( \6194 , \6192 , \6193 , RIaa97c20_13, RIaa97e00_17);
not \U$5525 ( \6195 , \6194 );
nand \U$5526 ( \6196 , \6195 , RIaa9c4c8_168);
not \U$5527 ( \6197 , RIaa97c20_13);
not \U$5528 ( \6198 , RIaa97e00_17);
nand \U$5529 ( \6199 , \6197 , \6198 , RIaa97c98_14, RIaa97d10_15);
not \U$5530 ( \6200 , \6199 );
nand \U$5531 ( \6201 , \6200 , RIaa9c540_169);
nand \U$5532 ( \6202 , RIaa97c20_13, RIaa97c98_14, RIaa97d10_15, RIaa97e00_17);
not \U$5533 ( \6203 , \6202 );
nand \U$5534 ( \6204 , \6203 , RIaa9c180_161);
nand \U$5535 ( \6205 , \6196 , \6201 , \6204 );
nor \U$5536 ( \6206 , \6191 , \6205 );
not \U$5537 ( \6207 , RIaa97e00_17);
nand \U$5538 ( \6208 , \6207 , \724 , \671 , RIaa97d10_15);
not \U$5539 ( \6209 , \6208 );
and \U$5540 ( \6210 , \6209 , RIaa9bf28_156);
nor \U$5541 ( \6211 , \6210 , \989 );
not \U$5542 ( \6212 , RIaa97c20_13);
nor \U$5543 ( \6213 , RIaa97d10_15, RIaa97e00_17);
nand \U$5544 ( \6214 , \6212 , \6213 , RIaa97c98_14);
not \U$5545 ( \6215 , \6214 );
nand \U$5546 ( \6216 , \6215 , RIaa9c2e8_164);
not \U$5547 ( \6217 , RIaa97d10_15);
nor \U$5548 ( \6218 , RIaa97c20_13, RIaa97c98_14);
nand \U$5549 ( \6219 , \6217 , \6218 , RIaa97e00_17);
not \U$5550 ( \6220 , \6219 );
nand \U$5551 ( \6221 , \6220 , RIaa9c018_158);
nand \U$5552 ( \6222 , \6211 , \6216 , \6221 );
not \U$5553 ( \6223 , RIaa9c090_159);
nor \U$5554 ( \6224 , RIaa97d10_15, RIaa97e00_17);
not \U$5555 ( \6225 , RIaa97d88_16);
and \U$5556 ( \6226 , \6224 , \6218 , \6225 );
not \U$5557 ( \6227 , \6226 );
or \U$5558 ( \6228 , \6223 , \6227 );
not \U$5559 ( \6229 , RIaa97e00_17);
nand \U$5560 ( \6230 , \6229 , RIaa97c20_13, RIaa97c98_14, RIaa97d10_15);
not \U$5561 ( \6231 , \6230 );
nand \U$5562 ( \6232 , \6231 , RIaa9c1f8_162);
nand \U$5563 ( \6233 , \6228 , \6232 );
nor \U$5564 ( \6234 , \6222 , \6233 );
not \U$5565 ( \6235 , RIaa9beb0_155);
not \U$5566 ( \6236 , RIaa97c20_13);
nand \U$5567 ( \6237 , \6236 , RIaa97d10_15, RIaa97e00_17, RIaa97c98_14);
not \U$5568 ( \6238 , \6237 );
not \U$5569 ( \6239 , \6238 );
or \U$5570 ( \6240 , \6235 , \6239 );
not \U$5571 ( \6241 , RIaa97c20_13);
not \U$5572 ( \6242 , RIaa97c98_14);
nand \U$5573 ( \6243 , \6241 , \6242 , RIaa97d10_15, RIaa97e00_17);
not \U$5574 ( \6244 , \6243 );
nand \U$5575 ( \6245 , \6244 , RIaa9bfa0_157);
nand \U$5576 ( \6246 , \6240 , \6245 );
not \U$5577 ( \6247 , RIaa9c3d8_166);
not \U$5578 ( \6248 , RIaa97c98_14);
nand \U$5579 ( \6249 , \6248 , RIaa97d10_15, RIaa97e00_17, RIaa97c20_13);
not \U$5580 ( \6250 , \6249 );
not \U$5581 ( \6251 , \6250 );
or \U$5582 ( \6252 , \6247 , \6251 );
not \U$5583 ( \6253 , RIaa97d10_15);
not \U$5584 ( \6254 , RIaa97e00_17);
nand \U$5585 ( \6255 , \6253 , \6254 , RIaa97c20_13, RIaa97c98_14);
not \U$5586 ( \6256 , \6255 );
nand \U$5587 ( \6257 , \6256 , RIaa9be38_154);
nand \U$5588 ( \6258 , \6252 , \6257 );
nor \U$5589 ( \6259 , \6246 , \6258 );
nand \U$5590 ( \6260 , \6206 , \6234 , \6259 );
not \U$5591 ( \6261 , \6260 );
not \U$5592 ( \6262 , \6261 );
and \U$5593 ( \6263 , \6113 , \6262 );
not \U$5594 ( \6264 , \6230 );
not \U$5595 ( \6265 , RIaa9c630_171);
not \U$5596 ( \6266 , \6265 );
and \U$5597 ( \6267 , \6264 , \6266 );
not \U$5598 ( \6268 , RIaa9c810_175);
nor \U$5599 ( \6269 , \6202 , \6268 );
nor \U$5600 ( \6270 , \6267 , \6269 );
not \U$5601 ( \6271 , \6214 );
not \U$5602 ( \6272 , RIaa9ccc0_185);
not \U$5603 ( \6273 , \6272 );
and \U$5604 ( \6274 , \6271 , \6273 );
not \U$5605 ( \6275 , RIaa9cc48_184);
nor \U$5606 ( \6276 , \6275 , \6188 );
nor \U$5607 ( \6277 , \6274 , \6276 );
nand \U$5608 ( \6278 , \6226 , RIaa9c798_174);
nand \U$5609 ( \6279 , \6270 , \6277 , \6278 );
not \U$5610 ( \6280 , \6199 );
not \U$5611 ( \6281 , RIaa9c900_177);
not \U$5612 ( \6282 , \6281 );
and \U$5613 ( \6283 , \6280 , \6282 );
and \U$5614 ( \6284 , \6250 , RIaa9cbd0_183);
nor \U$5615 ( \6285 , \6283 , \6284 );
not \U$5616 ( \6286 , \6255 );
not \U$5617 ( \6287 , RIaa9cd38_186);
not \U$5618 ( \6288 , \6287 );
and \U$5619 ( \6289 , \6286 , \6288 );
not \U$5620 ( \6290 , RIaa9c888_176);
nor \U$5621 ( \6291 , \6290 , \6172 );
nor \U$5622 ( \6292 , \6289 , \6291 );
nand \U$5623 ( \6293 , \6285 , \6292 );
nor \U$5624 ( \6294 , \6279 , \6293 );
not \U$5625 ( \6295 , \6219 );
not \U$5626 ( \6296 , RIaa9c6a8_172);
not \U$5627 ( \6297 , \6296 );
and \U$5628 ( \6298 , \6295 , \6297 );
nor \U$5629 ( \6299 , \6298 , \1030 );
nand \U$5630 ( \6300 , \6195 , RIaa9cb58_182);
nand \U$5631 ( \6301 , \6177 , RIaa9ca68_180);
nand \U$5632 ( \6302 , \6299 , \6300 , \6301 );
not \U$5633 ( \6303 , \6243 );
not \U$5634 ( \6304 , RIaa9c978_178);
not \U$5635 ( \6305 , \6304 );
and \U$5636 ( \6306 , \6303 , \6305 );
not \U$5637 ( \6307 , RIaa9cdb0_187);
nor \U$5638 ( \6308 , \6307 , \6237 );
nor \U$5639 ( \6309 , \6306 , \6308 );
not \U$5640 ( \6310 , \6208 );
not \U$5641 ( \6311 , RIaa9cae0_181);
not \U$5642 ( \6312 , \6311 );
and \U$5643 ( \6313 , \6310 , \6312 );
and \U$5644 ( \6314 , \6183 , RIaa9c9f0_179);
nor \U$5645 ( \6315 , \6313 , \6314 );
nand \U$5646 ( \6316 , \6309 , \6315 );
nor \U$5647 ( \6317 , \6302 , \6316 );
nand \U$5648 ( \6318 , \6294 , \6317 );
not \U$5649 ( \6319 , \6318 );
not \U$5650 ( \6320 , \6319 );
nor \U$5651 ( \6321 , \6263 , \3065 , \6320 );
nand \U$5652 ( \6322 , \6177 , RIaa9bd48_152);
nand \U$5653 ( \6323 , \6215 , RIaa9b6b8_138);
not \U$5654 ( \6324 , \6208 );
nand \U$5655 ( \6325 , \6324 , RIaa9bcd0_151);
nand \U$5656 ( \6326 , \6322 , \6323 , \6325 , \859 );
not \U$5657 ( \6327 , RIaa9b898_142);
not \U$5658 ( \6328 , \6226 );
or \U$5659 ( \6329 , \6327 , \6328 );
nand \U$5660 ( \6330 , \6231 , RIaa9b988_144);
nand \U$5661 ( \6331 , \6329 , \6330 );
nor \U$5662 ( \6332 , \6326 , \6331 );
not \U$5663 ( \6333 , RIaa9bbe0_149);
not \U$5664 ( \6334 , \6238 );
or \U$5665 ( \6335 , \6333 , \6334 );
not \U$5666 ( \6336 , \6255 );
nand \U$5667 ( \6337 , \6336 , RIaa9ba78_146);
nand \U$5668 ( \6338 , \6335 , \6337 );
not \U$5669 ( \6339 , RIaa9baf0_147);
not \U$5670 ( \6340 , \6250 );
or \U$5671 ( \6341 , \6339 , \6340 );
nand \U$5672 ( \6342 , \6244 , RIaa9bc58_150);
nand \U$5673 ( \6343 , \6341 , \6342 );
nor \U$5674 ( \6344 , \6338 , \6343 );
not \U$5675 ( \6345 , RIaa9b7a8_140);
not \U$5676 ( \6346 , \6200 );
or \U$5677 ( \6347 , \6345 , \6346 );
not \U$5678 ( \6348 , \6188 );
nand \U$5679 ( \6349 , \6348 , RIaa9b730_139);
nand \U$5680 ( \6350 , \6347 , \6349 );
not \U$5681 ( \6351 , RIaa9bdc0_153);
not \U$5682 ( \6352 , \6195 );
or \U$5683 ( \6353 , \6351 , \6352 );
nand \U$5684 ( \6354 , \6220 , RIaa9b820_141);
nand \U$5685 ( \6355 , \6353 , \6354 );
nor \U$5686 ( \6356 , \6350 , \6355 );
not \U$5687 ( \6357 , \6172 );
and \U$5688 ( \6358 , RIaa9b640_137, \6357 );
and \U$5689 ( \6359 , \6183 , RIaa9bb68_148);
nand \U$5690 ( \6360 , RIaa97c20_13, RIaa97c98_14, RIaa97d10_15, RIaa97e00_17);
not \U$5691 ( \6361 , \6360 );
not \U$5692 ( \6362 , \6361 );
not \U$5693 ( \6363 , RIaa9ba00_145);
nor \U$5694 ( \6364 , \6362 , \6363 );
nor \U$5695 ( \6365 , \6358 , \6359 , \6364 );
nand \U$5696 ( \6366 , \6332 , \6344 , \6356 , \6365 );
not \U$5697 ( \6367 , \6366 );
not \U$5698 ( \6368 , \6367 );
or \U$5699 ( \6369 , \6118 , \6368 );
or \U$5700 ( \6370 , \6113 , \6262 );
nand \U$5701 ( \6371 , \6369 , \6370 );
or \U$5702 ( \6372 , \6321 , \6371 );
not \U$5703 ( \6373 , \6120 );
nand \U$5704 ( \6374 , \6348 , RIaa9b190_127);
nand \U$5705 ( \6375 , \6215 , RIaa9b0a0_125);
nand \U$5706 ( \6376 , \6177 , RIaa9b460_133);
nand \U$5707 ( \6377 , \6250 , RIaa9b2f8_130);
nand \U$5708 ( \6378 , \6374 , \6375 , \6376 , \6377 );
not \U$5709 ( \6379 , \6219 );
not \U$5710 ( \6380 , \924 );
and \U$5711 ( \6381 , \6379 , \6380 );
and \U$5712 ( \6382 , \6183 , RIaa9b370_131);
nor \U$5713 ( \6383 , \6381 , \6382 );
not \U$5714 ( \6384 , \6194 );
not \U$5715 ( \6385 , RIaa9b4d8_134);
not \U$5716 ( \6386 , \6385 );
and \U$5717 ( \6387 , \6384 , \6386 );
and \U$5718 ( \6388 , \6324 , RIaa9b5c8_136);
nor \U$5719 ( \6389 , \6387 , \6388 );
nand \U$5720 ( \6390 , \6383 , \6389 );
nor \U$5721 ( \6391 , \6378 , \6390 );
and \U$5722 ( \6392 , \6231 , RIaa9afb0_123);
and \U$5723 ( \6393 , \6203 , RIaa9b028_124);
nor \U$5724 ( \6394 , \6392 , \6393 );
not \U$5725 ( \6395 , \6199 );
not \U$5726 ( \6396 , RIaa9b208_128);
not \U$5727 ( \6397 , \6396 );
and \U$5728 ( \6398 , \6395 , \6397 );
nor \U$5729 ( \6399 , \6398 , \944 );
nand \U$5730 ( \6400 , \6226 , RIaa9aec0_121);
nand \U$5731 ( \6401 , \6394 , \6399 , \6400 );
and \U$5732 ( \6402 , \6256 , RIaa9b280_129);
and \U$5733 ( \6403 , \6357 , RIaa9b118_126);
nor \U$5734 ( \6404 , \6402 , \6403 );
and \U$5735 ( \6405 , \6244 , RIaa9b550_135);
and \U$5736 ( \6406 , \6238 , RIaa9b3e8_132);
nor \U$5737 ( \6407 , \6405 , \6406 );
nand \U$5738 ( \6408 , \6404 , \6407 );
nor \U$5739 ( \6409 , \6401 , \6408 );
nand \U$5740 ( \6410 , \6391 , \6409 );
not \U$5741 ( \6411 , \6410 );
not \U$5742 ( \6412 , \6411 );
and \U$5743 ( \6413 , \6373 , \6412 );
and \U$5744 ( \6414 , \6118 , \6368 );
nor \U$5745 ( \6415 , \6413 , \6414 );
nand \U$5746 ( \6416 , \6372 , \6415 );
not \U$5747 ( \6417 , \1073 );
not \U$5748 ( \6418 , \6417 );
not \U$5749 ( \6419 , \6336 );
not \U$5750 ( \6420 , RIaa9d2d8_198);
or \U$5751 ( \6421 , \6419 , \6420 );
not \U$5752 ( \6422 , \6357 );
not \U$5753 ( \6423 , RIaa9d0f8_194);
or \U$5754 ( \6424 , \6422 , \6423 );
nand \U$5755 ( \6425 , \6421 , \6424 );
not \U$5756 ( \6426 , RIaa9d440_201);
not \U$5757 ( \6427 , \6237 );
not \U$5758 ( \6428 , \6427 );
or \U$5759 ( \6429 , \6426 , \6428 );
nand \U$5760 ( \6430 , \6244 , RIaa9d4b8_202);
nand \U$5761 ( \6431 , \6429 , \6430 );
nor \U$5762 ( \6432 , \6425 , \6431 );
and \U$5763 ( \6433 , RIaa9d260_197, \6200 );
and \U$5764 ( \6434 , \6183 , RIaa9d3c8_200);
not \U$5765 ( \6435 , RIaa9d170_195);
or \U$5766 ( \6436 , \6214 , \6435 );
nand \U$5767 ( \6437 , \6436 , \738 );
nor \U$5768 ( \6438 , \6433 , \6434 , \6437 );
not \U$5769 ( \6439 , \6231 );
not \U$5770 ( \6440 , \6439 );
not \U$5771 ( \6441 , RIaa9cf18_190);
not \U$5772 ( \6442 , \6441 );
and \U$5773 ( \6443 , \6440 , \6442 );
not \U$5774 ( \6444 , RIaa9cf90_191);
nor \U$5775 ( \6445 , \6444 , \6362 );
nor \U$5776 ( \6446 , \6443 , \6445 );
nand \U$5777 ( \6447 , \6432 , \6438 , \6446 );
buf \U$5778 ( \6448 , \6226 );
nand \U$5779 ( \6449 , \6448 , RIaa9d080_193);
nand \U$5780 ( \6450 , \6177 , RIaa9d5a8_204);
nand \U$5781 ( \6451 , \6195 , RIaa9d620_205);
and \U$5782 ( \6452 , \6449 , \6450 , \6451 );
not \U$5783 ( \6453 , RIaa9d350_199);
not \U$5784 ( \6454 , \6250 );
or \U$5785 ( \6455 , \6453 , \6454 );
nand \U$5786 ( \6456 , \6220 , RIaa9d008_192);
nand \U$5787 ( \6457 , \6455 , \6456 );
not \U$5788 ( \6458 , RIaa9d1e8_196);
not \U$5789 ( \6459 , \6348 );
or \U$5790 ( \6460 , \6458 , \6459 );
nand \U$5791 ( \6461 , \6324 , RIaa9d530_203);
nand \U$5792 ( \6462 , \6460 , \6461 );
nor \U$5793 ( \6463 , \6457 , \6462 );
nand \U$5794 ( \6464 , \6452 , \6463 );
nor \U$5795 ( \6465 , \6447 , \6464 );
not \U$5796 ( \6466 , \6465 );
not \U$5797 ( \6467 , \6466 );
and \U$5798 ( \6468 , \6418 , \6467 );
and \U$5799 ( \6469 , \6120 , \6411 );
nor \U$5800 ( \6470 , \6468 , \6469 );
and \U$5801 ( \6471 , \6416 , \6470 );
and \U$5802 ( \6472 , \6417 , \6466 );
and \U$5803 ( \6473 , \6427 , RIaa9abf0_115);
and \U$5804 ( \6474 , \6361 , RIaa9a830_107);
nor \U$5805 ( \6475 , \6473 , \6474 );
and \U$5806 ( \6476 , \6183 , RIaa9ab78_114);
not \U$5807 ( \6477 , \1109 );
nor \U$5808 ( \6478 , \6476 , \6477 );
nand \U$5809 ( \6479 , \6226 , RIaa9a6c8_104);
nand \U$5810 ( \6480 , \6475 , \6478 , \6479 );
nand \U$5811 ( \6481 , \6215 , RIaa9a8a8_108);
nand \U$5812 ( \6482 , \6220 , RIaa9a650_103);
nand \U$5813 ( \6483 , \6231 , RIaa9a7b8_106);
nand \U$5814 ( \6484 , \6348 , RIaa9a998_110);
nand \U$5815 ( \6485 , \6481 , \6482 , \6483 , \6484 );
nor \U$5816 ( \6486 , \6480 , \6485 );
nand \U$5817 ( \6487 , \6336 , RIaa9aa88_112);
nand \U$5818 ( \6488 , \6357 , RIaa9a920_109);
nand \U$5819 ( \6489 , \6250 , RIaa9ab00_113);
nand \U$5820 ( \6490 , \6244 , RIaa9ace0_117);
nand \U$5821 ( \6491 , \6487 , \6488 , \6489 , \6490 );
nand \U$5822 ( \6492 , \6177 , RIaa9ad58_118);
nand \U$5823 ( \6493 , \6195 , RIaa9add0_119);
nand \U$5824 ( \6494 , \6200 , RIaa9aa10_111);
nand \U$5825 ( \6495 , \6324 , RIaa9ac68_116);
nand \U$5826 ( \6496 , \6492 , \6493 , \6494 , \6495 );
nor \U$5827 ( \6497 , \6491 , \6496 );
nand \U$5828 ( \6498 , \6486 , \6497 );
buf \U$5829 ( \6499 , \6498 );
and \U$5830 ( \6500 , \1135 , \6499 );
nor \U$5831 ( \6501 , \6471 , \6472 , \6500 );
not \U$5832 ( \6502 , \6255 );
nand \U$5833 ( \6503 , \6502 , RIaa9a470_99);
nand \U$5834 ( \6504 , \6357 , RIaa9a308_96);
nand \U$5835 ( \6505 , \6244 , RIaa9a128_92);
nand \U$5836 ( \6506 , \6250 , RIaa9a560_101);
nand \U$5837 ( \6507 , \6503 , \6504 , \6505 , \6506 );
not \U$5838 ( \6508 , \6507 );
nand \U$5839 ( \6509 , \6348 , RIaa9a380_97);
nand \U$5840 ( \6510 , \6220 , RIaa99e58_86);
nand \U$5841 ( \6511 , \6177 , RIaa9a0b0_91);
nand \U$5842 ( \6512 , \6509 , \6510 , \6511 , \1216 );
not \U$5843 ( \6513 , RIaa99f48_88);
not \U$5844 ( \6514 , \6231 );
or \U$5845 ( \6515 , \6513 , \6514 );
nand \U$5846 ( \6516 , \6361 , RIaa9a038_90);
nand \U$5847 ( \6517 , \6515 , \6516 );
nor \U$5848 ( \6518 , \6512 , \6517 );
buf \U$5849 ( \6519 , \6226 );
and \U$5850 ( \6520 , \6519 , RIaa99fc0_89);
not \U$5851 ( \6521 , RIaa9a218_94);
not \U$5852 ( \6522 , \6195 );
or \U$5853 ( \6523 , \6521 , \6522 );
nand \U$5854 ( \6524 , \6324 , RIaa9a1a0_93);
nand \U$5855 ( \6525 , \6523 , \6524 );
nor \U$5856 ( \6526 , \6520 , \6525 );
not \U$5857 ( \6527 , RIaa9a290_95);
not \U$5858 ( \6528 , \6215 );
or \U$5859 ( \6529 , \6527 , \6528 );
nand \U$5860 ( \6530 , \6427 , RIaa9a5d8_102);
nand \U$5861 ( \6531 , \6529 , \6530 );
not \U$5862 ( \6532 , RIaa9a4e8_100);
not \U$5863 ( \6533 , \6183 );
or \U$5864 ( \6534 , \6532 , \6533 );
nand \U$5865 ( \6535 , \6200 , RIaa9a3f8_98);
nand \U$5866 ( \6536 , \6534 , \6535 );
nor \U$5867 ( \6537 , \6531 , \6536 );
nand \U$5868 ( \6538 , \6508 , \6518 , \6526 , \6537 );
buf \U$5869 ( \6539 , \6538 );
not \U$5870 ( \6540 , \1343 );
or \U$5871 ( \6541 , \6539 , \6540 );
not \U$5872 ( \6542 , \6103 );
not \U$5873 ( \6543 , RIaa99b88_80);
not \U$5874 ( \6544 , \6177 );
or \U$5875 ( \6545 , \6543 , \6544 );
nand \U$5876 ( \6546 , \6324 , RIaa99b10_79);
nand \U$5877 ( \6547 , \6545 , \6546 );
not \U$5878 ( \6548 , RIaa99750_71);
not \U$5879 ( \6549 , \6183 );
or \U$5880 ( \6550 , \6548 , \6549 );
nand \U$5881 ( \6551 , \6550 , \1273 );
nor \U$5882 ( \6552 , \6547 , \6551 );
not \U$5883 ( \6553 , \6439 );
not \U$5884 ( \6554 , \1268 );
and \U$5885 ( \6555 , \6553 , \6554 );
and \U$5886 ( \6556 , \6448 , RIaa998b8_74);
nor \U$5887 ( \6557 , \6555 , \6556 );
nand \U$5888 ( \6558 , \6552 , \6557 );
nand \U$5889 ( \6559 , \6195 , RIaa99c00_81);
nand \U$5890 ( \6560 , \6200 , RIaa996d8_70);
nand \U$5891 ( \6561 , \6220 , RIaa99840_73);
nand \U$5892 ( \6562 , \6348 , RIaa99660_69);
nand \U$5893 ( \6563 , \6559 , \6560 , \6561 , \6562 );
nor \U$5894 ( \6564 , \6558 , \6563 );
nand \U$5895 ( \6565 , \6336 , RIaa99cf0_83);
nand \U$5896 ( \6566 , \6427 , RIaa99de0_85);
nand \U$5897 ( \6567 , \6244 , RIaa99a98_78);
nand \U$5898 ( \6568 , \6250 , RIaa997c8_72);
nand \U$5899 ( \6569 , \6565 , \6566 , \6567 , \6568 );
nand \U$5900 ( \6570 , \6215 , RIaa99d68_84);
nand \U$5901 ( \6571 , \6357 , RIaa99c78_82);
nand \U$5902 ( \6572 , \6361 , RIaa99a20_77);
nand \U$5903 ( \6573 , \6570 , \6571 , \6572 );
nor \U$5904 ( \6574 , \6569 , \6573 );
nand \U$5905 ( \6575 , \6564 , \6574 );
buf \U$5906 ( \6576 , \6575 );
or \U$5907 ( \6577 , \6542 , \6576 );
or \U$5908 ( \6578 , \6499 , \1135 );
nand \U$5909 ( \6579 , \6541 , \6577 , \6578 );
or \U$5910 ( \6580 , \6501 , \6579 );
and \U$5911 ( \6581 , \6540 , \6576 , \6539 );
nor \U$5912 ( \6582 , \6581 , \6542 );
and \U$5913 ( \6583 , \6540 , \6539 );
nor \U$5914 ( \6584 , \6583 , \6576 );
or \U$5915 ( \6585 , \6582 , \6584 );
nand \U$5916 ( \6586 , \6580 , \6585 );
nand \U$5917 ( \6587 , \6519 , RIaa9df08_224);
buf \U$5918 ( \6588 , \6220 );
nand \U$5919 ( \6589 , \6588 , RIaa9de90_223);
and \U$5920 ( \6590 , \6587 , \6589 , \1732 );
and \U$5921 ( \6591 , \6195 , RIaa9e250_231);
and \U$5922 ( \6592 , \6231 , RIaa9e0e8_228);
nor \U$5923 ( \6593 , \6591 , \6592 );
and \U$5924 ( \6594 , \6177 , RIaa9e1d8_230);
buf \U$5925 ( \6595 , \6324 );
and \U$5926 ( \6596 , \6595 , RIaa9dff8_226);
nor \U$5927 ( \6597 , \6594 , \6596 );
buf \U$5928 ( \6598 , \6244 );
and \U$5929 ( \6599 , \6598 , RIaa9e070_227);
and \U$5930 ( \6600 , \6361 , RIaa9e160_229);
nor \U$5931 ( \6601 , \6599 , \6600 );
nand \U$5932 ( \6602 , \6590 , \6593 , \6597 , \6601 );
and \U$5933 ( \6603 , \6336 , RIaa9e2c8_232);
buf \U$5934 ( \6604 , \6357 );
and \U$5935 ( \6605 , \6604 , RIaa9e340_233);
nor \U$5936 ( \6606 , \6603 , \6605 );
and \U$5937 ( \6607 , \6250 , RIaa9e430_235);
buf \U$5938 ( \6608 , \6238 );
and \U$5939 ( \6609 , \6608 , RIaa9e610_239);
nor \U$5940 ( \6610 , \6607 , \6609 );
not \U$5941 ( \6611 , \6214 );
not \U$5942 ( \6612 , \1746 );
and \U$5943 ( \6613 , \6611 , \6612 );
buf \U$5944 ( \6614 , \6183 );
and \U$5945 ( \6615 , \6614 , RIaa9e3b8_234);
nor \U$5946 ( \6616 , \6613 , \6615 );
buf \U$5947 ( \6617 , \6200 );
and \U$5948 ( \6618 , \6617 , RIaa9e4a8_236);
and \U$5949 ( \6619 , \6348 , RIaa9e520_237);
nor \U$5950 ( \6620 , \6618 , \6619 );
nand \U$5951 ( \6621 , \6606 , \6610 , \6616 , \6620 );
nor \U$5952 ( \6622 , \6602 , \6621 );
and \U$5953 ( \6623 , \1768 , \6622 );
nand \U$5954 ( \6624 , \6519 , RIaa986e8_36);
nand \U$5955 ( \6625 , \6588 , RIaa98670_35);
and \U$5956 ( \6626 , \6624 , \6625 , \1857 );
and \U$5957 ( \6627 , \6195 , RIaa98a30_43);
and \U$5958 ( \6628 , \6231 , RIaa987d8_38);
nor \U$5959 ( \6629 , \6627 , \6628 );
and \U$5960 ( \6630 , \6177 , RIaa989b8_42);
and \U$5961 ( \6631 , \6595 , RIaa988c8_40);
nor \U$5962 ( \6632 , \6630 , \6631 );
and \U$5963 ( \6633 , \6598 , RIaa98940_41);
and \U$5964 ( \6634 , \6361 , RIaa98850_39);
nor \U$5965 ( \6635 , \6633 , \6634 );
nand \U$5966 ( \6636 , \6626 , \6629 , \6632 , \6635 );
not \U$5967 ( \6637 , \6419 );
and \U$5968 ( \6638 , \6637 , RIaa98c88_48);
and \U$5969 ( \6639 , \6348 , RIaa98df0_51);
nor \U$5970 ( \6640 , \6638 , \6639 );
and \U$5971 ( \6641 , \6250 , RIaa98c10_47);
and \U$5972 ( \6642 , \6608 , RIaa98d00_49);
nor \U$5973 ( \6643 , \6641 , \6642 );
and \U$5974 ( \6644 , \6215 , RIaa98b20_45);
and \U$5975 ( \6645 , \6604 , RIaa98aa8_44);
nor \U$5976 ( \6646 , \6644 , \6645 );
and \U$5977 ( \6647 , \6614 , RIaa98b98_46);
and \U$5978 ( \6648 , \6617 , RIaa98d78_50);
nor \U$5979 ( \6649 , \6647 , \6648 );
nand \U$5980 ( \6650 , \6640 , \6643 , \6646 , \6649 );
nor \U$5981 ( \6651 , \6636 , \6650 );
and \U$5982 ( \6652 , \1879 , \6651 );
nor \U$5983 ( \6653 , \6623 , \6652 );
nand \U$5984 ( \6654 , \6519 , RIaa9dad0_215);
nand \U$5985 ( \6655 , \6588 , RIaa9da58_214);
and \U$5986 ( \6656 , \6654 , \6655 , \1611 );
and \U$5987 ( \6657 , \6177 , RIaa9dcb0_219);
and \U$5988 ( \6658 , \6595 , RIaa9dbc0_217);
nor \U$5989 ( \6659 , \6657 , \6658 );
and \U$5990 ( \6660 , \6195 , RIaa9dd28_220);
and \U$5991 ( \6661 , \6231 , RIaa9dda0_221);
nor \U$5992 ( \6662 , \6660 , \6661 );
and \U$5993 ( \6663 , \6598 , RIaa9dc38_218);
not \U$5994 ( \6664 , \6362 );
and \U$5995 ( \6665 , \6664 , RIaa9de18_222);
nor \U$5996 ( \6666 , \6663 , \6665 );
and \U$5997 ( \6667 , \6656 , \6659 , \6662 , \6666 );
and \U$5998 ( \6668 , \6215 , RIaa9d788_208);
and \U$5999 ( \6669 , \6617 , RIaa9d968_212);
nor \U$6000 ( \6670 , \6668 , \6669 );
and \U$6001 ( \6671 , \6250 , RIaa9d8f0_211);
and \U$6002 ( \6672 , \6608 , RIaa9d800_209);
nor \U$6003 ( \6673 , \6671 , \6672 );
and \U$6004 ( \6674 , \6637 , RIaa9d698_206);
and \U$6005 ( \6675 , \6604 , RIaa9d710_207);
nor \U$6006 ( \6676 , \6674 , \6675 );
and \U$6007 ( \6677 , \6614 , RIaa9d878_210);
and \U$6008 ( \6678 , \6348 , RIaa9d9e0_213);
nor \U$6009 ( \6679 , \6677 , \6678 );
and \U$6010 ( \6680 , \6670 , \6673 , \6676 , \6679 );
nand \U$6011 ( \6681 , \6667 , \6680 );
not \U$6012 ( \6682 , \6681 );
nand \U$6013 ( \6683 , \1655 , \6682 );
nand \U$6014 ( \6684 , \6250 , RIaa99228_60);
nand \U$6015 ( \6685 , \6502 , RIaa99480_65);
nand \U$6016 ( \6686 , \6357 , RIaa990c0_57);
nand \U$6017 ( \6687 , \6324 , RIaa99318_62);
nand \U$6018 ( \6688 , \6684 , \6685 , \6686 , \6687 );
nand \U$6019 ( \6689 , \6177 , RIaa99390_63);
nand \U$6020 ( \6690 , \6195 , RIaa99408_64);
nand \U$6021 ( \6691 , \6200 , RIaa995e8_68);
nand \U$6022 ( \6692 , \6348 , RIaa99570_67);
nand \U$6023 ( \6693 , \6689 , \6690 , \6691 , \6692 );
nor \U$6024 ( \6694 , \6688 , \6693 );
and \U$6025 ( \6695 , \6427 , RIaa994f8_66);
and \U$6026 ( \6696 , \6361 , RIaa99048_56);
nor \U$6027 ( \6697 , \6695 , \6696 );
nand \U$6028 ( \6698 , \6448 , RIaa98ee0_53);
and \U$6029 ( \6699 , \6220 , RIaa98e68_52);
not \U$6030 ( \6700 , \1661 );
nor \U$6031 ( \6701 , \6699 , \6700 );
nand \U$6032 ( \6702 , \6697 , \6698 , \6701 );
nand \U$6033 ( \6703 , \6215 , RIaa99138_58);
nand \U$6034 ( \6704 , \6244 , RIaa992a0_61);
nand \U$6035 ( \6705 , \6231 , RIaa98fd0_55);
nand \U$6036 ( \6706 , \6183 , RIaa991b0_59);
nand \U$6037 ( \6707 , \6703 , \6704 , \6705 , \6706 );
nor \U$6038 ( \6708 , \6702 , \6707 );
nand \U$6039 ( \6709 , \6694 , \6708 );
buf \U$6040 ( \6710 , \6709 );
not \U$6041 ( \6711 , \6710 );
nand \U$6042 ( \6712 , \6711 , \6071 );
nand \U$6043 ( \6713 , \6586 , \6653 , \6683 , \6712 );
or \U$6044 ( \6714 , \1768 , \6622 );
or \U$6045 ( \6715 , \6682 , \1655 );
not \U$6046 ( \6716 , \6071 );
nand \U$6047 ( \6717 , \6716 , \6683 , \6710 );
nand \U$6048 ( \6718 , \6714 , \6715 , \6717 );
and \U$6049 ( \6719 , \6718 , \6653 );
or \U$6050 ( \6720 , \1879 , \6651 );
nand \U$6051 ( \6721 , \6519 , RIaa97e78_18);
nand \U$6052 ( \6722 , \6588 , RIaa97ef0_19);
and \U$6053 ( \6723 , \6721 , \6722 , \2057 );
and \U$6054 ( \6724 , \6195 , RIaa98238_26);
and \U$6055 ( \6725 , \6231 , RIaa980d0_23);
nor \U$6056 ( \6726 , \6724 , \6725 );
and \U$6057 ( \6727 , \6177 , RIaa981c0_25);
and \U$6058 ( \6728 , \6595 , RIaa97fe0_21);
nor \U$6059 ( \6729 , \6727 , \6728 );
and \U$6060 ( \6730 , \6598 , RIaa98058_22);
and \U$6061 ( \6731 , \6361 , RIaa98148_24);
nor \U$6062 ( \6732 , \6730 , \6731 );
nand \U$6063 ( \6733 , \6723 , \6726 , \6729 , \6732 );
and \U$6064 ( \6734 , \6617 , RIaa98490_31);
and \U$6065 ( \6735 , \6348 , RIaa98508_32);
nor \U$6066 ( \6736 , \6734 , \6735 );
and \U$6067 ( \6737 , \6250 , RIaa98418_30);
and \U$6068 ( \6738 , \6608 , RIaa985f8_34);
nor \U$6069 ( \6739 , \6737 , \6738 );
and \U$6070 ( \6740 , \6637 , RIaa982b0_27);
and \U$6071 ( \6741 , \6604 , RIaa98328_28);
nor \U$6072 ( \6742 , \6740 , \6741 );
and \U$6073 ( \6743 , \6215 , RIaa98580_33);
and \U$6074 ( \6744 , \6614 , RIaa983a0_29);
nor \U$6075 ( \6745 , \6743 , \6744 );
nand \U$6076 ( \6746 , \6736 , \6739 , \6742 , \6745 );
nor \U$6077 ( \6747 , \6733 , \6746 );
or \U$6078 ( \6748 , \2074 , \6747 );
nand \U$6079 ( \6749 , \6720 , \6748 );
nor \U$6080 ( \6750 , \6719 , \6749 );
not \U$6081 ( \6751 , \6160 );
not \U$6082 ( \6752 , RIaa97680_1);
and \U$6083 ( \6753 , \6751 , \6752 );
and \U$6084 ( \6754 , \6160 , RIaa97680_1);
nor \U$6085 ( \6755 , \6753 , \6754 );
not \U$6086 ( \6756 , \6755 );
nand \U$6087 ( \6757 , \6756 , \2074 );
and \U$6088 ( \6758 , \6713 , \6750 , \6757 );
and \U$6089 ( \6759 , \2074 , \6755 , \6747 );
nor \U$6090 ( \6760 , \6758 , \6759 );
nor \U$6091 ( \6761 , \6170 , \6760 );
and \U$6092 ( \6762 , \6713 , \6750 , \2073 , \6755 );
nor \U$6093 ( \6763 , \6761 , \6762 );
buf \U$6094 ( \6764 , \6763 );
not \U$6095 ( \6765 , \6764 );
nand \U$6096 ( \6766 , \6069 , \6070 , \6765 );
or \U$6097 ( \6767 , \6056 , \6766 );
not \U$6098 ( \6768 , \6765 );
buf \U$6099 ( \6769 , \6768 );
not \U$6100 ( \6770 , \6747 );
nand \U$6101 ( \6771 , \6770 , \2076 );
not \U$6102 ( \6772 , \6771 );
or \U$6103 ( \6773 , \1825 , \6651 );
not \U$6104 ( \6774 , \6773 );
not \U$6105 ( \6775 , \852 );
not \U$6106 ( \6776 , \6366 );
or \U$6107 ( \6777 , \6775 , \6776 );
not \U$6108 ( \6778 , RIaa977e8_4);
not \U$6109 ( \6779 , \6260 );
or \U$6110 ( \6780 , \6778 , \6779 );
nand \U$6111 ( \6781 , \6318 , \1017 );
nand \U$6112 ( \6782 , \6780 , \6781 );
nand \U$6113 ( \6783 , \6261 , \849 );
nand \U$6114 ( \6784 , \6782 , \6783 );
nand \U$6115 ( \6785 , \6777 , \6784 );
not \U$6116 ( \6786 , \6785 );
not \U$6117 ( \6787 , \6410 );
not \U$6118 ( \6788 , \960 );
and \U$6119 ( \6789 , \6787 , \6788 );
and \U$6120 ( \6790 , \6367 , \853 );
nor \U$6121 ( \6791 , \6789 , \6790 );
not \U$6122 ( \6792 , \6791 );
or \U$6123 ( \6793 , \6786 , \6792 );
nand \U$6124 ( \6794 , \6411 , \959 );
not \U$6125 ( \6795 , \6410 );
not \U$6126 ( \6796 , \959 );
and \U$6127 ( \6797 , \6795 , \6796 );
and \U$6128 ( \6798 , \6410 , \959 );
nor \U$6129 ( \6799 , \6797 , \6798 );
and \U$6130 ( \6800 , \6794 , \6799 );
nor \U$6131 ( \6801 , \6465 , \842 );
nor \U$6132 ( \6802 , \6800 , \6801 );
nand \U$6133 ( \6803 , \6793 , \6802 );
nand \U$6134 ( \6804 , \6709 , \1708 );
nand \U$6135 ( \6805 , \6575 , \1311 );
nand \U$6136 ( \6806 , \6498 , \1130 );
nand \U$6137 ( \6807 , \6538 , \1254 );
and \U$6138 ( \6808 , \6804 , \6805 , \6806 , \6807 );
not \U$6139 ( \6809 , \6808 );
or \U$6140 ( \6810 , \6803 , \6809 );
and \U$6141 ( \6811 , \6465 , \842 );
and \U$6142 ( \6812 , \6808 , \6811 );
nor \U$6143 ( \6813 , \6498 , \1130 );
and \U$6144 ( \6814 , \6813 , \6807 );
nor \U$6145 ( \6815 , \6538 , \1254 );
nor \U$6146 ( \6816 , \6814 , \6815 );
nand \U$6147 ( \6817 , \6804 , \6805 );
or \U$6148 ( \6818 , \6816 , \6817 );
nor \U$6149 ( \6819 , \6575 , \1311 );
and \U$6150 ( \6820 , \6819 , \6804 );
nor \U$6151 ( \6821 , \1708 , \6709 );
nor \U$6152 ( \6822 , \6820 , \6821 );
nand \U$6153 ( \6823 , \6818 , \6822 );
nor \U$6154 ( \6824 , \6812 , \6823 );
nand \U$6155 ( \6825 , \6810 , \6824 );
nor \U$6156 ( \6826 , \1604 , \6681 );
or \U$6157 ( \6827 , \6825 , \6826 );
nand \U$6158 ( \6828 , \1604 , \6681 );
nand \U$6159 ( \6829 , \6827 , \6828 );
not \U$6160 ( \6830 , \6622 );
nand \U$6161 ( \6831 , \6830 , \1774 );
not \U$6162 ( \6832 , \6831 );
or \U$6163 ( \6833 , \6829 , \6832 );
nand \U$6164 ( \6834 , \1773 , \6622 );
nand \U$6165 ( \6835 , \6833 , \6834 );
not \U$6166 ( \6836 , \6835 );
or \U$6167 ( \6837 , \6774 , \6836 );
nand \U$6168 ( \6838 , \1825 , \6651 );
nand \U$6169 ( \6839 , \6837 , \6838 );
not \U$6170 ( \6840 , \6839 );
or \U$6171 ( \6841 , \6772 , \6840 );
not \U$6172 ( \6842 , \2076 );
nand \U$6173 ( \6843 , \6842 , \6747 );
nand \U$6174 ( \6844 , \6841 , \6843 );
nand \U$6175 ( \6845 , \6844 , \2012 );
buf \U$6176 ( \6846 , \6845 );
not \U$6177 ( \6847 , \6846 );
not \U$6178 ( \6848 , \1861 );
not \U$6179 ( \6849 , \6848 );
not \U$6180 ( \6850 , RIaa9ec28_252);
not \U$6181 ( \6851 , \6850 );
and \U$6182 ( \6852 , \6849 , \6851 );
nor \U$6183 ( \6853 , \6852 , \1546 );
buf \U$6184 ( \6854 , \1874 );
and \U$6185 ( \6855 , \6854 , RIaa9ef70_259);
not \U$6186 ( \6856 , \1868 );
and \U$6187 ( \6857 , \6856 , RIaa9efe8_260);
nor \U$6188 ( \6858 , \6855 , \6857 );
and \U$6189 ( \6859 , \2061 , RIaa9eca0_253);
and \U$6190 ( \6860 , \2064 , RIaa9ee80_257);
nor \U$6191 ( \6861 , \6859 , \6860 );
buf \U$6192 ( \6862 , \1645 );
and \U$6193 ( \6863 , \6862 , RIaa9eac0_249);
and \U$6194 ( \6864 , \1372 , \6362 );
not \U$6195 ( \6865 , \1372 );
and \U$6196 ( \6866 , \6865 , \6439 );
or \U$6197 ( \6867 , \6864 , \6866 );
not \U$6198 ( \6868 , \6867 );
and \U$6199 ( \6869 , \6868 , RIaa9eb38_250);
nand \U$6200 ( \6870 , \6361 , \1373 );
nand \U$6201 ( \6871 , \6870 , \6225 );
and \U$6202 ( \6872 , \6871 , RIaa9ebb0_251);
nor \U$6203 ( \6873 , \6863 , \6869 , \6872 );
nand \U$6204 ( \6874 , \6853 , \6858 , \6861 , \6873 );
and \U$6205 ( \6875 , \1651 , RIaa9eef8_258);
not \U$6206 ( \6876 , \2020 );
and \U$6207 ( \6877 , \6876 , RIaa9f1c8_264);
nor \U$6208 ( \6878 , \6875 , \6877 );
and \U$6209 ( \6879 , \2023 , RIaa9ed18_254);
and \U$6210 ( \6880 , \1832 , RIaa9f0d8_262);
nor \U$6211 ( \6881 , \6879 , \6880 );
not \U$6212 ( \6882 , \1670 );
not \U$6213 ( \6883 , \6882 );
and \U$6214 ( \6884 , \6883 , RIaa9f150_263);
and \U$6215 ( \6885 , \1642 , RIaa9f060_261);
nor \U$6216 ( \6886 , \6884 , \6885 );
and \U$6217 ( \6887 , \1846 , RIaa9ee08_256);
not \U$6218 ( \6888 , \1647 );
not \U$6219 ( \6889 , \6888 );
and \U$6220 ( \6890 , \6889 , RIaa9ed90_255);
nor \U$6221 ( \6891 , \6887 , \6890 );
nand \U$6222 ( \6892 , \6878 , \6881 , \6886 , \6891 );
or \U$6223 ( \6893 , \6874 , \6892 );
buf \U$6224 ( \6894 , \6893 );
and \U$6225 ( \6895 , \6847 , \6894 );
nor \U$6226 ( \6896 , \6844 , \2012 );
not \U$6227 ( \6897 , \6896 );
nand \U$6228 ( \6898 , \6897 , \6845 );
not \U$6229 ( \6899 , \6839 );
nand \U$6230 ( \6900 , \6843 , \6771 );
not \U$6231 ( \6901 , \6900 );
and \U$6232 ( \6902 , \6899 , \6901 );
and \U$6233 ( \6903 , \6839 , \6900 );
nor \U$6234 ( \6904 , \6902 , \6903 );
not \U$6235 ( \6905 , \6904 );
nor \U$6236 ( \6906 , \6898 , \6905 );
not \U$6237 ( \6907 , \6906 );
nand \U$6238 ( \6908 , \6898 , \6905 );
not \U$6239 ( \6909 , \6835 );
nand \U$6240 ( \6910 , \6838 , \6773 );
not \U$6241 ( \6911 , \6910 );
and \U$6242 ( \6912 , \6909 , \6911 );
and \U$6243 ( \6913 , \6835 , \6910 );
nor \U$6244 ( \6914 , \6912 , \6913 );
buf \U$6245 ( \6915 , \6914 );
not \U$6246 ( \6916 , \6915 );
nand \U$6247 ( \6917 , \6905 , \6916 );
nand \U$6248 ( \6918 , \6904 , \6915 );
nand \U$6249 ( \6919 , \6917 , \6918 );
nand \U$6250 ( \6920 , \6907 , \6908 , \6919 );
not \U$6251 ( \6921 , \6920 );
buf \U$6252 ( \6922 , \6921 );
not \U$6253 ( \6923 , \6922 );
not \U$6254 ( \6924 , \6919 );
buf \U$6255 ( \6925 , \6924 );
not \U$6256 ( \6926 , \6925 );
and \U$6257 ( \6927 , \6923 , \6926 );
buf \U$6258 ( \6928 , \6898 );
buf \U$6259 ( \6929 , \6928 );
not \U$6260 ( \6930 , \6929 );
nor \U$6261 ( \6931 , \6895 , \6927 , \6930 );
and \U$6262 ( \6932 , \6854 , RIaa9f948_280);
and \U$6263 ( \6933 , \6856 , RIaa9f9c0_281);
nor \U$6264 ( \6934 , \6932 , \6933 );
not \U$6265 ( \6935 , \2026 );
not \U$6266 ( \6936 , \1416 );
and \U$6267 ( \6937 , \6935 , \6936 );
not \U$6268 ( \6938 , \1843 );
not \U$6269 ( \6939 , \6938 );
and \U$6270 ( \6940 , \6939 , RIaa9f8d0_279);
nor \U$6271 ( \6941 , \6937 , \6940 );
and \U$6272 ( \6942 , \1872 , RIaa9f330_267);
nor \U$6273 ( \6943 , \6942 , \1496 );
and \U$6274 ( \6944 , \1626 , RIaa9f3a8_268);
not \U$6275 ( \6945 , RIaa9f588_272);
not \U$6276 ( \6946 , \6871 );
or \U$6277 ( \6947 , \6945 , \6946 );
not \U$6278 ( \6948 , RIaa9f600_273);
or \U$6279 ( \6949 , \6867 , \6948 );
nand \U$6280 ( \6950 , \6947 , \6949 );
nor \U$6281 ( \6951 , \6944 , \6950 );
and \U$6282 ( \6952 , \6934 , \6941 , \6943 , \6951 );
and \U$6283 ( \6953 , \1832 , RIaa9f768_276);
and \U$6284 ( \6954 , \1642 , RIaa9f7e0_277);
nor \U$6285 ( \6955 , \6953 , \6954 );
and \U$6286 ( \6956 , \1861 , RIaa9f2b8_266);
and \U$6287 ( \6957 , \6883 , RIaa9f858_278);
nor \U$6288 ( \6958 , \6956 , \6957 );
nand \U$6289 ( \6959 , \6955 , \6958 );
not \U$6290 ( \6960 , \2063 );
not \U$6291 ( \6961 , RIaa9f678_274);
not \U$6292 ( \6962 , \6961 );
and \U$6293 ( \6963 , \6960 , \6962 );
and \U$6294 ( \6964 , \6862 , RIaa9f510_271);
nor \U$6295 ( \6965 , \6963 , \6964 );
not \U$6296 ( \6966 , \2052 );
not \U$6297 ( \6967 , RIaa9f420_269);
not \U$6298 ( \6968 , \6967 );
and \U$6299 ( \6969 , \6966 , \6968 );
and \U$6300 ( \6970 , \1755 , RIaa9f498_270);
nor \U$6301 ( \6971 , \6969 , \6970 );
nand \U$6302 ( \6972 , \6965 , \6971 );
nor \U$6303 ( \6973 , \6959 , \6972 );
and \U$6304 ( \6974 , \6952 , \6973 );
buf \U$6305 ( \6975 , \6974 );
not \U$6306 ( \6976 , \6975 );
buf \U$6307 ( \6977 , \6976 );
not \U$6308 ( \6978 , \6977 );
nor \U$6309 ( \6979 , \6846 , \6978 );
or \U$6310 ( \6980 , \6931 , \6979 );
nand \U$6311 ( \6981 , \6931 , \6979 );
nand \U$6312 ( \6982 , \6980 , \6981 );
not \U$6313 ( \6983 , \6982 );
not \U$6314 ( \6984 , \6928 );
nor \U$6315 ( \6985 , \6984 , \6920 );
buf \U$6316 ( \6986 , \6985 );
not \U$6317 ( \6987 , \6986 );
or \U$6318 ( \6988 , \6987 , \6894 );
not \U$6319 ( \6989 , \6928 );
and \U$6320 ( \6990 , \6921 , \6989 );
nand \U$6321 ( \6991 , \6990 , \6894 );
nand \U$6322 ( \6992 , \6928 , \6924 );
buf \U$6323 ( \6993 , \6992 );
nand \U$6324 ( \6994 , \6988 , \6991 , \6993 );
not \U$6325 ( \6995 , \6979 );
and \U$6326 ( \6996 , \6994 , \6995 );
not \U$6327 ( \6997 , \2026 );
not \U$6328 ( \6998 , RIaa9ffd8_294);
not \U$6329 ( \6999 , \6998 );
and \U$6330 ( \7000 , \6997 , \6999 );
and \U$6331 ( \7001 , \1755 , RIaaa00c8_296);
nor \U$6332 ( \7002 , \7000 , \7001 );
not \U$6333 ( \7003 , \1874 );
not \U$6334 ( \7004 , \7003 );
not \U$6335 ( \7005 , RIaa9fd08_288);
not \U$6336 ( \7006 , \7005 );
and \U$6337 ( \7007 , \7004 , \7006 );
and \U$6338 ( \7008 , \1846 , RIaa9fdf8_290);
nor \U$6339 ( \7009 , \7007 , \7008 );
nand \U$6340 ( \7010 , \7002 , \7009 );
nand \U$6341 ( \7011 , \1832 , RIaa9fe70_291);
nand \U$6342 ( \7012 , \1642 , RIaa9fee8_292);
not \U$6343 ( \7013 , \1622 );
not \U$6344 ( \7014 , \7013 );
nand \U$6345 ( \7015 , \7014 , RIaa9fd80_289);
nand \U$6346 ( \7016 , \7011 , \7012 , \7015 );
nor \U$6347 ( \7017 , \7010 , \7016 );
not \U$6348 ( \7018 , RIaa9ff60_293);
not \U$6349 ( \7019 , \2064 );
or \U$6350 ( \7020 , \7018 , \7019 );
nand \U$6351 ( \7021 , \7020 , \2264 );
nand \U$6352 ( \7022 , \6883 , RIaa9fa38_282);
not \U$6353 ( \7023 , \1316 );
not \U$6354 ( \7024 , \7023 );
nand \U$6355 ( \7025 , \7024 , RIaaa0140_297);
and \U$6356 ( \7026 , \6868 , RIaa9fc90_287);
and \U$6357 ( \7027 , \6871 , RIaa9fc18_286);
nor \U$6358 ( \7028 , \7026 , \7027 );
nand \U$6359 ( \7029 , \7022 , \7025 , \7028 );
nor \U$6360 ( \7030 , \7021 , \7029 );
and \U$6361 ( \7031 , \2023 , RIaaa0050_295);
and \U$6362 ( \7032 , \6939 , RIaa9fab0_283);
nor \U$6363 ( \7033 , \7031 , \7032 );
and \U$6364 ( \7034 , \6862 , RIaa9fba0_285);
and \U$6365 ( \7035 , \1861 , RIaaa01b8_298);
nor \U$6366 ( \7036 , \7034 , \7035 );
and \U$6367 ( \7037 , \7017 , \7030 , \7033 , \7036 );
buf \U$6368 ( \7038 , \7037 );
not \U$6369 ( \7039 , \7038 );
nand \U$6370 ( \7040 , \6847 , \7039 );
not \U$6371 ( \7041 , \6829 );
and \U$6372 ( \7042 , \6831 , \6834 );
not \U$6373 ( \7043 , \7042 );
and \U$6374 ( \7044 , \7041 , \7043 );
and \U$6375 ( \7045 , \6829 , \7042 );
nor \U$6376 ( \7046 , \7044 , \7045 );
or \U$6377 ( \7047 , \6914 , \7046 );
buf \U$6378 ( \7048 , \7046 );
nand \U$6379 ( \7049 , \6914 , \7048 );
not \U$6380 ( \7050 , \6826 );
nand \U$6381 ( \7051 , \7050 , \6828 );
not \U$6382 ( \7052 , \7051 );
buf \U$6383 ( \7053 , \6825 );
not \U$6384 ( \7054 , \7053 );
or \U$6385 ( \7055 , \7052 , \7054 );
or \U$6386 ( \7056 , \7053 , \7051 );
nand \U$6387 ( \7057 , \7055 , \7056 );
not \U$6388 ( \7058 , \7057 );
not \U$6389 ( \7059 , \7058 );
not \U$6390 ( \7060 , \7046 );
or \U$6391 ( \7061 , \7059 , \7060 );
or \U$6392 ( \7062 , \7058 , \7046 );
nand \U$6393 ( \7063 , \7061 , \7062 );
and \U$6394 ( \7064 , \7047 , \7049 , \7063 );
buf \U$6395 ( \7065 , \7064 );
not \U$6396 ( \7066 , \6915 );
nand \U$6397 ( \7067 , \7065 , \7066 );
not \U$6398 ( \7068 , \7063 );
nand \U$6399 ( \7069 , \7068 , \6916 );
not \U$6400 ( \7070 , \7069 );
not \U$6401 ( \7071 , \7070 );
and \U$6402 ( \7072 , \7040 , \7067 , \7071 );
not \U$6403 ( \7073 , \7072 );
not \U$6404 ( \7074 , \6977 );
not \U$6405 ( \7075 , \6990 );
or \U$6406 ( \7076 , \7074 , \7075 );
and \U$6407 ( \7077 , \6986 , \6978 );
not \U$6408 ( \7078 , \6928 );
nand \U$6409 ( \7079 , \7078 , \6924 );
buf \U$6410 ( \7080 , \7079 );
not \U$6411 ( \7081 , \7080 );
and \U$6412 ( \7082 , \7081 , \6894 );
not \U$6413 ( \7083 , \6993 );
not \U$6414 ( \7084 , \6894 );
and \U$6415 ( \7085 , \7083 , \7084 );
nor \U$6416 ( \7086 , \7077 , \7082 , \7085 );
nand \U$6417 ( \7087 , \7076 , \7086 );
not \U$6418 ( \7088 , \7087 );
or \U$6419 ( \7089 , \7073 , \7088 );
nand \U$6420 ( \7090 , \7089 , \7040 );
or \U$6421 ( \7091 , \6994 , \6979 );
nand \U$6422 ( \7092 , \7091 , \6981 );
and \U$6423 ( \7093 , \7090 , \7092 );
nor \U$6424 ( \7094 , \6996 , \7093 );
not \U$6425 ( \7095 , \7094 );
or \U$6426 ( \7096 , \6983 , \7095 );
or \U$6427 ( \7097 , \7094 , \6982 );
nand \U$6428 ( \7098 , \7096 , \7097 );
not \U$6429 ( \7099 , \7098 );
not \U$6430 ( \7100 , \7039 );
and \U$6431 ( \7101 , \7064 , \6915 );
buf \U$6432 ( \7102 , \7101 );
not \U$6433 ( \7103 , \7102 );
or \U$6434 ( \7104 , \7100 , \7103 );
not \U$6435 ( \7105 , \7063 );
nand \U$6436 ( \7106 , \7105 , \6915 );
not \U$6437 ( \7107 , \7106 );
and \U$6438 ( \7108 , \6976 , \7107 );
not \U$6439 ( \7109 , \6976 );
and \U$6440 ( \7110 , \7109 , \7070 );
nor \U$6441 ( \7111 , \7108 , \7110 );
nand \U$6442 ( \7112 , \7104 , \7111 );
nor \U$6443 ( \7113 , \7067 , \7039 );
or \U$6444 ( \7114 , \7112 , \7113 );
not \U$6445 ( \7115 , \7114 );
buf \U$6446 ( \7116 , \6805 );
not \U$6447 ( \7117 , \7116 );
not \U$6448 ( \7118 , \6807 );
not \U$6449 ( \7119 , \6806 );
not \U$6450 ( \7120 , \6811 );
nand \U$6451 ( \7121 , \6803 , \7120 );
not \U$6452 ( \7122 , \7121 );
or \U$6453 ( \7123 , \7119 , \7122 );
buf \U$6454 ( \7124 , \6813 );
not \U$6455 ( \7125 , \7124 );
nand \U$6456 ( \7126 , \7123 , \7125 );
not \U$6457 ( \7127 , \7126 );
or \U$6458 ( \7128 , \7118 , \7127 );
not \U$6459 ( \7129 , \6815 );
nand \U$6460 ( \7130 , \7128 , \7129 );
not \U$6461 ( \7131 , \7130 );
or \U$6462 ( \7132 , \7117 , \7131 );
not \U$6463 ( \7133 , \6819 );
nand \U$6464 ( \7134 , \7132 , \7133 );
not \U$6465 ( \7135 , \6821 );
nand \U$6466 ( \7136 , \7135 , \6804 );
and \U$6467 ( \7137 , \7134 , \7136 );
not \U$6468 ( \7138 , \7134 );
not \U$6469 ( \7139 , \7136 );
and \U$6470 ( \7140 , \7138 , \7139 );
nor \U$6471 ( \7141 , \7137 , \7140 );
not \U$6472 ( \7142 , \7141 );
nand \U$6473 ( \7143 , \7133 , \7116 );
not \U$6474 ( \7144 , \7143 );
not \U$6475 ( \7145 , \7130 );
or \U$6476 ( \7146 , \7144 , \7145 );
not \U$6477 ( \7147 , \7143 );
not \U$6478 ( \7148 , \7130 );
nand \U$6479 ( \7149 , \7147 , \7148 );
nand \U$6480 ( \7150 , \7146 , \7149 );
nand \U$6481 ( \7151 , \7142 , \7150 );
buf \U$6482 ( \7152 , \7058 );
not \U$6483 ( \7153 , \7152 );
nor \U$6484 ( \7154 , \7151 , \7153 );
buf \U$6485 ( \7155 , \7154 );
and \U$6486 ( \7156 , \7155 , \6894 );
not \U$6487 ( \7157 , \7058 );
buf \U$6488 ( \7158 , \7141 );
xnor \U$6489 ( \7159 , \7148 , \7143 );
nand \U$6490 ( \7160 , \7157 , \7158 , \7159 );
not \U$6491 ( \7161 , \7160 );
and \U$6492 ( \7162 , \7161 , \7084 );
not \U$6493 ( \7163 , \2014 );
not \U$6494 ( \7164 , RIaaa1dd8_358);
not \U$6495 ( \7165 , \7164 );
and \U$6496 ( \7166 , \7163 , \7165 );
and \U$6497 ( \7167 , \1626 , RIaaa1ce8_356);
nor \U$6498 ( \7168 , \7166 , \7167 );
nand \U$6499 ( \7169 , \2061 , RIaaa1c70_355);
nand \U$6500 ( \7170 , \7168 , \1932 , \7169 );
and \U$6501 ( \7171 , \1846 , RIaaa1d60_357);
and \U$6502 ( \7172 , \1861 , RIaaa1bf8_354);
nor \U$6503 ( \7173 , \7171 , \7172 );
not \U$6504 ( \7174 , \1852 );
and \U$6505 ( \7175 , \7174 , RIaaa1a90_351);
and \U$6506 ( \7176 , RIaaa1b80_353, \6868 );
and \U$6507 ( \7177 , \6871 , RIaaa1b08_352);
nor \U$6508 ( \7178 , \7175 , \7176 , \7177 );
nand \U$6509 ( \7179 , \7173 , \7178 );
nor \U$6510 ( \7180 , \7170 , \7179 );
not \U$6511 ( \7181 , RIaaa1e50_359);
nor \U$6512 ( \7182 , \2063 , \7181 );
not \U$6513 ( \7183 , \7182 );
not \U$6514 ( \7184 , \1842 );
not \U$6515 ( \7185 , \7184 );
not \U$6516 ( \7186 , \7185 );
nand \U$6517 ( \7187 , \7186 , RIaaa2198_366);
and \U$6518 ( \7188 , \6856 , RIaaa1fb8_362);
not \U$6519 ( \7189 , RIaaa1f40_361);
nor \U$6520 ( \7190 , \7189 , \2068 );
nor \U$6521 ( \7191 , \7188 , \7190 );
nand \U$6522 ( \7192 , \7183 , \7187 , \7191 );
and \U$6523 ( \7193 , \1832 , RIaaa2030_363);
and \U$6524 ( \7194 , \1642 , RIaaa20a8_364);
nor \U$6525 ( \7195 , \7193 , \7194 );
not \U$6526 ( \7196 , \6882 );
not \U$6527 ( \7197 , RIaaa2120_365);
not \U$6528 ( \7198 , \7197 );
and \U$6529 ( \7199 , \7196 , \7198 );
and \U$6530 ( \7200 , \1651 , RIaaa1ec8_360);
nor \U$6531 ( \7201 , \7199 , \7200 );
nand \U$6532 ( \7202 , \7195 , \7201 );
nor \U$6533 ( \7203 , \7192 , \7202 );
nand \U$6534 ( \7204 , \7180 , \7203 );
not \U$6535 ( \7205 , \7204 );
buf \U$6536 ( \7206 , \7205 );
not \U$6537 ( \7207 , \7206 );
and \U$6538 ( \7208 , \6847 , \7207 );
nor \U$6539 ( \7209 , \7156 , \7162 , \7208 );
not \U$6540 ( \7210 , \7142 );
not \U$6541 ( \7211 , \7159 );
or \U$6542 ( \7212 , \7210 , \7211 );
nand \U$6543 ( \7213 , \7141 , \7150 );
nand \U$6544 ( \7214 , \7212 , \7213 );
nand \U$6545 ( \7215 , \7214 , \7153 );
buf \U$6546 ( \7216 , \7215 );
nand \U$6547 ( \7217 , \7209 , \7216 );
nand \U$6548 ( \7218 , \7115 , \7217 );
not \U$6549 ( \7219 , \7218 );
not \U$6550 ( \7220 , \2026 );
not \U$6551 ( \7221 , RIaaa05f0_307);
not \U$6552 ( \7222 , \7221 );
and \U$6553 ( \7223 , \7220 , \7222 );
not \U$6554 ( \7224 , RIaaa0488_304);
nor \U$6555 ( \7225 , \7224 , \1838 );
nor \U$6556 ( \7226 , \7223 , \7225 );
not \U$6557 ( \7227 , RIaaa08c0_313);
nor \U$6558 ( \7228 , \7227 , \6938 );
not \U$6559 ( \7229 , RIaaa06e0_309);
nor \U$6560 ( \7230 , \7229 , \2036 );
nor \U$6561 ( \7231 , \7228 , \7230 );
nand \U$6562 ( \7232 , \7226 , \7231 );
not \U$6563 ( \7233 , RIaaa0668_308);
not \U$6564 ( \7234 , \2061 );
or \U$6565 ( \7235 , \7233 , \7234 );
and \U$6566 ( \7236 , \1640 , RIaaa0938_314);
not \U$6567 ( \7237 , RIaaa07d0_311);
not \U$6568 ( \7238 , \6871 );
or \U$6569 ( \7239 , \7237 , \7238 );
not \U$6570 ( \7240 , RIaaa0848_312);
or \U$6571 ( \7241 , \6867 , \7240 );
nand \U$6572 ( \7242 , \7239 , \7241 );
nor \U$6573 ( \7243 , \7236 , \7242 );
nand \U$6574 ( \7244 , \7235 , \7243 );
nor \U$6575 ( \7245 , \7232 , \7244 );
not \U$6576 ( \7246 , \6862 );
not \U$6577 ( \7247 , \7246 );
not \U$6578 ( \7248 , RIaaa0758_310);
not \U$6579 ( \7249 , \7248 );
and \U$6580 ( \7250 , \7247 , \7249 );
not \U$6581 ( \7251 , RIaaa0500_305);
nor \U$6582 ( \7252 , \7251 , \2014 );
nor \U$6583 ( \7253 , \7250 , \7252 );
nand \U$6584 ( \7254 , \2064 , RIaaa0578_306);
and \U$6585 ( \7255 , \7253 , \2354 , \7254 );
and \U$6586 ( \7256 , \6854 , RIaaa0320_301);
and \U$6587 ( \7257 , RIaaa0230_299, \1832 );
and \U$6588 ( \7258 , \1642 , RIaaa02a8_300);
nor \U$6589 ( \7259 , \7256 , \7257 , \7258 );
and \U$6590 ( \7260 , \1846 , RIaaa0410_303);
and \U$6591 ( \7261 , \2066 , RIaaa0398_302);
nor \U$6592 ( \7262 , \7260 , \7261 );
and \U$6593 ( \7263 , \7245 , \7255 , \7259 , \7262 );
not \U$6594 ( \7264 , \7263 );
buf \U$6595 ( \7265 , \7264 );
not \U$6596 ( \7266 , \7265 );
not \U$6597 ( \7267 , \6990 );
or \U$6598 ( \7268 , \7266 , \7267 );
not \U$6599 ( \7269 , \7265 );
and \U$6600 ( \7270 , \6986 , \7269 );
and \U$6601 ( \7271 , \7039 , \7080 );
not \U$6602 ( \7272 , \7039 );
and \U$6603 ( \7273 , \7272 , \6993 );
nor \U$6604 ( \7274 , \7271 , \7273 );
nor \U$6605 ( \7275 , \7270 , \7274 );
nand \U$6606 ( \7276 , \7268 , \7275 );
and \U$6607 ( \7277 , \1832 , RIaaa0cf8_322);
and \U$6608 ( \7278 , \1642 , RIaaa0d70_323);
nor \U$6609 ( \7279 , \7277 , \7278 );
and \U$6610 ( \7280 , \1872 , RIaaa0c08_320);
and \U$6611 ( \7281 , \1874 , RIaaa0de8_324);
nor \U$6612 ( \7282 , \7280 , \7281 );
nand \U$6613 ( \7283 , \2066 , RIaaa0e60_325);
nand \U$6614 ( \7284 , \7279 , \7282 , \7283 );
and \U$6615 ( \7285 , \6862 , RIaaa0f50_327);
and \U$6616 ( \7286 , \1861 , RIaaa0c80_321);
nor \U$6617 ( \7287 , \7285 , \7286 );
and \U$6618 ( \7288 , \1846 , RIaaa0ed8_326);
and \U$6619 ( \7289 , \2064 , RIaaa0b18_318);
nor \U$6620 ( \7290 , \7288 , \7289 );
nand \U$6621 ( \7291 , \7287 , \7290 );
nor \U$6622 ( \7292 , \7284 , \7291 );
and \U$6623 ( \7293 , \6889 , RIaaa0aa0_317);
and \U$6624 ( \7294 , \6876 , RIaaa10b8_330);
nor \U$6625 ( \7295 , \7293 , \7294 );
or \U$6626 ( \7296 , \1745 , \1946 );
and \U$6627 ( \7297 , \6868 , RIaaa1040_329);
and \U$6628 ( \7298 , \6871 , RIaaa0fc8_328);
nor \U$6629 ( \7299 , \7297 , \7298 );
nand \U$6630 ( \7300 , \7296 , \7299 );
nor \U$6631 ( \7301 , \7300 , \1975 );
and \U$6632 ( \7302 , \1626 , RIaaa0a28_316);
and \U$6633 ( \7303 , \1651 , RIaaa0b90_319);
nor \U$6634 ( \7304 , \7302 , \7303 );
and \U$6635 ( \7305 , \7295 , \7301 , \7304 );
nand \U$6636 ( \7306 , \7292 , \7305 );
not \U$6637 ( \7307 , \7306 );
buf \U$6638 ( \7308 , \7307 );
not \U$6639 ( \7309 , \7308 );
nand \U$6640 ( \7310 , \6847 , \7309 );
xor \U$6641 ( \7311 , \7276 , \7310 );
not \U$6642 ( \7312 , \7311 );
not \U$6643 ( \7313 , \7312 );
or \U$6644 ( \7314 , \7219 , \7313 );
not \U$6645 ( \7315 , \7218 );
nand \U$6646 ( \7316 , \7315 , \7311 );
nand \U$6647 ( \7317 , \7314 , \7316 );
not \U$6648 ( \7318 , \7317 );
and \U$6649 ( \7319 , \6930 , \7269 );
and \U$6650 ( \7320 , \6929 , \7265 );
nor \U$6651 ( \7321 , \7319 , \7320 );
or \U$6652 ( \7322 , \7321 , \6922 );
and \U$6653 ( \7323 , \7309 , \6930 );
not \U$6654 ( \7324 , \7309 );
and \U$6655 ( \7325 , \7324 , \6929 );
or \U$6656 ( \7326 , \7323 , \7325 );
or \U$6657 ( \7327 , \7326 , \6925 );
nor \U$6658 ( \7328 , \7309 , \7265 );
and \U$6659 ( \7329 , \7328 , \6930 );
nor \U$6660 ( \7330 , \7269 , \7308 );
and \U$6661 ( \7331 , \6929 , \7330 );
nor \U$6662 ( \7332 , \7329 , \7331 );
nand \U$6663 ( \7333 , \7322 , \7327 , \7332 );
nor \U$6664 ( \7334 , \7333 , \6927 );
not \U$6665 ( \7335 , \6894 );
and \U$6666 ( \7336 , \7214 , \7152 );
not \U$6667 ( \7337 , \7336 );
not \U$6668 ( \7338 , \7337 );
not \U$6669 ( \7339 , \7338 );
or \U$6670 ( \7340 , \7335 , \7339 );
not \U$6671 ( \7341 , \7161 );
not \U$6672 ( \7342 , \7341 );
not \U$6673 ( \7343 , \6977 );
and \U$6674 ( \7344 , \7342 , \7343 );
and \U$6675 ( \7345 , \7155 , \6977 );
nor \U$6676 ( \7346 , \7344 , \7345 );
nand \U$6677 ( \7347 , \7340 , \7346 );
nor \U$6678 ( \7348 , \7216 , \6894 );
nor \U$6679 ( \7349 , \7347 , \7348 );
buf \U$6680 ( \7350 , \7121 );
not \U$6681 ( \7351 , \7124 );
nand \U$6682 ( \7352 , \7351 , \6806 );
not \U$6683 ( \7353 , \7352 );
and \U$6684 ( \7354 , \7350 , \7353 );
not \U$6685 ( \7355 , \7350 );
and \U$6686 ( \7356 , \7355 , \7352 );
nor \U$6687 ( \7357 , \7354 , \7356 );
not \U$6688 ( \7358 , \7357 );
nand \U$6689 ( \7359 , \7129 , \6807 );
xnor \U$6690 ( \7360 , \7126 , \7359 );
not \U$6691 ( \7361 , \7360 );
not \U$6692 ( \7362 , \7361 );
or \U$6693 ( \7363 , \7358 , \7362 );
not \U$6694 ( \7364 , \7350 );
not \U$6695 ( \7365 , \7352 );
and \U$6696 ( \7366 , \7364 , \7365 );
and \U$6697 ( \7367 , \7350 , \7352 );
nor \U$6698 ( \7368 , \7366 , \7367 );
nand \U$6699 ( \7369 , \7360 , \7368 );
nand \U$6700 ( \7370 , \7363 , \7369 );
not \U$6701 ( \7371 , \7370 );
nand \U$6702 ( \7372 , \7371 , \7150 );
not \U$6703 ( \7373 , \7372 );
buf \U$6704 ( \7374 , \7360 );
not \U$6705 ( \7375 , \7374 );
nand \U$6706 ( \7376 , \7373 , \7375 );
nand \U$6707 ( \7377 , \7370 , \7150 );
buf \U$6708 ( \7378 , \7377 );
and \U$6709 ( \7379 , \7376 , \7378 );
and \U$6710 ( \7380 , \7102 , \7265 );
not \U$6711 ( \7381 , \7038 );
not \U$6712 ( \7382 , \7070 );
or \U$6713 ( \7383 , \7381 , \7382 );
nand \U$6714 ( \7384 , \7107 , \7039 );
nand \U$6715 ( \7385 , \7383 , \7384 );
nor \U$6716 ( \7386 , \7380 , \7385 );
not \U$6717 ( \7387 , \7064 );
nor \U$6718 ( \7388 , \7387 , \6915 );
buf \U$6719 ( \7389 , \7388 );
nand \U$6720 ( \7390 , \7389 , \7269 );
nand \U$6721 ( \7391 , \7386 , \7390 );
nor \U$6722 ( \7392 , \7379 , \7391 );
or \U$6723 ( \7393 , \7349 , \7392 );
nand \U$6724 ( \7394 , \7391 , \7379 );
nand \U$6725 ( \7395 , \7393 , \7394 );
xor \U$6726 ( \7396 , \7334 , \7395 );
not \U$6727 ( \7397 , \6927 );
and \U$6728 ( \7398 , \6929 , \7206 );
not \U$6729 ( \7399 , \6929 );
and \U$6730 ( \7400 , \7399 , \7207 );
or \U$6731 ( \7401 , \7398 , \7400 );
not \U$6732 ( \7402 , \7401 );
not \U$6733 ( \7403 , \6925 );
and \U$6734 ( \7404 , \7402 , \7403 );
nor \U$6735 ( \7405 , \7326 , \6922 );
nor \U$6736 ( \7406 , \7404 , \7405 );
nand \U$6737 ( \7407 , \7397 , \7406 );
not \U$6738 ( \7408 , \6846 );
not \U$6739 ( \7409 , \2066 );
not \U$6740 ( \7410 , \7409 );
not \U$6741 ( \7411 , RIaaa17c0_345);
not \U$6742 ( \7412 , \7411 );
and \U$6743 ( \7413 , \7410 , \7412 );
not \U$6744 ( \7414 , RIaaa1748_344);
not \U$6745 ( \7415 , \1874 );
nor \U$6746 ( \7416 , \7414 , \7415 );
nor \U$6747 ( \7417 , \7413 , \7416 );
not \U$6748 ( \7418 , RIaaa1478_338);
nor \U$6749 ( \7419 , \7418 , \7023 );
nor \U$6750 ( \7420 , \2191 , \7419 );
not \U$6751 ( \7421 , \2063 );
not \U$6752 ( \7422 , RIaaa1658_342);
not \U$6753 ( \7423 , \7422 );
and \U$6754 ( \7424 , \7421 , \7423 );
and \U$6755 ( \7425 , \1651 , RIaaa16d0_343);
nor \U$6756 ( \7426 , \7424 , \7425 );
not \U$6757 ( \7427 , \1852 );
not \U$6758 ( \7428 , RIaaa1298_334);
not \U$6759 ( \7429 , \7428 );
and \U$6760 ( \7430 , \7427 , \7429 );
not \U$6761 ( \7431 , RIaaa1568_340);
not \U$6762 ( \7432 , \1846 );
nor \U$6763 ( \7433 , \7431 , \7432 );
nor \U$6764 ( \7434 , \7430 , \7433 );
nand \U$6765 ( \7435 , \7417 , \7420 , \7426 , \7434 );
and \U$6766 ( \7436 , RIaaa1838_346, \1832 );
not \U$6767 ( \7437 , RIaaa18b0_347);
nor \U$6768 ( \7438 , \7437 , \1743 );
nor \U$6769 ( \7439 , \7436 , \7438 );
not \U$6770 ( \7440 , \1842 );
not \U$6771 ( \7441 , \7440 );
not \U$6772 ( \7442 , \7441 );
not \U$6773 ( \7443 , \2181 );
and \U$6774 ( \7444 , \7442 , \7443 );
and \U$6775 ( \7445 , \1640 , RIaaa1928_348);
nor \U$6776 ( \7446 , \7444 , \7445 );
not \U$6777 ( \7447 , \2036 );
not \U$6778 ( \7448 , RIaaa1400_337);
not \U$6779 ( \7449 , \7448 );
and \U$6780 ( \7450 , \7447 , \7449 );
and \U$6781 ( \7451 , \2023 , RIaaa14f0_339);
nor \U$6782 ( \7452 , \7450 , \7451 );
not \U$6783 ( \7453 , \6888 );
not \U$6784 ( \7454 , RIaaa15e0_341);
not \U$6785 ( \7455 , \7454 );
and \U$6786 ( \7456 , \7453 , \7455 );
not \U$6787 ( \7457 , RIaaa1388_336);
not \U$6788 ( \7458 , \6868 );
or \U$6789 ( \7459 , \7457 , \7458 );
nand \U$6790 ( \7460 , \6871 , RIaaa1310_335);
nand \U$6791 ( \7461 , \7459 , \7460 );
nor \U$6792 ( \7462 , \7456 , \7461 );
nand \U$6793 ( \7463 , \7439 , \7446 , \7452 , \7462 );
nor \U$6794 ( \7464 , \7435 , \7463 );
buf \U$6795 ( \7465 , \7464 );
buf \U$6796 ( \7466 , \7465 );
not \U$6797 ( \7467 , \7466 );
and \U$6798 ( \7468 , \7408 , \7467 );
and \U$6799 ( \7469 , \7102 , \7309 );
or \U$6800 ( \7470 , \7071 , \7265 );
not \U$6801 ( \7471 , \7107 );
not \U$6802 ( \7472 , \7471 );
nand \U$6803 ( \7473 , \7472 , \7265 );
nand \U$6804 ( \7474 , \7470 , \7473 );
nor \U$6805 ( \7475 , \7469 , \7474 );
nand \U$6806 ( \7476 , \7389 , \7308 );
nand \U$6807 ( \7477 , \7475 , \7476 );
nor \U$6808 ( \7478 , \7468 , \7477 );
nor \U$6809 ( \7479 , \7407 , \7478 );
and \U$6810 ( \7480 , \7396 , \7479 );
and \U$6811 ( \7481 , \7334 , \7395 );
or \U$6812 ( \7482 , \7480 , \7481 );
not \U$6813 ( \7483 , \6978 );
not \U$6814 ( \7484 , \7389 );
or \U$6815 ( \7485 , \7483 , \7484 );
and \U$6816 ( \7486 , \7102 , \6977 );
and \U$6817 ( \7487 , \7107 , \6894 );
and \U$6818 ( \7488 , \7070 , \7084 );
nor \U$6819 ( \7489 , \7486 , \7487 , \7488 );
nand \U$6820 ( \7490 , \7485 , \7489 );
and \U$6821 ( \7491 , \7490 , \7114 );
not \U$6822 ( \7492 , \7490 );
and \U$6823 ( \7493 , \7492 , \7115 );
nor \U$6824 ( \7494 , \7491 , \7493 );
not \U$6825 ( \7495 , \7151 );
not \U$6826 ( \7496 , \7495 );
nand \U$6827 ( \7497 , \7496 , \7153 );
xor \U$6828 ( \7498 , \7494 , \7497 );
or \U$6829 ( \7499 , \7482 , \7498 );
not \U$6830 ( \7500 , \7499 );
or \U$6831 ( \7501 , \7318 , \7500 );
nand \U$6832 ( \7502 , \7482 , \7498 );
nand \U$6833 ( \7503 , \7501 , \7502 );
not \U$6834 ( \7504 , \7503 );
not \U$6835 ( \7505 , \7218 );
nand \U$6836 ( \7506 , \7505 , \7312 );
not \U$6837 ( \7507 , \7310 );
nand \U$6838 ( \7508 , \7507 , \7276 );
and \U$6839 ( \7509 , \7506 , \7508 );
and \U$6840 ( \7510 , \7494 , \7497 );
and \U$6841 ( \7511 , \7490 , \7114 );
nor \U$6842 ( \7512 , \7510 , \7511 );
xor \U$6843 ( \7513 , \7509 , \7512 );
or \U$6844 ( \7514 , \7067 , \6894 );
and \U$6845 ( \7515 , \7102 , \6894 );
or \U$6846 ( \7516 , \6846 , \7269 );
nand \U$6847 ( \7517 , \7516 , \7071 );
nor \U$6848 ( \7518 , \7515 , \7517 );
nand \U$6849 ( \7519 , \7514 , \7518 );
not \U$6850 ( \7520 , \7519 );
not \U$6851 ( \7521 , \7039 );
not \U$6852 ( \7522 , \6990 );
or \U$6853 ( \7523 , \7521 , \7522 );
and \U$6854 ( \7524 , \6986 , \7038 );
or \U$6855 ( \7525 , \7080 , \6978 );
or \U$6856 ( \7526 , \6993 , \6977 );
nand \U$6857 ( \7527 , \7525 , \7526 );
nor \U$6858 ( \7528 , \7524 , \7527 );
nand \U$6859 ( \7529 , \7523 , \7528 );
not \U$6860 ( \7530 , \7529 );
or \U$6861 ( \7531 , \7520 , \7530 );
or \U$6862 ( \7532 , \7529 , \7519 );
nand \U$6863 ( \7533 , \7531 , \7532 );
not \U$6864 ( \7534 , \7533 );
xor \U$6865 ( \7535 , \7513 , \7534 );
nand \U$6866 ( \7536 , \7504 , \7535 );
nand \U$6867 ( \7537 , \6367 , \853 );
nand \U$6868 ( \7538 , \6785 , \7537 );
buf \U$6869 ( \7539 , \6799 );
xnor \U$6870 ( \7540 , \7538 , \7539 );
not \U$6871 ( \7541 , \7539 );
not \U$6872 ( \7542 , \7541 );
not \U$6873 ( \7543 , \7538 );
or \U$6874 ( \7544 , \7542 , \7543 );
nand \U$6875 ( \7545 , \7544 , \6794 );
not \U$6876 ( \7546 , \6801 );
nand \U$6877 ( \7547 , \7546 , \7120 );
not \U$6878 ( \7548 , \7547 );
and \U$6879 ( \7549 , \7545 , \7548 );
not \U$6880 ( \7550 , \7545 );
and \U$6881 ( \7551 , \7550 , \7547 );
nor \U$6882 ( \7552 , \7549 , \7551 );
xnor \U$6883 ( \7553 , \7540 , \7552 );
buf \U$6884 ( \7554 , \7553 );
not \U$6885 ( \7555 , \7554 );
not \U$6886 ( \7556 , \7357 );
not \U$6887 ( \7557 , \7556 );
nand \U$6888 ( \7558 , \7555 , \7557 );
buf \U$6889 ( \7559 , \7558 );
buf \U$6890 ( \7560 , \7554 );
buf \U$6891 ( \7561 , \7552 );
nand \U$6892 ( \7562 , \7561 , \7357 );
not \U$6893 ( \7563 , \7561 );
nand \U$6894 ( \7564 , \7563 , \7368 );
nand \U$6895 ( \7565 , \7560 , \7562 , \7564 );
nand \U$6896 ( \7566 , \7559 , \7565 );
and \U$6897 ( \7567 , \6893 , \7560 , \7557 );
not \U$6898 ( \7568 , \6893 );
not \U$6899 ( \7569 , \7368 );
not \U$6900 ( \7570 , \7569 );
and \U$6901 ( \7571 , \7568 , \7570 );
nor \U$6902 ( \7572 , \7567 , \7571 );
and \U$6903 ( \7573 , \7566 , \7572 );
not \U$6904 ( \7574 , \7573 );
not \U$6905 ( \7575 , \7574 );
and \U$6906 ( \7576 , \7554 , \7562 , \7564 , \7557 );
buf \U$6907 ( \7577 , \7576 );
not \U$6908 ( \7578 , \7577 );
nand \U$6909 ( \7579 , \7578 , \7559 );
not \U$6910 ( \7580 , \7579 );
or \U$6911 ( \7581 , \7575 , \7580 );
xor \U$6912 ( \7582 , \7579 , \7573 );
not \U$6913 ( \7583 , \7582 );
not \U$6914 ( \7584 , \7066 );
not \U$6915 ( \7585 , \7308 );
not \U$6916 ( \7586 , \7585 );
and \U$6917 ( \7587 , \7584 , \7586 );
and \U$6918 ( \7588 , \7066 , \7309 );
nor \U$6919 ( \7589 , \7587 , \7588 );
or \U$6920 ( \7590 , \7589 , \7065 );
xnor \U$6921 ( \7591 , \7206 , \7066 );
not \U$6922 ( \7592 , \7591 );
not \U$6923 ( \7593 , \7065 );
or \U$6924 ( \7594 , \7592 , \7593 );
nand \U$6925 ( \7595 , \7594 , \7063 );
nand \U$6926 ( \7596 , \7590 , \7595 );
nand \U$6927 ( \7597 , \7583 , \7596 );
nand \U$6928 ( \7598 , \7581 , \7597 );
xor \U$6929 ( \7599 , \7477 , \7598 );
not \U$6930 ( \7600 , \7466 );
and \U$6931 ( \7601 , \7600 , \6930 );
not \U$6932 ( \7602 , \7600 );
and \U$6933 ( \7603 , \7602 , \6929 );
nor \U$6934 ( \7604 , \7601 , \7603 );
not \U$6935 ( \7605 , \7604 );
or \U$6936 ( \7606 , \7605 , \6925 );
or \U$6937 ( \7607 , \7401 , \6922 );
nand \U$6938 ( \7608 , \7606 , \7607 );
or \U$6939 ( \7609 , \7608 , \6927 );
and \U$6940 ( \7610 , \7599 , \7609 );
and \U$6941 ( \7611 , \7477 , \7598 );
nor \U$6942 ( \7612 , \7610 , \7611 );
not \U$6943 ( \7613 , \7612 );
not \U$6944 ( \7614 , \7394 );
nor \U$6945 ( \7615 , \7614 , \7392 );
xor \U$6946 ( \7616 , \7615 , \7349 );
or \U$6947 ( \7617 , \7153 , \6976 );
or \U$6948 ( \7618 , \7152 , \6975 );
nand \U$6949 ( \7619 , \7617 , \7618 );
not \U$6950 ( \7620 , \7619 );
not \U$6951 ( \7621 , \7155 );
nand \U$6952 ( \7622 , \7621 , \7160 );
not \U$6953 ( \7623 , \7622 );
not \U$6954 ( \7624 , \7623 );
or \U$6955 ( \7625 , \7620 , \7624 );
not \U$6956 ( \7626 , \7214 );
or \U$6957 ( \7627 , \7038 , \7152 );
nand \U$6958 ( \7628 , \7038 , \7152 );
nand \U$6959 ( \7629 , \7627 , \7628 );
and \U$6960 ( \7630 , \7626 , \7629 );
not \U$6961 ( \7631 , \7628 );
and \U$6962 ( \7632 , \7631 , \6975 );
nor \U$6963 ( \7633 , \7630 , \7632 );
nand \U$6964 ( \7634 , \7625 , \7633 );
not \U$6965 ( \7635 , \7634 );
nand \U$6966 ( \7636 , \7623 , \7626 );
nand \U$6967 ( \7637 , \7635 , \7636 );
not \U$6968 ( \7638 , \7637 );
not \U$6969 ( \7639 , \7376 );
and \U$6970 ( \7640 , \7371 , \7159 , \7374 );
nor \U$6971 ( \7641 , \7639 , \7640 );
not \U$6972 ( \7642 , \7641 );
not \U$6973 ( \7643 , \7378 );
or \U$6974 ( \7644 , \7642 , \7643 );
and \U$6975 ( \7645 , \7373 , \6894 );
buf \U$6976 ( \7646 , \7159 );
and \U$6977 ( \7647 , \7646 , \7084 );
nor \U$6978 ( \7648 , \7645 , \7647 );
nand \U$6979 ( \7649 , \7644 , \7648 );
not \U$6980 ( \7650 , \7637 );
xor \U$6981 ( \7651 , \7649 , \7650 );
nand \U$6982 ( \7652 , \7638 , \7651 );
xor \U$6983 ( \7653 , \7616 , \7652 );
not \U$6984 ( \7654 , \7653 );
or \U$6985 ( \7655 , \7613 , \7654 );
or \U$6986 ( \7656 , \7653 , \7612 );
nand \U$6987 ( \7657 , \7655 , \7656 );
not \U$6988 ( \7658 , \7657 );
not \U$6989 ( \7659 , \6923 );
not \U$6990 ( \7660 , \7604 );
or \U$6991 ( \7661 , \7659 , \7660 );
not \U$6992 ( \7662 , \1852 );
not \U$6993 ( \7663 , RIaaa3020_397);
not \U$6994 ( \7664 , \7663 );
and \U$6995 ( \7665 , \7662 , \7664 );
not \U$6996 ( \7666 , \2020 );
and \U$6997 ( \7667 , \7666 , RIaaa2f30_395);
nor \U$6998 ( \7668 , \7665 , \7667 );
and \U$6999 ( \7669 , \1640 , RIaaa2fa8_396);
and \U$7000 ( \7670 , \1642 , RIaaa2cd8_390);
nor \U$7001 ( \7671 , \7669 , \7670 );
not \U$7002 ( \7672 , RIaaa2eb8_394);
or \U$7003 ( \7673 , \7432 , \7672 );
not \U$7004 ( \7674 , RIaaa2be8_388);
or \U$7005 ( \7675 , \6848 , \7674 );
nand \U$7006 ( \7676 , \7673 , \7675 );
not \U$7007 ( \7677 , RIaaa2a08_384);
or \U$7008 ( \7678 , \2026 , \7677 );
and \U$7009 ( \7679 , \6868 , RIaaa3098_398);
and \U$7010 ( \7680 , \6871 , RIaaa3110_399);
nor \U$7011 ( \7681 , \7679 , \7680 );
nand \U$7012 ( \7682 , \7678 , \7681 );
nor \U$7013 ( \7683 , \7676 , \7682 );
not \U$7014 ( \7684 , \7013 );
not \U$7015 ( \7685 , RIaaa2dc8_392);
not \U$7016 ( \7686 , \7685 );
and \U$7017 ( \7687 , \7684 , \7686 );
not \U$7018 ( \7688 , RIaaa2e40_393);
nor \U$7019 ( \7689 , \7688 , \2068 );
nor \U$7020 ( \7690 , \7687 , \7689 );
nand \U$7021 ( \7691 , \7668 , \7671 , \7683 , \7690 );
not \U$7022 ( \7692 , \2061 );
not \U$7023 ( \7693 , \7692 );
not \U$7024 ( \7694 , RIaaa2c60_389);
not \U$7025 ( \7695 , \7694 );
and \U$7026 ( \7696 , \7693 , \7695 );
and \U$7027 ( \7697 , \1832 , RIaaa2d50_391);
nor \U$7028 ( \7698 , \7696 , \7697 );
not \U$7029 ( \7699 , \2014 );
not \U$7030 ( \7700 , RIaaa2af8_386);
not \U$7031 ( \7701 , \7700 );
and \U$7032 ( \7702 , \7699 , \7701 );
and \U$7033 ( \7703 , \2023 , RIaaa2b70_387);
nor \U$7034 ( \7704 , \7702 , \7703 );
nand \U$7035 ( \7705 , \2064 , RIaaa2a80_385);
nand \U$7036 ( \7706 , \7698 , \7704 , \2118 , \7705 );
nor \U$7037 ( \7707 , \7691 , \7706 );
buf \U$7038 ( \7708 , \7707 );
not \U$7039 ( \7709 , \7708 );
not \U$7040 ( \7710 , \7709 );
not \U$7041 ( \7711 , \7710 );
not \U$7042 ( \7712 , \7711 );
not \U$7043 ( \7713 , \6929 );
or \U$7044 ( \7714 , \7712 , \7713 );
or \U$7045 ( \7715 , \6929 , \7711 );
nand \U$7046 ( \7716 , \7714 , \7715 );
and \U$7047 ( \7717 , \7716 , \6926 );
or \U$7048 ( \7718 , \6929 , \7711 , \7600 );
nor \U$7049 ( \7719 , \7466 , \7710 );
nand \U$7050 ( \7720 , \6929 , \7719 );
nand \U$7051 ( \7721 , \7718 , \7720 );
nor \U$7052 ( \7722 , \7717 , \7721 );
nand \U$7053 ( \7723 , \7661 , \7722 );
nor \U$7054 ( \7724 , \7723 , \6927 );
not \U$7055 ( \7725 , \7724 );
not \U$7056 ( \7726 , \7725 );
xor \U$7057 ( \7727 , \7596 , \7582 );
not \U$7058 ( \7728 , \7727 );
not \U$7059 ( \7729 , \7038 );
not \U$7060 ( \7730 , \7639 );
or \U$7061 ( \7731 , \7729 , \7730 );
nor \U$7062 ( \7732 , \7150 , \7375 );
nand \U$7063 ( \7733 , \7732 , \7371 );
not \U$7064 ( \7734 , \7733 );
not \U$7065 ( \7735 , \7038 );
and \U$7066 ( \7736 , \7734 , \7735 );
and \U$7067 ( \7737 , \6975 , \7378 );
not \U$7068 ( \7738 , \6975 );
nand \U$7069 ( \7739 , \7370 , \7159 );
not \U$7070 ( \7740 , \7739 );
not \U$7071 ( \7741 , \7740 );
and \U$7072 ( \7742 , \7738 , \7741 );
nor \U$7073 ( \7743 , \7737 , \7742 );
nor \U$7074 ( \7744 , \7736 , \7743 );
nand \U$7075 ( \7745 , \7731 , \7744 );
nand \U$7076 ( \7746 , \7745 , \7574 );
not \U$7077 ( \7747 , \7746 );
not \U$7078 ( \7748 , \7600 );
not \U$7079 ( \7749 , \7102 );
or \U$7080 ( \7750 , \7748 , \7749 );
and \U$7081 ( \7751 , \7207 , \7472 );
not \U$7082 ( \7752 , \7207 );
and \U$7083 ( \7753 , \7752 , \7070 );
nor \U$7084 ( \7754 , \7751 , \7753 );
nand \U$7085 ( \7755 , \7750 , \7754 );
nor \U$7086 ( \7756 , \7067 , \7600 );
nor \U$7087 ( \7757 , \7755 , \7756 );
not \U$7088 ( \7758 , \7757 );
or \U$7089 ( \7759 , \7747 , \7758 );
not \U$7090 ( \7760 , \7745 );
nand \U$7091 ( \7761 , \7760 , \7573 );
nand \U$7092 ( \7762 , \7759 , \7761 );
not \U$7093 ( \7763 , \7762 );
or \U$7094 ( \7764 , \7728 , \7763 );
or \U$7095 ( \7765 , \7762 , \7727 );
nand \U$7096 ( \7766 , \7764 , \7765 );
not \U$7097 ( \7767 , \7766 );
or \U$7098 ( \7768 , \7726 , \7767 );
not \U$7099 ( \7769 , \7727 );
nand \U$7100 ( \7770 , \7769 , \7762 );
nand \U$7101 ( \7771 , \7768 , \7770 );
not \U$7102 ( \7772 , \7771 );
and \U$7103 ( \7773 , \7623 , \7629 );
not \U$7104 ( \7774 , \7626 );
and \U$7105 ( \7775 , \7265 , \7153 );
not \U$7106 ( \7776 , \7265 );
and \U$7107 ( \7777 , \7776 , \7152 );
nor \U$7108 ( \7778 , \7775 , \7777 );
or \U$7109 ( \7779 , \7774 , \7778 );
or \U$7110 ( \7780 , \7628 , \7265 );
nand \U$7111 ( \7781 , \7779 , \7780 );
nor \U$7112 ( \7782 , \7773 , \7781 );
nand \U$7113 ( \7783 , \7782 , \7636 );
not \U$7114 ( \7784 , \7783 );
not \U$7115 ( \7785 , \7639 );
nor \U$7116 ( \7786 , \7785 , \6976 );
not \U$7117 ( \7787 , \6976 );
not \U$7118 ( \7788 , \7640 );
or \U$7119 ( \7789 , \7787 , \7788 );
and \U$7120 ( \7790 , \7370 , \7150 );
and \U$7121 ( \7791 , \7084 , \7790 );
not \U$7122 ( \7792 , \7084 );
and \U$7123 ( \7793 , \7792 , \7740 );
nor \U$7124 ( \7794 , \7791 , \7793 );
nand \U$7125 ( \7795 , \7789 , \7794 );
nor \U$7126 ( \7796 , \7786 , \7795 );
not \U$7127 ( \7797 , \7796 );
nand \U$7128 ( \7798 , \7784 , \7797 );
not \U$7129 ( \7799 , \7798 );
nand \U$7130 ( \7800 , \6847 , \7711 );
nand \U$7131 ( \7801 , \7651 , \7800 );
not \U$7132 ( \7802 , \7801 );
or \U$7133 ( \7803 , \7799 , \7802 );
or \U$7134 ( \7804 , \7801 , \7798 );
nand \U$7135 ( \7805 , \7803 , \7804 );
not \U$7136 ( \7806 , \7805 );
or \U$7137 ( \7807 , \7772 , \7806 );
not \U$7138 ( \7808 , \7801 );
nand \U$7139 ( \7809 , \7808 , \7798 );
nand \U$7140 ( \7810 , \7807 , \7809 );
and \U$7141 ( \7811 , \7407 , \7478 );
nor \U$7142 ( \7812 , \7811 , \7479 );
and \U$7143 ( \7813 , \7810 , \7812 );
not \U$7144 ( \7814 , \7810 );
not \U$7145 ( \7815 , \7812 );
and \U$7146 ( \7816 , \7814 , \7815 );
or \U$7147 ( \7817 , \7813 , \7816 );
not \U$7148 ( \7818 , \7817 );
or \U$7149 ( \7819 , \7658 , \7818 );
nand \U$7150 ( \7820 , \7810 , \7815 );
nand \U$7151 ( \7821 , \7819 , \7820 );
not \U$7152 ( \7822 , \7612 );
not \U$7153 ( \7823 , \7822 );
not \U$7154 ( \7824 , \7653 );
or \U$7155 ( \7825 , \7823 , \7824 );
nand \U$7156 ( \7826 , \7652 , \7616 );
nand \U$7157 ( \7827 , \7825 , \7826 );
not \U$7158 ( \7828 , \7114 );
not \U$7159 ( \7829 , \7217 );
and \U$7160 ( \7830 , \7828 , \7829 );
and \U$7161 ( \7831 , \7114 , \7217 );
nor \U$7162 ( \7832 , \7830 , \7831 );
buf \U$7163 ( \7833 , \7832 );
not \U$7164 ( \7834 , \7833 );
xor \U$7165 ( \7835 , \7334 , \7395 );
xor \U$7166 ( \7836 , \7835 , \7479 );
not \U$7167 ( \7837 , \7836 );
or \U$7168 ( \7838 , \7834 , \7837 );
or \U$7169 ( \7839 , \7836 , \7833 );
nand \U$7170 ( \7840 , \7838 , \7839 );
xor \U$7171 ( \7841 , \7827 , \7840 );
nand \U$7172 ( \7842 , \7821 , \7841 );
xor \U$7173 ( \7843 , \7498 , \7482 );
xnor \U$7174 ( \7844 , \7843 , \7317 );
not \U$7175 ( \7845 , \7840 );
not \U$7176 ( \7846 , \7827 );
or \U$7177 ( \7847 , \7845 , \7846 );
not \U$7178 ( \7848 , \7836 );
nand \U$7179 ( \7849 , \7848 , \7833 );
nand \U$7180 ( \7850 , \7847 , \7849 );
nand \U$7181 ( \7851 , \7844 , \7850 );
nand \U$7182 ( \7852 , \7536 , \7842 , \7851 );
not \U$7183 ( \7853 , \7852 );
not \U$7184 ( \7854 , \7853 );
nor \U$7185 ( \7855 , \7554 , \7557 );
buf \U$7186 ( \7856 , \7855 );
not \U$7187 ( \7857 , \7856 );
not \U$7188 ( \7858 , \6893 );
or \U$7189 ( \7859 , \7857 , \7858 );
or \U$7190 ( \7860 , \7559 , \6894 );
nand \U$7191 ( \7861 , \7859 , \7860 );
not \U$7192 ( \7862 , \7861 );
and \U$7193 ( \7863 , \7554 , \7562 , \7564 , \7368 );
not \U$7194 ( \7864 , \7863 );
not \U$7195 ( \7865 , \7864 );
and \U$7196 ( \7866 , \6976 , \7865 );
not \U$7197 ( \7867 , \6976 );
and \U$7198 ( \7868 , \7867 , \7577 );
nor \U$7199 ( \7869 , \7866 , \7868 );
nand \U$7200 ( \7870 , \7862 , \7869 );
not \U$7201 ( \7871 , \7870 );
buf \U$7202 ( \7872 , \7540 );
xnor \U$7203 ( \7873 , \853 , \6367 );
buf \U$7204 ( \7874 , \6784 );
xor \U$7205 ( \7875 , \7873 , \7874 );
not \U$7206 ( \7876 , \7875 );
buf \U$7207 ( \7877 , \6781 );
and \U$7208 ( \7878 , \6262 , RIaa977e8_4);
not \U$7209 ( \7879 , \6262 );
and \U$7210 ( \7880 , \7879 , \849 );
nor \U$7211 ( \7881 , \7878 , \7880 );
xor \U$7212 ( \7882 , \7877 , \7881 );
nand \U$7213 ( \7883 , \7876 , \7882 );
and \U$7214 ( \7884 , \7872 , \7883 );
not \U$7215 ( \7885 , \7884 );
nor \U$7216 ( \7886 , \7554 , \7570 );
buf \U$7217 ( \7887 , \7886 );
not \U$7218 ( \7888 , \7887 );
not \U$7219 ( \7889 , \6974 );
or \U$7220 ( \7890 , \7888 , \7889 );
not \U$7221 ( \7891 , \7856 );
not \U$7222 ( \7892 , \6974 );
not \U$7223 ( \7893 , \7892 );
or \U$7224 ( \7894 , \7891 , \7893 );
nand \U$7225 ( \7895 , \7890 , \7894 );
not \U$7226 ( \7896 , \7895 );
and \U$7227 ( \7897 , \7039 , \7865 );
not \U$7228 ( \7898 , \7039 );
and \U$7229 ( \7899 , \7898 , \7577 );
nor \U$7230 ( \7900 , \7897 , \7899 );
nand \U$7231 ( \7901 , \7896 , \7900 );
not \U$7232 ( \7902 , \7901 );
or \U$7233 ( \7903 , \7885 , \7902 );
or \U$7234 ( \7904 , \7901 , \7884 );
nand \U$7235 ( \7905 , \7903 , \7904 );
not \U$7236 ( \7906 , \7905 );
or \U$7237 ( \7907 , \7871 , \7906 );
not \U$7238 ( \7908 , \7884 );
and \U$7239 ( \7909 , \7901 , \7908 );
nand \U$7240 ( \7910 , \1872 , RIaaa3f20_429);
not \U$7241 ( \7911 , RIaaa3d40_425);
nor \U$7242 ( \7912 , \7911 , \7013 );
not \U$7243 ( \7913 , RIaaa3cc8_424);
nor \U$7244 ( \7914 , \7913 , \2068 );
nor \U$7245 ( \7915 , \7912 , \7914 );
nand \U$7246 ( \7916 , \7910 , \2662 , \7915 );
not \U$7247 ( \7917 , \2063 );
not \U$7248 ( \7918 , RIaaa39f8_418);
not \U$7249 ( \7919 , \7918 );
and \U$7250 ( \7920 , \7917 , \7919 );
and \U$7251 ( \7921 , \2023 , RIaaa3ea8_428);
nor \U$7252 ( \7922 , \7920 , \7921 );
not \U$7253 ( \7923 , \2026 );
not \U$7254 ( \7924 , RIaaa3a70_419);
not \U$7255 ( \7925 , \7924 );
and \U$7256 ( \7926 , \7923 , \7925 );
and \U$7257 ( \7927 , \1861 , RIaaa3e30_427);
nor \U$7258 ( \7928 , \7926 , \7927 );
nand \U$7259 ( \7929 , \7922 , \7928 );
nor \U$7260 ( \7930 , \7916 , \7929 );
not \U$7261 ( \7931 , \6882 );
not \U$7262 ( \7932 , \2680 );
and \U$7263 ( \7933 , \7931 , \7932 );
not \U$7264 ( \7934 , RIaaa3b60_421);
nor \U$7265 ( \7935 , \7934 , \1743 );
nor \U$7266 ( \7936 , \7933 , \7935 );
and \U$7267 ( \7937 , \1832 , RIaaa3ae8_420);
and \U$7268 ( \7938 , \6868 , RIaaa4178_434);
and \U$7269 ( \7939 , \6871 , RIaaa4100_433);
nor \U$7270 ( \7940 , \7938 , \7939 );
not \U$7271 ( \7941 , \7940 );
nor \U$7272 ( \7942 , \7937 , \7941 );
nand \U$7273 ( \7943 , \7936 , \7942 );
not \U$7274 ( \7944 , RIaaa3c50_423);
nor \U$7275 ( \7945 , \7944 , \2020 );
not \U$7276 ( \7946 , RIaaa3f98_430);
nor \U$7277 ( \7947 , \7946 , \2052 );
nor \U$7278 ( \7948 , \7945 , \7947 );
not \U$7279 ( \7949 , \2014 );
not \U$7280 ( \7950 , RIaaa4010_431);
not \U$7281 ( \7951 , \7950 );
and \U$7282 ( \7952 , \7949 , \7951 );
not \U$7283 ( \7953 , RIaaa4088_432);
nor \U$7284 ( \7954 , \1852 , \7953 );
nor \U$7285 ( \7955 , \7952 , \7954 );
nand \U$7286 ( \7956 , \7948 , \7955 );
nor \U$7287 ( \7957 , \7943 , \7956 );
nand \U$7288 ( \7958 , \7930 , \7957 );
not \U$7289 ( \7959 , \7958 );
buf \U$7290 ( \7960 , \7959 );
not \U$7291 ( \7961 , \7960 );
and \U$7292 ( \7962 , \6847 , \7961 );
nor \U$7293 ( \7963 , \7909 , \7962 );
nand \U$7294 ( \7964 , \7907 , \7963 );
and \U$7295 ( \7965 , \7338 , \7265 );
and \U$7296 ( \7966 , \7309 , \7155 );
not \U$7297 ( \7967 , \7309 );
and \U$7298 ( \7968 , \7967 , \7161 );
or \U$7299 ( \7969 , \7966 , \7968 );
nor \U$7300 ( \7970 , \7965 , \7969 );
not \U$7301 ( \7971 , \7216 );
nand \U$7302 ( \7972 , \7971 , \7269 );
nand \U$7303 ( \7973 , \7970 , \7972 );
nand \U$7304 ( \7974 , \7964 , \7973 );
not \U$7305 ( \7975 , \7974 );
and \U$7306 ( \7976 , \7174 , RIaaa2828_380);
and \U$7307 ( \7977 , \7666 , RIaaa27b0_379);
nor \U$7308 ( \7978 , \7976 , \7977 );
and \U$7309 ( \7979 , \1626 , RIaaa2558_374);
and \U$7310 ( \7980 , \6889 , RIaaa25d0_375);
nor \U$7311 ( \7981 , \7979 , \7980 );
and \U$7312 ( \7982 , \6883 , RIaaa2738_378);
and \U$7313 ( \7983 , RIaaa28a0_381, \6871 );
and \U$7314 ( \7984 , \6868 , RIaaa2918_382);
nor \U$7315 ( \7985 , \7982 , \7983 , \7984 );
nand \U$7316 ( \7986 , \7978 , \7981 , \7985 , \2480 );
not \U$7317 ( \7987 , \7986 );
not \U$7318 ( \7988 , \2026 );
not \U$7319 ( \7989 , RIaaa24e0_373);
not \U$7320 ( \7990 , \7989 );
and \U$7321 ( \7991 , \7988 , \7990 );
and \U$7322 ( \7992 , \1861 , RIaaa26c0_377);
nor \U$7323 ( \7993 , \7991 , \7992 );
and \U$7324 ( \7994 , \2064 , RIaaa2468_372);
not \U$7325 ( \7995 , RIaaa23f0_371);
nor \U$7326 ( \7996 , \7995 , \2052 );
nor \U$7327 ( \7997 , \7994 , \7996 );
nand \U$7328 ( \7998 , \7993 , \7997 );
nand \U$7329 ( \7999 , \1832 , RIaaa2300_369);
nand \U$7330 ( \8000 , \1642 , RIaaa2378_370);
not \U$7331 ( \8001 , \7415 );
nand \U$7332 ( \8002 , \8001 , RIaaa2288_368);
nand \U$7333 ( \8003 , \7999 , \8000 , \8002 );
not \U$7334 ( \8004 , RIaaa2210_367);
not \U$7335 ( \8005 , \7014 );
or \U$7336 ( \8006 , \8004 , \8005 );
not \U$7337 ( \8007 , \7692 );
nand \U$7338 ( \8008 , \8007 , RIaaa2648_376);
nand \U$7339 ( \8009 , \8006 , \8008 );
nor \U$7340 ( \8010 , \7998 , \8003 , \8009 );
nand \U$7341 ( \8011 , \7987 , \8010 );
not \U$7342 ( \8012 , \8011 );
not \U$7343 ( \8013 , \8012 );
not \U$7344 ( \8014 , \8013 );
not \U$7345 ( \8015 , \6847 );
or \U$7346 ( \8016 , \8014 , \8015 );
not \U$7347 ( \8017 , \7783 );
not \U$7348 ( \8018 , \7796 );
or \U$7349 ( \8019 , \8017 , \8018 );
nand \U$7350 ( \8020 , \8019 , \7798 );
nand \U$7351 ( \8021 , \8016 , \8020 );
not \U$7352 ( \8022 , \8021 );
or \U$7353 ( \8023 , \7975 , \8022 );
or \U$7354 ( \8024 , \8021 , \7974 );
nand \U$7355 ( \8025 , \8023 , \8024 );
not \U$7356 ( \8026 , \8025 );
not \U$7357 ( \8027 , \7724 );
not \U$7358 ( \8028 , \7766 );
or \U$7359 ( \8029 , \8027 , \8028 );
or \U$7360 ( \8030 , \7766 , \7724 );
nand \U$7361 ( \8031 , \8029 , \8030 );
not \U$7362 ( \8032 , \8031 );
or \U$7363 ( \8033 , \8026 , \8032 );
or \U$7364 ( \8034 , \8031 , \8025 );
nand \U$7365 ( \8035 , \8033 , \8034 );
not \U$7366 ( \8036 , \8035 );
xor \U$7367 ( \8037 , \7574 , \7745 );
xnor \U$7368 ( \8038 , \8037 , \7757 );
not \U$7369 ( \8039 , \8013 );
and \U$7370 ( \8040 , \6986 , \8039 );
and \U$7371 ( \8041 , \7711 , \7080 );
not \U$7372 ( \8042 , \7711 );
and \U$7373 ( \8043 , \8042 , \6993 );
nor \U$7374 ( \8044 , \8041 , \8043 );
nor \U$7375 ( \8045 , \8040 , \8044 );
nand \U$7376 ( \8046 , \6990 , \8013 );
nand \U$7377 ( \8047 , \8045 , \8046 );
xor \U$7378 ( \8048 , \8038 , \8047 );
or \U$7379 ( \8049 , \7337 , \7308 );
not \U$7380 ( \8050 , \7155 );
not \U$7381 ( \8051 , \8050 );
not \U$7382 ( \8052 , \7206 );
and \U$7383 ( \8053 , \8051 , \8052 );
and \U$7384 ( \8054 , \7161 , \7206 );
nor \U$7385 ( \8055 , \8053 , \8054 );
nand \U$7386 ( \8056 , \8049 , \8055 );
nor \U$7387 ( \8057 , \7216 , \7309 );
nor \U$7388 ( \8058 , \8056 , \8057 );
not \U$7389 ( \8059 , \8058 );
not \U$7390 ( \8060 , \7269 );
not \U$7391 ( \8061 , \7376 );
not \U$7392 ( \8062 , \8061 );
or \U$7393 ( \8063 , \8060 , \8062 );
not \U$7394 ( \8064 , \7733 );
not \U$7395 ( \8065 , \7269 );
and \U$7396 ( \8066 , \8064 , \8065 );
and \U$7397 ( \8067 , \7039 , \7741 );
not \U$7398 ( \8068 , \7039 );
and \U$7399 ( \8069 , \8068 , \7378 );
nor \U$7400 ( \8070 , \8067 , \8069 );
nor \U$7401 ( \8071 , \8066 , \8070 );
nand \U$7402 ( \8072 , \8063 , \8071 );
not \U$7403 ( \8073 , \7710 );
not \U$7404 ( \8074 , \7389 );
or \U$7405 ( \8075 , \8073 , \8074 );
and \U$7406 ( \8076 , \7102 , \7711 );
or \U$7407 ( \8077 , \7071 , \7600 );
nand \U$7408 ( \8078 , \7472 , \7600 );
nand \U$7409 ( \8079 , \8077 , \8078 );
nor \U$7410 ( \8080 , \8076 , \8079 );
nand \U$7411 ( \8081 , \8075 , \8080 );
xor \U$7412 ( \8082 , \8072 , \8081 );
and \U$7413 ( \8083 , \8059 , \8082 );
and \U$7414 ( \8084 , \8072 , \8081 );
nor \U$7415 ( \8085 , \8083 , \8084 );
not \U$7416 ( \8086 , \8085 );
and \U$7417 ( \8087 , \8048 , \8086 );
and \U$7418 ( \8088 , \8038 , \8047 );
nor \U$7419 ( \8089 , \8087 , \8088 );
not \U$7420 ( \8090 , \8089 );
and \U$7421 ( \8091 , \8036 , \8090 );
and \U$7422 ( \8092 , \8035 , \8089 );
nor \U$7423 ( \8093 , \8091 , \8092 );
not \U$7424 ( \8094 , \8093 );
xor \U$7425 ( \8095 , \8082 , \8058 );
not \U$7426 ( \8096 , \8095 );
not \U$7427 ( \8097 , \8096 );
and \U$7428 ( \8098 , \7038 , \7887 );
not \U$7429 ( \8099 , \7038 );
and \U$7430 ( \8100 , \8099 , \7856 );
or \U$7431 ( \8101 , \8098 , \8100 );
not \U$7432 ( \8102 , \8101 );
and \U$7433 ( \8103 , \7265 , \7865 );
not \U$7434 ( \8104 , \7265 );
and \U$7435 ( \8105 , \8104 , \7577 );
nor \U$7436 ( \8106 , \8103 , \8105 );
nand \U$7437 ( \8107 , \8102 , \8106 );
not \U$7438 ( \8108 , \7882 );
nor \U$7439 ( \8109 , \8107 , \8108 );
buf \U$7440 ( \8110 , \8109 );
not \U$7441 ( \8111 , \8110 );
not \U$7442 ( \8112 , \8111 );
not \U$7443 ( \8113 , \6894 );
xnor \U$7444 ( \8114 , \7540 , \7875 );
not \U$7445 ( \8115 , \7882 );
nand \U$7446 ( \8116 , \8115 , \7875 );
nand \U$7447 ( \8117 , \7883 , \8116 );
nand \U$7448 ( \8118 , \8114 , \8117 );
not \U$7449 ( \8119 , \8118 );
not \U$7450 ( \8120 , \7872 );
nand \U$7451 ( \8121 , \8119 , \8120 );
not \U$7452 ( \8122 , \8121 );
not \U$7453 ( \8123 , \8122 );
or \U$7454 ( \8124 , \8113 , \8123 );
buf \U$7455 ( \8125 , \8118 );
nor \U$7456 ( \8126 , \8125 , \8120 );
buf \U$7457 ( \8127 , \8126 );
and \U$7458 ( \8128 , \8127 , \7568 );
not \U$7459 ( \8129 , \8117 );
nand \U$7460 ( \8130 , \8129 , \7872 );
not \U$7461 ( \8131 , \8130 );
nor \U$7462 ( \8132 , \8128 , \8131 );
nand \U$7463 ( \8133 , \8124 , \8132 );
and \U$7464 ( \8134 , \8133 , \7901 );
not \U$7465 ( \8135 , \8133 );
not \U$7466 ( \8136 , \7901 );
and \U$7467 ( \8137 , \8135 , \8136 );
or \U$7468 ( \8138 , \8134 , \8137 );
not \U$7469 ( \8139 , \8138 );
or \U$7470 ( \8140 , \8112 , \8139 );
nand \U$7471 ( \8141 , \8136 , \8133 );
nand \U$7472 ( \8142 , \8140 , \8141 );
or \U$7473 ( \8143 , \7216 , \7207 );
nand \U$7474 ( \8144 , \7338 , \7207 );
and \U$7475 ( \8145 , \7161 , \7466 );
and \U$7476 ( \8146 , \7155 , \7600 );
nor \U$7477 ( \8147 , \8145 , \8146 );
nand \U$7478 ( \8148 , \8143 , \8144 , \8147 );
not \U$7479 ( \8149 , \8148 );
not \U$7480 ( \8150 , \7308 );
not \U$7481 ( \8151 , \8061 );
or \U$7482 ( \8152 , \8150 , \8151 );
not \U$7483 ( \8153 , \7308 );
not \U$7484 ( \8154 , \7733 );
and \U$7485 ( \8155 , \8153 , \8154 );
and \U$7486 ( \8156 , \7265 , \7741 );
not \U$7487 ( \8157 , \7265 );
and \U$7488 ( \8158 , \8157 , \7378 );
nor \U$7489 ( \8159 , \8156 , \8158 );
nor \U$7490 ( \8160 , \8155 , \8159 );
nand \U$7491 ( \8161 , \8152 , \8160 );
not \U$7492 ( \8162 , \8039 );
not \U$7493 ( \8163 , \7389 );
or \U$7494 ( \8164 , \8162 , \8163 );
and \U$7495 ( \8165 , \7102 , \8013 );
or \U$7496 ( \8166 , \7069 , \7711 );
nand \U$7497 ( \8167 , \7107 , \7711 );
nand \U$7498 ( \8168 , \8166 , \8167 );
nor \U$7499 ( \8169 , \8165 , \8168 );
nand \U$7500 ( \8170 , \8164 , \8169 );
xor \U$7501 ( \8171 , \8161 , \8170 );
not \U$7502 ( \8172 , \8171 );
or \U$7503 ( \8173 , \8149 , \8172 );
nand \U$7504 ( \8174 , \8170 , \8161 );
nand \U$7505 ( \8175 , \8173 , \8174 );
xor \U$7506 ( \8176 , \8142 , \8175 );
not \U$7507 ( \8177 , \8176 );
or \U$7508 ( \8178 , \8097 , \8177 );
nand \U$7509 ( \8179 , \8175 , \8142 );
nand \U$7510 ( \8180 , \8178 , \8179 );
not \U$7511 ( \8181 , \8180 );
or \U$7512 ( \8182 , \7080 , \8039 );
not \U$7513 ( \8183 , \6992 );
nand \U$7514 ( \8184 , \8183 , \8039 );
nand \U$7515 ( \8185 , \8182 , \8184 );
not \U$7516 ( \8186 , \8185 );
not \U$7517 ( \8187 , \7961 );
nand \U$7518 ( \8188 , \8187 , \6986 );
nand \U$7519 ( \8189 , \6990 , \7961 );
nand \U$7520 ( \8190 , \8186 , \8188 , \8189 );
xor \U$7521 ( \8191 , \7870 , \7905 );
buf \U$7522 ( \8192 , \8191 );
xor \U$7523 ( \8193 , \8190 , \8192 );
nand \U$7524 ( \8194 , \2023 , RIaaa32f0_403);
nand \U$7525 ( \8195 , \6889 , RIaaa3458_406);
nand \U$7526 ( \8196 , \8007 , RIaaa3368_404);
nand \U$7527 ( \8197 , \2901 , \8194 , \8195 , \8196 );
not \U$7528 ( \8198 , \1852 );
not \U$7529 ( \8199 , RIaaa34d0_407);
not \U$7530 ( \8200 , \8199 );
and \U$7531 ( \8201 , \8198 , \8200 );
not \U$7532 ( \8202 , \2036 );
and \U$7533 ( \8203 , \8202 , RIaaa3278_402);
nor \U$7534 ( \8204 , \8201 , \8203 );
and \U$7535 ( \8205 , \1846 , RIaaa33e0_405);
and \U$7536 ( \8206 , RIaaa35c0_409, \6868 );
and \U$7537 ( \8207 , \6871 , RIaaa3548_408);
nor \U$7538 ( \8208 , \8205 , \8206 , \8207 );
nand \U$7539 ( \8209 , \8204 , \8208 );
nor \U$7540 ( \8210 , \8197 , \8209 );
and \U$7541 ( \8211 , \1832 , RIaaa3728_412);
and \U$7542 ( \8212 , \1642 , RIaaa37a0_413);
nor \U$7543 ( \8213 , \8211 , \8212 );
not \U$7544 ( \8214 , \2046 );
not \U$7545 ( \8215 , RIaaa3638_410);
not \U$7546 ( \8216 , \8215 );
and \U$7547 ( \8217 , \8214 , \8216 );
and \U$7548 ( \8218 , \6939 , RIaaa36b0_411);
nor \U$7549 ( \8219 , \8217 , \8218 );
nand \U$7550 ( \8220 , \8213 , \8219 );
nand \U$7551 ( \8221 , \2064 , RIaaa3818_414);
nand \U$7552 ( \8222 , \2069 , RIaaa3908_416);
nand \U$7553 ( \8223 , \6856 , RIaaa3980_417);
not \U$7554 ( \8224 , \2026 );
nand \U$7555 ( \8225 , \8224 , RIaaa3890_415);
nand \U$7556 ( \8226 , \8221 , \8222 , \8223 , \8225 );
nor \U$7557 ( \8227 , \8220 , \8226 );
nand \U$7558 ( \8228 , \8210 , \8227 );
buf \U$7559 ( \8229 , \8228 );
not \U$7560 ( \8230 , \8229 );
not \U$7561 ( \8231 , \8230 );
not \U$7562 ( \8232 , \8231 );
not \U$7563 ( \8233 , \8232 );
and \U$7564 ( \8234 , \6847 , \8233 );
and \U$7565 ( \8235 , \8193 , \8234 );
and \U$7566 ( \8236 , \8190 , \8192 );
nor \U$7567 ( \8237 , \8235 , \8236 );
not \U$7568 ( \8238 , \8237 );
not \U$7569 ( \8239 , \7974 );
nor \U$7570 ( \8240 , \7964 , \7973 );
nor \U$7571 ( \8241 , \8239 , \8240 );
not \U$7572 ( \8242 , \8241 );
or \U$7573 ( \8243 , \8238 , \8242 );
or \U$7574 ( \8244 , \8237 , \8241 );
nand \U$7575 ( \8245 , \8243 , \8244 );
not \U$7576 ( \8246 , \8245 );
or \U$7577 ( \8247 , \8181 , \8246 );
not \U$7578 ( \8248 , \8237 );
nand \U$7579 ( \8249 , \8248 , \8241 );
nand \U$7580 ( \8250 , \8247 , \8249 );
nand \U$7581 ( \8251 , \8094 , \8250 );
xor \U$7582 ( \8252 , \7771 , \7805 );
not \U$7583 ( \8253 , \7974 );
nand \U$7584 ( \8254 , \8021 , \8253 );
not \U$7585 ( \8255 , \8254 );
not \U$7586 ( \8256 , \8031 );
or \U$7587 ( \8257 , \8255 , \8256 );
or \U$7588 ( \8258 , \8021 , \8253 );
nand \U$7589 ( \8259 , \8257 , \8258 );
not \U$7590 ( \8260 , \8259 );
xnor \U$7591 ( \8261 , \7609 , \7599 );
not \U$7592 ( \8262 , \8261 );
and \U$7593 ( \8263 , \8260 , \8262 );
and \U$7594 ( \8264 , \8259 , \8261 );
nor \U$7595 ( \8265 , \8263 , \8264 );
not \U$7596 ( \8266 , \8265 );
xor \U$7597 ( \8267 , \8252 , \8266 );
not \U$7598 ( \8268 , \8089 );
nand \U$7599 ( \8269 , \8268 , \8035 );
nand \U$7600 ( \8270 , \8251 , \8267 , \8269 );
not \U$7601 ( \8271 , \8245 );
not \U$7602 ( \8272 , \8180 );
not \U$7603 ( \8273 , \8272 );
and \U$7604 ( \8274 , \8271 , \8273 );
and \U$7605 ( \8275 , \8245 , \8272 );
nor \U$7606 ( \8276 , \8274 , \8275 );
not \U$7607 ( \8277 , \8276 );
xnor \U$7608 ( \8278 , \8085 , \8048 );
not \U$7609 ( \8279 , \8278 );
and \U$7610 ( \8280 , \8138 , \8110 );
not \U$7611 ( \8281 , \8138 );
and \U$7612 ( \8282 , \8281 , \8111 );
or \U$7613 ( \8283 , \8280 , \8282 );
nor \U$7614 ( \8284 , \7216 , \7600 );
not \U$7615 ( \8285 , \8284 );
nand \U$7616 ( \8286 , \7336 , \7600 );
and \U$7617 ( \8287 , \7155 , \7711 );
nor \U$7618 ( \8288 , \7160 , \7711 );
nor \U$7619 ( \8289 , \8287 , \8288 );
nand \U$7620 ( \8290 , \8285 , \8286 , \8289 );
not \U$7621 ( \8291 , \8290 );
not \U$7622 ( \8292 , \7067 );
not \U$7623 ( \8293 , \7961 );
and \U$7624 ( \8294 , \8292 , \8293 );
not \U$7625 ( \8295 , \7961 );
not \U$7626 ( \8296 , \7101 );
or \U$7627 ( \8297 , \8295 , \8296 );
and \U$7628 ( \8298 , \8013 , \7107 );
not \U$7629 ( \8299 , \8013 );
and \U$7630 ( \8300 , \8299 , \7070 );
nor \U$7631 ( \8301 , \8298 , \8300 );
nand \U$7632 ( \8302 , \8297 , \8301 );
nor \U$7633 ( \8303 , \8294 , \8302 );
not \U$7634 ( \8304 , \8303 );
not \U$7635 ( \8305 , \8304 );
not \U$7636 ( \8306 , \8109 );
nand \U$7637 ( \8307 , \8107 , \8108 );
nand \U$7638 ( \8308 , \8306 , \8307 );
not \U$7639 ( \8309 , \8308 );
not \U$7640 ( \8310 , \8309 );
or \U$7641 ( \8311 , \8305 , \8310 );
nand \U$7642 ( \8312 , \8303 , \8308 );
nand \U$7643 ( \8313 , \8311 , \8312 );
not \U$7644 ( \8314 , \8313 );
or \U$7645 ( \8315 , \8291 , \8314 );
nand \U$7646 ( \8316 , \8304 , \8308 );
nand \U$7647 ( \8317 , \8315 , \8316 );
xor \U$7648 ( \8318 , \8283 , \8317 );
xor \U$7649 ( \8319 , \8148 , \8171 );
and \U$7650 ( \8320 , \8318 , \8319 );
and \U$7651 ( \8321 , \8283 , \8317 );
nor \U$7652 ( \8322 , \8320 , \8321 );
not \U$7653 ( \8323 , \8322 );
not \U$7654 ( \8324 , \8323 );
xor \U$7655 ( \8325 , \8234 , \8191 );
xnor \U$7656 ( \8326 , \8325 , \8190 );
not \U$7657 ( \8327 , \8326 );
not \U$7658 ( \8328 , \8327 );
or \U$7659 ( \8329 , \8324 , \8328 );
not \U$7660 ( \8330 , \8326 );
not \U$7661 ( \8331 , \8322 );
or \U$7662 ( \8332 , \8330 , \8331 );
not \U$7663 ( \8333 , \8233 );
not \U$7664 ( \8334 , \6990 );
or \U$7665 ( \8335 , \8333 , \8334 );
and \U$7666 ( \8336 , \6986 , \8232 );
and \U$7667 ( \8337 , \7960 , \6993 );
not \U$7668 ( \8338 , \7960 );
and \U$7669 ( \8339 , \8338 , \7080 );
nor \U$7670 ( \8340 , \8337 , \8339 );
nor \U$7671 ( \8341 , \8336 , \8340 );
nand \U$7672 ( \8342 , \8335 , \8341 );
not \U$7673 ( \8343 , RIaa9ce28_188);
not \U$7674 ( \8344 , \6319 );
or \U$7675 ( \8345 , \8343 , \8344 );
nand \U$7676 ( \8346 , \8345 , \6781 );
not \U$7677 ( \8347 , \8346 );
and \U$7678 ( \8348 , \7882 , \8347 );
not \U$7679 ( \8349 , \8348 );
not \U$7680 ( \8350 , \6893 );
or \U$7681 ( \8351 , \8349 , \8350 );
nand \U$7682 ( \8352 , \8351 , \7882 );
not \U$7683 ( \8353 , \8352 );
not \U$7684 ( \8354 , \8353 );
not \U$7685 ( \8355 , \7039 );
not \U$7686 ( \8356 , \8122 );
or \U$7687 ( \8357 , \8355 , \8356 );
and \U$7688 ( \8358 , \8126 , \7038 );
not \U$7689 ( \8359 , \8117 );
nand \U$7690 ( \8360 , \8359 , \8120 );
not \U$7691 ( \8361 , \8360 );
not \U$7692 ( \8362 , \8361 );
or \U$7693 ( \8363 , \8362 , \6974 );
nand \U$7694 ( \8364 , \8131 , \6974 );
nand \U$7695 ( \8365 , \8363 , \8364 );
nor \U$7696 ( \8366 , \8358 , \8365 );
nand \U$7697 ( \8367 , \8357 , \8366 );
not \U$7698 ( \8368 , \8367 );
or \U$7699 ( \8369 , \8354 , \8368 );
not \U$7700 ( \8370 , \6974 );
not \U$7701 ( \8371 , \8127 );
or \U$7702 ( \8372 , \8370 , \8371 );
and \U$7703 ( \8373 , \7568 , \8131 );
not \U$7704 ( \8374 , \7568 );
and \U$7705 ( \8375 , \8374 , \8361 );
nor \U$7706 ( \8376 , \8373 , \8375 );
nand \U$7707 ( \8377 , \8372 , \8376 );
and \U$7708 ( \8378 , \8122 , \7892 );
nor \U$7709 ( \8379 , \8377 , \8378 );
nand \U$7710 ( \8380 , \8369 , \8379 );
not \U$7711 ( \8381 , \8380 );
not \U$7712 ( \8382 , \7785 );
not \U$7713 ( \8383 , \7207 );
and \U$7714 ( \8384 , \8382 , \8383 );
not \U$7715 ( \8385 , \7207 );
not \U$7716 ( \8386 , \7640 );
or \U$7717 ( \8387 , \8385 , \8386 );
and \U$7718 ( \8388 , \7585 , \7740 );
not \U$7719 ( \8389 , \7585 );
and \U$7720 ( \8390 , \8389 , \7790 );
nor \U$7721 ( \8391 , \8388 , \8390 );
nand \U$7722 ( \8392 , \8387 , \8391 );
nor \U$7723 ( \8393 , \8384 , \8392 );
not \U$7724 ( \8394 , \8393 );
not \U$7725 ( \8395 , \8394 );
or \U$7726 ( \8396 , \8381 , \8395 );
not \U$7727 ( \8397 , \6888 );
not \U$7728 ( \8398 , \3138 );
and \U$7729 ( \8399 , \8397 , \8398 );
and \U$7730 ( \8400 , \1626 , RIaaa44c0_441);
nor \U$7731 ( \8401 , \8399 , \8400 );
nand \U$7732 ( \8402 , \2061 , RIaaa4448_440);
nand \U$7733 ( \8403 , \8401 , \3129 , \8402 );
not \U$7734 ( \8404 , \2052 );
not \U$7735 ( \8405 , RIaaa4538_442);
not \U$7736 ( \8406 , \8405 );
and \U$7737 ( \8407 , \8404 , \8406 );
not \U$7738 ( \8408 , RIaaa43d0_439);
nor \U$7739 ( \8409 , \8408 , \2036 );
nor \U$7740 ( \8410 , \8407 , \8409 );
and \U$7741 ( \8411 , \7174 , RIaaa4268_436);
and \U$7742 ( \8412 , \6868 , RIaaa4358_438);
and \U$7743 ( \8413 , \6871 , RIaaa42e0_437);
nor \U$7744 ( \8414 , \8412 , \8413 );
not \U$7745 ( \8415 , \8414 );
nor \U$7746 ( \8416 , \8411 , \8415 );
nand \U$7747 ( \8417 , \8410 , \8416 );
nor \U$7748 ( \8418 , \8403 , \8417 );
and \U$7749 ( \8419 , \7440 , RIaaa4970_451);
and \U$7750 ( \8420 , \1642 , RIaaa4880_449);
nor \U$7751 ( \8421 , \8419 , \8420 );
not \U$7752 ( \8422 , \1745 );
not \U$7753 ( \8423 , RIaaa48f8_450);
not \U$7754 ( \8424 , \8423 );
and \U$7755 ( \8425 , \8422 , \8424 );
and \U$7756 ( \8426 , \1832 , RIaaa4808_448);
nor \U$7757 ( \8427 , \8425 , \8426 );
nand \U$7758 ( \8428 , \8421 , \8427 );
nand \U$7759 ( \8429 , \6856 , RIaaa4790_447);
nand \U$7760 ( \8430 , \1874 , RIaaa4718_446);
not \U$7761 ( \8431 , \1735 );
nand \U$7762 ( \8432 , \8431 , RIaaa4628_444);
not \U$7763 ( \8433 , \2026 );
nand \U$7764 ( \8434 , \8433 , RIaaa46a0_445);
nand \U$7765 ( \8435 , \8429 , \8430 , \8432 , \8434 );
nor \U$7766 ( \8436 , \8428 , \8435 );
nand \U$7767 ( \8437 , \8418 , \8436 );
buf \U$7768 ( \8438 , \8437 );
buf \U$7769 ( \8439 , \8438 );
not \U$7770 ( \8440 , \8439 );
not \U$7771 ( \8441 , \8440 );
and \U$7772 ( \8442 , \6847 , \8441 );
not \U$7773 ( \8443 , \8379 );
nand \U$7774 ( \8444 , \8443 , \8367 , \8353 );
not \U$7775 ( \8445 , \8444 );
nor \U$7776 ( \8446 , \8442 , \8445 );
nand \U$7777 ( \8447 , \8396 , \8446 );
nand \U$7778 ( \8448 , \8342 , \8447 );
not \U$7779 ( \8449 , \8448 );
nand \U$7780 ( \8450 , \8332 , \8449 );
nand \U$7781 ( \8451 , \8329 , \8450 );
not \U$7782 ( \8452 , \8451 );
not \U$7783 ( \8453 , \8452 );
or \U$7784 ( \8454 , \8279 , \8453 );
not \U$7785 ( \8455 , \8278 );
nand \U$7786 ( \8456 , \8455 , \8451 );
nand \U$7787 ( \8457 , \8454 , \8456 );
nand \U$7788 ( \8458 , \8277 , \8457 );
not \U$7789 ( \8459 , \8250 );
not \U$7790 ( \8460 , \8093 );
and \U$7791 ( \8461 , \8459 , \8460 );
and \U$7792 ( \8462 , \8250 , \8093 );
nor \U$7793 ( \8463 , \8461 , \8462 );
nand \U$7794 ( \8464 , \8451 , \8278 );
and \U$7795 ( \8465 , \8458 , \8463 , \8464 );
xnor \U$7796 ( \8466 , \8276 , \8457 );
xor \U$7797 ( \8467 , \8448 , \8323 );
xnor \U$7798 ( \8468 , \8467 , \8326 );
not \U$7799 ( \8469 , \8468 );
not \U$7800 ( \8470 , \8469 );
not \U$7801 ( \8471 , \8352 );
not \U$7802 ( \8472 , \8367 );
or \U$7803 ( \8473 , \8471 , \8472 );
or \U$7804 ( \8474 , \8367 , \8352 );
nand \U$7805 ( \8475 , \8473 , \8474 );
not \U$7806 ( \8476 , \8475 );
buf \U$7807 ( \8477 , \8126 );
buf \U$7808 ( \8478 , \7263 );
and \U$7809 ( \8479 , \8477 , \8478 );
not \U$7810 ( \8480 , \8131 );
not \U$7811 ( \8481 , \7037 );
or \U$7812 ( \8482 , \8480 , \8481 );
or \U$7813 ( \8483 , \8360 , \7038 );
nand \U$7814 ( \8484 , \8482 , \8483 );
nor \U$7815 ( \8485 , \8479 , \8484 );
nand \U$7816 ( \8486 , \8122 , \7264 );
nand \U$7817 ( \8487 , \8485 , \8486 );
not \U$7818 ( \8488 , \8348 );
not \U$7819 ( \8489 , \6974 );
or \U$7820 ( \8490 , \8488 , \8489 );
and \U$7821 ( \8491 , \7882 , \8346 );
and \U$7822 ( \8492 , \7568 , \8491 );
and \U$7823 ( \8493 , \8108 , \8346 );
and \U$7824 ( \8494 , \6893 , \8493 );
nor \U$7825 ( \8495 , \8492 , \8494 );
nand \U$7826 ( \8496 , \8490 , \8495 );
nand \U$7827 ( \8497 , \8487 , \8496 );
not \U$7828 ( \8498 , \8497 );
not \U$7829 ( \8499 , \7308 );
not \U$7830 ( \8500 , \7577 );
or \U$7831 ( \8501 , \8499 , \8500 );
buf \U$7832 ( \8502 , \7863 );
and \U$7833 ( \8503 , \8502 , \7585 );
not \U$7834 ( \8504 , \7264 );
not \U$7835 ( \8505 , \7856 );
or \U$7836 ( \8506 , \8504 , \8505 );
not \U$7837 ( \8507 , \7559 );
nand \U$7838 ( \8508 , \8507 , \8478 );
nand \U$7839 ( \8509 , \8506 , \8508 );
nor \U$7840 ( \8510 , \8503 , \8509 );
nand \U$7841 ( \8511 , \8501 , \8510 );
not \U$7842 ( \8512 , \8511 );
or \U$7843 ( \8513 , \8498 , \8512 );
not \U$7844 ( \8514 , \8511 );
not \U$7845 ( \8515 , \8497 );
nand \U$7846 ( \8516 , \8514 , \8515 );
nand \U$7847 ( \8517 , \8513 , \8516 );
not \U$7848 ( \8518 , \8517 );
or \U$7849 ( \8519 , \8476 , \8518 );
not \U$7850 ( \8520 , \6846 );
not \U$7851 ( \8521 , \1735 );
not \U$7852 ( \8522 , RIaaa6860_517);
not \U$7853 ( \8523 , \8522 );
and \U$7854 ( \8524 , \8521 , \8523 );
not \U$7855 ( \8525 , RIaaa68d8_518);
nor \U$7856 ( \8526 , \8525 , \7003 );
nor \U$7857 ( \8527 , \8524 , \8526 );
not \U$7858 ( \8528 , \8527 );
not \U$7859 ( \8529 , \2066 );
not \U$7860 ( \8530 , RIaaa6950_519);
or \U$7861 ( \8531 , \8529 , \8530 );
nand \U$7862 ( \8532 , \8531 , \3204 );
and \U$7863 ( \8533 , \6862 , RIaaa6248_504);
not \U$7864 ( \8534 , RIaaa62c0_505);
not \U$7865 ( \8535 , \6871 );
or \U$7866 ( \8536 , \8534 , \8535 );
not \U$7867 ( \8537 , RIaaa6338_506);
or \U$7868 ( \8538 , \6867 , \8537 );
nand \U$7869 ( \8539 , \8536 , \8538 );
nor \U$7870 ( \8540 , \8533 , \8539 );
and \U$7871 ( \8541 , RIaaa6428_508, \2061 );
not \U$7872 ( \8542 , RIaaa63b0_507);
nor \U$7873 ( \8543 , \8542 , \6848 );
nor \U$7874 ( \8544 , \8541 , \8543 );
nand \U$7875 ( \8545 , \8540 , \8544 );
nor \U$7876 ( \8546 , \8528 , \8532 , \8545 );
nand \U$7877 ( \8547 , \1832 , RIaaa6680_513);
nand \U$7878 ( \8548 , \1642 , RIaaa6608_512);
nand \U$7879 ( \8549 , \1755 , RIaaa6518_510);
nand \U$7880 ( \8550 , \1640 , RIaaa66f8_514);
nand \U$7881 ( \8551 , \8547 , \8548 , \8549 , \8550 );
and \U$7882 ( \8552 , \7184 , RIaaa6770_515);
not \U$7883 ( \8553 , RIaaa6590_511);
nor \U$7884 ( \8554 , \8553 , \2052 );
nor \U$7885 ( \8555 , \8552 , \8554 );
and \U$7886 ( \8556 , \1626 , RIaaa64a0_509);
and \U$7887 ( \8557 , \1651 , RIaaa67e8_516);
nor \U$7888 ( \8558 , \8556 , \8557 );
nand \U$7889 ( \8559 , \8555 , \8558 );
nor \U$7890 ( \8560 , \8551 , \8559 );
nand \U$7891 ( \8561 , \8546 , \8560 );
not \U$7892 ( \8562 , \8561 );
not \U$7893 ( \8563 , \8562 );
buf \U$7894 ( \8564 , \8563 );
not \U$7895 ( \8565 , \8564 );
not \U$7896 ( \8566 , \8565 );
and \U$7897 ( \8567 , \8520 , \8566 );
and \U$7898 ( \8568 , \8511 , \8515 );
nor \U$7899 ( \8569 , \8567 , \8568 );
nand \U$7900 ( \8570 , \8519 , \8569 );
not \U$7901 ( \8571 , \8441 );
and \U$7902 ( \8572 , \6921 , \6989 );
not \U$7903 ( \8573 , \8572 );
or \U$7904 ( \8574 , \8571 , \8573 );
not \U$7905 ( \8575 , \8441 );
and \U$7906 ( \8576 , \6985 , \8575 );
and \U$7907 ( \8577 , \8233 , \7079 );
not \U$7908 ( \8578 , \8233 );
and \U$7909 ( \8579 , \8578 , \6992 );
nor \U$7910 ( \8580 , \8577 , \8579 );
nor \U$7911 ( \8581 , \8576 , \8580 );
nand \U$7912 ( \8582 , \8574 , \8581 );
and \U$7913 ( \8583 , \8570 , \8582 );
nand \U$7914 ( \8584 , \8380 , \8444 );
xor \U$7915 ( \8585 , \8393 , \8584 );
not \U$7916 ( \8586 , \7466 );
not \U$7917 ( \8587 , \7639 );
or \U$7918 ( \8588 , \8586 , \8587 );
and \U$7919 ( \8589 , \7206 , \7378 );
not \U$7920 ( \8590 , \7206 );
and \U$7921 ( \8591 , \8590 , \7741 );
nor \U$7922 ( \8592 , \8589 , \8591 );
nor \U$7923 ( \8593 , \7466 , \7733 );
nor \U$7924 ( \8594 , \8592 , \8593 );
nand \U$7925 ( \8595 , \8588 , \8594 );
not \U$7926 ( \8596 , \8232 );
not \U$7927 ( \8597 , \7389 );
or \U$7928 ( \8598 , \8596 , \8597 );
and \U$7929 ( \8599 , \7101 , \8233 );
and \U$7930 ( \8600 , \7961 , \7106 );
not \U$7931 ( \8601 , \7961 );
buf \U$7932 ( \8602 , \7069 );
and \U$7933 ( \8603 , \8601 , \8602 );
nor \U$7934 ( \8604 , \8600 , \8603 );
nor \U$7935 ( \8605 , \8599 , \8604 );
nand \U$7936 ( \8606 , \8598 , \8605 );
xor \U$7937 ( \8607 , \8595 , \8606 );
not \U$7938 ( \8608 , \7710 );
not \U$7939 ( \8609 , \7971 );
or \U$7940 ( \8610 , \8608 , \8609 );
not \U$7941 ( \8611 , \7161 );
not \U$7942 ( \8612 , \8012 );
or \U$7943 ( \8613 , \8611 , \8612 );
or \U$7944 ( \8614 , \8039 , \8050 );
nand \U$7945 ( \8615 , \8613 , \8614 );
nor \U$7946 ( \8616 , \7337 , \7710 );
nor \U$7947 ( \8617 , \8615 , \8616 );
nand \U$7948 ( \8618 , \8610 , \8617 );
and \U$7949 ( \8619 , \8607 , \8618 );
and \U$7950 ( \8620 , \8595 , \8606 );
or \U$7951 ( \8621 , \8619 , \8620 );
xor \U$7952 ( \8622 , \8585 , \8621 );
xor \U$7953 ( \8623 , \8290 , \8313 );
and \U$7954 ( \8624 , \8622 , \8623 );
and \U$7955 ( \8625 , \8585 , \8621 );
or \U$7956 ( \8626 , \8624 , \8625 );
xor \U$7957 ( \8627 , \8583 , \8626 );
xor \U$7958 ( \8628 , \8447 , \8342 );
and \U$7959 ( \8629 , \8627 , \8628 );
and \U$7960 ( \8630 , \8583 , \8626 );
nor \U$7961 ( \8631 , \8629 , \8630 );
not \U$7962 ( \8632 , \8631 );
not \U$7963 ( \8633 , \8095 );
not \U$7964 ( \8634 , \8176 );
or \U$7965 ( \8635 , \8633 , \8634 );
or \U$7966 ( \8636 , \8176 , \8095 );
nand \U$7967 ( \8637 , \8635 , \8636 );
not \U$7968 ( \8638 , \8637 );
or \U$7969 ( \8639 , \8632 , \8638 );
or \U$7970 ( \8640 , \8631 , \8637 );
nand \U$7971 ( \8641 , \8639 , \8640 );
not \U$7972 ( \8642 , \8641 );
or \U$7973 ( \8643 , \8470 , \8642 );
not \U$7974 ( \8644 , \8631 );
nand \U$7975 ( \8645 , \8644 , \8637 );
nand \U$7976 ( \8646 , \8643 , \8645 );
nand \U$7977 ( \8647 , \8466 , \8646 );
or \U$7978 ( \8648 , \8465 , \8647 );
not \U$7979 ( \8649 , \8464 );
not \U$7980 ( \8650 , \8458 );
or \U$7981 ( \8651 , \8649 , \8650 );
not \U$7982 ( \8652 , \8463 );
nand \U$7983 ( \8653 , \8651 , \8652 );
nand \U$7984 ( \8654 , \8648 , \8653 );
and \U$7985 ( \8655 , \8270 , \8654 );
not \U$7986 ( \8656 , \8269 );
not \U$7987 ( \8657 , \8251 );
or \U$7988 ( \8658 , \8656 , \8657 );
not \U$7989 ( \8659 , \8267 );
nand \U$7990 ( \8660 , \8658 , \8659 );
not \U$7991 ( \8661 , \8265 );
and \U$7992 ( \8662 , \8661 , \8252 );
not \U$7993 ( \8663 , \8259 );
nor \U$7994 ( \8664 , \8663 , \8261 );
nor \U$7995 ( \8665 , \8662 , \8664 );
not \U$7996 ( \8666 , \7657 );
and \U$7997 ( \8667 , \7817 , \8666 );
not \U$7998 ( \8668 , \7817 );
and \U$7999 ( \8669 , \8668 , \7657 );
nor \U$8000 ( \8670 , \8667 , \8669 );
nand \U$8001 ( \8671 , \8665 , \8670 );
nand \U$8002 ( \8672 , \8660 , \8671 );
nor \U$8003 ( \8673 , \8655 , \8672 );
or \U$8004 ( \8674 , \8665 , \8670 );
not \U$8005 ( \8675 , \8674 );
nor \U$8006 ( \8676 , \8673 , \8675 );
not \U$8007 ( \8677 , \8676 );
or \U$8008 ( \8678 , \7854 , \8677 );
not \U$8009 ( \8679 , \7851 );
nor \U$8010 ( \8680 , \7821 , \7841 );
not \U$8011 ( \8681 , \8680 );
or \U$8012 ( \8682 , \8679 , \8681 );
or \U$8013 ( \8683 , \7844 , \7850 );
nand \U$8014 ( \8684 , \8682 , \8683 );
not \U$8015 ( \8685 , \7503 );
nor \U$8016 ( \8686 , \7535 , \8685 );
or \U$8017 ( \8687 , \8684 , \8686 );
nand \U$8018 ( \8688 , \7535 , \8685 );
nand \U$8019 ( \8689 , \8687 , \8688 );
xor \U$8020 ( \8690 , \7509 , \7512 );
not \U$8021 ( \8691 , \7533 );
and \U$8022 ( \8692 , \8690 , \8691 );
and \U$8023 ( \8693 , \7509 , \7512 );
or \U$8024 ( \8694 , \8692 , \8693 );
not \U$8025 ( \8695 , \8694 );
xor \U$8026 ( \8696 , \7087 , \7072 );
xor \U$8027 ( \8697 , \7532 , \8696 );
nand \U$8028 ( \8698 , \8695 , \8697 );
and \U$8029 ( \8699 , \8689 , \8698 );
nand \U$8030 ( \8700 , \8678 , \8699 );
not \U$8031 ( \8701 , \8700 );
nor \U$8032 ( \8702 , \8695 , \8697 );
not \U$8033 ( \8703 , \8702 );
not \U$8034 ( \8704 , \8703 );
or \U$8035 ( \8705 , \8701 , \8704 );
not \U$8036 ( \8706 , RIaaa5f78_498);
nor \U$8037 ( \8707 , \8706 , \7409 );
not \U$8038 ( \8708 , \8707 );
nor \U$8039 ( \8709 , \7003 , \4179 );
not \U$8040 ( \8710 , \8709 );
nand \U$8041 ( \8711 , \2061 , RIaaa5c30_491);
nand \U$8042 ( \8712 , \8708 , \8710 , \4172 , \8711 );
not \U$8043 ( \8713 , \2063 );
not \U$8044 ( \8714 , \4144 );
and \U$8045 ( \8715 , \8713 , \8714 );
and \U$8046 ( \8716 , \7174 , RIaaa5e10_495);
nor \U$8047 ( \8717 , \8715 , \8716 );
not \U$8048 ( \8718 , RIaaa5bb8_490);
nor \U$8049 ( \8719 , \8718 , \6848 );
not \U$8050 ( \8720 , RIaaa5a50_487);
nor \U$8051 ( \8721 , \8720 , \2026 );
nor \U$8052 ( \8722 , \8719 , \8721 );
nand \U$8053 ( \8723 , \8717 , \8722 );
nor \U$8054 ( \8724 , \8712 , \8723 );
not \U$8055 ( \8725 , \1832 );
nor \U$8056 ( \8726 , \8725 , \4148 );
not \U$8057 ( \8727 , RIaaa6158_502);
nor \U$8058 ( \8728 , \8727 , \1743 );
nor \U$8059 ( \8729 , \8726 , \8728 );
and \U$8060 ( \8730 , \6883 , RIaaa5ca8_492);
and \U$8061 ( \8731 , RIaaa5e88_496, \6871 );
and \U$8062 ( \8732 , \6868 , RIaaa5f00_497);
nor \U$8063 ( \8733 , \8730 , \8731 , \8732 );
nand \U$8064 ( \8734 , \8729 , \8733 );
not \U$8065 ( \8735 , RIaaa6068_500);
nor \U$8066 ( \8736 , \8735 , \7432 );
not \U$8067 ( \8737 , \8736 );
not \U$8068 ( \8738 , \7185 );
nand \U$8069 ( \8739 , \8738 , RIaaa5d20_493);
not \U$8070 ( \8740 , \2014 );
not \U$8071 ( \8741 , RIaaa5ac8_488);
not \U$8072 ( \8742 , \8741 );
and \U$8073 ( \8743 , \8740 , \8742 );
and \U$8074 ( \8744 , \2023 , RIaaa5b40_489);
nor \U$8075 ( \8745 , \8743 , \8744 );
nand \U$8076 ( \8746 , \8737 , \8739 , \8745 );
nor \U$8077 ( \8747 , \8734 , \8746 );
nand \U$8078 ( \8748 , \8724 , \8747 );
not \U$8079 ( \8749 , \8748 );
buf \U$8080 ( \8750 , \8749 );
not \U$8081 ( \8751 , \8750 );
not \U$8082 ( \8752 , \8751 );
and \U$8083 ( \8753 , \6986 , \8752 );
not \U$8084 ( \8754 , RIaaa4e98_462);
nor \U$8085 ( \8755 , \8754 , \2063 );
not \U$8086 ( \8756 , RIaaa4d30_459);
nor \U$8087 ( \8757 , \8756 , \7415 );
nor \U$8088 ( \8758 , \8755 , \8757 );
nand \U$8089 ( \8759 , \2061 , RIaaa5078_466);
nand \U$8090 ( \8760 , \8758 , \3901 , \8759 );
not \U$8091 ( \8761 , \6848 );
not \U$8092 ( \8762 , RIaaa5000_465);
not \U$8093 ( \8763 , \8762 );
and \U$8094 ( \8764 , \8761 , \8763 );
and \U$8095 ( \8765 , \1622 , RIaaa4cb8_458);
nor \U$8096 ( \8766 , \8764 , \8765 );
not \U$8097 ( \8767 , \1852 );
not \U$8098 ( \8768 , RIaaa4b50_455);
not \U$8099 ( \8769 , \8768 );
and \U$8100 ( \8770 , \8767 , \8769 );
not \U$8101 ( \8771 , RIaaa4e20_461);
nor \U$8102 ( \8772 , \2026 , \8771 );
nor \U$8103 ( \8773 , \8770 , \8772 );
nand \U$8104 ( \8774 , \8766 , \8773 );
nor \U$8105 ( \8775 , \8760 , \8774 );
not \U$8106 ( \8776 , \6882 );
not \U$8107 ( \8777 , \3879 );
and \U$8108 ( \8778 , \8776 , \8777 );
and \U$8109 ( \8779 , \6868 , RIaaa4c40_457);
and \U$8110 ( \8780 , \6871 , RIaaa4bc8_456);
nor \U$8111 ( \8781 , \8779 , \8780 );
not \U$8112 ( \8782 , \8781 );
nor \U$8113 ( \8783 , \8778 , \8782 );
nand \U$8114 ( \8784 , \1832 , RIaaa50f0_467);
nand \U$8115 ( \8785 , \1642 , RIaaa5168_468);
nand \U$8116 ( \8786 , \8783 , \8784 , \8785 );
not \U$8117 ( \8787 , RIaaa4f10_463);
nor \U$8118 ( \8788 , \8787 , \2014 );
not \U$8119 ( \8789 , \8788 );
not \U$8120 ( \8790 , \2020 );
nand \U$8121 ( \8791 , \8790 , RIaaa4a60_453);
not \U$8122 ( \8792 , \7432 );
not \U$8123 ( \8793 , RIaaa4da8_460);
not \U$8124 ( \8794 , \8793 );
and \U$8125 ( \8795 , \8792 , \8794 );
and \U$8126 ( \8796 , \1626 , RIaaa4f88_464);
nor \U$8127 ( \8797 , \8795 , \8796 );
nand \U$8128 ( \8798 , \8789 , \8791 , \8797 );
nor \U$8129 ( \8799 , \8786 , \8798 );
nand \U$8130 ( \8800 , \8775 , \8799 );
not \U$8131 ( \8801 , \8800 );
not \U$8132 ( \8802 , \8801 );
buf \U$8133 ( \8803 , \8802 );
not \U$8134 ( \8804 , \8803 );
or \U$8135 ( \8805 , \7080 , \8804 );
nand \U$8136 ( \8806 , \8183 , \8804 );
nand \U$8137 ( \8807 , \8805 , \8806 );
nor \U$8138 ( \8808 , \8753 , \8807 );
nand \U$8139 ( \8809 , \8572 , \8751 );
nand \U$8140 ( \8810 , \8808 , \8809 );
not \U$8141 ( \8811 , \8126 );
not \U$8142 ( \8812 , \7465 );
or \U$8143 ( \8813 , \8811 , \8812 );
nand \U$8144 ( \8814 , \8122 , \8812 );
and \U$8145 ( \8815 , \7205 , \8131 );
not \U$8146 ( \8816 , \7205 );
and \U$8147 ( \8817 , \8816 , \8361 );
nor \U$8148 ( \8818 , \8815 , \8817 );
nand \U$8149 ( \8819 , \8813 , \8814 , \8818 );
buf \U$8150 ( \8820 , \8819 );
not \U$8151 ( \8821 , \8820 );
not \U$8152 ( \8822 , \8493 );
not \U$8153 ( \8823 , \7264 );
or \U$8154 ( \8824 , \8822 , \8823 );
and \U$8155 ( \8825 , \7307 , \8348 );
and \U$8156 ( \8826 , \7263 , \8491 );
nor \U$8157 ( \8827 , \8825 , \8826 );
nand \U$8158 ( \8828 , \8824 , \8827 );
not \U$8159 ( \8829 , \8828 );
not \U$8160 ( \8830 , \8829 );
and \U$8161 ( \8831 , \8821 , \8830 );
and \U$8162 ( \8832 , \8820 , \8829 );
nor \U$8163 ( \8833 , \8831 , \8832 );
not \U$8164 ( \8834 , \8833 );
not \U$8165 ( \8835 , \8834 );
not \U$8166 ( \8836 , \8039 );
not \U$8167 ( \8837 , \7577 );
or \U$8168 ( \8838 , \8836 , \8837 );
and \U$8169 ( \8839 , \8502 , \8013 );
and \U$8170 ( \8840 , \7709 , \7856 );
not \U$8171 ( \8841 , \7709 );
and \U$8172 ( \8842 , \8841 , \7887 );
or \U$8173 ( \8843 , \8840 , \8842 );
nor \U$8174 ( \8844 , \8839 , \8843 );
nand \U$8175 ( \8845 , \8838 , \8844 );
not \U$8176 ( \8846 , \8845 );
and \U$8177 ( \8847 , \7205 , \8348 );
and \U$8178 ( \8848 , \7307 , \8491 );
nor \U$8179 ( \8849 , \8847 , \8848 );
nand \U$8180 ( \8850 , \7306 , \8493 );
and \U$8181 ( \8851 , \8849 , \8850 );
not \U$8182 ( \8852 , \8851 );
or \U$8183 ( \8853 , \8362 , \7465 );
nand \U$8184 ( \8854 , \8131 , \7465 );
nand \U$8185 ( \8855 , \8853 , \8854 );
not \U$8186 ( \8856 , \8855 );
not \U$8187 ( \8857 , \7709 );
nand \U$8188 ( \8858 , \8857 , \8127 );
nand \U$8189 ( \8859 , \7709 , \8122 );
nand \U$8190 ( \8860 , \8856 , \8858 , \8859 );
nand \U$8191 ( \8861 , \8852 , \8860 );
not \U$8192 ( \8862 , \8861 );
or \U$8193 ( \8863 , \8846 , \8862 );
or \U$8194 ( \8864 , \8845 , \8861 );
nand \U$8195 ( \8865 , \8863 , \8864 );
not \U$8196 ( \8866 , \8865 );
or \U$8197 ( \8867 , \8835 , \8866 );
not \U$8198 ( \8868 , \6846 );
and \U$8199 ( \8869 , \1832 , RIaaa6d88_528);
and \U$8200 ( \8870 , \1642 , RIaaa6e00_529);
nor \U$8201 ( \8871 , \8869 , \8870 );
not \U$8202 ( \8872 , \2068 );
not \U$8203 ( \8873 , \4324 );
and \U$8204 ( \8874 , \8872 , \8873 );
not \U$8205 ( \8875 , RIaaa6ba8_524);
nor \U$8206 ( \8876 , \8875 , \7692 );
nor \U$8207 ( \8877 , \8874 , \8876 );
nand \U$8208 ( \8878 , \7014 , RIaaa6d10_527);
nand \U$8209 ( \8879 , \8871 , \8877 , \8878 );
and \U$8210 ( \8880 , \1651 , RIaaa6ab8_522);
and \U$8211 ( \8881 , \8202 , RIaaa6c20_525);
nor \U$8212 ( \8882 , \8880 , \8881 );
and \U$8213 ( \8883 , \1846 , RIaaa6e78_530);
and \U$8214 ( \8884 , \8431 , RIaaa6b30_523);
nor \U$8215 ( \8885 , \8883 , \8884 );
nand \U$8216 ( \8886 , \8882 , \8885 );
nor \U$8217 ( \8887 , \8879 , \8886 );
not \U$8218 ( \8888 , \1852 );
not \U$8219 ( \8889 , RIaaa6fe0_533);
not \U$8220 ( \8890 , \8889 );
and \U$8221 ( \8891 , \8888 , \8890 );
and \U$8222 ( \8892 , \7666 , RIaaa6f68_532);
nor \U$8223 ( \8893 , \8891 , \8892 );
and \U$8224 ( \8894 , \2023 , RIaaa69c8_520);
and \U$8225 ( \8895 , \6889 , RIaaa6a40_521);
nor \U$8226 ( \8896 , \8894 , \8895 );
nand \U$8227 ( \8897 , \8893 , \8896 );
and \U$8228 ( \8898 , \6883 , RIaaa6ef0_531);
not \U$8229 ( \8899 , RIaaa7058_534);
not \U$8230 ( \8900 , \6871 );
or \U$8231 ( \8901 , \8899 , \8900 );
or \U$8232 ( \8902 , \6867 , \4334 );
nand \U$8233 ( \8903 , \8901 , \8902 );
nor \U$8234 ( \8904 , \8898 , \8903 );
nand \U$8235 ( \8905 , \8904 , \4315 );
nor \U$8236 ( \8906 , \8897 , \8905 );
nand \U$8237 ( \8907 , \8887 , \8906 );
not \U$8238 ( \8908 , \8907 );
not \U$8239 ( \8909 , \8908 );
not \U$8240 ( \8910 , \8909 );
not \U$8241 ( \8911 , \8910 );
and \U$8242 ( \8912 , \8868 , \8911 );
not \U$8243 ( \8913 , \8861 );
and \U$8244 ( \8914 , \8845 , \8913 );
nor \U$8245 ( \8915 , \8912 , \8914 );
nand \U$8246 ( \8916 , \8867 , \8915 );
nand \U$8247 ( \8917 , \8810 , \8916 );
not \U$8248 ( \8918 , \8804 );
and \U$8249 ( \8919 , \6990 , \8918 );
not \U$8250 ( \8920 , \6985 );
not \U$8251 ( \8921 , \8804 );
or \U$8252 ( \8922 , \8920 , \8921 );
not \U$8253 ( \8923 , \1832 );
not \U$8254 ( \8924 , \8923 );
not \U$8255 ( \8925 , RIaaa5708_480);
not \U$8256 ( \8926 , \8925 );
and \U$8257 ( \8927 , \8924 , \8926 );
and \U$8258 ( \8928 , \1642 , RIaaa5780_481);
nor \U$8259 ( \8929 , \8927 , \8928 );
not \U$8260 ( \8930 , \1745 );
not \U$8261 ( \8931 , RIaaa57f8_482);
not \U$8262 ( \8932 , \8931 );
and \U$8263 ( \8933 , \8930 , \8932 );
and \U$8264 ( \8934 , \7666 , RIaaa5870_483);
nor \U$8265 ( \8935 , \8933 , \8934 );
not \U$8266 ( \8936 , \2068 );
not \U$8267 ( \8937 , RIaaa5960_485);
not \U$8268 ( \8938 , \8937 );
and \U$8269 ( \8939 , \8936 , \8938 );
and \U$8270 ( \8940 , \8431 , RIaaa5618_478);
nor \U$8271 ( \8941 , \8939 , \8940 );
not \U$8272 ( \8942 , \7013 );
not \U$8273 ( \8943 , RIaaa58e8_484);
not \U$8274 ( \8944 , \8943 );
and \U$8275 ( \8945 , \8942 , \8944 );
and \U$8276 ( \8946 , \1651 , RIaaa5690_479);
nor \U$8277 ( \8947 , \8945 , \8946 );
nand \U$8278 ( \8948 , \8929 , \8935 , \8941 , \8947 );
not \U$8279 ( \8949 , RIaaa5348_472);
nor \U$8280 ( \8950 , \8949 , \1871 );
nor \U$8281 ( \8951 , \3671 , \8950 );
not \U$8282 ( \8952 , \6888 );
not \U$8283 ( \8953 , RIaaa5438_474);
not \U$8284 ( \8954 , \8953 );
and \U$8285 ( \8955 , \8952 , \8954 );
and \U$8286 ( \8956 , \2023 , RIaaa52d0_471);
nor \U$8287 ( \8957 , \8955 , \8956 );
not \U$8288 ( \8958 , \1852 );
not \U$8289 ( \8959 , \3643 );
and \U$8290 ( \8960 , \8958 , \8959 );
and \U$8291 ( \8961 , \1861 , RIaaa5258_470);
nor \U$8292 ( \8962 , \8960 , \8961 );
and \U$8293 ( \8963 , \1846 , RIaaa53c0_473);
and \U$8294 ( \8964 , \6868 , RIaaa5528_476);
and \U$8295 ( \8965 , \6871 , RIaaa55a0_477);
nor \U$8296 ( \8966 , \8963 , \8964 , \8965 );
nand \U$8297 ( \8967 , \8951 , \8957 , \8962 , \8966 );
nor \U$8298 ( \8968 , \8948 , \8967 );
buf \U$8299 ( \8969 , \8968 );
not \U$8300 ( \8970 , \8969 );
not \U$8301 ( \8971 , \7079 );
and \U$8302 ( \8972 , \8970 , \8971 );
not \U$8303 ( \8973 , \8970 );
and \U$8304 ( \8974 , \8973 , \8183 );
nor \U$8305 ( \8975 , \8972 , \8974 );
nand \U$8306 ( \8976 , \8922 , \8975 );
nor \U$8307 ( \8977 , \8919 , \8976 );
not \U$8308 ( \8978 , \8977 );
and \U$8309 ( \8979 , \8502 , \7711 );
and \U$8310 ( \8980 , \7465 , \7887 );
not \U$8311 ( \8981 , \7465 );
and \U$8312 ( \8982 , \8981 , \7856 );
or \U$8313 ( \8983 , \8980 , \8982 );
nor \U$8314 ( \8984 , \8979 , \8983 );
nand \U$8315 ( \8985 , \8819 , \8828 );
nand \U$8316 ( \8986 , \7577 , \7710 );
nand \U$8317 ( \8987 , \8984 , \8985 , \8986 );
not \U$8318 ( \8988 , \8987 );
not \U$8319 ( \8989 , \8985 );
nand \U$8320 ( \8990 , \8986 , \8984 );
nand \U$8321 ( \8991 , \8989 , \8990 );
not \U$8322 ( \8992 , \7207 );
buf \U$8323 ( \8993 , \8122 );
not \U$8324 ( \8994 , \8993 );
or \U$8325 ( \8995 , \8992 , \8994 );
and \U$8326 ( \8996 , \8477 , \7206 );
not \U$8327 ( \8997 , \8131 );
not \U$8328 ( \8998 , \7307 );
or \U$8329 ( \8999 , \8997 , \8998 );
or \U$8330 ( \9000 , \8362 , \7307 );
nand \U$8331 ( \9001 , \8999 , \9000 );
nor \U$8332 ( \9002 , \8996 , \9001 );
nand \U$8333 ( \9003 , \8995 , \9002 );
not \U$8334 ( \9004 , \9003 );
and \U$8335 ( \9005 , \7037 , \8491 );
not \U$8336 ( \9006 , \7037 );
and \U$8337 ( \9007 , \9006 , \8493 );
nor \U$8338 ( \9008 , \9005 , \9007 );
nand \U$8339 ( \9009 , \7263 , \8348 );
and \U$8340 ( \9010 , \9008 , \9009 );
not \U$8341 ( \9011 , \9010 );
and \U$8342 ( \9012 , \9004 , \9011 );
and \U$8343 ( \9013 , \9003 , \9010 );
nor \U$8344 ( \9014 , \9012 , \9013 );
nand \U$8345 ( \9015 , \8991 , \9014 );
not \U$8346 ( \9016 , \9015 );
or \U$8347 ( \9017 , \8988 , \9016 );
nand \U$8348 ( \9018 , \6847 , \8751 );
nand \U$8349 ( \9019 , \9017 , \9018 );
not \U$8350 ( \9020 , \9019 );
and \U$8351 ( \9021 , \8978 , \9020 );
and \U$8352 ( \9022 , \8977 , \9019 );
nor \U$8353 ( \9023 , \9021 , \9022 );
xor \U$8354 ( \9024 , \8917 , \9023 );
not \U$8355 ( \9025 , \8230 );
not \U$8356 ( \9026 , \7639 );
or \U$8357 ( \9027 , \9025 , \9026 );
or \U$8358 ( \9028 , \7961 , \7378 );
nand \U$8359 ( \9029 , \7740 , \7961 );
nand \U$8360 ( \9030 , \9028 , \9029 );
nor \U$8361 ( \9031 , \7733 , \8232 );
nor \U$8362 ( \9032 , \9030 , \9031 );
nand \U$8363 ( \9033 , \9027 , \9032 );
not \U$8364 ( \9034 , \8804 );
not \U$8365 ( \9035 , \7388 );
or \U$8366 ( \9036 , \9034 , \9035 );
not \U$8367 ( \9037 , \6915 );
nor \U$8368 ( \9038 , \9037 , \7387 );
not \U$8369 ( \9039 , \8803 );
not \U$8370 ( \9040 , \9039 );
and \U$8371 ( \9041 , \9038 , \9040 );
not \U$8372 ( \9042 , \8968 );
buf \U$8373 ( \9043 , \9042 );
or \U$8374 ( \9044 , \7069 , \9043 );
nand \U$8375 ( \9045 , \7107 , \9043 );
nand \U$8376 ( \9046 , \9044 , \9045 );
nor \U$8377 ( \9047 , \9041 , \9046 );
nand \U$8378 ( \9048 , \9036 , \9047 );
xor \U$8379 ( \9049 , \9033 , \9048 );
not \U$8380 ( \9050 , \8564 );
or \U$8381 ( \9051 , \7153 , \9050 );
or \U$8382 ( \9052 , \7152 , \8564 );
nand \U$8383 ( \9053 , \9051 , \9052 );
not \U$8384 ( \9054 , \9053 );
not \U$8385 ( \9055 , \7622 );
or \U$8386 ( \9056 , \9054 , \9055 );
and \U$8387 ( \9057 , \8441 , \7336 );
not \U$8388 ( \9058 , \8441 );
not \U$8389 ( \9059 , \7215 );
and \U$8390 ( \9060 , \9058 , \9059 );
nor \U$8391 ( \9061 , \9057 , \9060 );
nand \U$8392 ( \9062 , \9056 , \9061 );
and \U$8393 ( \9063 , \9049 , \9062 );
and \U$8394 ( \9064 , \9033 , \9048 );
nor \U$8395 ( \9065 , \9063 , \9064 );
not \U$8396 ( \9066 , \9065 );
nand \U$8397 ( \9067 , \8991 , \8987 );
xor \U$8398 ( \9068 , \9067 , \9014 );
not \U$8399 ( \9069 , \9068 );
not \U$8400 ( \9070 , \9069 );
and \U$8401 ( \9071 , \9066 , \9070 );
not \U$8402 ( \9072 , \9068 );
not \U$8403 ( \9073 , \9065 );
or \U$8404 ( \9074 , \9072 , \9073 );
or \U$8405 ( \9075 , \9065 , \9068 );
nand \U$8406 ( \9076 , \9074 , \9075 );
not \U$8407 ( \9077 , \7960 );
not \U$8408 ( \9078 , \8061 );
or \U$8409 ( \9079 , \9077 , \9078 );
not \U$8410 ( \9080 , \7960 );
not \U$8411 ( \9081 , \7733 );
and \U$8412 ( \9082 , \9080 , \9081 );
and \U$8413 ( \9083 , \8013 , \7741 );
not \U$8414 ( \9084 , \8013 );
and \U$8415 ( \9085 , \9084 , \7378 );
nor \U$8416 ( \9086 , \9083 , \9085 );
nor \U$8417 ( \9087 , \9082 , \9086 );
nand \U$8418 ( \9088 , \9079 , \9087 );
not \U$8419 ( \9089 , \8970 );
not \U$8420 ( \9090 , \9089 );
not \U$8421 ( \9091 , \7389 );
or \U$8422 ( \9092 , \9090 , \9091 );
and \U$8423 ( \9093 , \7101 , \8970 );
and \U$8424 ( \9094 , \8564 , \7471 );
not \U$8425 ( \9095 , \8564 );
and \U$8426 ( \9096 , \9095 , \8602 );
nor \U$8427 ( \9097 , \9094 , \9096 );
nor \U$8428 ( \9098 , \9093 , \9097 );
nand \U$8429 ( \9099 , \9092 , \9098 );
xor \U$8430 ( \9100 , \9088 , \9099 );
or \U$8431 ( \9101 , \7216 , \8233 );
nand \U$8432 ( \9102 , \7336 , \8233 );
and \U$8433 ( \9103 , \7155 , \8441 );
nor \U$8434 ( \9104 , \7341 , \8441 );
nor \U$8435 ( \9105 , \9103 , \9104 );
nand \U$8436 ( \9106 , \9101 , \9102 , \9105 );
xor \U$8437 ( \9107 , \9100 , \9106 );
and \U$8438 ( \9108 , \9076 , \9107 );
nor \U$8439 ( \9109 , \9071 , \9108 );
xor \U$8440 ( \9110 , \9024 , \9109 );
not \U$8441 ( \9111 , \9110 );
not \U$8442 ( \9112 , \8910 );
not \U$8443 ( \9113 , \9112 );
not \U$8444 ( \9114 , \6990 );
or \U$8445 ( \9115 , \9113 , \9114 );
and \U$8446 ( \9116 , \6985 , \8910 );
and \U$8447 ( \9117 , \8751 , \7080 );
not \U$8448 ( \9118 , \8751 );
and \U$8449 ( \9119 , \9118 , \6992 );
nor \U$8450 ( \9120 , \9117 , \9119 );
nor \U$8451 ( \9121 , \9116 , \9120 );
nand \U$8452 ( \9122 , \9115 , \9121 );
not \U$8453 ( \9123 , \8851 );
not \U$8454 ( \9124 , \8860 );
or \U$8455 ( \9125 , \9123 , \9124 );
or \U$8456 ( \9126 , \8860 , \8851 );
nand \U$8457 ( \9127 , \9125 , \9126 );
not \U$8458 ( \9128 , \9127 );
not \U$8459 ( \9129 , \7960 );
not \U$8460 ( \9130 , \7577 );
or \U$8461 ( \9131 , \9129 , \9130 );
and \U$8462 ( \9132 , \7865 , \7961 );
and \U$8463 ( \9133 , \8013 , \7856 );
and \U$8464 ( \9134 , \7887 , \8012 );
nor \U$8465 ( \9135 , \9132 , \9133 , \9134 );
nand \U$8466 ( \9136 , \9131 , \9135 );
not \U$8467 ( \9137 , \9136 );
or \U$8468 ( \9138 , \9128 , \9137 );
nand \U$8469 ( \9139 , \2066 , RIaaa7760_549);
nand \U$8470 ( \9140 , \2064 , RIaaa75f8_546);
nand \U$8471 ( \9141 , \1874 , RIaaa76e8_548);
nand \U$8472 ( \9142 , \4560 , \9139 , \9140 , \9141 );
nand \U$8473 ( \9143 , \6862 , RIaaa7238_538);
nand \U$8474 ( \9144 , \1861 , RIaaa73a0_541);
nand \U$8475 ( \9145 , \1872 , RIaaa7418_542);
and \U$8476 ( \9146 , \6868 , RIaaa7328_540);
and \U$8477 ( \9147 , \6871 , RIaaa72b0_539);
nor \U$8478 ( \9148 , \9146 , \9147 );
nand \U$8479 ( \9149 , \9143 , \9144 , \9145 , \9148 );
nor \U$8480 ( \9150 , \9142 , \9149 );
not \U$8481 ( \9151 , \6882 );
not \U$8482 ( \9152 , \4543 );
and \U$8483 ( \9153 , \9151 , \9152 );
and \U$8484 ( \9154 , \1832 , RIaaa77d8_550);
nor \U$8485 ( \9155 , \9153 , \9154 );
not \U$8486 ( \9156 , \2052 );
not \U$8487 ( \9157 , \4566 );
and \U$8488 ( \9158 , \9156 , \9157 );
and \U$8489 ( \9159 , \1642 , RIaaa7850_551);
nor \U$8490 ( \9160 , \9158 , \9159 );
nand \U$8491 ( \9161 , \9155 , \9160 );
and \U$8492 ( \9162 , \6876 , RIaaa7940_553);
not \U$8493 ( \9163 , RIaaa7580_545);
nor \U$8494 ( \9164 , \9163 , \2014 );
nor \U$8495 ( \9165 , \9162 , \9164 );
and \U$8496 ( \9166 , \2023 , RIaaa7490_543);
and \U$8497 ( \9167 , \1651 , RIaaa7670_547);
nor \U$8498 ( \9168 , \9166 , \9167 );
nand \U$8499 ( \9169 , \9165 , \9168 );
nor \U$8500 ( \9170 , \9161 , \9169 );
nand \U$8501 ( \9171 , \9150 , \9170 );
not \U$8502 ( \9172 , \9171 );
not \U$8503 ( \9173 , \9172 );
nand \U$8504 ( \9174 , \6847 , \9173 );
nand \U$8505 ( \9175 , \9138 , \9174 );
and \U$8506 ( \9176 , \9122 , \9175 );
not \U$8507 ( \9177 , \9176 );
xor \U$8508 ( \9178 , \9049 , \9062 );
not \U$8509 ( \9179 , \9178 );
not \U$8510 ( \9180 , \8865 );
not \U$8511 ( \9181 , \8833 );
and \U$8512 ( \9182 , \9180 , \9181 );
and \U$8513 ( \9183 , \8865 , \8833 );
nor \U$8514 ( \9184 , \9182 , \9183 );
not \U$8515 ( \9185 , \9184 );
not \U$8516 ( \9186 , \8752 );
not \U$8517 ( \9187 , \7389 );
or \U$8518 ( \9188 , \9186 , \9187 );
and \U$8519 ( \9189 , \9038 , \8751 );
or \U$8520 ( \9190 , \8602 , \9040 );
not \U$8521 ( \9191 , \9039 );
nand \U$8522 ( \9192 , \9191 , \7107 );
nand \U$8523 ( \9193 , \9190 , \9192 );
nor \U$8524 ( \9194 , \9189 , \9193 );
nand \U$8525 ( \9195 , \9188 , \9194 );
not \U$8526 ( \9196 , \9195 );
nor \U$8527 ( \9197 , \7376 , \8441 );
not \U$8528 ( \9198 , \8441 );
not \U$8529 ( \9199 , \7640 );
or \U$8530 ( \9200 , \9198 , \9199 );
and \U$8531 ( \9201 , \7370 , \7159 );
and \U$8532 ( \9202 , \8231 , \9201 );
not \U$8533 ( \9203 , \8231 );
and \U$8534 ( \9204 , \9203 , \7790 );
nor \U$8535 ( \9205 , \9202 , \9204 );
nand \U$8536 ( \9206 , \9200 , \9205 );
nor \U$8537 ( \9207 , \9197 , \9206 );
not \U$8538 ( \9208 , \9207 );
not \U$8539 ( \9209 , \8012 );
nor \U$8540 ( \9210 , \8125 , \8120 );
not \U$8541 ( \9211 , \9210 );
or \U$8542 ( \9212 , \9209 , \9211 );
and \U$8543 ( \9213 , \7707 , \8131 );
not \U$8544 ( \9214 , \7707 );
and \U$8545 ( \9215 , \9214 , \8361 );
nor \U$8546 ( \9216 , \9213 , \9215 );
nand \U$8547 ( \9217 , \9212 , \9216 );
and \U$8548 ( \9218 , \8122 , \8011 );
nor \U$8549 ( \9219 , \9217 , \9218 );
nand \U$8550 ( \9220 , \7205 , \8491 );
nand \U$8551 ( \9221 , \7204 , \8493 );
nand \U$8552 ( \9222 , \7464 , \8348 );
nand \U$8553 ( \9223 , \9220 , \9221 , \9222 );
not \U$8554 ( \9224 , \9223 );
and \U$8555 ( \9225 , \9219 , \9224 );
not \U$8556 ( \9226 , \9219 );
and \U$8557 ( \9227 , \9226 , \9223 );
nor \U$8558 ( \9228 , \9225 , \9227 );
not \U$8559 ( \9229 , \9228 );
and \U$8560 ( \9230 , \7554 , \7562 , \7564 , \7368 );
and \U$8561 ( \9231 , \9230 , \8231 );
buf \U$8562 ( \9232 , \7958 );
nor \U$8563 ( \9233 , \7554 , \7557 );
not \U$8564 ( \9234 , \9233 );
and \U$8565 ( \9235 , \9232 , \9234 );
not \U$8566 ( \9236 , \9232 );
and \U$8567 ( \9237 , \9236 , \7558 );
nor \U$8568 ( \9238 , \9235 , \9237 );
nor \U$8569 ( \9239 , \9231 , \9238 );
and \U$8570 ( \9240 , \7554 , \7562 , \7564 , \7557 );
nand \U$8571 ( \9241 , \9240 , \8230 );
nand \U$8572 ( \9242 , \9239 , \9241 );
not \U$8573 ( \9243 , \9242 );
or \U$8574 ( \9244 , \9229 , \9243 );
or \U$8575 ( \9245 , \9217 , \9218 );
nand \U$8576 ( \9246 , \9245 , \9223 );
nand \U$8577 ( \9247 , \9244 , \9246 );
not \U$8578 ( \9248 , \9247 );
or \U$8579 ( \9249 , \9208 , \9248 );
or \U$8580 ( \9250 , \9247 , \9207 );
nand \U$8581 ( \9251 , \9249 , \9250 );
not \U$8582 ( \9252 , \9251 );
or \U$8583 ( \9253 , \9196 , \9252 );
not \U$8584 ( \9254 , \9207 );
nand \U$8585 ( \9255 , \9254 , \9247 );
nand \U$8586 ( \9256 , \9253 , \9255 );
not \U$8587 ( \9257 , \9256 );
or \U$8588 ( \9258 , \9185 , \9257 );
or \U$8589 ( \9259 , \9256 , \9184 );
nand \U$8590 ( \9260 , \9258 , \9259 );
not \U$8591 ( \9261 , \9260 );
or \U$8592 ( \9262 , \9179 , \9261 );
not \U$8593 ( \9263 , \9184 );
nand \U$8594 ( \9264 , \9263 , \9256 );
nand \U$8595 ( \9265 , \9262 , \9264 );
not \U$8596 ( \9266 , \9265 );
or \U$8597 ( \9267 , \9177 , \9266 );
nor \U$8598 ( \9268 , \8810 , \8916 );
not \U$8599 ( \9269 , \9268 );
nand \U$8600 ( \9270 , \9269 , \8917 );
nand \U$8601 ( \9271 , \9267 , \9270 );
not \U$8602 ( \9272 , \9176 );
not \U$8603 ( \9273 , \9265 );
nand \U$8604 ( \9274 , \9272 , \9273 );
nand \U$8605 ( \9275 , \9271 , \9274 );
not \U$8606 ( \9276 , \7585 );
not \U$8607 ( \9277 , \8993 );
or \U$8608 ( \9278 , \9276 , \9277 );
and \U$8609 ( \9279 , \8127 , \7308 );
or \U$8610 ( \9280 , \7264 , \8130 );
nand \U$8611 ( \9281 , \8361 , \7264 );
nand \U$8612 ( \9282 , \9280 , \9281 );
nor \U$8613 ( \9283 , \9279 , \9282 );
nand \U$8614 ( \9284 , \9278 , \9283 );
not \U$8615 ( \9285 , \8348 );
not \U$8616 ( \9286 , \7038 );
or \U$8617 ( \9287 , \9285 , \9286 );
and \U$8618 ( \9288 , \6974 , \8491 );
not \U$8619 ( \9289 , \6974 );
and \U$8620 ( \9290 , \9289 , \8493 );
nor \U$8621 ( \9291 , \9288 , \9290 );
nand \U$8622 ( \9292 , \9287 , \9291 );
xor \U$8623 ( \9293 , \9284 , \9292 );
not \U$8624 ( \9294 , \9010 );
nand \U$8625 ( \9295 , \9294 , \9003 );
not \U$8626 ( \9296 , \9295 );
and \U$8627 ( \9297 , \7865 , \7600 );
or \U$8628 ( \9298 , \7559 , \7207 );
nand \U$8629 ( \9299 , \7856 , \7207 );
nand \U$8630 ( \9300 , \9298 , \9299 );
nor \U$8631 ( \9301 , \9297 , \9300 );
nand \U$8632 ( \9302 , \7577 , \7466 );
nand \U$8633 ( \9303 , \9301 , \9302 );
not \U$8634 ( \9304 , \9303 );
or \U$8635 ( \9305 , \9296 , \9304 );
or \U$8636 ( \9306 , \9295 , \9303 );
nand \U$8637 ( \9307 , \9305 , \9306 );
xor \U$8638 ( \9308 , \9293 , \9307 );
xor \U$8639 ( \9309 , \9088 , \9099 );
and \U$8640 ( \9310 , \9309 , \9106 );
and \U$8641 ( \9311 , \9088 , \9099 );
or \U$8642 ( \9312 , \9310 , \9311 );
xor \U$8643 ( \9313 , \9308 , \9312 );
not \U$8644 ( \9314 , \9313 );
not \U$8645 ( \9315 , \8039 );
not \U$8646 ( \9316 , \8061 );
or \U$8647 ( \9317 , \9315 , \9316 );
and \U$8648 ( \9318 , \7711 , \7739 );
not \U$8649 ( \9319 , \7711 );
and \U$8650 ( \9320 , \9319 , \7378 );
nor \U$8651 ( \9321 , \9318 , \9320 );
nor \U$8652 ( \9322 , \7733 , \8012 );
nor \U$8653 ( \9323 , \9321 , \9322 );
nand \U$8654 ( \9324 , \9317 , \9323 );
and \U$8655 ( \9325 , \7102 , \8564 );
or \U$8656 ( \9326 , \7069 , \8441 );
nand \U$8657 ( \9327 , \7107 , \8441 );
nand \U$8658 ( \9328 , \9326 , \9327 );
nor \U$8659 ( \9329 , \9325 , \9328 );
nand \U$8660 ( \9330 , \7389 , \8565 );
nand \U$8661 ( \9331 , \9329 , \9330 );
xor \U$8662 ( \9332 , \9324 , \9331 );
not \U$8663 ( \9333 , \7774 );
and \U$8664 ( \9334 , \8232 , \7152 );
and \U$8665 ( \9335 , \8231 , \7153 );
nor \U$8666 ( \9336 , \9334 , \9335 );
not \U$8667 ( \9337 , \9336 );
and \U$8668 ( \9338 , \9333 , \9337 );
nor \U$8669 ( \9339 , \7960 , \7152 );
and \U$8670 ( \9340 , \7623 , \9339 );
nor \U$8671 ( \9341 , \9338 , \9340 );
not \U$8672 ( \9342 , \8233 );
not \U$8673 ( \9343 , \7622 );
or \U$8674 ( \9344 , \9342 , \9343 );
nor \U$8675 ( \9345 , \7153 , \7961 );
nand \U$8676 ( \9346 , \9344 , \9345 );
and \U$8677 ( \9347 , \9341 , \9346 , \7636 );
xor \U$8678 ( \9348 , \9332 , \9347 );
not \U$8679 ( \9349 , \9348 );
or \U$8680 ( \9350 , \9314 , \9349 );
or \U$8681 ( \9351 , \9348 , \9313 );
nand \U$8682 ( \9352 , \9350 , \9351 );
xor \U$8683 ( \9353 , \9275 , \9352 );
not \U$8684 ( \9354 , \9353 );
not \U$8685 ( \9355 , \9354 );
or \U$8686 ( \9356 , \9111 , \9355 );
not \U$8687 ( \9357 , \9110 );
nand \U$8688 ( \9358 , \9357 , \9353 );
nand \U$8689 ( \9359 , \9356 , \9358 );
xnor \U$8690 ( \9360 , \9076 , \9107 );
xor \U$8691 ( \9361 , \9127 , \9136 );
xor \U$8692 ( \9362 , \9251 , \9195 );
not \U$8693 ( \9363 , \9362 );
and \U$8694 ( \9364 , \9361 , \9363 );
not \U$8695 ( \9365 , \9361 );
and \U$8696 ( \9366 , \9365 , \9362 );
nor \U$8697 ( \9367 , \9364 , \9366 );
not \U$8698 ( \9368 , \9367 );
and \U$8699 ( \9369 , \8061 , \8565 );
not \U$8700 ( \9370 , \8564 );
not \U$8701 ( \9371 , \7640 );
or \U$8702 ( \9372 , \9370 , \9371 );
and \U$8703 ( \9373 , \8575 , \7790 );
not \U$8704 ( \9374 , \8575 );
and \U$8705 ( \9375 , \9374 , \7740 );
nor \U$8706 ( \9376 , \9373 , \9375 );
nand \U$8707 ( \9377 , \9372 , \9376 );
nor \U$8708 ( \9378 , \9369 , \9377 );
not \U$8709 ( \9379 , \9378 );
not \U$8710 ( \9380 , \7464 );
or \U$8711 ( \9381 , \9380 , \8347 );
nor \U$8712 ( \9382 , \8348 , \8493 );
nand \U$8713 ( \9383 , \9381 , \9382 );
nand \U$8714 ( \9384 , \7709 , \8348 );
or \U$8715 ( \9385 , \7464 , \8347 );
nand \U$8716 ( \9386 , \9385 , \8108 );
and \U$8717 ( \9387 , \9383 , \9384 , \9386 );
and \U$8718 ( \9388 , \8477 , \7960 );
or \U$8719 ( \9389 , \8362 , \8012 );
nand \U$8720 ( \9390 , \8131 , \8012 );
nand \U$8721 ( \9391 , \9389 , \9390 );
nor \U$8722 ( \9392 , \9388 , \9391 );
nand \U$8723 ( \9393 , \8993 , \7961 );
nand \U$8724 ( \9394 , \9392 , \9393 );
and \U$8725 ( \9395 , \9387 , \9394 );
nand \U$8726 ( \9396 , \9379 , \9395 );
not \U$8727 ( \9397 , \9396 );
and \U$8728 ( \9398 , \9368 , \9397 );
and \U$8729 ( \9399 , \9362 , \9361 );
nor \U$8730 ( \9400 , \9398 , \9399 );
and \U$8731 ( \9401 , \6990 , \9173 );
not \U$8732 ( \9402 , \9172 );
not \U$8733 ( \9403 , \6986 );
or \U$8734 ( \9404 , \9402 , \9403 );
and \U$8735 ( \9405 , \9112 , \8971 );
not \U$8736 ( \9406 , \9112 );
and \U$8737 ( \9407 , \9406 , \8183 );
nor \U$8738 ( \9408 , \9405 , \9407 );
nand \U$8739 ( \9409 , \9404 , \9408 );
nor \U$8740 ( \9410 , \9401 , \9409 );
not \U$8741 ( \9411 , \9410 );
not \U$8742 ( \9412 , \7341 );
not \U$8743 ( \9413 , \8970 );
and \U$8744 ( \9414 , \9412 , \9413 );
and \U$8745 ( \9415 , \7155 , \8970 );
nor \U$8746 ( \9416 , \9414 , \9415 );
and \U$8747 ( \9417 , \7774 , \9053 );
not \U$8748 ( \9418 , RIaaa8480_577);
nor \U$8749 ( \9419 , \9418 , \1871 );
nor \U$8750 ( \9420 , \4488 , \9419 );
and \U$8751 ( \9421 , \6862 , RIaaa8228_572);
and \U$8752 ( \9422 , \1846 , RIaaa84f8_578);
nor \U$8753 ( \9423 , \9421 , \9422 );
and \U$8754 ( \9424 , \2023 , RIaaa8408_576);
and \U$8755 ( \9425 , \8202 , RIaaa8390_575);
nor \U$8756 ( \9426 , \9424 , \9425 );
and \U$8757 ( \9427 , \6889 , RIaaa8570_579);
and \U$8758 ( \9428 , \6868 , RIaaa8318_574);
and \U$8759 ( \9429 , \6871 , RIaaa82a0_573);
nor \U$8760 ( \9430 , \9427 , \9428 , \9429 );
nand \U$8761 ( \9431 , \9420 , \9423 , \9426 , \9430 );
not \U$8762 ( \9432 , \1745 );
not \U$8763 ( \9433 , RIaaa88b8_586);
not \U$8764 ( \9434 , \9433 );
and \U$8765 ( \9435 , \9432 , \9434 );
and \U$8766 ( \9436 , \1832 , RIaaa87c8_584);
nor \U$8767 ( \9437 , \9435 , \9436 );
and \U$8768 ( \9438 , \7440 , RIaaa8930_587);
and \U$8769 ( \9439 , \1642 , RIaaa8840_585);
nor \U$8770 ( \9440 , \9438 , \9439 );
and \U$8771 ( \9441 , \2064 , RIaaa85e8_580);
and \U$8772 ( \9442 , \7014 , RIaaa8750_583);
nor \U$8773 ( \9443 , \9441 , \9442 );
and \U$8774 ( \9444 , \1651 , RIaaa8660_581);
and \U$8775 ( \9445 , \1874 , RIaaa86d8_582);
nor \U$8776 ( \9446 , \9444 , \9445 );
nand \U$8777 ( \9447 , \9437 , \9440 , \9443 , \9446 );
or \U$8778 ( \9448 , \9431 , \9447 );
buf \U$8779 ( \9449 , \9448 );
and \U$8780 ( \9450 , \6847 , \9449 );
nor \U$8781 ( \9451 , \9417 , \9450 );
nand \U$8782 ( \9452 , \9416 , \9451 );
nand \U$8783 ( \9453 , \9411 , \9452 );
nand \U$8784 ( \9454 , \9400 , \9453 );
xor \U$8785 ( \9455 , \9122 , \9175 );
and \U$8786 ( \9456 , \9454 , \9455 );
nor \U$8787 ( \9457 , \9400 , \9453 );
nor \U$8788 ( \9458 , \9456 , \9457 );
xor \U$8789 ( \9459 , \9360 , \9458 );
xor \U$8790 ( \9460 , \9176 , \9270 );
xnor \U$8791 ( \9461 , \9460 , \9273 );
and \U$8792 ( \9462 , \9459 , \9461 );
and \U$8793 ( \9463 , \9360 , \9458 );
or \U$8794 ( \9464 , \9462 , \9463 );
nand \U$8795 ( \9465 , \9359 , \9464 );
not \U$8796 ( \9466 , \9271 );
not \U$8797 ( \9467 , \9274 );
or \U$8798 ( \9468 , \9466 , \9467 );
nand \U$8799 ( \9469 , \9468 , \9352 );
not \U$8800 ( \9470 , \9469 );
nand \U$8801 ( \9471 , \9353 , \9110 );
not \U$8802 ( \9472 , \9471 );
or \U$8803 ( \9473 , \9470 , \9472 );
xor \U$8804 ( \9474 , \8917 , \9023 );
and \U$8805 ( \9475 , \9474 , \9109 );
and \U$8806 ( \9476 , \8917 , \9023 );
or \U$8807 ( \9477 , \9475 , \9476 );
nand \U$8808 ( \9478 , \7338 , \8013 );
nand \U$8809 ( \9479 , \7971 , \8039 );
and \U$8810 ( \9480 , \7155 , \7961 );
nor \U$8811 ( \9481 , \7341 , \7961 );
nor \U$8812 ( \9482 , \9480 , \9481 );
nand \U$8813 ( \9483 , \9478 , \9479 , \9482 );
not \U$8814 ( \9484 , \7710 );
not \U$8815 ( \9485 , \8061 );
or \U$8816 ( \9486 , \9484 , \9485 );
nor \U$8817 ( \9487 , \7733 , \7710 );
or \U$8818 ( \9488 , \7741 , \7466 );
or \U$8819 ( \9489 , \7378 , \7600 );
nand \U$8820 ( \9490 , \9488 , \9489 );
nor \U$8821 ( \9491 , \9487 , \9490 );
nand \U$8822 ( \9492 , \9486 , \9491 );
not \U$8823 ( \9493 , \8575 );
not \U$8824 ( \9494 , \7389 );
or \U$8825 ( \9495 , \9493 , \9494 );
and \U$8826 ( \9496 , \8441 , \7102 );
or \U$8827 ( \9497 , \7071 , \8231 );
nand \U$8828 ( \9498 , \7107 , \8233 );
nand \U$8829 ( \9499 , \9497 , \9498 );
nor \U$8830 ( \9500 , \9496 , \9499 );
nand \U$8831 ( \9501 , \9495 , \9500 );
xor \U$8832 ( \9502 , \9492 , \9501 );
xor \U$8833 ( \9503 , \9483 , \9502 );
nand \U$8834 ( \9504 , \9284 , \9292 );
xor \U$8835 ( \9505 , \8487 , \8496 );
xor \U$8836 ( \9506 , \9504 , \9505 );
or \U$8837 ( \9507 , \7585 , \7559 );
nand \U$8838 ( \9508 , \7856 , \7585 );
nand \U$8839 ( \9509 , \9507 , \9508 );
not \U$8840 ( \9510 , \9509 );
and \U$8841 ( \9511 , \7207 , \7865 );
not \U$8842 ( \9512 , \7207 );
and \U$8843 ( \9513 , \9512 , \7577 );
nor \U$8844 ( \9514 , \9511 , \9513 );
nand \U$8845 ( \9515 , \9510 , \9514 );
xnor \U$8846 ( \9516 , \9506 , \9515 );
xor \U$8847 ( \9517 , \9324 , \9331 );
and \U$8848 ( \9518 , \9517 , \9347 );
and \U$8849 ( \9519 , \9324 , \9331 );
or \U$8850 ( \9520 , \9518 , \9519 );
xor \U$8851 ( \9521 , \9516 , \9520 );
not \U$8852 ( \9522 , \9521 );
and \U$8853 ( \9523 , \9503 , \9522 );
not \U$8854 ( \9524 , \9503 );
and \U$8855 ( \9525 , \9524 , \9521 );
nor \U$8856 ( \9526 , \9523 , \9525 );
xor \U$8857 ( \9527 , \9477 , \9526 );
not \U$8858 ( \9528 , \8977 );
nand \U$8859 ( \9529 , \9528 , \9019 );
not \U$8860 ( \9530 , \8970 );
not \U$8861 ( \9531 , \6990 );
or \U$8862 ( \9532 , \9530 , \9531 );
and \U$8863 ( \9533 , \6986 , \9089 );
or \U$8864 ( \9534 , \7080 , \8565 );
nand \U$8865 ( \9535 , \8183 , \8565 );
nand \U$8866 ( \9536 , \9534 , \9535 );
nor \U$8867 ( \9537 , \9533 , \9536 );
nand \U$8868 ( \9538 , \9532 , \9537 );
not \U$8869 ( \9539 , \9293 );
not \U$8870 ( \9540 , \9307 );
or \U$8871 ( \9541 , \9539 , \9540 );
not \U$8872 ( \9542 , \6846 );
not \U$8873 ( \9543 , \8804 );
and \U$8874 ( \9544 , \9542 , \9543 );
not \U$8875 ( \9545 , \9295 );
and \U$8876 ( \9546 , \9303 , \9545 );
nor \U$8877 ( \9547 , \9544 , \9546 );
nand \U$8878 ( \9548 , \9541 , \9547 );
xnor \U$8879 ( \9549 , \9538 , \9548 );
xor \U$8880 ( \9550 , \9529 , \9549 );
or \U$8881 ( \9551 , \9308 , \9312 );
and \U$8882 ( \9552 , \9348 , \9551 );
and \U$8883 ( \9553 , \9308 , \9312 );
nor \U$8884 ( \9554 , \9552 , \9553 );
xor \U$8885 ( \9555 , \9550 , \9554 );
xor \U$8886 ( \9556 , \9527 , \9555 );
nand \U$8887 ( \9557 , \9473 , \9556 );
xor \U$8888 ( \9558 , \9360 , \9458 );
xor \U$8889 ( \9559 , \9558 , \9461 );
xor \U$8890 ( \9560 , \9260 , \9178 );
not \U$8891 ( \9561 , \9452 );
not \U$8892 ( \9562 , \9561 );
not \U$8893 ( \9563 , \9411 );
or \U$8894 ( \9564 , \9562 , \9563 );
nand \U$8895 ( \9565 , \9410 , \9452 );
nand \U$8896 ( \9566 , \9564 , \9565 );
not \U$8897 ( \9567 , \9566 );
not \U$8898 ( \9568 , \8910 );
not \U$8899 ( \9569 , \7389 );
or \U$8900 ( \9570 , \9568 , \9569 );
and \U$8901 ( \9571 , \7102 , \9112 );
or \U$8902 ( \9572 , \7071 , \8751 );
nand \U$8903 ( \9573 , \7107 , \8751 );
nand \U$8904 ( \9574 , \9572 , \9573 );
nor \U$8905 ( \9575 , \9571 , \9574 );
nand \U$8906 ( \9576 , \9570 , \9575 );
buf \U$8907 ( \9577 , \9228 );
xnor \U$8908 ( \9578 , \9242 , \9577 );
not \U$8909 ( \9579 , \9578 );
xor \U$8910 ( \9580 , \9576 , \9579 );
not \U$8911 ( \9581 , \9089 );
not \U$8912 ( \9582 , \7971 );
or \U$8913 ( \9583 , \9581 , \9582 );
and \U$8914 ( \9584 , \7336 , \8970 );
or \U$8915 ( \9585 , \7160 , \8918 );
nand \U$8916 ( \9586 , \7155 , \8918 );
nand \U$8917 ( \9587 , \9585 , \9586 );
nor \U$8918 ( \9588 , \9584 , \9587 );
nand \U$8919 ( \9589 , \9583 , \9588 );
and \U$8920 ( \9590 , \9580 , \9589 );
and \U$8921 ( \9591 , \9576 , \9579 );
nor \U$8922 ( \9592 , \9590 , \9591 );
nand \U$8923 ( \9593 , \9567 , \9592 );
not \U$8924 ( \9594 , \9593 );
xor \U$8925 ( \9595 , \9387 , \9394 );
and \U$8926 ( \9596 , \7865 , \8441 );
or \U$8927 ( \9597 , \7559 , \8231 );
nand \U$8928 ( \9598 , \7856 , \8231 );
nand \U$8929 ( \9599 , \9597 , \9598 );
nor \U$8930 ( \9600 , \9596 , \9599 );
nand \U$8931 ( \9601 , \7577 , \8575 );
nand \U$8932 ( \9602 , \9600 , \9601 );
xor \U$8933 ( \9603 , \9595 , \9602 );
not \U$8934 ( \9604 , \6918 );
or \U$8935 ( \9605 , \1745 , \4761 );
not \U$8936 ( \9606 , \1832 );
or \U$8937 ( \9607 , \9606 , \4799 );
and \U$8938 ( \9608 , \1642 , RIaaa8138_570);
and \U$8939 ( \9609 , RIaaa7df0_563, \6868 );
and \U$8940 ( \9610 , \6871 , RIaaa7e68_564);
nor \U$8941 ( \9611 , \9608 , \9609 , \9610 );
nand \U$8942 ( \9612 , \9605 , \9607 , \9611 );
not \U$8943 ( \9613 , \9612 );
not \U$8944 ( \9614 , RIaaa7fd0_567);
not \U$8945 ( \9615 , \7014 );
or \U$8946 ( \9616 , \9614 , \9615 );
nand \U$8947 ( \9617 , \9616 , \4783 );
not \U$8948 ( \9618 , \9617 );
not \U$8949 ( \9619 , \1838 );
not \U$8950 ( \9620 , \4802 );
and \U$8951 ( \9621 , \9619 , \9620 );
not \U$8952 ( \9622 , RIaaa7a30_555);
nor \U$8953 ( \9623 , \9622 , \2026 );
nor \U$8954 ( \9624 , \9621 , \9623 );
and \U$8955 ( \9625 , \6889 , RIaaa7b20_557);
and \U$8956 ( \9626 , \1861 , RIaaa7b98_558);
nor \U$8957 ( \9627 , \9625 , \9626 );
nand \U$8958 ( \9628 , \9624 , \9627 );
not \U$8959 ( \9629 , RIaaa79b8_554);
not \U$8960 ( \9630 , \2064 );
or \U$8961 ( \9631 , \9629 , \9630 );
not \U$8962 ( \9632 , RIaaa7c10_559);
not \U$8963 ( \9633 , \9632 );
nand \U$8964 ( \9634 , \9633 , \7024 );
nand \U$8965 ( \9635 , \9631 , \9634 );
nor \U$8966 ( \9636 , \9628 , \9635 );
not \U$8967 ( \9637 , RIaaa8048_568);
not \U$8968 ( \9638 , \1846 );
or \U$8969 ( \9639 , \9637 , \9638 );
nand \U$8970 ( \9640 , \6862 , RIaaa7d78_562);
nand \U$8971 ( \9641 , \9639 , \9640 );
not \U$8972 ( \9642 , RIaaa7c88_560);
not \U$8973 ( \9643 , \7184 );
or \U$8974 ( \9644 , \9642 , \9643 );
nand \U$8975 ( \9645 , \1874 , RIaaa7f58_566);
nand \U$8976 ( \9646 , \9644 , \9645 );
nor \U$8977 ( \9647 , \9641 , \9646 );
nand \U$8978 ( \9648 , \9613 , \9618 , \9636 , \9647 );
buf \U$8979 ( \9649 , \9648 );
not \U$8980 ( \9650 , \9649 );
or \U$8981 ( \9651 , \9604 , \9650 );
nand \U$8982 ( \9652 , \9651 , \6917 );
nor \U$8983 ( \9653 , \6989 , \9652 );
and \U$8984 ( \9654 , \9603 , \9653 );
and \U$8985 ( \9655 , \9595 , \9602 );
or \U$8986 ( \9656 , \9654 , \9655 );
not \U$8987 ( \9657 , \9449 );
and \U$8988 ( \9658 , \6985 , \9657 );
and \U$8989 ( \9659 , \9173 , \7079 );
not \U$8990 ( \9660 , \9173 );
and \U$8991 ( \9661 , \9660 , \6992 );
nor \U$8992 ( \9662 , \9659 , \9661 );
nor \U$8993 ( \9663 , \9658 , \9662 );
nand \U$8994 ( \9664 , \6990 , \9449 );
nand \U$8995 ( \9665 , \9663 , \9664 );
xor \U$8996 ( \9666 , \9656 , \9665 );
not \U$8997 ( \9667 , \9089 );
not \U$8998 ( \9668 , \7639 );
or \U$8999 ( \9669 , \9667 , \9668 );
and \U$9000 ( \9670 , \9050 , \7378 );
not \U$9001 ( \9671 , \9050 );
and \U$9002 ( \9672 , \9671 , \7739 );
nor \U$9003 ( \9673 , \9670 , \9672 );
nor \U$9004 ( \9674 , \7733 , \9089 );
nor \U$9005 ( \9675 , \9673 , \9674 );
nand \U$9006 ( \9676 , \9669 , \9675 );
not \U$9007 ( \9677 , \8229 );
not \U$9008 ( \9678 , \9677 );
not \U$9009 ( \9679 , \8126 );
or \U$9010 ( \9680 , \9678 , \9679 );
and \U$9011 ( \9681 , \7959 , \8131 );
not \U$9012 ( \9682 , \7959 );
and \U$9013 ( \9683 , \9682 , \8361 );
nor \U$9014 ( \9684 , \9681 , \9683 );
nand \U$9015 ( \9685 , \9680 , \9684 );
and \U$9016 ( \9686 , \8122 , \8229 );
nor \U$9017 ( \9687 , \9685 , \9686 );
not \U$9018 ( \9688 , \9687 );
not \U$9019 ( \9689 , \8493 );
not \U$9020 ( \9690 , \7709 );
or \U$9021 ( \9691 , \9689 , \9690 );
and \U$9022 ( \9692 , \8012 , \8348 );
and \U$9023 ( \9693 , \7708 , \8491 );
nor \U$9024 ( \9694 , \9692 , \9693 );
nand \U$9025 ( \9695 , \9691 , \9694 );
not \U$9026 ( \9696 , \9695 );
and \U$9027 ( \9697 , \9688 , \9696 );
and \U$9028 ( \9698 , \9687 , \9695 );
nor \U$9029 ( \9699 , \9697 , \9698 );
not \U$9030 ( \9700 , \9699 );
not \U$9031 ( \9701 , \9700 );
and \U$9032 ( \9702 , \8502 , \8564 );
not \U$9033 ( \9703 , \7886 );
not \U$9034 ( \9704 , \8439 );
not \U$9035 ( \9705 , \9704 );
or \U$9036 ( \9706 , \9703 , \9705 );
or \U$9037 ( \9707 , \7891 , \8440 );
nand \U$9038 ( \9708 , \9706 , \9707 );
nor \U$9039 ( \9709 , \9702 , \9708 );
nand \U$9040 ( \9710 , \7577 , \9050 );
nand \U$9041 ( \9711 , \9709 , \9710 );
not \U$9042 ( \9712 , \9711 );
or \U$9043 ( \9713 , \9701 , \9712 );
not \U$9044 ( \9714 , \9687 );
nand \U$9045 ( \9715 , \9714 , \9695 );
nand \U$9046 ( \9716 , \9713 , \9715 );
xor \U$9047 ( \9717 , \9676 , \9716 );
not \U$9048 ( \9718 , \9172 );
not \U$9049 ( \9719 , \7389 );
or \U$9050 ( \9720 , \9718 , \9719 );
and \U$9051 ( \9721 , \7102 , \9173 );
or \U$9052 ( \9722 , \7106 , \8910 );
nand \U$9053 ( \9723 , \7070 , \8910 );
nand \U$9054 ( \9724 , \9722 , \9723 );
nor \U$9055 ( \9725 , \9721 , \9724 );
nand \U$9056 ( \9726 , \9720 , \9725 );
and \U$9057 ( \9727 , \9717 , \9726 );
and \U$9058 ( \9728 , \9676 , \9716 );
or \U$9059 ( \9729 , \9727 , \9728 );
and \U$9060 ( \9730 , \9666 , \9729 );
and \U$9061 ( \9731 , \9656 , \9665 );
nor \U$9062 ( \9732 , \9730 , \9731 );
not \U$9063 ( \9733 , \9732 );
not \U$9064 ( \9734 , \9733 );
or \U$9065 ( \9735 , \9594 , \9734 );
not \U$9066 ( \9736 , \9592 );
nand \U$9067 ( \9737 , \9736 , \9566 );
nand \U$9068 ( \9738 , \9735 , \9737 );
xor \U$9069 ( \9739 , \9560 , \9738 );
xor \U$9070 ( \9740 , \9455 , \9453 );
xor \U$9071 ( \9741 , \9740 , \9400 );
and \U$9072 ( \9742 , \9739 , \9741 );
and \U$9073 ( \9743 , \9560 , \9738 );
nor \U$9074 ( \9744 , \9742 , \9743 );
nand \U$9075 ( \9745 , \9559 , \9744 );
and \U$9076 ( \9746 , \9465 , \9557 , \9745 );
not \U$9077 ( \9747 , \9739 );
and \U$9078 ( \9748 , \9741 , \9747 );
not \U$9079 ( \9749 , \9741 );
and \U$9080 ( \9750 , \9749 , \9739 );
nor \U$9081 ( \9751 , \9748 , \9750 );
xor \U$9082 ( \9752 , \9361 , \9396 );
xor \U$9083 ( \9753 , \9752 , \9362 );
not \U$9084 ( \9754 , \9395 );
not \U$9085 ( \9755 , \9754 );
not \U$9086 ( \9756 , \9379 );
or \U$9087 ( \9757 , \9755 , \9756 );
and \U$9088 ( \9758 , \9378 , \9395 );
not \U$9089 ( \9759 , \9650 );
and \U$9090 ( \9760 , \6847 , \9759 );
nor \U$9091 ( \9761 , \9758 , \9760 );
nand \U$9092 ( \9762 , \9757 , \9761 );
xor \U$9093 ( \9763 , \9578 , \9576 );
xnor \U$9094 ( \9764 , \9763 , \9589 );
xor \U$9095 ( \9765 , \9762 , \9764 );
not \U$9096 ( \9766 , \9765 );
not \U$9097 ( \9767 , \9766 );
not \U$9098 ( \9768 , \9729 );
and \U$9099 ( \9769 , \9666 , \9768 );
not \U$9100 ( \9770 , \9666 );
and \U$9101 ( \9771 , \9770 , \9729 );
nor \U$9102 ( \9772 , \9769 , \9771 );
not \U$9103 ( \9773 , \9772 );
and \U$9104 ( \9774 , \9767 , \9773 );
and \U$9105 ( \9775 , \9762 , \9764 );
nor \U$9106 ( \9776 , \9774 , \9775 );
xor \U$9107 ( \9777 , \9753 , \9776 );
xor \U$9108 ( \9778 , \9592 , \9566 );
xnor \U$9109 ( \9779 , \9778 , \9732 );
and \U$9110 ( \9780 , \9777 , \9779 );
and \U$9111 ( \9781 , \9753 , \9776 );
or \U$9112 ( \9782 , \9780 , \9781 );
or \U$9113 ( \9783 , \9751 , \9782 );
not \U$9114 ( \9784 , \9559 );
not \U$9115 ( \9785 , \9744 );
nand \U$9116 ( \9786 , \9784 , \9785 );
nand \U$9117 ( \9787 , \9783 , \9786 );
and \U$9118 ( \9788 , \9746 , \9787 );
not \U$9119 ( \9789 , \9464 );
not \U$9120 ( \9790 , \9359 );
nand \U$9121 ( \9791 , \9789 , \9790 );
not \U$9122 ( \9792 , \9557 );
or \U$9123 ( \9793 , \9791 , \9792 );
not \U$9124 ( \9794 , \9556 );
nand \U$9125 ( \9795 , \9794 , \9471 , \9469 );
nand \U$9126 ( \9796 , \9793 , \9795 );
nor \U$9127 ( \9797 , \9788 , \9796 );
xor \U$9128 ( \9798 , \8627 , \8628 );
not \U$9129 ( \9799 , \9798 );
xnor \U$9130 ( \9800 , \8318 , \8319 );
not \U$9131 ( \9801 , \9800 );
nand \U$9132 ( \9802 , \8572 , \8564 );
not \U$9133 ( \9803 , \9802 );
not \U$9134 ( \9804 , \8565 );
not \U$9135 ( \9805 , \6985 );
or \U$9136 ( \9806 , \9804 , \9805 );
and \U$9137 ( \9807 , \8183 , \8575 );
nor \U$9138 ( \9808 , \7079 , \8575 );
nor \U$9139 ( \9809 , \9807 , \9808 );
nand \U$9140 ( \9810 , \9806 , \9809 );
not \U$9141 ( \9811 , \9810 );
not \U$9142 ( \9812 , \9811 );
or \U$9143 ( \9813 , \9803 , \9812 );
not \U$9144 ( \9814 , \9505 );
not \U$9145 ( \9815 , \9504 );
not \U$9146 ( \9816 , \9515 );
or \U$9147 ( \9817 , \9815 , \9816 );
or \U$9148 ( \9818 , \9504 , \9515 );
nand \U$9149 ( \9819 , \9817 , \9818 );
not \U$9150 ( \9820 , \9819 );
or \U$9151 ( \9821 , \9814 , \9820 );
not \U$9152 ( \9822 , \6846 );
not \U$9153 ( \9823 , \9089 );
and \U$9154 ( \9824 , \9822 , \9823 );
not \U$9155 ( \9825 , \9504 );
and \U$9156 ( \9826 , \9515 , \9825 );
nor \U$9157 ( \9827 , \9824 , \9826 );
nand \U$9158 ( \9828 , \9821 , \9827 );
nand \U$9159 ( \9829 , \9813 , \9828 );
not \U$9160 ( \9830 , \9829 );
xor \U$9161 ( \9831 , \8570 , \8582 );
not \U$9162 ( \9832 , \9831 );
or \U$9163 ( \9833 , \9830 , \9832 );
or \U$9164 ( \9834 , \9831 , \9829 );
nand \U$9165 ( \9835 , \9833 , \9834 );
not \U$9166 ( \9836 , \9835 );
xor \U$9167 ( \9837 , \8475 , \8517 );
xor \U$9168 ( \9838 , \8595 , \8606 );
xor \U$9169 ( \9839 , \9838 , \8618 );
xor \U$9170 ( \9840 , \9837 , \9839 );
not \U$9171 ( \9841 , \9483 );
not \U$9172 ( \9842 , \9502 );
or \U$9173 ( \9843 , \9841 , \9842 );
nand \U$9174 ( \9844 , \9501 , \9492 );
nand \U$9175 ( \9845 , \9843 , \9844 );
and \U$9176 ( \9846 , \9840 , \9845 );
and \U$9177 ( \9847 , \9837 , \9839 );
nor \U$9178 ( \9848 , \9846 , \9847 );
not \U$9179 ( \9849 , \9848 );
not \U$9180 ( \9850 , \9849 );
or \U$9181 ( \9851 , \9836 , \9850 );
not \U$9182 ( \9852 , \9829 );
nand \U$9183 ( \9853 , \9852 , \9831 );
nand \U$9184 ( \9854 , \9851 , \9853 );
not \U$9185 ( \9855 , \9854 );
or \U$9186 ( \9856 , \9801 , \9855 );
or \U$9187 ( \9857 , \9854 , \9800 );
nand \U$9188 ( \9858 , \9856 , \9857 );
not \U$9189 ( \9859 , \9858 );
nand \U$9190 ( \9860 , \9799 , \9859 );
nand \U$9191 ( \9861 , \9858 , \9798 );
and \U$9192 ( \9862 , \9860 , \9861 );
xor \U$9193 ( \9863 , \8585 , \8621 );
xor \U$9194 ( \9864 , \9863 , \8623 );
not \U$9195 ( \9865 , \9864 );
xnor \U$9196 ( \9866 , \9848 , \9835 );
not \U$9197 ( \9867 , \9866 );
or \U$9198 ( \9868 , \9865 , \9867 );
or \U$9199 ( \9869 , \9864 , \9866 );
not \U$9200 ( \9870 , \9802 );
nor \U$9201 ( \9871 , \9870 , \9810 );
xor \U$9202 ( \9872 , \9871 , \9828 );
not \U$9203 ( \9873 , \9872 );
and \U$9204 ( \9874 , \9538 , \9548 );
not \U$9205 ( \9875 , \9874 );
or \U$9206 ( \9876 , \9873 , \9875 );
or \U$9207 ( \9877 , \9874 , \9872 );
nand \U$9208 ( \9878 , \9876 , \9877 );
not \U$9209 ( \9879 , \9878 );
and \U$9210 ( \9880 , \9521 , \9503 );
and \U$9211 ( \9881 , \9516 , \9520 );
nor \U$9212 ( \9882 , \9880 , \9881 );
not \U$9213 ( \9883 , \9882 );
not \U$9214 ( \9884 , \9883 );
or \U$9215 ( \9885 , \9879 , \9884 );
not \U$9216 ( \9886 , \9872 );
nand \U$9217 ( \9887 , \9886 , \9874 );
nand \U$9218 ( \9888 , \9885 , \9887 );
nand \U$9219 ( \9889 , \9869 , \9888 );
nand \U$9220 ( \9890 , \9868 , \9889 );
nor \U$9221 ( \9891 , \9862 , \9890 );
not \U$9222 ( \9892 , \9891 );
not \U$9223 ( \9893 , \8468 );
not \U$9224 ( \9894 , \8641 );
or \U$9225 ( \9895 , \9893 , \9894 );
or \U$9226 ( \9896 , \8468 , \8641 );
nand \U$9227 ( \9897 , \9895 , \9896 );
not \U$9228 ( \9898 , \9800 );
not \U$9229 ( \9899 , \9898 );
not \U$9230 ( \9900 , \9854 );
or \U$9231 ( \9901 , \9899 , \9900 );
nand \U$9232 ( \9902 , \9901 , \9861 );
nand \U$9233 ( \9903 , \9897 , \9902 );
not \U$9234 ( \9904 , \9903 );
or \U$9235 ( \9905 , \9892 , \9904 );
xor \U$9236 ( \9906 , \9864 , \9866 );
xnor \U$9237 ( \9907 , \9906 , \9888 );
xnor \U$9238 ( \9908 , \9840 , \9845 );
xor \U$9239 ( \9909 , \9529 , \9549 );
and \U$9240 ( \9910 , \9909 , \9554 );
and \U$9241 ( \9911 , \9529 , \9549 );
or \U$9242 ( \9912 , \9910 , \9911 );
xor \U$9243 ( \9913 , \9908 , \9912 );
not \U$9244 ( \9914 , \9882 );
not \U$9245 ( \9915 , \9878 );
and \U$9246 ( \9916 , \9914 , \9915 );
and \U$9247 ( \9917 , \9878 , \9882 );
nor \U$9248 ( \9918 , \9916 , \9917 );
and \U$9249 ( \9919 , \9913 , \9918 );
and \U$9250 ( \9920 , \9908 , \9912 );
or \U$9251 ( \9921 , \9919 , \9920 );
nand \U$9252 ( \9922 , \9907 , \9921 );
xor \U$9253 ( \9923 , \9908 , \9912 );
xor \U$9254 ( \9924 , \9923 , \9918 );
xor \U$9255 ( \9925 , \9477 , \9526 );
and \U$9256 ( \9926 , \9925 , \9555 );
and \U$9257 ( \9927 , \9477 , \9526 );
or \U$9258 ( \9928 , \9926 , \9927 );
nand \U$9259 ( \9929 , \9924 , \9928 );
nand \U$9260 ( \9930 , \9922 , \9929 );
not \U$9261 ( \9931 , \9930 );
nand \U$9262 ( \9932 , \9905 , \9931 );
or \U$9263 ( \9933 , \9797 , \9932 );
nor \U$9264 ( \9934 , \9924 , \9928 );
nand \U$9265 ( \9935 , \9922 , \9934 );
not \U$9266 ( \9936 , \9907 );
not \U$9267 ( \9937 , \9921 );
nand \U$9268 ( \9938 , \9936 , \9937 );
and \U$9269 ( \9939 , \9935 , \9938 );
nand \U$9270 ( \9940 , \9860 , \9861 , \9890 );
nand \U$9271 ( \9941 , \9939 , \9903 , \9940 );
nand \U$9272 ( \9942 , \9903 , \9891 );
nand \U$9273 ( \9943 , \9941 , \9942 );
nand \U$9274 ( \9944 , \9933 , \9943 );
xor \U$9275 ( \9945 , \9595 , \9602 );
xor \U$9276 ( \9946 , \9945 , \9653 );
not \U$9277 ( \9947 , \9946 );
not \U$9278 ( \9948 , \9657 );
not \U$9279 ( \9949 , \7389 );
or \U$9280 ( \9950 , \9948 , \9949 );
and \U$9281 ( \9951 , \9038 , \9449 );
and \U$9282 ( \9952 , \9173 , \7106 );
not \U$9283 ( \9953 , \9173 );
and \U$9284 ( \9954 , \9953 , \8602 );
nor \U$9285 ( \9955 , \9952 , \9954 );
nor \U$9286 ( \9956 , \9951 , \9955 );
nand \U$9287 ( \9957 , \9950 , \9956 );
not \U$9288 ( \9958 , \9957 );
not \U$9289 ( \9959 , \9958 );
not \U$9290 ( \9960 , \9700 );
not \U$9291 ( \9961 , \9711 );
not \U$9292 ( \9962 , \9961 );
or \U$9293 ( \9963 , \9960 , \9962 );
nand \U$9294 ( \9964 , \9699 , \9711 );
nand \U$9295 ( \9965 , \9963 , \9964 );
not \U$9296 ( \9966 , \9965 );
not \U$9297 ( \9967 , \9966 );
or \U$9298 ( \9968 , \9959 , \9967 );
not \U$9299 ( \9969 , \9957 );
not \U$9300 ( \9970 , \9965 );
or \U$9301 ( \9971 , \9969 , \9970 );
not \U$9302 ( \9972 , \8752 );
not \U$9303 ( \9973 , \9059 );
or \U$9304 ( \9974 , \9972 , \9973 );
and \U$9305 ( \9975 , \7214 , \7152 );
and \U$9306 ( \9976 , \9975 , \8751 );
not \U$9307 ( \9977 , \8909 );
not \U$9308 ( \9978 , \7154 );
or \U$9309 ( \9979 , \9977 , \9978 );
or \U$9310 ( \9980 , \7160 , \8909 );
nand \U$9311 ( \9981 , \9979 , \9980 );
nor \U$9312 ( \9982 , \9976 , \9981 );
nand \U$9313 ( \9983 , \9974 , \9982 );
not \U$9314 ( \9984 , \9983 );
nand \U$9315 ( \9985 , \9971 , \9984 );
nand \U$9316 ( \9986 , \9968 , \9985 );
not \U$9317 ( \9987 , \9986 );
or \U$9318 ( \9988 , \9947 , \9987 );
or \U$9319 ( \9989 , \9986 , \9946 );
nand \U$9320 ( \9990 , \9988 , \9989 );
not \U$9321 ( \9991 , \9990 );
xor \U$9322 ( \9992 , \9676 , \9716 );
xor \U$9323 ( \9993 , \9992 , \9726 );
not \U$9324 ( \9994 , \9993 );
and \U$9325 ( \9995 , \9991 , \9994 );
and \U$9326 ( \9996 , \9990 , \9993 );
nor \U$9327 ( \9997 , \9995 , \9996 );
not \U$9328 ( \9998 , \9997 );
not \U$9329 ( \9999 , \9998 );
buf \U$9330 ( \10000 , \7150 );
nand \U$9331 ( \10001 , \10000 , \8970 );
not \U$9332 ( \10002 , \10001 );
not \U$9333 ( \10003 , \9043 );
and \U$9334 ( \10004 , \7646 , \10003 );
nor \U$9335 ( \10005 , \10004 , \7371 );
not \U$9336 ( \10006 , \10005 );
or \U$9337 ( \10007 , \10002 , \10006 );
nand \U$9338 ( \10008 , \10007 , \7641 );
not \U$9339 ( \10009 , \7373 );
nor \U$9340 ( \10010 , \10009 , \8804 );
and \U$9341 ( \10011 , \7646 , \7371 , \9039 );
nor \U$9342 ( \10012 , \10010 , \10011 );
nand \U$9343 ( \10013 , \10008 , \10012 );
not \U$9344 ( \10014 , \10013 );
nand \U$9345 ( \10015 , \7048 , \7058 );
and \U$9346 ( \10016 , \9649 , \10015 );
nor \U$9347 ( \10017 , \7048 , \7058 );
nor \U$9348 ( \10018 , \10016 , \10017 );
nand \U$9349 ( \10019 , \6916 , \10018 );
not \U$9350 ( \10020 , \8348 );
not \U$9351 ( \10021 , \7959 );
or \U$9352 ( \10022 , \10020 , \10021 );
nand \U$9353 ( \10023 , \8012 , \8491 );
nand \U$9354 ( \10024 , \10022 , \10023 );
not \U$9355 ( \10025 , \8493 );
nor \U$9356 ( \10026 , \10025 , \8012 );
nor \U$9357 ( \10027 , \10024 , \10026 );
nor \U$9358 ( \10028 , \10019 , \10027 );
not \U$9359 ( \10029 , \10028 );
not \U$9360 ( \10030 , \10029 );
nor \U$9361 ( \10031 , \6919 , \9650 );
not \U$9362 ( \10032 , \10031 );
or \U$9363 ( \10033 , \10030 , \10032 );
or \U$9364 ( \10034 , \10031 , \10029 );
nand \U$9365 ( \10035 , \10033 , \10034 );
not \U$9366 ( \10036 , \10035 );
or \U$9367 ( \10037 , \10014 , \10036 );
not \U$9368 ( \10038 , \10031 );
nand \U$9369 ( \10039 , \10038 , \10029 );
nand \U$9370 ( \10040 , \10037 , \10039 );
or \U$9371 ( \10041 , \7337 , \8804 );
not \U$9372 ( \10042 , \8050 );
not \U$9373 ( \10043 , \8752 );
and \U$9374 ( \10044 , \10042 , \10043 );
and \U$9375 ( \10045 , \7161 , \8752 );
nor \U$9376 ( \10046 , \10044 , \10045 );
nand \U$9377 ( \10047 , \10041 , \10046 );
nor \U$9378 ( \10048 , \7216 , \8918 );
nor \U$9379 ( \10049 , \10047 , \10048 );
nor \U$9380 ( \10050 , \10040 , \10049 );
not \U$9381 ( \10051 , \10050 );
nand \U$9382 ( \10052 , \10040 , \10049 );
nand \U$9383 ( \10053 , \10051 , \10052 );
not \U$9384 ( \10054 , \10053 );
xor \U$9385 ( \10055 , \6929 , \9650 );
not \U$9386 ( \10056 , \10055 );
not \U$9387 ( \10057 , \6923 );
and \U$9388 ( \10058 , \10056 , \10057 );
or \U$9389 ( \10059 , \7079 , \9657 );
nand \U$9390 ( \10060 , \8183 , \9657 );
nand \U$9391 ( \10061 , \10059 , \10060 );
nor \U$9392 ( \10062 , \10058 , \10061 );
not \U$9393 ( \10063 , \10062 );
and \U$9394 ( \10064 , \10054 , \10063 );
and \U$9395 ( \10065 , \10053 , \10062 );
nor \U$9396 ( \10066 , \10064 , \10065 );
not \U$9397 ( \10067 , \10066 );
not \U$9398 ( \10068 , \10067 );
buf \U$9399 ( \10069 , \10013 );
buf \U$9400 ( \10070 , \10035 );
xor \U$9401 ( \10071 , \10069 , \10070 );
not \U$9402 ( \10072 , \10071 );
not \U$9403 ( \10073 , \8752 );
not \U$9404 ( \10074 , \8061 );
or \U$9405 ( \10075 , \10073 , \10074 );
or \U$9406 ( \10076 , \7378 , \8803 );
nand \U$9407 ( \10077 , \9201 , \8803 );
nand \U$9408 ( \10078 , \10076 , \10077 );
and \U$9409 ( \10079 , \7640 , \8751 );
nor \U$9410 ( \10080 , \10078 , \10079 );
nand \U$9411 ( \10081 , \10075 , \10080 );
not \U$9412 ( \10082 , \10081 );
not \U$9413 ( \10083 , \10082 );
nor \U$9414 ( \10084 , \7063 , \9650 );
not \U$9415 ( \10085 , \10084 );
not \U$9416 ( \10086 , \8348 );
not \U$9417 ( \10087 , \9677 );
or \U$9418 ( \10088 , \10086 , \10087 );
not \U$9419 ( \10089 , \7958 );
not \U$9420 ( \10090 , \8491 );
not \U$9421 ( \10091 , \10090 );
and \U$9422 ( \10092 , \10089 , \10091 );
and \U$9423 ( \10093 , \9232 , \8493 );
nor \U$9424 ( \10094 , \10092 , \10093 );
nand \U$9425 ( \10095 , \10088 , \10094 );
not \U$9426 ( \10096 , \8563 );
not \U$9427 ( \10097 , \8122 );
or \U$9428 ( \10098 , \10096 , \10097 );
and \U$9429 ( \10099 , \9210 , \8562 );
and \U$9430 ( \10100 , \8437 , \8360 );
not \U$9431 ( \10101 , \8437 );
and \U$9432 ( \10102 , \10101 , \8130 );
nor \U$9433 ( \10103 , \10100 , \10102 );
nor \U$9434 ( \10104 , \10099 , \10103 );
nand \U$9435 ( \10105 , \10098 , \10104 );
xor \U$9436 ( \10106 , \10095 , \10105 );
not \U$9437 ( \10107 , \10106 );
or \U$9438 ( \10108 , \10085 , \10107 );
nand \U$9439 ( \10109 , \10105 , \10095 );
nand \U$9440 ( \10110 , \10108 , \10109 );
not \U$9441 ( \10111 , \10110 );
not \U$9442 ( \10112 , \10111 );
or \U$9443 ( \10113 , \10083 , \10112 );
not \U$9444 ( \10114 , \10081 );
not \U$9445 ( \10115 , \10110 );
or \U$9446 ( \10116 , \10114 , \10115 );
not \U$9447 ( \10117 , \9759 );
not \U$9448 ( \10118 , \9038 );
or \U$9449 ( \10119 , \10117 , \10118 );
and \U$9450 ( \10120 , \9448 , \7107 );
not \U$9451 ( \10121 , \9448 );
and \U$9452 ( \10122 , \10121 , \7070 );
nor \U$9453 ( \10123 , \10120 , \10122 );
nand \U$9454 ( \10124 , \10119 , \10123 );
and \U$9455 ( \10125 , \7388 , \9650 );
nor \U$9456 ( \10126 , \10124 , \10125 );
nand \U$9457 ( \10127 , \10116 , \10126 );
nand \U$9458 ( \10128 , \10113 , \10127 );
not \U$9459 ( \10129 , \10128 );
and \U$9460 ( \10130 , \8477 , \8440 );
or \U$9461 ( \10131 , \8362 , \8230 );
nand \U$9462 ( \10132 , \8131 , \8230 );
nand \U$9463 ( \10133 , \10131 , \10132 );
nor \U$9464 ( \10134 , \10130 , \10133 );
nand \U$9465 ( \10135 , \8122 , \8439 );
nand \U$9466 ( \10136 , \10134 , \10135 );
and \U$9467 ( \10137 , \8502 , \9043 );
or \U$9468 ( \10138 , \7559 , \8563 );
nand \U$9469 ( \10139 , \7856 , \8563 );
nand \U$9470 ( \10140 , \10138 , \10139 );
nor \U$9471 ( \10141 , \10137 , \10140 );
nand \U$9472 ( \10142 , \7577 , \8969 );
nand \U$9473 ( \10143 , \10141 , \10142 );
xor \U$9474 ( \10144 , \10136 , \10143 );
nand \U$9475 ( \10145 , \10019 , \10027 );
not \U$9476 ( \10146 , \10145 );
nor \U$9477 ( \10147 , \10146 , \10028 );
and \U$9478 ( \10148 , \10144 , \10147 );
and \U$9479 ( \10149 , \10136 , \10143 );
or \U$9480 ( \10150 , \10148 , \10149 );
not \U$9481 ( \10151 , \10150 );
and \U$9482 ( \10152 , \10129 , \10151 );
and \U$9483 ( \10153 , \10128 , \10150 );
nor \U$9484 ( \10154 , \10152 , \10153 );
not \U$9485 ( \10155 , \10154 );
not \U$9486 ( \10156 , \10155 );
or \U$9487 ( \10157 , \10072 , \10156 );
not \U$9488 ( \10158 , \10150 );
nand \U$9489 ( \10159 , \10158 , \10128 );
nand \U$9490 ( \10160 , \10157 , \10159 );
not \U$9491 ( \10161 , \10160 );
not \U$9492 ( \10162 , \10161 );
or \U$9493 ( \10163 , \10068 , \10162 );
nand \U$9494 ( \10164 , \10160 , \10066 );
nand \U$9495 ( \10165 , \10163 , \10164 );
not \U$9496 ( \10166 , \10165 );
or \U$9497 ( \10167 , \9999 , \10166 );
not \U$9498 ( \10168 , \10066 );
nand \U$9499 ( \10169 , \10168 , \10160 );
nand \U$9500 ( \10170 , \10167 , \10169 );
not \U$9501 ( \10171 , \10062 );
and \U$9502 ( \10172 , \10052 , \10171 );
nor \U$9503 ( \10173 , \10172 , \10050 );
not \U$9504 ( \10174 , \9993 );
not \U$9505 ( \10175 , \10174 );
not \U$9506 ( \10176 , \9990 );
or \U$9507 ( \10177 , \10175 , \10176 );
not \U$9508 ( \10178 , \9946 );
nand \U$9509 ( \10179 , \10178 , \9986 );
nand \U$9510 ( \10180 , \10177 , \10179 );
xor \U$9511 ( \10181 , \10173 , \10180 );
not \U$9512 ( \10182 , \9772 );
not \U$9513 ( \10183 , \9765 );
and \U$9514 ( \10184 , \10182 , \10183 );
and \U$9515 ( \10185 , \9765 , \9772 );
nor \U$9516 ( \10186 , \10184 , \10185 );
xor \U$9517 ( \10187 , \10181 , \10186 );
xor \U$9518 ( \10188 , \10170 , \10187 );
xor \U$9519 ( \10189 , \10106 , \10084 );
or \U$9520 ( \10190 , \7215 , \9173 );
nand \U$9521 ( \10191 , \9975 , \9173 );
and \U$9522 ( \10192 , \7161 , \9657 );
and \U$9523 ( \10193 , \7155 , \9448 );
nor \U$9524 ( \10194 , \10192 , \10193 );
nand \U$9525 ( \10195 , \10190 , \10191 , \10194 );
and \U$9526 ( \10196 , \7158 , \7646 );
nor \U$9527 ( \10197 , \10196 , \9650 );
nor \U$9528 ( \10198 , \10197 , \7497 );
not \U$9529 ( \10199 , \10198 );
not \U$9530 ( \10200 , \9210 );
not \U$9531 ( \10201 , \8968 );
or \U$9532 ( \10202 , \10200 , \10201 );
and \U$9533 ( \10203 , \8561 , \8361 );
not \U$9534 ( \10204 , \8561 );
and \U$9535 ( \10205 , \10204 , \8131 );
nor \U$9536 ( \10206 , \10203 , \10205 );
nand \U$9537 ( \10207 , \10202 , \10206 );
not \U$9538 ( \10208 , \10207 );
nand \U$9539 ( \10209 , \9042 , \8122 );
nand \U$9540 ( \10210 , \10208 , \10209 );
not \U$9541 ( \10211 , \10210 );
not \U$9542 ( \10212 , \8438 );
nand \U$9543 ( \10213 , \10212 , \8348 );
not \U$9544 ( \10214 , \8228 );
nand \U$9545 ( \10215 , \10214 , \8491 );
nand \U$9546 ( \10216 , \8228 , \8493 );
and \U$9547 ( \10217 , \10213 , \10215 , \10216 );
not \U$9548 ( \10218 , \10217 );
and \U$9549 ( \10219 , \10211 , \10218 );
and \U$9550 ( \10220 , \10210 , \10217 );
nor \U$9551 ( \10221 , \10219 , \10220 );
not \U$9552 ( \10222 , \10221 );
not \U$9553 ( \10223 , \8750 );
not \U$9554 ( \10224 , \9240 );
or \U$9555 ( \10225 , \10223 , \10224 );
not \U$9556 ( \10226 , \8750 );
and \U$9557 ( \10227 , \9230 , \10226 );
or \U$9558 ( \10228 , \9234 , \8801 );
nand \U$9559 ( \10229 , \7886 , \8801 );
nand \U$9560 ( \10230 , \10228 , \10229 );
nor \U$9561 ( \10231 , \10227 , \10230 );
nand \U$9562 ( \10232 , \10225 , \10231 );
not \U$9563 ( \10233 , \10232 );
or \U$9564 ( \10234 , \10222 , \10233 );
or \U$9565 ( \10235 , \10232 , \10221 );
nand \U$9566 ( \10236 , \10234 , \10235 );
not \U$9567 ( \10237 , \10236 );
or \U$9568 ( \10238 , \10199 , \10237 );
not \U$9569 ( \10239 , \10221 );
nand \U$9570 ( \10240 , \10239 , \10232 );
nand \U$9571 ( \10241 , \10238 , \10240 );
xor \U$9572 ( \10242 , \10195 , \10241 );
xor \U$9573 ( \10243 , \10189 , \10242 );
not \U$9574 ( \10244 , \10243 );
not \U$9575 ( \10245 , \9059 );
not \U$9576 ( \10246 , \9657 );
or \U$9577 ( \10247 , \10245 , \10246 );
not \U$9578 ( \10248 , \9448 );
not \U$9579 ( \10249 , \7214 );
or \U$9580 ( \10250 , \10248 , \10249 );
nand \U$9581 ( \10251 , \7495 , \9649 );
nand \U$9582 ( \10252 , \10250 , \10251 );
and \U$9583 ( \10253 , \10252 , \7152 );
and \U$9584 ( \10254 , \7161 , \9650 );
nor \U$9585 ( \10255 , \10253 , \10254 );
nand \U$9586 ( \10256 , \10247 , \10255 );
and \U$9587 ( \10257 , \7640 , \9173 );
not \U$9588 ( \10258 , \10257 );
not \U$9589 ( \10259 , \9173 );
nand \U$9590 ( \10260 , \10259 , \7639 );
and \U$9591 ( \10261 , \8909 , \7740 );
not \U$9592 ( \10262 , \8909 );
and \U$9593 ( \10263 , \10262 , \7790 );
nor \U$9594 ( \10264 , \10261 , \10263 );
nand \U$9595 ( \10265 , \10258 , \10260 , \10264 );
xor \U$9596 ( \10266 , \10256 , \10265 );
not \U$9597 ( \10267 , \8125 );
and \U$9598 ( \10268 , \7872 , \8968 );
not \U$9599 ( \10269 , \7872 );
and \U$9600 ( \10270 , \10269 , \9042 );
nor \U$9601 ( \10271 , \10268 , \10270 );
not \U$9602 ( \10272 , \10271 );
or \U$9603 ( \10273 , \10267 , \10272 );
not \U$9604 ( \10274 , \8120 );
and \U$9605 ( \10275 , \8800 , \10274 );
not \U$9606 ( \10276 , \8800 );
and \U$9607 ( \10277 , \10276 , \8120 );
nor \U$9608 ( \10278 , \10275 , \10277 );
not \U$9609 ( \10279 , \8125 );
nand \U$9610 ( \10280 , \10278 , \10279 );
nand \U$9611 ( \10281 , \10280 , \8117 );
nand \U$9612 ( \10282 , \10273 , \10281 );
and \U$9613 ( \10283 , \8439 , \8493 );
not \U$9614 ( \10284 , \8348 );
or \U$9615 ( \10285 , \8563 , \10284 );
or \U$9616 ( \10286 , \8438 , \10090 );
nand \U$9617 ( \10287 , \10285 , \10286 );
nor \U$9618 ( \10288 , \10283 , \10287 );
nand \U$9619 ( \10289 , \10282 , \10288 );
not \U$9620 ( \10290 , \10289 );
and \U$9621 ( \10291 , \7865 , \9112 );
and \U$9622 ( \10292 , \10226 , \7891 );
not \U$9623 ( \10293 , \10226 );
and \U$9624 ( \10294 , \10293 , \7559 );
nor \U$9625 ( \10295 , \10292 , \10294 );
nor \U$9626 ( \10296 , \10291 , \10295 );
nand \U$9627 ( \10297 , \7577 , \8910 );
nand \U$9628 ( \10298 , \10296 , \10297 );
not \U$9629 ( \10299 , \10298 );
or \U$9630 ( \10300 , \10290 , \10299 );
or \U$9631 ( \10301 , \10282 , \10288 );
nand \U$9632 ( \10302 , \10300 , \10301 );
and \U$9633 ( \10303 , \10266 , \10302 );
and \U$9634 ( \10304 , \10256 , \10265 );
nor \U$9635 ( \10305 , \10303 , \10304 );
not \U$9636 ( \10306 , \10217 );
and \U$9637 ( \10307 , \10210 , \10306 );
not \U$9638 ( \10308 , \10307 );
not \U$9639 ( \10309 , \8800 );
not \U$9640 ( \10310 , \9230 );
or \U$9641 ( \10311 , \10309 , \10310 );
and \U$9642 ( \10312 , \8969 , \7887 );
not \U$9643 ( \10313 , \8969 );
and \U$9644 ( \10314 , \10313 , \7856 );
nor \U$9645 ( \10315 , \10312 , \10314 );
nand \U$9646 ( \10316 , \10311 , \10315 );
not \U$9647 ( \10317 , \9240 );
nor \U$9648 ( \10318 , \10317 , \8803 );
nor \U$9649 ( \10319 , \10316 , \10318 );
not \U$9650 ( \10320 , \10319 );
or \U$9651 ( \10321 , \10308 , \10320 );
or \U$9652 ( \10322 , \10319 , \10307 );
nand \U$9653 ( \10323 , \10321 , \10322 );
not \U$9654 ( \10324 , \8910 );
not \U$9655 ( \10325 , \7639 );
or \U$9656 ( \10326 , \10324 , \10325 );
or \U$9657 ( \10327 , \7378 , \8751 );
nand \U$9658 ( \10328 , \9201 , \8751 );
nand \U$9659 ( \10329 , \10327 , \10328 );
not \U$9660 ( \10330 , \8909 );
nor \U$9661 ( \10331 , \10330 , \7733 );
nor \U$9662 ( \10332 , \10329 , \10331 );
nand \U$9663 ( \10333 , \10326 , \10332 );
xor \U$9664 ( \10334 , \10323 , \10333 );
xor \U$9665 ( \10335 , \10305 , \10334 );
not \U$9666 ( \10336 , \10335 );
or \U$9667 ( \10337 , \10244 , \10336 );
or \U$9668 ( \10338 , \10335 , \10243 );
nand \U$9669 ( \10339 , \10337 , \10338 );
not \U$9670 ( \10340 , \10339 );
not \U$9671 ( \10341 , \10340 );
xor \U$9672 ( \10342 , \10236 , \10198 );
not \U$9673 ( \10343 , \10342 );
not \U$9674 ( \10344 , \8811 );
and \U$9675 ( \10345 , \10344 , \8750 );
not \U$9676 ( \10346 , \8131 );
and \U$9677 ( \10347 , \8801 , \10346 );
not \U$9678 ( \10348 , \8801 );
and \U$9679 ( \10349 , \10348 , \8362 );
nor \U$9680 ( \10350 , \10347 , \10349 );
nor \U$9681 ( \10351 , \10345 , \10350 );
nand \U$9682 ( \10352 , \8122 , \10226 );
nand \U$9683 ( \10353 , \10351 , \10352 );
not \U$9684 ( \10354 , \9649 );
and \U$9685 ( \10355 , \10354 , \7570 );
nor \U$9686 ( \10356 , \10355 , \7375 );
nor \U$9687 ( \10357 , \10354 , \7570 );
nor \U$9688 ( \10358 , \10356 , \10357 );
and \U$9689 ( \10359 , \10000 , \10358 );
nand \U$9690 ( \10360 , \10353 , \10359 );
not \U$9691 ( \10361 , \9650 );
nand \U$9692 ( \10362 , \10361 , \7774 );
xor \U$9693 ( \10363 , \10360 , \10362 );
and \U$9694 ( \10364 , \9173 , \7740 );
not \U$9695 ( \10365 , \9173 );
and \U$9696 ( \10366 , \10365 , \7790 );
nor \U$9697 ( \10367 , \10364 , \10366 );
nand \U$9698 ( \10368 , \7640 , \9449 );
nand \U$9699 ( \10369 , \10367 , \10368 );
nor \U$9700 ( \10370 , \7376 , \9448 );
nor \U$9701 ( \10371 , \10369 , \10370 );
and \U$9702 ( \10372 , \10363 , \10371 );
and \U$9703 ( \10373 , \10360 , \10362 );
or \U$9704 ( \10374 , \10372 , \10373 );
not \U$9705 ( \10375 , \10374 );
or \U$9706 ( \10376 , \10343 , \10375 );
or \U$9707 ( \10377 , \10374 , \10342 );
nand \U$9708 ( \10378 , \10376 , \10377 );
not \U$9709 ( \10379 , \10378 );
xnor \U$9710 ( \10380 , \10266 , \10302 );
not \U$9711 ( \10381 , \10380 );
not \U$9712 ( \10382 , \10381 );
or \U$9713 ( \10383 , \10379 , \10382 );
not \U$9714 ( \10384 , \10374 );
nand \U$9715 ( \10385 , \10384 , \10342 );
nand \U$9716 ( \10386 , \10383 , \10385 );
not \U$9717 ( \10387 , \10386 );
not \U$9718 ( \10388 , \10387 );
and \U$9719 ( \10389 , \10341 , \10388 );
and \U$9720 ( \10390 , \10339 , \10387 );
not \U$9721 ( \10391 , \10339 );
and \U$9722 ( \10392 , \10391 , \10386 );
or \U$9723 ( \10393 , \10390 , \10392 );
and \U$9724 ( \10394 , \8562 , \8491 );
and \U$9725 ( \10395 , \8563 , \8493 );
nor \U$9726 ( \10396 , \10394 , \10395 );
nand \U$9727 ( \10397 , \8969 , \8348 );
and \U$9728 ( \10398 , \10396 , \10397 );
not \U$9729 ( \10399 , \10398 );
and \U$9730 ( \10400 , \8909 , \9233 );
not \U$9731 ( \10401 , \8909 );
and \U$9732 ( \10402 , \10401 , \7886 );
nor \U$9733 ( \10403 , \10400 , \10402 );
not \U$9734 ( \10404 , \10403 );
and \U$9735 ( \10405 , \9173 , \9230 );
not \U$9736 ( \10406 , \9173 );
and \U$9737 ( \10407 , \10406 , \9240 );
or \U$9738 ( \10408 , \10405 , \10407 );
nor \U$9739 ( \10409 , \10404 , \10408 );
not \U$9740 ( \10410 , \10409 );
nand \U$9741 ( \10411 , \10399 , \10410 );
not \U$9742 ( \10412 , \10411 );
xnor \U$9743 ( \10413 , \10353 , \10359 );
not \U$9744 ( \10414 , \10413 );
or \U$9745 ( \10415 , \10412 , \10414 );
nand \U$9746 ( \10416 , \10409 , \10398 );
nand \U$9747 ( \10417 , \10415 , \10416 );
nand \U$9748 ( \10418 , \10301 , \10289 );
xor \U$9749 ( \10419 , \10418 , \10298 );
xor \U$9750 ( \10420 , \10417 , \10419 );
xor \U$9751 ( \10421 , \10360 , \10362 );
xor \U$9752 ( \10422 , \10421 , \10371 );
xor \U$9753 ( \10423 , \10420 , \10422 );
nor \U$9754 ( \10424 , \7371 , \10354 );
not \U$9755 ( \10425 , \10424 );
not \U$9756 ( \10426 , \10425 );
and \U$9757 ( \10427 , \8122 , \8909 );
not \U$9758 ( \10428 , \8908 );
not \U$9759 ( \10429 , \8126 );
or \U$9760 ( \10430 , \10428 , \10429 );
and \U$9761 ( \10431 , \8749 , \8131 );
not \U$9762 ( \10432 , \8749 );
and \U$9763 ( \10433 , \10432 , \8361 );
nor \U$9764 ( \10434 , \10431 , \10433 );
nand \U$9765 ( \10435 , \10430 , \10434 );
nor \U$9766 ( \10436 , \10427 , \10435 );
not \U$9767 ( \10437 , \10436 );
not \U$9768 ( \10438 , \10437 );
or \U$9769 ( \10439 , \10426 , \10438 );
nand \U$9770 ( \10440 , \10436 , \10424 );
nand \U$9771 ( \10441 , \10439 , \10440 );
not \U$9772 ( \10442 , \10441 );
or \U$9773 ( \10443 , \7559 , \9173 );
nand \U$9774 ( \10444 , \9233 , \9173 );
nand \U$9775 ( \10445 , \10443 , \10444 );
not \U$9776 ( \10446 , \10445 );
not \U$9777 ( \10447 , \9448 );
not \U$9778 ( \10448 , \10447 );
nand \U$9779 ( \10449 , \10448 , \8502 );
nand \U$9780 ( \10450 , \7577 , \10447 );
nand \U$9781 ( \10451 , \10446 , \10449 , \10450 );
not \U$9782 ( \10452 , \10451 );
or \U$9783 ( \10453 , \10442 , \10452 );
nand \U$9784 ( \10454 , \10437 , \10424 );
nand \U$9785 ( \10455 , \10453 , \10454 );
not \U$9786 ( \10456 , \10455 );
and \U$9787 ( \10457 , \7639 , \9650 );
not \U$9788 ( \10458 , \9649 );
not \U$9789 ( \10459 , \7640 );
or \U$9790 ( \10460 , \10458 , \10459 );
and \U$9791 ( \10461 , \10447 , \7790 );
not \U$9792 ( \10462 , \10447 );
and \U$9793 ( \10463 , \10462 , \7740 );
nor \U$9794 ( \10464 , \10461 , \10463 );
nand \U$9795 ( \10465 , \10460 , \10464 );
nor \U$9796 ( \10466 , \10457 , \10465 );
not \U$9797 ( \10467 , \10466 );
and \U$9798 ( \10468 , \10456 , \10467 );
and \U$9799 ( \10469 , \10455 , \10466 );
nor \U$9800 ( \10470 , \10468 , \10469 );
not \U$9801 ( \10471 , \10470 );
nand \U$9802 ( \10472 , \10411 , \10416 );
and \U$9803 ( \10473 , \10472 , \10413 );
not \U$9804 ( \10474 , \10472 );
not \U$9805 ( \10475 , \10413 );
and \U$9806 ( \10476 , \10474 , \10475 );
nor \U$9807 ( \10477 , \10473 , \10476 );
and \U$9808 ( \10478 , \10471 , \10477 );
not \U$9809 ( \10479 , \10455 );
nor \U$9810 ( \10480 , \10479 , \10466 );
nor \U$9811 ( \10481 , \10478 , \10480 );
nand \U$9812 ( \10482 , \10423 , \10481 );
not \U$9813 ( \10483 , \10482 );
xor \U$9814 ( \10484 , \10470 , \10477 );
not \U$9815 ( \10485 , \9173 );
not \U$9816 ( \10486 , \8122 );
or \U$9817 ( \10487 , \10485 , \10486 );
and \U$9818 ( \10488 , \8477 , \9172 );
and \U$9819 ( \10489 , \8908 , \8130 );
not \U$9820 ( \10490 , \8908 );
and \U$9821 ( \10491 , \10490 , \8362 );
nor \U$9822 ( \10492 , \10489 , \10491 );
nor \U$9823 ( \10493 , \10488 , \10492 );
nand \U$9824 ( \10494 , \10487 , \10493 );
nand \U$9825 ( \10495 , \7563 , \8120 );
nand \U$9826 ( \10496 , \9649 , \10495 );
nand \U$9827 ( \10497 , \7561 , \10274 );
and \U$9828 ( \10498 , \10496 , \7557 , \10497 );
nand \U$9829 ( \10499 , \10494 , \10498 );
not \U$9830 ( \10500 , \10499 );
not \U$9831 ( \10501 , \8348 );
not \U$9832 ( \10502 , \9039 );
or \U$9833 ( \10503 , \10501 , \10502 );
and \U$9834 ( \10504 , \10003 , \8491 );
and \U$9835 ( \10505 , \9043 , \8493 );
nor \U$9836 ( \10506 , \10504 , \10505 );
nand \U$9837 ( \10507 , \10503 , \10506 );
not \U$9838 ( \10508 , \10507 );
and \U$9839 ( \10509 , \10500 , \10508 );
and \U$9840 ( \10510 , \10499 , \10507 );
nor \U$9841 ( \10511 , \10509 , \10510 );
not \U$9842 ( \10512 , \10511 );
xor \U$9843 ( \10513 , \10441 , \10451 );
and \U$9844 ( \10514 , \10512 , \10513 );
not \U$9845 ( \10515 , \10507 );
nor \U$9846 ( \10516 , \10515 , \10499 );
nor \U$9847 ( \10517 , \10514 , \10516 );
nand \U$9848 ( \10518 , \10484 , \10517 );
not \U$9849 ( \10519 , \10518 );
not \U$9850 ( \10520 , \7578 );
not \U$9851 ( \10521 , \9649 );
and \U$9852 ( \10522 , \10520 , \10521 );
not \U$9853 ( \10523 , \9759 );
not \U$9854 ( \10524 , \7863 );
or \U$9855 ( \10525 , \10523 , \10524 );
and \U$9856 ( \10526 , \10447 , \7887 );
not \U$9857 ( \10527 , \10447 );
and \U$9858 ( \10528 , \10527 , \7856 );
nor \U$9859 ( \10529 , \10526 , \10528 );
nand \U$9860 ( \10530 , \10525 , \10529 );
nor \U$9861 ( \10531 , \10522 , \10530 );
and \U$9862 ( \10532 , \10226 , \8348 );
and \U$9863 ( \10533 , \8801 , \8108 );
nor \U$9864 ( \10534 , \10532 , \10533 );
or \U$9865 ( \10535 , \8802 , \8347 );
nand \U$9866 ( \10536 , \10535 , \9382 );
nand \U$9867 ( \10537 , \10534 , \10536 );
nand \U$9868 ( \10538 , \10531 , \10537 );
not \U$9869 ( \10539 , \10538 );
xor \U$9870 ( \10540 , \10498 , \10494 );
not \U$9871 ( \10541 , \10540 );
or \U$9872 ( \10542 , \10539 , \10541 );
not \U$9873 ( \10543 , \10537 );
not \U$9874 ( \10544 , \10531 );
nand \U$9875 ( \10545 , \10543 , \10544 );
nand \U$9876 ( \10546 , \10542 , \10545 );
not \U$9877 ( \10547 , \10546 );
not \U$9878 ( \10548 , \10547 );
not \U$9879 ( \10549 , \10513 );
not \U$9880 ( \10550 , \10511 );
and \U$9881 ( \10551 , \10549 , \10550 );
and \U$9882 ( \10552 , \10513 , \10511 );
nor \U$9883 ( \10553 , \10551 , \10552 );
not \U$9884 ( \10554 , \10553 );
or \U$9885 ( \10555 , \10548 , \10554 );
and \U$9886 ( \10556 , \8748 , \8493 );
not \U$9887 ( \10557 , \8748 );
and \U$9888 ( \10558 , \10557 , \8491 );
nor \U$9889 ( \10559 , \10556 , \10558 );
nand \U$9890 ( \10560 , \8908 , \8348 );
nand \U$9891 ( \10561 , \10559 , \10560 );
nor \U$9892 ( \10562 , \7560 , \10354 );
or \U$9893 ( \10563 , \10561 , \10562 );
nand \U$9894 ( \10564 , \10562 , \10561 );
nand \U$9895 ( \10565 , \10563 , \10564 );
not \U$9896 ( \10566 , \9448 );
not \U$9897 ( \10567 , \8122 );
or \U$9898 ( \10568 , \10566 , \10567 );
and \U$9899 ( \10569 , \8127 , \10447 );
or \U$9900 ( \10570 , \8360 , \9172 );
nand \U$9901 ( \10571 , \8131 , \9172 );
nand \U$9902 ( \10572 , \10570 , \10571 );
nor \U$9903 ( \10573 , \10569 , \10572 );
nand \U$9904 ( \10574 , \10568 , \10573 );
nor \U$9905 ( \10575 , \10565 , \10574 );
not \U$9906 ( \10576 , \10575 );
not \U$9907 ( \10577 , \8116 );
not \U$9908 ( \10578 , \9648 );
or \U$9909 ( \10579 , \10577 , \10578 );
nand \U$9910 ( \10580 , \10579 , \7884 );
not \U$9911 ( \10581 , \10580 );
not \U$9912 ( \10582 , \8348 );
not \U$9913 ( \10583 , \9172 );
or \U$9914 ( \10584 , \10582 , \10583 );
and \U$9915 ( \10585 , \8907 , \8493 );
not \U$9916 ( \10586 , \8907 );
and \U$9917 ( \10587 , \10586 , \8491 );
nor \U$9918 ( \10588 , \10585 , \10587 );
nand \U$9919 ( \10589 , \10584 , \10588 );
nand \U$9920 ( \10590 , \10581 , \10589 );
nand \U$9921 ( \10591 , \10565 , \10574 );
nand \U$9922 ( \10592 , \10576 , \10590 , \10591 );
not \U$9923 ( \10593 , \8493 );
nand \U$9924 ( \10594 , \10593 , \9171 );
nand \U$9925 ( \10595 , \9172 , \10090 );
nand \U$9926 ( \10596 , \10594 , \10595 , \9649 );
nand \U$9927 ( \10597 , \10596 , \9448 );
and \U$9928 ( \10598 , \9649 , \8117 );
not \U$9929 ( \10599 , \9649 );
and \U$9930 ( \10600 , \10599 , \8108 );
nor \U$9931 ( \10601 , \10598 , \10600 );
nand \U$9932 ( \10602 , \10595 , \10594 );
nand \U$9933 ( \10603 , \10602 , \10284 );
nand \U$9934 ( \10604 , \10597 , \10601 , \10603 );
not \U$9935 ( \10605 , \10589 );
not \U$9936 ( \10606 , \10580 );
and \U$9937 ( \10607 , \10605 , \10606 );
and \U$9938 ( \10608 , \10589 , \10580 );
nor \U$9939 ( \10609 , \10607 , \10608 );
or \U$9940 ( \10610 , \10604 , \10609 );
and \U$9941 ( \10611 , \8811 , \9650 );
nor \U$9942 ( \10612 , \8122 , \9650 );
nor \U$9943 ( \10613 , \10611 , \10612 );
and \U$9944 ( \10614 , \8360 , \9448 );
and \U$9945 ( \10615 , \8130 , \10447 );
nor \U$9946 ( \10616 , \10614 , \10615 );
or \U$9947 ( \10617 , \10613 , \10616 );
nand \U$9948 ( \10618 , \10609 , \10604 );
nand \U$9949 ( \10619 , \10617 , \10618 );
nand \U$9950 ( \10620 , \10610 , \10619 );
and \U$9951 ( \10621 , \10592 , \10620 );
not \U$9952 ( \10622 , \10575 );
and \U$9953 ( \10623 , \10622 , \10591 );
nor \U$9954 ( \10624 , \10623 , \10590 );
nor \U$9955 ( \10625 , \10621 , \10624 );
not \U$9956 ( \10626 , \10574 );
nand \U$9957 ( \10627 , \10626 , \10564 );
nand \U$9958 ( \10628 , \10627 , \10563 );
and \U$9959 ( \10629 , \10625 , \10628 );
nand \U$9960 ( \10630 , \10545 , \10538 );
and \U$9961 ( \10631 , \10630 , \10540 );
not \U$9962 ( \10632 , \10630 );
not \U$9963 ( \10633 , \10540 );
and \U$9964 ( \10634 , \10632 , \10633 );
nor \U$9965 ( \10635 , \10631 , \10634 );
or \U$9966 ( \10636 , \10629 , \10635 );
buf \U$9967 ( \10637 , \10625 );
or \U$9968 ( \10638 , \10637 , \10628 );
nand \U$9969 ( \10639 , \10636 , \10638 );
nand \U$9970 ( \10640 , \10555 , \10639 );
not \U$9971 ( \10641 , \10553 );
nand \U$9972 ( \10642 , \10546 , \10641 );
nand \U$9973 ( \10643 , \10640 , \10642 );
not \U$9974 ( \10644 , \10643 );
or \U$9975 ( \10645 , \10519 , \10644 );
or \U$9976 ( \10646 , \10484 , \10517 );
nand \U$9977 ( \10647 , \10645 , \10646 );
not \U$9978 ( \10648 , \10647 );
or \U$9979 ( \10649 , \10483 , \10648 );
not \U$9980 ( \10650 , \10423 );
not \U$9981 ( \10651 , \10481 );
nand \U$9982 ( \10652 , \10650 , \10651 );
nand \U$9983 ( \10653 , \10649 , \10652 );
not \U$9984 ( \10654 , \10653 );
xor \U$9985 ( \10655 , \10417 , \10419 );
and \U$9986 ( \10656 , \10655 , \10422 );
and \U$9987 ( \10657 , \10417 , \10419 );
or \U$9988 ( \10658 , \10656 , \10657 );
not \U$9989 ( \10659 , \10658 );
not \U$9990 ( \10660 , \10659 );
not \U$9991 ( \10661 , \10378 );
not \U$9992 ( \10662 , \10661 );
not \U$9993 ( \10663 , \10381 );
or \U$9994 ( \10664 , \10662 , \10663 );
nand \U$9995 ( \10665 , \10380 , \10378 );
nand \U$9996 ( \10666 , \10664 , \10665 );
not \U$9997 ( \10667 , \10666 );
not \U$9998 ( \10668 , \10667 );
or \U$9999 ( \10669 , \10660 , \10668 );
nand \U$10000 ( \10670 , \10666 , \10658 );
nand \U$10001 ( \10671 , \10669 , \10670 );
not \U$10002 ( \10672 , \10671 );
or \U$10003 ( \10673 , \10654 , \10672 );
nand \U$10004 ( \10674 , \10666 , \10659 );
nand \U$10005 ( \10675 , \10673 , \10674 );
and \U$10006 ( \10676 , \10393 , \10675 );
nor \U$10007 ( \10677 , \10389 , \10676 );
not \U$10008 ( \10678 , \10243 );
not \U$10009 ( \10679 , \10335 );
not \U$10010 ( \10680 , \10679 );
or \U$10011 ( \10681 , \10678 , \10680 );
not \U$10012 ( \10682 , \10305 );
nand \U$10013 ( \10683 , \10682 , \10334 );
nand \U$10014 ( \10684 , \10681 , \10683 );
and \U$10015 ( \10685 , \10242 , \10189 );
and \U$10016 ( \10686 , \10195 , \10241 );
nor \U$10017 ( \10687 , \10685 , \10686 );
and \U$10018 ( \10688 , \10111 , \10081 );
not \U$10019 ( \10689 , \10111 );
and \U$10020 ( \10690 , \10689 , \10082 );
or \U$10021 ( \10691 , \10688 , \10690 );
buf \U$10022 ( \10692 , \10126 );
xor \U$10023 ( \10693 , \10691 , \10692 );
nor \U$10024 ( \10694 , \10687 , \10693 );
not \U$10025 ( \10695 , \10694 );
nand \U$10026 ( \10696 , \10687 , \10693 );
nand \U$10027 ( \10697 , \10695 , \10696 );
not \U$10028 ( \10698 , \10333 );
not \U$10029 ( \10699 , \10323 );
or \U$10030 ( \10700 , \10698 , \10699 );
not \U$10031 ( \10701 , \10319 );
nand \U$10032 ( \10702 , \10701 , \10307 );
nand \U$10033 ( \10703 , \10700 , \10702 );
not \U$10034 ( \10704 , \10703 );
xor \U$10035 ( \10705 , \10136 , \10143 );
xor \U$10036 ( \10706 , \10705 , \10147 );
not \U$10037 ( \10707 , \10706 );
nand \U$10038 ( \10708 , \10704 , \10707 );
nand \U$10039 ( \10709 , \10703 , \10706 );
nand \U$10040 ( \10710 , \10708 , \10709 );
not \U$10041 ( \10711 , \10710 );
or \U$10042 ( \10712 , \7337 , \8910 );
nand \U$10043 ( \10713 , \7971 , \8910 );
not \U$10044 ( \10714 , \7341 );
not \U$10045 ( \10715 , \9173 );
and \U$10046 ( \10716 , \10714 , \10715 );
and \U$10047 ( \10717 , \7155 , \9173 );
nor \U$10048 ( \10718 , \10716 , \10717 );
nand \U$10049 ( \10719 , \10712 , \10713 , \10718 );
buf \U$10050 ( \10720 , \10719 );
not \U$10051 ( \10721 , \10720 );
and \U$10052 ( \10722 , \10711 , \10721 );
and \U$10053 ( \10723 , \10710 , \10720 );
nor \U$10054 ( \10724 , \10722 , \10723 );
and \U$10055 ( \10725 , \10697 , \10724 );
not \U$10056 ( \10726 , \10697 );
not \U$10057 ( \10727 , \10724 );
and \U$10058 ( \10728 , \10726 , \10727 );
nor \U$10059 ( \10729 , \10725 , \10728 );
xor \U$10060 ( \10730 , \10684 , \10729 );
not \U$10061 ( \10731 , \10694 );
nand \U$10062 ( \10732 , \10731 , \10724 );
and \U$10063 ( \10733 , \10732 , \10696 );
not \U$10064 ( \10734 , \10719 );
nand \U$10065 ( \10735 , \10734 , \10709 );
nand \U$10066 ( \10736 , \10735 , \10708 );
not \U$10067 ( \10737 , \10736 );
not \U$10068 ( \10738 , \9984 );
not \U$10069 ( \10739 , \9965 );
or \U$10070 ( \10740 , \10738 , \10739 );
or \U$10071 ( \10741 , \9965 , \9984 );
nand \U$10072 ( \10742 , \10740 , \10741 );
and \U$10073 ( \10743 , \10742 , \9957 );
not \U$10074 ( \10744 , \10742 );
and \U$10075 ( \10745 , \10744 , \9958 );
nor \U$10076 ( \10746 , \10743 , \10745 );
nand \U$10077 ( \10747 , \10737 , \10746 );
not \U$10078 ( \10748 , \10746 );
nand \U$10079 ( \10749 , \10748 , \10736 );
nand \U$10080 ( \10750 , \10747 , \10749 );
not \U$10081 ( \10751 , \10750 );
not \U$10082 ( \10752 , \10071 );
not \U$10083 ( \10753 , \10154 );
or \U$10084 ( \10754 , \10752 , \10753 );
or \U$10085 ( \10755 , \10071 , \10154 );
nand \U$10086 ( \10756 , \10754 , \10755 );
not \U$10087 ( \10757 , \10756 );
and \U$10088 ( \10758 , \10751 , \10757 );
and \U$10089 ( \10759 , \10756 , \10750 );
nor \U$10090 ( \10760 , \10758 , \10759 );
nor \U$10091 ( \10761 , \10733 , \10760 );
not \U$10092 ( \10762 , \10761 );
nand \U$10093 ( \10763 , \10730 , \10762 );
nor \U$10094 ( \10764 , \10677 , \10763 );
not \U$10095 ( \10765 , \9997 );
not \U$10096 ( \10766 , \10165 );
or \U$10097 ( \10767 , \10765 , \10766 );
or \U$10098 ( \10768 , \10165 , \9997 );
nand \U$10099 ( \10769 , \10767 , \10768 );
not \U$10100 ( \10770 , \10756 );
and \U$10101 ( \10771 , \10770 , \10749 );
not \U$10102 ( \10772 , \10747 );
nor \U$10103 ( \10773 , \10771 , \10772 );
nand \U$10104 ( \10774 , \10769 , \10773 );
and \U$10105 ( \10775 , \10764 , \10774 );
nand \U$10106 ( \10776 , \10729 , \10684 );
or \U$10107 ( \10777 , \10776 , \10761 );
nand \U$10108 ( \10778 , \10760 , \10733 );
nand \U$10109 ( \10779 , \10777 , \10778 );
not \U$10110 ( \10780 , \10779 );
not \U$10111 ( \10781 , \10774 );
or \U$10112 ( \10782 , \10780 , \10781 );
not \U$10113 ( \10783 , \10769 );
not \U$10114 ( \10784 , \10773 );
nand \U$10115 ( \10785 , \10783 , \10784 );
nand \U$10116 ( \10786 , \10782 , \10785 );
nor \U$10117 ( \10787 , \10775 , \10786 );
and \U$10118 ( \10788 , \10188 , \10787 );
and \U$10119 ( \10789 , \10170 , \10187 );
or \U$10120 ( \10790 , \10788 , \10789 );
xor \U$10121 ( \10791 , \9753 , \9776 );
xor \U$10122 ( \10792 , \10791 , \9779 );
xor \U$10123 ( \10793 , \10173 , \10180 );
and \U$10124 ( \10794 , \10793 , \10186 );
and \U$10125 ( \10795 , \10173 , \10180 );
or \U$10126 ( \10796 , \10794 , \10795 );
or \U$10127 ( \10797 , \10792 , \10796 );
and \U$10128 ( \10798 , \10790 , \10797 );
nand \U$10129 ( \10799 , \10792 , \10796 );
nand \U$10130 ( \10800 , \9751 , \9782 );
nand \U$10131 ( \10801 , \10799 , \10800 );
nor \U$10132 ( \10802 , \10798 , \10801 );
nor \U$10133 ( \10803 , \9930 , \9891 );
and \U$10134 ( \10804 , \10802 , \10803 , \9746 );
or \U$10135 ( \10805 , \9944 , \10804 );
or \U$10136 ( \10806 , \9897 , \9902 );
nand \U$10137 ( \10807 , \10805 , \10806 );
not \U$10138 ( \10808 , \10807 );
not \U$10139 ( \10809 , \8465 );
or \U$10140 ( \10810 , \8466 , \8646 );
nand \U$10141 ( \10811 , \10809 , \10810 , \8270 , \8674 );
not \U$10142 ( \10812 , \10811 );
nor \U$10143 ( \10813 , \7852 , \8702 );
nand \U$10144 ( \10814 , \10808 , \10812 , \10813 );
nand \U$10145 ( \10815 , \8705 , \10814 );
and \U$10146 ( \10816 , \7532 , \8696 );
xor \U$10147 ( \10817 , \7090 , \7092 );
xor \U$10148 ( \10818 , \10816 , \10817 );
and \U$10149 ( \10819 , \10815 , \10818 );
and \U$10150 ( \10820 , \10816 , \10817 );
nor \U$10151 ( \10821 , \10819 , \10820 );
not \U$10152 ( \10822 , \10821 );
or \U$10153 ( \10823 , \7099 , \10822 );
or \U$10154 ( \10824 , \10821 , \7098 );
nand \U$10155 ( \10825 , \10823 , \10824 );
nand \U$10156 ( \10826 , \6769 , \10825 );
nand \U$10157 ( \10827 , \6767 , \10826 );
buf \U$10158 ( \10828 , \10827 );
buf \U$10159 ( \10829 , \5994 );
not \U$10160 ( \10830 , \6055 );
nand \U$10161 ( \10831 , \10830 , \6070 );
nand \U$10162 ( \10832 , \10831 , \6765 );
or \U$10163 ( \10833 , \10829 , \10832 );
not \U$10164 ( \10834 , \6036 );
not \U$10165 ( \10835 , \10834 );
nor \U$10166 ( \10836 , \10831 , \6768 );
nand \U$10167 ( \10837 , \10835 , \10829 , \10836 );
xnor \U$10168 ( \10838 , \10815 , \10818 );
not \U$10169 ( \10839 , \10838 );
not \U$10170 ( \10840 , \6765 );
and \U$10171 ( \10841 , \10839 , \10840 );
not \U$10172 ( \10842 , \10832 );
and \U$10173 ( \10843 , \10834 , \10842 );
nor \U$10174 ( \10844 , \10841 , \10843 );
nand \U$10175 ( \10845 , \10833 , \10837 , \10844 );
buf \U$10176 ( \10846 , \10845 );
not \U$10177 ( \10847 , \3581 );
not \U$10178 ( \10848 , \5974 );
nand \U$10179 ( \10849 , \5482 , \10848 );
not \U$10180 ( \10850 , \10849 );
not \U$10181 ( \10851 , \4445 );
or \U$10182 ( \10852 , \10850 , \10851 );
nand \U$10183 ( \10853 , \10852 , \5992 );
nand \U$10184 ( \10854 , \10853 , \3432 );
and \U$10185 ( \10855 , \5958 , \4444 );
nor \U$10186 ( \10856 , \4004 , \4222 );
and \U$10187 ( \10857 , \10855 , \10856 , \3431 );
not \U$10188 ( \10858 , \5479 );
nand \U$10189 ( \10859 , \5486 , \5952 , \5218 , \5480 );
not \U$10190 ( \10860 , \10859 );
not \U$10191 ( \10861 , \10860 );
or \U$10192 ( \10862 , \10858 , \10861 );
buf \U$10193 ( \10863 , \5965 );
not \U$10194 ( \10864 , \10863 );
nand \U$10195 ( \10865 , \10862 , \10864 );
and \U$10196 ( \10866 , \10857 , \10865 );
nor \U$10197 ( \10867 , \10866 , \6019 );
nand \U$10198 ( \10868 , \10854 , \10867 );
not \U$10199 ( \10869 , \10868 );
or \U$10200 ( \10870 , \10847 , \10869 );
nand \U$10201 ( \10871 , \10870 , \6032 );
not \U$10202 ( \10872 , \3618 );
nor \U$10203 ( \10873 , \10872 , \6035 );
nand \U$10204 ( \10874 , \10873 , \6765 );
or \U$10205 ( \10875 , \10871 , \10874 );
nor \U$10206 ( \10876 , \10873 , \6768 );
nand \U$10207 ( \10877 , \10871 , \10876 );
nand \U$10208 ( \10878 , \8703 , \8698 );
not \U$10209 ( \10879 , \10878 );
not \U$10210 ( \10880 , \7853 );
not \U$10211 ( \10881 , \10807 );
not \U$10212 ( \10882 , \10811 );
and \U$10213 ( \10883 , \10881 , \10882 );
nor \U$10214 ( \10884 , \10883 , \8676 );
not \U$10215 ( \10885 , \10884 );
not \U$10216 ( \10886 , \10885 );
or \U$10217 ( \10887 , \10880 , \10886 );
nand \U$10218 ( \10888 , \10887 , \8689 );
not \U$10219 ( \10889 , \10888 );
or \U$10220 ( \10890 , \10879 , \10889 );
or \U$10221 ( \10891 , \10888 , \10878 );
nand \U$10222 ( \10892 , \10890 , \10891 );
nand \U$10223 ( \10893 , \10892 , \6764 );
nand \U$10224 ( \10894 , \10875 , \10877 , \10893 );
buf \U$10225 ( \10895 , \10894 );
not \U$10226 ( \10896 , \3549 );
not \U$10227 ( \10897 , \10896 );
not \U$10228 ( \10898 , \10868 );
or \U$10229 ( \10899 , \10897 , \10898 );
not \U$10230 ( \10900 , \6027 );
nand \U$10231 ( \10901 , \10899 , \10900 );
not \U$10232 ( \10902 , \6030 );
nor \U$10233 ( \10903 , \10902 , \3580 );
nand \U$10234 ( \10904 , \10903 , \6765 );
or \U$10235 ( \10905 , \10901 , \10904 );
nor \U$10236 ( \10906 , \10903 , \6764 );
nand \U$10237 ( \10907 , \10901 , \10906 );
not \U$10238 ( \10908 , \6765 );
not \U$10239 ( \10909 , \7535 );
not \U$10240 ( \10910 , \7503 );
and \U$10241 ( \10911 , \10909 , \10910 );
and \U$10242 ( \10912 , \7535 , \7503 );
nor \U$10243 ( \10913 , \10911 , \10912 );
not \U$10244 ( \10914 , \10913 );
not \U$10245 ( \10915 , \7851 );
not \U$10246 ( \10916 , \7842 );
nor \U$10247 ( \10917 , \10884 , \10916 );
not \U$10248 ( \10918 , \10917 );
or \U$10249 ( \10919 , \10915 , \10918 );
not \U$10250 ( \10920 , \8684 );
nand \U$10251 ( \10921 , \10919 , \10920 );
not \U$10252 ( \10922 , \10921 );
or \U$10253 ( \10923 , \10914 , \10922 );
or \U$10254 ( \10924 , \10921 , \10913 );
nand \U$10255 ( \10925 , \10923 , \10924 );
nand \U$10256 ( \10926 , \10908 , \10925 );
nand \U$10257 ( \10927 , \10905 , \10907 , \10926 );
buf \U$10258 ( \10928 , \10927 );
not \U$10259 ( \10929 , \3548 );
not \U$10260 ( \10930 , \10868 );
or \U$10261 ( \10931 , \10929 , \10930 );
nand \U$10262 ( \10932 , \10931 , \6024 );
xor \U$10263 ( \10933 , \3484 , \3535 );
nand \U$10264 ( \10934 , \10933 , \6765 );
or \U$10265 ( \10935 , \10932 , \10934 );
not \U$10266 ( \10936 , \7842 );
not \U$10267 ( \10937 , \10885 );
or \U$10268 ( \10938 , \10936 , \10937 );
not \U$10269 ( \10939 , \8680 );
nand \U$10270 ( \10940 , \10938 , \10939 );
nand \U$10271 ( \10941 , \7851 , \8683 );
and \U$10272 ( \10942 , \10940 , \10941 );
not \U$10273 ( \10943 , \10940 );
not \U$10274 ( \10944 , \10941 );
and \U$10275 ( \10945 , \10943 , \10944 );
nor \U$10276 ( \10946 , \10942 , \10945 );
or \U$10277 ( \10947 , \10946 , \6765 );
nor \U$10278 ( \10948 , \10933 , \6769 );
nand \U$10279 ( \10949 , \10932 , \10948 );
nand \U$10280 ( \10950 , \10935 , \10947 , \10949 );
buf \U$10281 ( \10951 , \10950 );
nand \U$10282 ( \10952 , \6024 , \3548 );
xor \U$10283 ( \10953 , \10952 , \10868 );
or \U$10284 ( \10954 , \10953 , \6764 );
nand \U$10285 ( \10955 , \10939 , \7842 );
xor \U$10286 ( \10956 , \10955 , \10885 );
or \U$10287 ( \10957 , \10956 , \6765 );
nand \U$10288 ( \10958 , \10954 , \10957 );
buf \U$10289 ( \10959 , \10958 );
buf \U$10290 ( \10960 , \2979 );
not \U$10291 ( \10961 , \10960 );
not \U$10292 ( \10962 , \3430 );
and \U$10293 ( \10963 , \10962 , \4223 , \4444 , \4005 );
not \U$10294 ( \10964 , \10963 );
not \U$10295 ( \10965 , \5976 );
or \U$10296 ( \10966 , \10964 , \10965 );
and \U$10297 ( \10967 , \5991 , \10962 );
not \U$10298 ( \10968 , \6002 );
nor \U$10299 ( \10969 , \10967 , \10968 );
nand \U$10300 ( \10970 , \10966 , \10969 );
not \U$10301 ( \10971 , \10970 );
or \U$10302 ( \10972 , \10961 , \10971 );
nand \U$10303 ( \10973 , \10972 , \6013 );
nand \U$10304 ( \10974 , \6018 , \2714 );
xor \U$10305 ( \10975 , \10973 , \10974 );
and \U$10306 ( \10976 , \6765 , \10975 );
not \U$10307 ( \10977 , \6765 );
buf \U$10308 ( \10978 , \8270 );
not \U$10309 ( \10979 , \10978 );
not \U$10310 ( \10980 , \10808 );
not \U$10311 ( \10981 , \8465 );
nand \U$10312 ( \10982 , \10981 , \10810 );
or \U$10313 ( \10983 , \10980 , \10982 );
not \U$10314 ( \10984 , \8654 );
nand \U$10315 ( \10985 , \10983 , \10984 );
not \U$10316 ( \10986 , \10985 );
or \U$10317 ( \10987 , \10979 , \10986 );
nand \U$10318 ( \10988 , \10987 , \8660 );
nand \U$10319 ( \10989 , \8674 , \8671 );
xor \U$10320 ( \10990 , \10988 , \10989 );
and \U$10321 ( \10991 , \10977 , \10990 );
nor \U$10322 ( \10992 , \10976 , \10991 );
buf \U$10323 ( \10993 , \10992 );
not \U$10324 ( \10994 , \10985 );
nand \U$10325 ( \10995 , \8660 , \10978 );
not \U$10326 ( \10996 , \10995 );
and \U$10327 ( \10997 , \10994 , \10996 );
and \U$10328 ( \10998 , \10995 , \10985 );
nor \U$10329 ( \10999 , \10997 , \10998 );
and \U$10330 ( \11000 , \6769 , \10999 );
not \U$10331 ( \11001 , \6769 );
nand \U$10332 ( \11002 , \10960 , \6013 );
and \U$10333 ( \11003 , \10970 , \11002 );
not \U$10334 ( \11004 , \10970 );
not \U$10335 ( \11005 , \11002 );
and \U$10336 ( \11006 , \11004 , \11005 );
nor \U$10337 ( \11007 , \11003 , \11006 );
and \U$10338 ( \11008 , \11001 , \11007 );
nor \U$10339 ( \11009 , \11000 , \11008 );
buf \U$10340 ( \11010 , \11009 );
not \U$10341 ( \11011 , \8466 );
not \U$10342 ( \11012 , \8646 );
or \U$10343 ( \11013 , \11011 , \11012 );
not \U$10344 ( \11014 , \10810 );
or \U$10345 ( \11015 , \10980 , \11014 );
nand \U$10346 ( \11016 , \11013 , \11015 );
not \U$10347 ( \11017 , \11016 );
nand \U$10348 ( \11018 , \10981 , \8653 );
not \U$10349 ( \11019 , \11018 );
and \U$10350 ( \11020 , \11017 , \11019 );
and \U$10351 ( \11021 , \11016 , \11018 );
nor \U$10352 ( \11022 , \11020 , \11021 );
and \U$10353 ( \11023 , \6764 , \11022 );
not \U$10354 ( \11024 , \6764 );
not \U$10355 ( \11025 , \3422 );
not \U$10356 ( \11026 , \5993 );
or \U$10357 ( \11027 , \11025 , \11026 );
buf \U$10358 ( \11028 , \6000 );
buf \U$10359 ( \11029 , \11028 );
nand \U$10360 ( \11030 , \11027 , \11029 );
nand \U$10361 ( \11031 , \5999 , \3429 );
xor \U$10362 ( \11032 , \11030 , \11031 );
and \U$10363 ( \11033 , \11024 , \11032 );
nor \U$10364 ( \11034 , \11023 , \11033 );
buf \U$10365 ( \11035 , \11034 );
nand \U$10366 ( \11036 , \3422 , \11028 );
xor \U$10367 ( \11037 , \5993 , \11036 );
or \U$10368 ( \11038 , \11037 , \6764 );
nand \U$10369 ( \11039 , \8647 , \10810 );
xnor \U$10370 ( \11040 , \10980 , \11039 );
or \U$10371 ( \11041 , \11040 , \6765 );
nand \U$10372 ( \11042 , \11038 , \11041 );
buf \U$10373 ( \11043 , \11042 );
not \U$10374 ( \11044 , \4223 );
not \U$10375 ( \11045 , \5481 );
not \U$10376 ( \11046 , \5446 );
or \U$10377 ( \11047 , \11045 , \11046 );
nand \U$10378 ( \11048 , \11047 , \10859 );
nand \U$10379 ( \11049 , \11048 , \5479 );
not \U$10380 ( \11050 , \10855 );
or \U$10381 ( \11051 , \11049 , \11050 );
and \U$10382 ( \11052 , \10855 , \10863 );
not \U$10383 ( \11053 , \4444 );
or \U$10384 ( \11054 , \10848 , \11053 );
not \U$10385 ( \11055 , \5979 );
nand \U$10386 ( \11056 , \11054 , \11055 );
nor \U$10387 ( \11057 , \11052 , \11056 );
nand \U$10388 ( \11058 , \11051 , \11057 );
not \U$10389 ( \11059 , \11058 );
or \U$10390 ( \11060 , \11044 , \11059 );
not \U$10391 ( \11061 , \5982 );
nand \U$10392 ( \11062 , \11060 , \11061 );
buf \U$10393 ( \11063 , \3992 );
nand \U$10394 ( \11064 , \11062 , \11063 );
xnor \U$10395 ( \11065 , \5989 , \5988 );
buf \U$10396 ( \11066 , \5983 );
not \U$10397 ( \11067 , \11066 );
nand \U$10398 ( \11068 , \11067 , \6765 );
nor \U$10399 ( \11069 , \11065 , \11068 );
and \U$10400 ( \11070 , \11064 , \11069 );
and \U$10401 ( \11071 , \11065 , \11066 , \6765 );
nor \U$10402 ( \11072 , \11070 , \11071 );
and \U$10403 ( \11073 , \11065 , \6765 );
and \U$10404 ( \11074 , \11062 , \11073 , \11063 );
not \U$10405 ( \11075 , \9891 );
not \U$10406 ( \11076 , \11075 );
not \U$10407 ( \11077 , \9931 );
not \U$10408 ( \11078 , \9746 );
not \U$10409 ( \11079 , \10802 );
or \U$10410 ( \11080 , \11078 , \11079 );
buf \U$10411 ( \11081 , \9745 );
and \U$10412 ( \11082 , \9787 , \11081 );
and \U$10413 ( \11083 , \9465 , \9557 );
and \U$10414 ( \11084 , \11082 , \11083 );
nor \U$10415 ( \11085 , \11084 , \9796 );
nand \U$10416 ( \11086 , \11080 , \11085 );
not \U$10417 ( \11087 , \11086 );
or \U$10418 ( \11088 , \11077 , \11087 );
nand \U$10419 ( \11089 , \11088 , \9939 );
not \U$10420 ( \11090 , \11089 );
or \U$10421 ( \11091 , \11076 , \11090 );
buf \U$10422 ( \11092 , \9940 );
nand \U$10423 ( \11093 , \11091 , \11092 );
nand \U$10424 ( \11094 , \9903 , \10806 );
xor \U$10425 ( \11095 , \11093 , \11094 );
buf \U$10426 ( \11096 , \6765 );
nor \U$10427 ( \11097 , \11095 , \11096 );
nor \U$10428 ( \11098 , \11074 , \11097 );
nand \U$10429 ( \11099 , \11072 , \11098 );
buf \U$10430 ( \11100 , \11099 );
nand \U$10431 ( \11101 , \11092 , \11075 );
xor \U$10432 ( \11102 , \11089 , \11101 );
and \U$10433 ( \11103 , \6764 , \11102 );
not \U$10434 ( \11104 , \6764 );
not \U$10435 ( \11105 , \11062 );
nand \U$10436 ( \11106 , \11063 , \11067 );
not \U$10437 ( \11107 , \11106 );
and \U$10438 ( \11108 , \11105 , \11107 );
and \U$10439 ( \11109 , \11062 , \11106 );
nor \U$10440 ( \11110 , \11108 , \11109 );
and \U$10441 ( \11111 , \11104 , \11110 );
nor \U$10442 ( \11112 , \11103 , \11111 );
buf \U$10443 ( \11113 , \11112 );
buf \U$10444 ( \11114 , \4220 );
not \U$10445 ( \11115 , \4007 );
xor \U$10446 ( \11116 , \11114 , \11115 );
buf \U$10447 ( \11117 , \11058 );
xor \U$10448 ( \11118 , \11116 , \11117 );
or \U$10449 ( \11119 , \11118 , \6769 );
not \U$10450 ( \11120 , \9929 );
not \U$10451 ( \11121 , \11086 );
or \U$10452 ( \11122 , \11120 , \11121 );
not \U$10453 ( \11123 , \9934 );
nand \U$10454 ( \11124 , \11122 , \11123 );
nand \U$10455 ( \11125 , \9922 , \9938 );
xor \U$10456 ( \11126 , \11124 , \11125 );
or \U$10457 ( \11127 , \11126 , \6765 );
nand \U$10458 ( \11128 , \11119 , \11127 );
buf \U$10459 ( \11129 , \11128 );
nand \U$10460 ( \11130 , \11123 , \9929 );
xor \U$10461 ( \11131 , \11086 , \11130 );
and \U$10462 ( \11132 , \6768 , \11131 );
not \U$10463 ( \11133 , \6768 );
xnor \U$10464 ( \11134 , \4229 , \4443 );
xor \U$10465 ( \11135 , \11134 , \5976 );
and \U$10466 ( \11136 , \11133 , \11135 );
nor \U$10467 ( \11137 , \11132 , \11136 );
buf \U$10468 ( \11138 , \11137 );
not \U$10469 ( \11139 , \5479 );
not \U$10470 ( \11140 , \11048 );
or \U$10471 ( \11141 , \11139 , \11140 );
nand \U$10472 ( \11142 , \11141 , \10864 );
buf \U$10473 ( \11143 , \4731 );
and \U$10474 ( \11144 , \11142 , \11143 );
buf \U$10475 ( \11145 , \5967 );
nor \U$10476 ( \11146 , \11144 , \11145 );
nand \U$10477 ( \11147 , \5973 , \4746 );
not \U$10478 ( \11148 , \11147 );
and \U$10479 ( \11149 , \11146 , \11148 );
not \U$10480 ( \11150 , \11146 );
and \U$10481 ( \11151 , \11150 , \11147 );
nor \U$10482 ( \11152 , \11149 , \11151 );
or \U$10483 ( \11153 , \11152 , \6769 );
and \U$10484 ( \11154 , \9795 , \9557 );
not \U$10485 ( \11155 , \11154 );
not \U$10486 ( \11156 , \11081 );
buf \U$10487 ( \11157 , \10802 );
not \U$10488 ( \11158 , \11157 );
or \U$10489 ( \11159 , \11156 , \11158 );
not \U$10490 ( \11160 , \11082 );
nand \U$10491 ( \11161 , \11159 , \11160 );
and \U$10492 ( \11162 , \11161 , \9465 );
not \U$10493 ( \11163 , \9791 );
nor \U$10494 ( \11164 , \11162 , \11163 );
not \U$10495 ( \11165 , \11164 );
and \U$10496 ( \11166 , \11155 , \11165 );
and \U$10497 ( \11167 , \11164 , \11154 );
nor \U$10498 ( \11168 , \11166 , \11167 );
or \U$10499 ( \11169 , \11168 , \6765 );
nand \U$10500 ( \11170 , \11153 , \11169 );
buf \U$10501 ( \11171 , \11170 );
not \U$10502 ( \11172 , \11161 );
xor \U$10503 ( \11173 , \9790 , \9464 );
not \U$10504 ( \11174 , \11173 );
and \U$10505 ( \11175 , \11172 , \11174 );
and \U$10506 ( \11176 , \11161 , \11173 );
nor \U$10507 ( \11177 , \11175 , \11176 );
and \U$10508 ( \11178 , \6764 , \11177 );
not \U$10509 ( \11179 , \6764 );
not \U$10510 ( \11180 , \11145 );
nand \U$10511 ( \11181 , \11180 , \11143 );
and \U$10512 ( \11182 , \11142 , \11181 );
not \U$10513 ( \11183 , \11142 );
not \U$10514 ( \11184 , \11181 );
and \U$10515 ( \11185 , \11183 , \11184 );
nor \U$10516 ( \11186 , \11182 , \11185 );
and \U$10517 ( \11187 , \11179 , \11186 );
nor \U$10518 ( \11188 , \11178 , \11187 );
buf \U$10519 ( \11189 , \11188 );
buf \U$10520 ( \11190 , \11048 );
buf \U$10521 ( \11191 , \5477 );
and \U$10522 ( \11192 , \11190 , \11191 );
not \U$10523 ( \11193 , \5962 );
nor \U$10524 ( \11194 , \11192 , \11193 );
nand \U$10525 ( \11195 , \5960 , \5469 );
not \U$10526 ( \11196 , \11195 );
and \U$10527 ( \11197 , \11194 , \11196 );
not \U$10528 ( \11198 , \11194 );
and \U$10529 ( \11199 , \11198 , \11195 );
nor \U$10530 ( \11200 , \11197 , \11199 );
or \U$10531 ( \11201 , \11200 , \6764 );
not \U$10532 ( \11202 , \11157 );
nand \U$10533 ( \11203 , \11202 , \9783 );
nand \U$10534 ( \11204 , \9786 , \11081 );
xor \U$10535 ( \11205 , \11203 , \11204 );
or \U$10536 ( \11206 , \11205 , \6765 );
nand \U$10537 ( \11207 , \11201 , \11206 );
buf \U$10538 ( \11208 , \11207 );
buf \U$10539 ( \11209 , \10790 );
not \U$10540 ( \11210 , \11209 );
and \U$10541 ( \11211 , \11210 , \10799 );
not \U$10542 ( \11212 , \10797 );
nor \U$10543 ( \11213 , \11211 , \11212 );
not \U$10544 ( \11214 , \11213 );
and \U$10545 ( \11215 , \9783 , \10800 );
not \U$10546 ( \11216 , \11215 );
and \U$10547 ( \11217 , \11214 , \11216 );
and \U$10548 ( \11218 , \11213 , \11215 );
nor \U$10549 ( \11219 , \11217 , \11218 );
and \U$10550 ( \11220 , \6764 , \11219 );
not \U$10551 ( \11221 , \6764 );
nand \U$10552 ( \11222 , \5962 , \11191 );
and \U$10553 ( \11223 , \11190 , \11222 );
not \U$10554 ( \11224 , \11190 );
not \U$10555 ( \11225 , \11222 );
and \U$10556 ( \11226 , \11224 , \11225 );
nor \U$10557 ( \11227 , \11223 , \11226 );
and \U$10558 ( \11228 , \11221 , \11227 );
nor \U$10559 ( \11229 , \11220 , \11228 );
buf \U$10560 ( \11230 , \11229 );
not \U$10561 ( \11231 , \5218 );
not \U$10562 ( \11232 , \5952 );
not \U$10563 ( \11233 , \5486 );
or \U$10564 ( \11234 , \11232 , \11233 );
nand \U$10565 ( \11235 , \11234 , \5404 );
not \U$10566 ( \11236 , \11235 );
or \U$10567 ( \11237 , \11231 , \11236 );
not \U$10568 ( \11238 , \5444 );
nand \U$10569 ( \11239 , \11237 , \11238 );
not \U$10570 ( \11240 , \5443 );
nand \U$10571 ( \11241 , \11240 , \5481 );
xor \U$10572 ( \11242 , \11239 , \11241 );
and \U$10573 ( \11243 , \6765 , \11242 );
not \U$10574 ( \11244 , \6765 );
not \U$10575 ( \11245 , \11209 );
not \U$10576 ( \11246 , \10799 );
nor \U$10577 ( \11247 , \11246 , \11212 );
not \U$10578 ( \11248 , \11247 );
and \U$10579 ( \11249 , \11245 , \11248 );
and \U$10580 ( \11250 , \11209 , \11247 );
nor \U$10581 ( \11251 , \11249 , \11250 );
and \U$10582 ( \11252 , \11244 , \11251 );
nor \U$10583 ( \11253 , \11243 , \11252 );
buf \U$10584 ( \11254 , \11253 );
nand \U$10585 ( \11255 , \11238 , \5218 );
and \U$10586 ( \11256 , \11235 , \11255 );
not \U$10587 ( \11257 , \11235 );
not \U$10588 ( \11258 , \11255 );
and \U$10589 ( \11259 , \11257 , \11258 );
nor \U$10590 ( \11260 , \11256 , \11259 );
or \U$10591 ( \11261 , \11260 , \6768 );
xor \U$10592 ( \11262 , \10170 , \10187 );
xor \U$10593 ( \11263 , \11262 , \10787 );
or \U$10594 ( \11264 , \11263 , \6765 );
nand \U$10595 ( \11265 , \11261 , \11264 );
buf \U$10596 ( \11266 , \11265 );
buf \U$10597 ( \11267 , \10677 );
not \U$10598 ( \11268 , \10730 );
or \U$10599 ( \11269 , \11267 , \11268 );
nand \U$10600 ( \11270 , \11269 , \10776 );
and \U$10601 ( \11271 , \11270 , \10762 );
not \U$10602 ( \11272 , \10778 );
nor \U$10603 ( \11273 , \11271 , \11272 );
nand \U$10604 ( \11274 , \10785 , \10774 );
xnor \U$10605 ( \11275 , \11273 , \11274 );
and \U$10606 ( \11276 , \6764 , \11275 );
not \U$10607 ( \11277 , \6764 );
buf \U$10608 ( \11278 , \5401 );
not \U$10609 ( \11279 , \11278 );
not \U$10610 ( \11280 , \5402 );
and \U$10611 ( \11281 , \11279 , \11280 );
and \U$10612 ( \11282 , \11278 , \5402 );
nor \U$10613 ( \11283 , \11281 , \11282 );
not \U$10614 ( \11284 , \5485 );
not \U$10615 ( \11285 , \5952 );
or \U$10616 ( \11286 , \11284 , \11285 );
buf \U$10617 ( \11287 , \5399 );
nand \U$10618 ( \11288 , \11286 , \11287 );
not \U$10619 ( \11289 , \11288 );
and \U$10620 ( \11290 , \11283 , \11289 );
not \U$10621 ( \11291 , \11283 );
and \U$10622 ( \11292 , \11291 , \11288 );
nor \U$10623 ( \11293 , \11290 , \11292 );
and \U$10624 ( \11294 , \11277 , \11293 );
nor \U$10625 ( \11295 , \11276 , \11294 );
buf \U$10626 ( \11296 , \11295 );
and \U$10627 ( \11297 , \5399 , \5485 );
xnor \U$10628 ( \11298 , \11297 , \5952 );
or \U$10629 ( \11299 , \11298 , \6764 );
not \U$10630 ( \11300 , \11270 );
nand \U$10631 ( \11301 , \10778 , \10762 );
not \U$10632 ( \11302 , \11301 );
and \U$10633 ( \11303 , \11300 , \11302 );
and \U$10634 ( \11304 , \11270 , \11301 );
nor \U$10635 ( \11305 , \11303 , \11304 );
or \U$10636 ( \11306 , \11305 , \6765 );
nand \U$10637 ( \11307 , \11299 , \11306 );
buf \U$10638 ( \11308 , \11307 );
nand \U$10639 ( \11309 , \5951 , \5566 );
buf \U$10640 ( \11310 , \5946 );
and \U$10641 ( \11311 , \11309 , \11310 );
not \U$10642 ( \11312 , \11309 );
not \U$10643 ( \11313 , \11310 );
and \U$10644 ( \11314 , \11312 , \11313 );
nor \U$10645 ( \11315 , \11311 , \11314 );
or \U$10646 ( \11316 , \11315 , \6764 );
xnor \U$10647 ( \11317 , \11268 , \11267 );
or \U$10648 ( \11318 , \11317 , \6765 );
nand \U$10649 ( \11319 , \11316 , \11318 );
buf \U$10650 ( \11320 , \11319 );
nand \U$10651 ( \11321 , \5945 , \5633 );
xor \U$10652 ( \11322 , \11321 , \5939 );
or \U$10653 ( \11323 , \11322 , \6764 );
xnor \U$10654 ( \11324 , \10675 , \10393 );
or \U$10655 ( \11325 , \11324 , \6765 );
nand \U$10656 ( \11326 , \11323 , \11325 );
buf \U$10657 ( \11327 , \11326 );
xnor \U$10658 ( \11328 , \5918 , \5934 );
or \U$10659 ( \11329 , \11328 , \6764 );
buf \U$10660 ( \11330 , \10653 );
xnor \U$10661 ( \11331 , \10671 , \11330 );
or \U$10662 ( \11332 , \11331 , \6765 );
nand \U$10663 ( \11333 , \11329 , \11332 );
buf \U$10664 ( \11334 , \11333 );
not \U$10665 ( \11335 , \10647 );
nand \U$10666 ( \11336 , \10482 , \10652 );
not \U$10667 ( \11337 , \11336 );
and \U$10668 ( \11338 , \11335 , \11337 );
and \U$10669 ( \11339 , \10647 , \11336 );
nor \U$10670 ( \11340 , \11338 , \11339 );
and \U$10671 ( \11341 , \6763 , \11340 );
not \U$10672 ( \11342 , \6763 );
nand \U$10673 ( \11343 , \5713 , \5917 );
and \U$10674 ( \11344 , \11343 , \5912 );
not \U$10675 ( \11345 , \11343 );
not \U$10676 ( \11346 , \5912 );
and \U$10677 ( \11347 , \11345 , \11346 );
nor \U$10678 ( \11348 , \11344 , \11347 );
and \U$10679 ( \11349 , \11342 , \11348 );
nor \U$10680 ( \11350 , \11341 , \11349 );
buf \U$10681 ( \11351 , \11350 );
nand \U$10682 ( \11352 , \10646 , \10518 );
xor \U$10683 ( \11353 , \11352 , \10643 );
and \U$10684 ( \11354 , \6763 , \11353 );
not \U$10685 ( \11355 , \6763 );
and \U$10686 ( \11356 , \5765 , \5910 );
not \U$10687 ( \11357 , \5765 );
and \U$10688 ( \11358 , \11357 , \5758 );
nor \U$10689 ( \11359 , \11356 , \11358 );
xor \U$10690 ( \11360 , \5907 , \11359 );
and \U$10691 ( \11361 , \11355 , \11360 );
nor \U$10692 ( \11362 , \11354 , \11361 );
buf \U$10693 ( \11363 , \11362 );
nand \U$10694 ( \11364 , RIaaa9218_606, RIaaa90b0_603, RIaaa9128_604, RIaaa91a0_605);
not \U$10695 ( \11365 , \11364 );
and \U$10696 ( \11366 , \11365 , RIaaa9380_609, RIaaa9308_608, RIaaa9290_607);
not \U$10697 ( \11367 , \11366 );
nand \U$10698 ( \11368 , RIaaa9038_602, RIaaa93f8_610, RIaaa9470_611, RIaaa94e8_612);
nor \U$10699 ( \11369 , \11367 , \11368 );
and \U$10700 ( \11370 , RIaaa95d8_614, \11369 );
not \U$10701 ( \11371 , RIaa9b0a0_125);
nor \U$10702 ( \11372 , RIaaa8c78_594, RIaaa8cf0_595);
nor \U$10703 ( \11373 , RIaaa8a98_590, RIaaa8b10_591);
not \U$10704 ( \11374 , RIaaa8a20_589);
nand \U$10705 ( \11375 , \11372 , \11373 , \11374 );
not \U$10706 ( \11376 , \11375 );
nor \U$10707 ( \11377 , RIaaa8b88_592, RIaaa8c00_593);
nor \U$10708 ( \11378 , RIaaa8d68_596, RIaaa8de0_597);
nand \U$10709 ( \11379 , \11377 , \11378 );
not \U$10710 ( \11380 , \11379 );
and \U$10711 ( \11381 , RIaaa8e58_598, RIaaa8ed0_599);
nand \U$10712 ( \11382 , RIaaa8f48_600, RIaaa8fc0_601);
nor \U$10713 ( \11383 , \11381 , \11382 );
nand \U$10714 ( \11384 , \11376 , \11380 , \11383 );
and \U$10715 ( \11385 , \11384 , RIaaa8ed0_599);
not \U$10716 ( \11386 , \11384 );
not \U$10717 ( \11387 , RIaaa8ed0_599);
and \U$10718 ( \11388 , \11386 , \11387 );
or \U$10719 ( \11389 , \11385 , \11388 );
not \U$10720 ( \11390 , \11389 );
not \U$10721 ( \11391 , \11390 );
not \U$10722 ( \11392 , RIaaa8ed0_599);
not \U$10723 ( \11393 , \11384 );
not \U$10724 ( \11394 , \11393 );
or \U$10725 ( \11395 , \11392 , \11394 );
not \U$10726 ( \11396 , RIaaa8e58_598);
nand \U$10727 ( \11397 , \11395 , \11396 );
buf \U$10728 ( \11398 , \11397 );
buf \U$10729 ( \11399 , \11398 );
not \U$10730 ( \11400 , \11399 );
buf \U$10731 ( \11401 , \11393 );
not \U$10732 ( \11402 , \11401 );
not \U$10733 ( \11403 , RIaaa8f48_600);
not \U$10734 ( \11404 , RIaaa8fc0_601);
nand \U$10735 ( \11405 , RIaaa8ed0_599, RIaaa8f48_600);
not \U$10736 ( \11406 , \11405 );
or \U$10737 ( \11407 , \11404 , \11406 );
not \U$10738 ( \11408 , RIaaa8e58_598);
nand \U$10739 ( \11409 , \11408 , RIaaa8fc0_601);
nand \U$10740 ( \11410 , \11407 , \11409 );
and \U$10741 ( \11411 , \11376 , \11410 , \11380 );
not \U$10742 ( \11412 , \11411 );
nand \U$10743 ( \11413 , \11403 , \11412 );
nand \U$10744 ( \11414 , \11402 , \11413 );
buf \U$10745 ( \11415 , \11414 );
buf \U$10746 ( \11416 , \11376 );
nand \U$10747 ( \11417 , \11416 , \11380 );
not \U$10748 ( \11418 , RIaaa8fc0_601);
nand \U$10749 ( \11419 , \11417 , \11418 );
nand \U$10750 ( \11420 , \11412 , \11419 );
buf \U$10751 ( \11421 , \11420 );
nand \U$10752 ( \11422 , \11391 , \11400 , \11415 , \11421 );
not \U$10753 ( \11423 , \11422 );
not \U$10754 ( \11424 , \11423 );
or \U$10755 ( \11425 , \11371 , \11424 );
not \U$10756 ( \11426 , \11389 );
not \U$10757 ( \11427 , \11426 );
not \U$10758 ( \11428 , \11398 );
not \U$10759 ( \11429 , \11428 );
buf \U$10760 ( \11430 , \11414 );
nand \U$10761 ( \11431 , \11427 , \11429 , \11430 , \11421 );
not \U$10762 ( \11432 , \11431 );
nand \U$10763 ( \11433 , \11432 , RIaa9b280_129);
nand \U$10764 ( \11434 , \11425 , \11433 );
not \U$10765 ( \11435 , RIaa9b3e8_132);
not \U$10766 ( \11436 , \11389 );
not \U$10767 ( \11437 , \11436 );
not \U$10768 ( \11438 , \11398 );
not \U$10769 ( \11439 , \11438 );
not \U$10770 ( \11440 , \11439 );
not \U$10771 ( \11441 , \11411 );
not \U$10772 ( \11442 , RIaaa8f48_600);
and \U$10773 ( \11443 , \11441 , \11442 );
nor \U$10774 ( \11444 , \11443 , \11401 );
buf \U$10775 ( \11445 , \11444 );
and \U$10776 ( \11446 , \11412 , \11419 );
buf \U$10777 ( \11447 , \11446 );
nand \U$10778 ( \11448 , \11437 , \11440 , \11445 , \11447 );
not \U$10779 ( \11449 , \11448 );
not \U$10780 ( \11450 , \11449 );
or \U$10781 ( \11451 , \11435 , \11450 );
not \U$10782 ( \11452 , \11398 );
not \U$10783 ( \11453 , \11452 );
buf \U$10784 ( \11454 , \11389 );
not \U$10785 ( \11455 , \11454 );
nand \U$10786 ( \11456 , \11453 , \11455 , \11415 , \11447 );
not \U$10787 ( \11457 , \11456 );
nand \U$10788 ( \11458 , \11457 , RIaa9b4d8_134);
nand \U$10789 ( \11459 , \11451 , \11458 );
nor \U$10790 ( \11460 , \11434 , \11459 );
buf \U$10791 ( \11461 , \11446 );
nand \U$10792 ( \11462 , \11461 , \11454 , \11445 , \11399 );
not \U$10793 ( \11463 , \11462 );
nand \U$10794 ( \11464 , \11463 , RIaa9b028_124);
not \U$10795 ( \11465 , \11380 );
and \U$10796 ( \11466 , \11373 , \11372 );
not \U$10797 ( \11467 , \11466 );
or \U$10798 ( \11468 , \11465 , \11467 );
nor \U$10799 ( \11469 , RIaaa8ed0_599, RIaaa8fc0_601);
nor \U$10800 ( \11470 , RIaaa8e58_598, RIaaa8f48_600);
and \U$10801 ( \11471 , \11374 , \11469 , \11470 );
nand \U$10802 ( \11472 , \11468 , \11471 );
not \U$10803 ( \11473 , \11472 );
nand \U$10804 ( \11474 , \11473 , RIaa9aec0_121);
nand \U$10805 ( \11475 , RIaa9af38_122, RIaaa8a20_589);
nand \U$10806 ( \11476 , \11464 , \11474 , \11475 );
not \U$10807 ( \11477 , RIaa9b208_128);
not \U$10808 ( \11478 , \11399 );
nand \U$10809 ( \11479 , \11454 , \11478 , \11445 , \11421 );
not \U$10810 ( \11480 , \11479 );
not \U$10811 ( \11481 , \11480 );
or \U$10812 ( \11482 , \11477 , \11481 );
and \U$10813 ( \11483 , \11390 , \11439 );
and \U$10814 ( \11484 , \11414 , \11421 );
nand \U$10815 ( \11485 , \11483 , \11484 );
not \U$10816 ( \11486 , \11485 );
nand \U$10817 ( \11487 , \11486 , RIaa9b460_133);
nand \U$10818 ( \11488 , \11482 , \11487 );
nor \U$10819 ( \11489 , \11476 , \11488 );
not \U$10820 ( \11490 , RIaa9afb0_123);
not \U$10821 ( \11491 , \11390 );
nand \U$10822 ( \11492 , \11491 , \11399 , \11445 , \11421 );
not \U$10823 ( \11493 , \11492 );
not \U$10824 ( \11494 , \11493 );
or \U$10825 ( \11495 , \11490 , \11494 );
not \U$10826 ( \11496 , \11454 );
nand \U$10827 ( \11497 , \11439 , \11496 , \11445 , \11421 );
not \U$10828 ( \11498 , \11497 );
nand \U$10829 ( \11499 , \11498 , RIaa9b370_131);
nand \U$10830 ( \11500 , \11495 , \11499 );
not \U$10831 ( \11501 , RIaa9b118_126);
not \U$10832 ( \11502 , \11399 );
not \U$10833 ( \11503 , \11502 );
nand \U$10834 ( \11504 , \11503 , \11454 , \11430 , \11447 );
not \U$10835 ( \11505 , \11504 );
not \U$10836 ( \11506 , \11505 );
or \U$10837 ( \11507 , \11501 , \11506 );
not \U$10838 ( \11508 , \11428 );
nand \U$10839 ( \11509 , \11508 , \11461 , \11445 , \11436 );
not \U$10840 ( \11510 , \11509 );
nand \U$10841 ( \11511 , \11510 , RIaa9b2f8_130);
nand \U$10842 ( \11512 , \11507 , \11511 );
nor \U$10843 ( \11513 , \11500 , \11512 );
not \U$10844 ( \11514 , RIaa9b190_127);
not \U$10845 ( \11515 , \11426 );
not \U$10846 ( \11516 , \11439 );
nand \U$10847 ( \11517 , \11515 , \11516 , \11430 , \11447 );
not \U$10848 ( \11518 , \11517 );
not \U$10849 ( \11519 , \11518 );
or \U$10850 ( \11520 , \11514 , \11519 );
not \U$10851 ( \11521 , \11399 );
and \U$10852 ( \11522 , \11436 , \11521 , \11445 , \11421 );
nand \U$10853 ( \11523 , \11522 , RIaa9b5c8_136);
nand \U$10854 ( \11524 , \11520 , \11523 );
not \U$10855 ( \11525 , RIaa9b550_135);
nand \U$10856 ( \11526 , \11502 , \11426 , \11445 , \11461 );
not \U$10857 ( \11527 , \11526 );
not \U$10858 ( \11528 , \11527 );
or \U$10859 ( \11529 , \11525 , \11528 );
not \U$10860 ( \11530 , \11445 );
not \U$10861 ( \11531 , \11454 );
nand \U$10862 ( \11532 , \11530 , \11531 , \11452 , \11447 );
not \U$10863 ( \11533 , \11532 );
nand \U$10864 ( \11534 , \11533 , RIaa9ae48_120);
nand \U$10865 ( \11535 , \11529 , \11534 );
nor \U$10866 ( \11536 , \11524 , \11535 );
nand \U$10867 ( \11537 , \11460 , \11489 , \11513 , \11536 );
not \U$10868 ( \11538 , \11537 );
nand \U$10869 ( \11539 , RIaaa9128_604, RIaaa91a0_605);
not \U$10870 ( \11540 , \11539 );
nand \U$10871 ( \11541 , \11540 , RIaaa90b0_603);
not \U$10872 ( \11542 , RIaaa90b0_603);
nand \U$10873 ( \11543 , \11542 , \11539 );
nand \U$10874 ( \11544 , \11541 , \11543 );
not \U$10875 ( \11545 , \11544 );
nor \U$10876 ( \11546 , \11538 , \11545 );
buf \U$10877 ( \11547 , \11462 );
not \U$10878 ( \11548 , RIaa99a20_77);
or \U$10879 ( \11549 , \11547 , \11548 );
nand \U$10880 ( \11550 , \11473 , RIaa998b8_74);
nand \U$10881 ( \11551 , RIaa99930_75, RIaaa8a20_589);
nand \U$10882 ( \11552 , \11549 , \11550 , \11551 );
not \U$10883 ( \11553 , RIaa997c8_72);
not \U$10884 ( \11554 , \11510 );
or \U$10885 ( \11555 , \11553 , \11554 );
and \U$10886 ( \11556 , \11461 , \11452 , \11445 , \11426 );
nand \U$10887 ( \11557 , \11556 , RIaa99a98_78);
nand \U$10888 ( \11558 , \11555 , \11557 );
nor \U$10889 ( \11559 , \11552 , \11558 );
not \U$10890 ( \11560 , RIaa99cf0_83);
not \U$10891 ( \11561 , \11432 );
or \U$10892 ( \11562 , \11560 , \11561 );
not \U$10893 ( \11563 , \11454 );
not \U$10894 ( \11564 , \11438 );
nand \U$10895 ( \11565 , \11563 , \11564 , \11415 , \11421 );
not \U$10896 ( \11566 , \11565 );
nand \U$10897 ( \11567 , \11566 , RIaa99b88_80);
nand \U$10898 ( \11568 , \11562 , \11567 );
not \U$10899 ( \11569 , RIaa99d68_84);
not \U$10900 ( \11570 , \11422 );
not \U$10901 ( \11571 , \11570 );
or \U$10902 ( \11572 , \11569 , \11571 );
not \U$10903 ( \11573 , \11436 );
nand \U$10904 ( \11574 , \11573 , \11429 , \11415 , \11447 );
not \U$10905 ( \11575 , \11574 );
nand \U$10906 ( \11576 , \11575 , RIaa99c78_82);
nand \U$10907 ( \11577 , \11572 , \11576 );
nor \U$10908 ( \11578 , \11568 , \11577 );
not \U$10909 ( \11579 , \11492 );
not \U$10910 ( \11580 , \11579 );
or \U$10911 ( \11581 , \11580 , \1268 );
not \U$10912 ( \11582 , RIaa99c00_81);
or \U$10913 ( \11583 , \11582 , \11456 );
nand \U$10914 ( \11584 , \11581 , \11583 );
not \U$10915 ( \11585 , \11399 );
nand \U$10916 ( \11586 , \11454 , \11585 , \11445 , \11461 );
not \U$10917 ( \11587 , RIaa99de0_85);
or \U$10918 ( \11588 , \11586 , \11587 );
not \U$10919 ( \11589 , RIaa996d8_70);
or \U$10920 ( \11590 , \11589 , \11479 );
nand \U$10921 ( \11591 , \11588 , \11590 );
nor \U$10922 ( \11592 , \11584 , \11591 );
not \U$10923 ( \11593 , RIaa99660_69);
not \U$10924 ( \11594 , \11399 );
nand \U$10925 ( \11595 , \11594 , \11491 , \11414 , \11461 );
not \U$10926 ( \11596 , \11595 );
not \U$10927 ( \11597 , \11596 );
or \U$10928 ( \11598 , \11593 , \11597 );
not \U$10929 ( \11599 , \11452 );
nand \U$10930 ( \11600 , \11599 , \11563 , \11445 , \11421 );
not \U$10931 ( \11601 , \11600 );
nand \U$10932 ( \11602 , \11601 , RIaa99750_71);
nand \U$10933 ( \11603 , \11598 , \11602 );
not \U$10934 ( \11604 , RIaa99b10_79);
not \U$10935 ( \11605 , \11522 );
or \U$10936 ( \11606 , \11604 , \11605 );
nand \U$10937 ( \11607 , \11415 , \11400 , \11455 , \11447 );
not \U$10938 ( \11608 , \11607 );
nand \U$10939 ( \11609 , \11608 , RIaa99840_73);
nand \U$10940 ( \11610 , \11606 , \11609 );
nor \U$10941 ( \11611 , \11603 , \11610 );
nand \U$10942 ( \11612 , \11559 , \11578 , \11592 , \11611 );
not \U$10943 ( \11613 , RIaaa9290_607);
nor \U$10944 ( \11614 , \11364 , \11613 );
and \U$10945 ( \11615 , RIaaa9308_608, \11614 );
nor \U$10946 ( \11616 , \11615 , RIaaa9380_609);
not \U$10947 ( \11617 , \11616 );
nand \U$10948 ( \11618 , \11617 , \11367 );
buf \U$10949 ( \11619 , \11618 );
nand \U$10950 ( \11620 , \11612 , \11619 );
not \U$10951 ( \11621 , \11620 );
nor \U$10952 ( \11622 , \11546 , \11621 );
nand \U$10953 ( \11623 , \11391 , \11400 , \11415 , \11421 );
not \U$10954 ( \11624 , \11623 );
not \U$10955 ( \11625 , \6435 );
and \U$10956 ( \11626 , \11624 , \11625 );
and \U$10957 ( \11627 , \11445 , \11428 , \11390 , \11421 );
and \U$10958 ( \11628 , \11627 , RIaa9d530_203);
nor \U$10959 ( \11629 , \11626 , \11628 );
not \U$10960 ( \11630 , \11462 );
and \U$10961 ( \11631 , \11630 , RIaa9cf90_191);
and \U$10962 ( \11632 , RIaa9cea0_189, RIaaa8a20_589);
nor \U$10963 ( \11633 , \11631 , \11632 );
nand \U$10964 ( \11634 , \11486 , RIaa9d5a8_204);
nand \U$10965 ( \11635 , \11629 , \11633 , \11634 );
not \U$10966 ( \11636 , \11479 );
not \U$10967 ( \11637 , RIaa9d260_197);
not \U$10968 ( \11638 , \11637 );
and \U$10969 ( \11639 , \11636 , \11638 );
not \U$10970 ( \11640 , RIaa9d440_201);
nor \U$10971 ( \11641 , \11586 , \11640 );
nor \U$10972 ( \11642 , \11639 , \11641 );
and \U$10973 ( \11643 , \11556 , RIaa9d4b8_202);
and \U$10974 ( \11644 , \11510 , RIaa9d350_199);
nor \U$10975 ( \11645 , \11643 , \11644 );
nand \U$10976 ( \11646 , \11642 , \11645 );
nor \U$10977 ( \11647 , \11635 , \11646 );
and \U$10978 ( \11648 , \11575 , RIaa9d0f8_194);
and \U$10979 ( \11649 , \11473 , RIaa9d080_193);
nor \U$10980 ( \11650 , \11648 , \11649 );
not \U$10981 ( \11651 , \11607 );
not \U$10982 ( \11652 , RIaa9d008_192);
not \U$10983 ( \11653 , \11652 );
and \U$10984 ( \11654 , \11651 , \11653 );
and \U$10985 ( \11655 , \11493 , RIaa9cf18_190);
nor \U$10986 ( \11656 , \11654 , \11655 );
nand \U$10987 ( \11657 , \11650 , \11656 );
not \U$10988 ( \11658 , \11454 );
nand \U$10989 ( \11659 , \11658 , \11564 , \11415 , \11461 );
not \U$10990 ( \11660 , \11659 );
nand \U$10991 ( \11661 , \11660 , RIaa9d620_205);
nand \U$10992 ( \11662 , \11601 , RIaa9d3c8_200);
nand \U$10993 ( \11663 , \11596 , RIaa9d1e8_196);
nand \U$10994 ( \11664 , \11454 , \11439 , \11415 , \11421 );
not \U$10995 ( \11665 , \11664 );
nand \U$10996 ( \11666 , \11665 , RIaa9d2d8_198);
nand \U$10997 ( \11667 , \11661 , \11662 , \11663 , \11666 );
nor \U$10998 ( \11668 , \11657 , \11667 );
nand \U$10999 ( \11669 , \11647 , \11668 );
not \U$11000 ( \11670 , RIaaa9218_606);
not \U$11001 ( \11671 , \11670 );
not \U$11002 ( \11672 , \11541 );
or \U$11003 ( \11673 , \11671 , \11672 );
nand \U$11004 ( \11674 , \11673 , \11364 );
nand \U$11005 ( \11675 , \11669 , \11674 );
not \U$11006 ( \11676 , \11509 );
not \U$11007 ( \11677 , RIaa9ab00_113);
not \U$11008 ( \11678 , \11677 );
and \U$11009 ( \11679 , \11676 , \11678 );
and \U$11010 ( \11680 , \11473 , RIaa9a6c8_104);
nor \U$11011 ( \11681 , \11679 , \11680 );
and \U$11012 ( \11682 , RIaa9a830_107, \11463 );
and \U$11013 ( \11683 , RIaa9a740_105, RIaaa8a20_589);
nor \U$11014 ( \11684 , \11682 , \11683 );
nand \U$11015 ( \11685 , \11486 , RIaa9ad58_118);
nand \U$11016 ( \11686 , \11681 , \11684 , \11685 );
not \U$11017 ( \11687 , \11659 );
not \U$11018 ( \11688 , RIaa9add0_119);
not \U$11019 ( \11689 , \11688 );
and \U$11020 ( \11690 , \11687 , \11689 );
not \U$11021 ( \11691 , RIaa9a998_110);
nor \U$11022 ( \11692 , \11595 , \11691 );
nor \U$11023 ( \11693 , \11690 , \11692 );
not \U$11024 ( \11694 , \11623 );
not \U$11025 ( \11695 , RIaa9a8a8_108);
not \U$11026 ( \11696 , \11695 );
and \U$11027 ( \11697 , \11694 , \11696 );
and \U$11028 ( \11698 , \11533 , RIaa9a650_103);
nor \U$11029 ( \11699 , \11697 , \11698 );
nand \U$11030 ( \11700 , \11693 , \11699 );
nor \U$11031 ( \11701 , \11686 , \11700 );
not \U$11032 ( \11702 , RIaa9aa88_112);
or \U$11033 ( \11703 , \11664 , \11702 );
not \U$11034 ( \11704 , RIaa9a920_109);
or \U$11035 ( \11705 , \11574 , \11704 );
not \U$11036 ( \11706 , \11600 );
not \U$11037 ( \11707 , RIaa9ab78_114);
not \U$11038 ( \11708 , \11707 );
and \U$11039 ( \11709 , \11706 , \11708 );
not \U$11040 ( \11710 , RIaa9aa10_111);
nor \U$11041 ( \11711 , \11479 , \11710 );
nor \U$11042 ( \11712 , \11709 , \11711 );
nand \U$11043 ( \11713 , \11703 , \11705 , \11712 );
nand \U$11044 ( \11714 , \11493 , RIaa9a7b8_106);
not \U$11045 ( \11715 , \11586 );
nand \U$11046 ( \11716 , \11715 , RIaa9abf0_115);
nand \U$11047 ( \11717 , \11627 , RIaa9ac68_116);
nand \U$11048 ( \11718 , \11556 , RIaa9ace0_117);
nand \U$11049 ( \11719 , \11714 , \11716 , \11717 , \11718 );
nor \U$11050 ( \11720 , \11713 , \11719 );
nand \U$11051 ( \11721 , \11701 , \11720 );
not \U$11052 ( \11722 , \11614 );
nand \U$11053 ( \11723 , \11364 , \11613 );
nand \U$11054 ( \11724 , \11722 , \11723 );
nand \U$11055 ( \11725 , \11721 , \11724 );
and \U$11056 ( \11726 , \11675 , \11725 );
and \U$11057 ( \11727 , \11518 , RIaa9a380_97);
and \U$11058 ( \11728 , \11473 , RIaa99fc0_89);
nor \U$11059 ( \11729 , \11727 , \11728 );
not \U$11060 ( \11730 , \11547 );
and \U$11061 ( \11731 , \11730 , RIaa9a038_90);
and \U$11062 ( \11732 , RIaa99ed0_87, RIaaa8a20_589);
nor \U$11063 ( \11733 , \11731 , \11732 );
nand \U$11064 ( \11734 , \11579 , RIaa99f48_88);
nand \U$11065 ( \11735 , \11729 , \11733 , \11734 );
nand \U$11066 ( \11736 , \11423 , RIaa9a290_95);
nand \U$11067 ( \11737 , \11505 , RIaa9a308_96);
nand \U$11068 ( \11738 , \11449 , RIaa9a5d8_102);
nand \U$11069 ( \11739 , \11498 , RIaa9a4e8_100);
nand \U$11070 ( \11740 , \11736 , \11737 , \11738 , \11739 );
nor \U$11071 ( \11741 , \11735 , \11740 );
nand \U$11072 ( \11742 , \11486 , RIaa9a0b0_91);
nand \U$11073 ( \11743 , \11432 , RIaa9a470_99);
nand \U$11074 ( \11744 , \11480 , RIaa9a3f8_98);
not \U$11075 ( \11745 , \11456 );
nand \U$11076 ( \11746 , \11745 , RIaa9a218_94);
nand \U$11077 ( \11747 , \11742 , \11743 , \11744 , \11746 );
nand \U$11078 ( \11748 , \11510 , RIaa9a560_101);
nand \U$11079 ( \11749 , \11522 , RIaa9a1a0_93);
nand \U$11080 ( \11750 , \11533 , RIaa99e58_86);
nand \U$11081 ( \11751 , \11527 , RIaa9a128_92);
nand \U$11082 ( \11752 , \11748 , \11749 , \11750 , \11751 );
nor \U$11083 ( \11753 , \11747 , \11752 );
nand \U$11084 ( \11754 , \11741 , \11753 );
and \U$11085 ( \11755 , \11614 , RIaaa9308_608);
not \U$11086 ( \11756 , \11614 );
not \U$11087 ( \11757 , RIaaa9308_608);
and \U$11088 ( \11758 , \11756 , \11757 );
or \U$11089 ( \11759 , \11755 , \11758 );
nand \U$11090 ( \11760 , \11754 , \11759 );
nand \U$11091 ( \11761 , \11622 , \11726 , \11760 );
not \U$11092 ( \11762 , RIaa9beb0_155);
not \U$11093 ( \11763 , \11449 );
or \U$11094 ( \11764 , \11762 , \11763 );
nand \U$11095 ( \11765 , \11480 , RIaa9c540_169);
nand \U$11096 ( \11766 , \11764 , \11765 );
nand \U$11097 ( \11767 , \11463 , RIaa9c180_161);
nand \U$11098 ( \11768 , \11473 , RIaa9c090_159);
nand \U$11099 ( \11769 , RIaa9c108_160, RIaaa8a20_589);
nand \U$11100 ( \11770 , \11767 , \11768 , \11769 );
nor \U$11101 ( \11771 , \11766 , \11770 );
not \U$11102 ( \11772 , RIaa9c3d8_166);
not \U$11103 ( \11773 , \11510 );
or \U$11104 ( \11774 , \11772 , \11773 );
nand \U$11105 ( \11775 , \11601 , RIaa9c360_165);
nand \U$11106 ( \11776 , \11774 , \11775 );
not \U$11107 ( \11777 , RIaa9c2e8_164);
not \U$11108 ( \11778 , \11570 );
or \U$11109 ( \11779 , \11777 , \11778 );
nand \U$11110 ( \11780 , \11665 , RIaa9be38_154);
nand \U$11111 ( \11781 , \11779 , \11780 );
nor \U$11112 ( \11782 , \11776 , \11781 );
not \U$11113 ( \11783 , RIaa9c5b8_170);
not \U$11114 ( \11784 , \11575 );
or \U$11115 ( \11785 , \11783 , \11784 );
nand \U$11116 ( \11786 , \11566 , RIaa9c450_167);
nand \U$11117 ( \11787 , \11785 , \11786 );
not \U$11118 ( \11788 , RIaa9c270_163);
not \U$11119 ( \11789 , \11596 );
or \U$11120 ( \11790 , \11788 , \11789 );
nand \U$11121 ( \11791 , \11579 , RIaa9c1f8_162);
nand \U$11122 ( \11792 , \11790 , \11791 );
nor \U$11123 ( \11793 , \11787 , \11792 );
not \U$11124 ( \11794 , RIaa9c4c8_168);
not \U$11125 ( \11795 , \11456 );
not \U$11126 ( \11796 , \11795 );
or \U$11127 ( \11797 , \11794 , \11796 );
nand \U$11128 ( \11798 , \11533 , RIaa9c018_158);
nand \U$11129 ( \11799 , \11797 , \11798 );
not \U$11130 ( \11800 , RIaa9bfa0_157);
not \U$11131 ( \11801 , \11527 );
or \U$11132 ( \11802 , \11800 , \11801 );
nand \U$11133 ( \11803 , \11627 , RIaa9bf28_156);
nand \U$11134 ( \11804 , \11802 , \11803 );
nor \U$11135 ( \11805 , \11799 , \11804 );
nand \U$11136 ( \11806 , \11771 , \11782 , \11793 , \11805 );
not \U$11137 ( \11807 , \11806 );
not \U$11138 ( \11808 , RIaaa91a0_605);
and \U$11139 ( \11809 , \11807 , \11808 );
not \U$11140 ( \11810 , RIaaa9128_604);
not \U$11141 ( \11811 , \11810 );
not \U$11142 ( \11812 , \11808 );
or \U$11143 ( \11813 , \11811 , \11812 );
nand \U$11144 ( \11814 , \11813 , \11539 );
nand \U$11145 ( \11815 , \11463 , RIaa9ba00_145);
nand \U$11146 ( \11816 , \11473 , RIaa9b898_142);
nand \U$11147 ( \11817 , RIaa9b910_143, RIaaa8a20_589);
nand \U$11148 ( \11818 , \11815 , \11816 , \11817 );
not \U$11149 ( \11819 , RIaa9b640_137);
not \U$11150 ( \11820 , \11505 );
or \U$11151 ( \11821 , \11819 , \11820 );
nand \U$11152 ( \11822 , \11510 , RIaa9baf0_147);
nand \U$11153 ( \11823 , \11821 , \11822 );
nor \U$11154 ( \11824 , \11818 , \11823 );
not \U$11155 ( \11825 , RIaa9b988_144);
not \U$11156 ( \11826 , \11493 );
or \U$11157 ( \11827 , \11825 , \11826 );
nand \U$11158 ( \11828 , \11498 , RIaa9bb68_148);
nand \U$11159 ( \11829 , \11827 , \11828 );
not \U$11160 ( \11830 , RIaa9b730_139);
not \U$11161 ( \11831 , \11518 );
or \U$11162 ( \11832 , \11830 , \11831 );
not \U$11163 ( \11833 , \11623 );
nand \U$11164 ( \11834 , \11833 , RIaa9b6b8_138);
nand \U$11165 ( \11835 , \11832 , \11834 );
nor \U$11166 ( \11836 , \11829 , \11835 );
not \U$11167 ( \11837 , RIaa9ba78_146);
not \U$11168 ( \11838 , \11432 );
or \U$11169 ( \11839 , \11837 , \11838 );
nand \U$11170 ( \11840 , \11566 , RIaa9bd48_152);
nand \U$11171 ( \11841 , \11839 , \11840 );
not \U$11172 ( \11842 , RIaa9b7a8_140);
not \U$11173 ( \11843 , \11480 );
or \U$11174 ( \11844 , \11842 , \11843 );
nand \U$11175 ( \11845 , \11556 , RIaa9bc58_150);
nand \U$11176 ( \11846 , \11844 , \11845 );
nor \U$11177 ( \11847 , \11841 , \11846 );
not \U$11178 ( \11848 , RIaa9bbe0_149);
not \U$11179 ( \11849 , \11715 );
or \U$11180 ( \11850 , \11848 , \11849 );
not \U$11181 ( \11851 , \11659 );
nand \U$11182 ( \11852 , \11851 , RIaa9bdc0_153);
nand \U$11183 ( \11853 , \11850 , \11852 );
not \U$11184 ( \11854 , RIaa9bcd0_151);
not \U$11185 ( \11855 , \11522 );
or \U$11186 ( \11856 , \11854 , \11855 );
nand \U$11187 ( \11857 , \11608 , RIaa9b820_141);
nand \U$11188 ( \11858 , \11856 , \11857 );
nor \U$11189 ( \11859 , \11853 , \11858 );
nand \U$11190 ( \11860 , \11824 , \11836 , \11847 , \11859 );
nor \U$11191 ( \11861 , \11814 , \11860 );
nor \U$11192 ( \11862 , \11809 , \11861 );
not \U$11193 ( \11863 , \11862 );
not \U$11194 ( \11864 , RIaaa91a0_605);
not \U$11195 ( \11865 , \11806 );
or \U$11196 ( \11866 , \11864 , \11865 );
nand \U$11197 ( \11867 , \11630 , RIaa9c810_175);
nand \U$11198 ( \11868 , \11473 , RIaa9c798_174);
nand \U$11199 ( \11869 , RIaa9c720_173, RIaaa8a20_589);
nand \U$11200 ( \11870 , \11867 , \11868 , \11869 );
not \U$11201 ( \11871 , RIaa9c9f0_179);
not \U$11202 ( \11872 , \11498 );
or \U$11203 ( \11873 , \11871 , \11872 );
nand \U$11204 ( \11874 , \11660 , RIaa9cb58_182);
nand \U$11205 ( \11875 , \11873 , \11874 );
nor \U$11206 ( \11876 , \11870 , \11875 );
not \U$11207 ( \11877 , RIaa9c888_176);
not \U$11208 ( \11878 , \11505 );
or \U$11209 ( \11879 , \11877 , \11878 );
nand \U$11210 ( \11880 , \11665 , RIaa9cd38_186);
nand \U$11211 ( \11881 , \11879 , \11880 );
not \U$11212 ( \11882 , RIaa9cdb0_187);
not \U$11213 ( \11883 , \11449 );
or \U$11214 ( \11884 , \11882 , \11883 );
nand \U$11215 ( \11885 , \11510 , RIaa9cbd0_183);
nand \U$11216 ( \11886 , \11884 , \11885 );
nor \U$11217 ( \11887 , \11881 , \11886 );
not \U$11218 ( \11888 , RIaa9cc48_184);
not \U$11219 ( \11889 , \11518 );
or \U$11220 ( \11890 , \11888 , \11889 );
nand \U$11221 ( \11891 , \11493 , RIaa9c630_171);
nand \U$11222 ( \11892 , \11890 , \11891 );
not \U$11223 ( \11893 , RIaa9ccc0_185);
not \U$11224 ( \11894 , \11833 );
or \U$11225 ( \11895 , \11893 , \11894 );
nand \U$11226 ( \11896 , \11627 , RIaa9cae0_181);
nand \U$11227 ( \11897 , \11895 , \11896 );
nor \U$11228 ( \11898 , \11892 , \11897 );
not \U$11229 ( \11899 , RIaa9c900_177);
not \U$11230 ( \11900 , \11480 );
or \U$11231 ( \11901 , \11899 , \11900 );
nand \U$11232 ( \11902 , \11566 , RIaa9ca68_180);
nand \U$11233 ( \11903 , \11901 , \11902 );
not \U$11234 ( \11904 , RIaa9c978_178);
not \U$11235 ( \11905 , \11527 );
or \U$11236 ( \11906 , \11904 , \11905 );
nand \U$11237 ( \11907 , \11608 , RIaa9c6a8_172);
nand \U$11238 ( \11908 , \11906 , \11907 );
nor \U$11239 ( \11909 , \11903 , \11908 );
nand \U$11240 ( \11910 , \11876 , \11887 , \11898 , \11909 );
not \U$11241 ( \11911 , RIaaa9560_613);
nand \U$11242 ( \11912 , \11910 , \11911 );
nand \U$11243 ( \11913 , \11866 , \11912 );
not \U$11244 ( \11914 , \11913 );
or \U$11245 ( \11915 , \11863 , \11914 );
not \U$11246 ( \11916 , \11860 );
not \U$11247 ( \11917 , \11814 );
nor \U$11248 ( \11918 , \11916 , \11917 );
not \U$11249 ( \11919 , \11918 );
nand \U$11250 ( \11920 , \11915 , \11919 );
or \U$11251 ( \11921 , \11761 , \11920 );
not \U$11252 ( \11922 , \11754 );
not \U$11253 ( \11923 , \11759 );
nor \U$11254 ( \11924 , \11922 , \11923 );
nand \U$11255 ( \11925 , \11620 , \11725 );
nor \U$11256 ( \11926 , \11924 , \11925 );
nand \U$11257 ( \11927 , \11675 , \11538 , \11545 );
not \U$11258 ( \11928 , \11669 );
not \U$11259 ( \11929 , \11674 );
nand \U$11260 ( \11930 , \11928 , \11929 );
not \U$11261 ( \11931 , \11721 );
not \U$11262 ( \11932 , \11724 );
nand \U$11263 ( \11933 , \11931 , \11932 );
nand \U$11264 ( \11934 , \11927 , \11930 , \11933 );
and \U$11265 ( \11935 , \11926 , \11934 );
not \U$11266 ( \11936 , \11754 );
nand \U$11267 ( \11937 , \11936 , \11923 );
not \U$11268 ( \11938 , \11619 );
not \U$11269 ( \11939 , \11612 );
nand \U$11270 ( \11940 , \11938 , \11939 );
and \U$11271 ( \11941 , \11937 , \11940 );
not \U$11272 ( \11942 , \11620 );
nor \U$11273 ( \11943 , \11941 , \11942 );
nor \U$11274 ( \11944 , \11935 , \11943 );
nand \U$11275 ( \11945 , \11921 , \11944 );
buf \U$11276 ( \11946 , \11945 );
buf \U$11277 ( \11947 , \11498 );
buf \U$11278 ( \11948 , \11947 );
nand \U$11279 ( \11949 , \11948 , RIaa9e3b8_234);
not \U$11280 ( \11950 , \11510 );
not \U$11281 ( \11951 , \11950 );
nand \U$11282 ( \11952 , \11951 , RIaa9e430_235);
buf \U$11283 ( \11953 , \11505 );
nand \U$11284 ( \11954 , \11953 , RIaa9e340_233);
buf \U$11285 ( \11955 , \11527 );
nand \U$11286 ( \11956 , \11955 , RIaa9e070_227);
nand \U$11287 ( \11957 , \11949 , \11952 , \11954 , \11956 );
not \U$11288 ( \11958 , \11957 );
buf \U$11289 ( \11959 , \11547 );
not \U$11290 ( \11960 , \11959 );
nand \U$11291 ( \11961 , \11960 , RIaa9e160_229);
nand \U$11292 ( \11962 , \11473 , RIaa9df08_224);
nand \U$11293 ( \11963 , RIaa9df80_225, RIaaa8a20_589);
nand \U$11294 ( \11964 , \11961 , \11962 , \11963 );
not \U$11295 ( \11965 , RIaa9e4a8_236);
buf \U$11296 ( \11966 , \11480 );
not \U$11297 ( \11967 , \11966 );
or \U$11298 ( \11968 , \11965 , \11967 );
buf \U$11299 ( \11969 , \11518 );
nand \U$11300 ( \11970 , \11969 , RIaa9e520_237);
nand \U$11301 ( \11971 , \11968 , \11970 );
nor \U$11302 ( \11972 , \11964 , \11971 );
not \U$11303 ( \11973 , RIaa9e250_231);
not \U$11304 ( \11974 , \11745 );
not \U$11305 ( \11975 , \11974 );
not \U$11306 ( \11976 , \11975 );
or \U$11307 ( \11977 , \11973 , \11976 );
not \U$11308 ( \11978 , \11431 );
nand \U$11309 ( \11979 , \11978 , RIaa9e2c8_232);
nand \U$11310 ( \11980 , \11977 , \11979 );
not \U$11311 ( \11981 , RIaa9e598_238);
buf \U$11312 ( \11982 , \11423 );
not \U$11313 ( \11983 , \11982 );
or \U$11314 ( \11984 , \11981 , \11983 );
buf \U$11315 ( \11985 , \11486 );
nand \U$11316 ( \11986 , \11985 , RIaa9e1d8_230);
nand \U$11317 ( \11987 , \11984 , \11986 );
nor \U$11318 ( \11988 , \11980 , \11987 );
not \U$11319 ( \11989 , RIaa9e610_239);
not \U$11320 ( \11990 , \11448 );
not \U$11321 ( \11991 , \11990 );
or \U$11322 ( \11992 , \11989 , \11991 );
buf \U$11323 ( \11993 , \11580 );
not \U$11324 ( \11994 , \11993 );
nand \U$11325 ( \11995 , \11994 , RIaa9e0e8_228);
nand \U$11326 ( \11996 , \11992 , \11995 );
not \U$11327 ( \11997 , RIaa9de90_223);
buf \U$11328 ( \11998 , \11533 );
not \U$11329 ( \11999 , \11998 );
or \U$11330 ( \12000 , \11997 , \11999 );
buf \U$11331 ( \12001 , \11522 );
nand \U$11332 ( \12002 , \12001 , RIaa9dff8_226);
nand \U$11333 ( \12003 , \12000 , \12002 );
nor \U$11334 ( \12004 , \11996 , \12003 );
nand \U$11335 ( \12005 , \11958 , \11972 , \11988 , \12004 );
nand \U$11336 ( \12006 , \11366 , RIaaa93f8_610);
not \U$11337 ( \12007 , \12006 );
nand \U$11338 ( \12008 , \12007 , RIaaa9038_602);
not \U$11339 ( \12009 , \12008 );
nor \U$11340 ( \12010 , \12009 , RIaaa9470_611);
not \U$11341 ( \12011 , \12010 );
nand \U$11342 ( \12012 , \12009 , RIaaa9470_611);
nand \U$11343 ( \12013 , \12011 , \12012 );
buf \U$11344 ( \12014 , \12013 );
nand \U$11345 ( \12015 , \12005 , \12014 );
not \U$11346 ( \12016 , RIaaa94e8_612);
nand \U$11347 ( \12017 , \12016 , \12012 );
not \U$11348 ( \12018 , \11369 );
and \U$11349 ( \12019 , \12017 , \12018 );
not \U$11350 ( \12020 , \12019 );
nand \U$11351 ( \12021 , \11960 , RIaa98850_39);
nand \U$11352 ( \12022 , \11473 , RIaa986e8_36);
nand \U$11353 ( \12023 , RIaa98760_37, RIaaa8a20_589);
nand \U$11354 ( \12024 , \12021 , \12022 , \12023 );
not \U$11355 ( \12025 , RIaa98b98_46);
not \U$11356 ( \12026 , \11948 );
or \U$11357 ( \12027 , \12025 , \12026 );
nand \U$11358 ( \12028 , \11975 , RIaa98a30_43);
nand \U$11359 ( \12029 , \12027 , \12028 );
nor \U$11360 ( \12030 , \12024 , \12029 );
not \U$11361 ( \12031 , RIaa987d8_38);
not \U$11362 ( \12032 , \11994 );
or \U$11363 ( \12033 , \12031 , \12032 );
nand \U$11364 ( \12034 , \11985 , RIaa989b8_42);
nand \U$11365 ( \12035 , \12033 , \12034 );
not \U$11366 ( \12036 , RIaa98b20_45);
not \U$11367 ( \12037 , \11982 );
or \U$11368 ( \12038 , \12036 , \12037 );
nand \U$11369 ( \12039 , \11953 , RIaa98aa8_44);
nand \U$11370 ( \12040 , \12038 , \12039 );
nor \U$11371 ( \12041 , \12035 , \12040 );
not \U$11372 ( \12042 , RIaa98df0_51);
not \U$11373 ( \12043 , \11969 );
or \U$11374 ( \12044 , \12042 , \12043 );
nand \U$11375 ( \12045 , \11951 , RIaa98c10_47);
nand \U$11376 ( \12046 , \12044 , \12045 );
not \U$11377 ( \12047 , RIaa98d00_49);
not \U$11378 ( \12048 , \11990 );
or \U$11379 ( \12049 , \12047 , \12048 );
not \U$11380 ( \12050 , \11431 );
nand \U$11381 ( \12051 , \12050 , RIaa98c88_48);
nand \U$11382 ( \12052 , \12049 , \12051 );
nor \U$11383 ( \12053 , \12046 , \12052 );
not \U$11384 ( \12054 , RIaa98d78_50);
not \U$11385 ( \12055 , \11966 );
or \U$11386 ( \12056 , \12054 , \12055 );
buf \U$11387 ( \12057 , \11998 );
nand \U$11388 ( \12058 , \12057 , RIaa98670_35);
nand \U$11389 ( \12059 , \12056 , \12058 );
not \U$11390 ( \12060 , RIaa98940_41);
not \U$11391 ( \12061 , \11955 );
or \U$11392 ( \12062 , \12060 , \12061 );
nand \U$11393 ( \12063 , \12001 , RIaa988c8_40);
nand \U$11394 ( \12064 , \12062 , \12063 );
nor \U$11395 ( \12065 , \12059 , \12064 );
nand \U$11396 ( \12066 , \12030 , \12041 , \12053 , \12065 );
nand \U$11397 ( \12067 , \12020 , \12066 );
nand \U$11398 ( \12068 , \11960 , RIaa9de18_222);
nand \U$11399 ( \12069 , \11473 , RIaa9dad0_215);
nand \U$11400 ( \12070 , RIaa9db48_216, RIaaa8a20_589);
nand \U$11401 ( \12071 , \12068 , \12069 , \12070 );
not \U$11402 ( \12072 , RIaa9d878_210);
not \U$11403 ( \12073 , \11947 );
or \U$11404 ( \12074 , \12072 , \12073 );
not \U$11405 ( \12075 , \11974 );
nand \U$11406 ( \12076 , \12075 , RIaa9dd28_220);
nand \U$11407 ( \12077 , \12074 , \12076 );
nor \U$11408 ( \12078 , \12071 , \12077 );
not \U$11409 ( \12079 , RIaa9d788_208);
not \U$11410 ( \12080 , \11982 );
or \U$11411 ( \12081 , \12079 , \12080 );
nand \U$11412 ( \12082 , \11985 , RIaa9dcb0_219);
nand \U$11413 ( \12083 , \12081 , \12082 );
not \U$11414 ( \12084 , RIaa9d968_212);
not \U$11415 ( \12085 , \11966 );
or \U$11416 ( \12086 , \12084 , \12085 );
nand \U$11417 ( \12087 , \11951 , RIaa9d8f0_211);
nand \U$11418 ( \12088 , \12086 , \12087 );
nor \U$11419 ( \12089 , \12083 , \12088 );
not \U$11420 ( \12090 , RIaa9d9e0_213);
not \U$11421 ( \12091 , \11969 );
or \U$11422 ( \12092 , \12090 , \12091 );
nand \U$11423 ( \12093 , \11953 , RIaa9d710_207);
nand \U$11424 ( \12094 , \12092 , \12093 );
not \U$11425 ( \12095 , RIaa9d800_209);
not \U$11426 ( \12096 , \11990 );
or \U$11427 ( \12097 , \12095 , \12096 );
nand \U$11428 ( \12098 , \11994 , RIaa9dda0_221);
nand \U$11429 ( \12099 , \12097 , \12098 );
nor \U$11430 ( \12100 , \12094 , \12099 );
not \U$11431 ( \12101 , RIaa9d698_206);
not \U$11432 ( \12102 , \11978 );
or \U$11433 ( \12103 , \12101 , \12102 );
nand \U$11434 ( \12104 , \11998 , RIaa9da58_214);
nand \U$11435 ( \12105 , \12103 , \12104 );
not \U$11436 ( \12106 , \11955 );
not \U$11437 ( \12107 , RIaa9dc38_218);
or \U$11438 ( \12108 , \12106 , \12107 );
not \U$11439 ( \12109 , \12001 );
or \U$11440 ( \12110 , \12109 , \1619 );
nand \U$11441 ( \12111 , \12108 , \12110 );
nor \U$11442 ( \12112 , \12105 , \12111 );
nand \U$11443 ( \12113 , \12078 , \12089 , \12100 , \12112 );
nor \U$11444 ( \12114 , \12007 , RIaaa9038_602);
not \U$11445 ( \12115 , \12114 );
nand \U$11446 ( \12116 , \12115 , \12008 );
buf \U$11447 ( \12117 , \12116 );
nand \U$11448 ( \12118 , \12113 , \12117 );
buf \U$11449 ( \12119 , \12118 );
or \U$11450 ( \12120 , \11366 , RIaaa93f8_610);
nand \U$11451 ( \12121 , \12120 , \12006 );
not \U$11452 ( \12122 , \12121 );
not \U$11453 ( \12123 , \12122 );
not \U$11454 ( \12124 , RIaa991b0_59);
not \U$11455 ( \12125 , \11947 );
or \U$11456 ( \12126 , \12124 , \12125 );
nand \U$11457 ( \12127 , \12075 , RIaa99408_64);
nand \U$11458 ( \12128 , \12126 , \12127 );
not \U$11459 ( \12129 , RIaa995e8_68);
not \U$11460 ( \12130 , \11966 );
or \U$11461 ( \12131 , \12129 , \12130 );
nand \U$11462 ( \12132 , \11969 , RIaa99570_67);
nand \U$11463 ( \12133 , \12131 , \12132 );
nor \U$11464 ( \12134 , \12128 , \12133 );
nand \U$11465 ( \12135 , \11960 , RIaa99048_56);
nand \U$11466 ( \12136 , \11473 , RIaa98ee0_53);
nand \U$11467 ( \12137 , RIaa98f58_54, RIaaa8a20_589);
nand \U$11468 ( \12138 , \12135 , \12136 , \12137 );
not \U$11469 ( \12139 , RIaa990c0_57);
not \U$11470 ( \12140 , \11953 );
or \U$11471 ( \12141 , \12139 , \12140 );
nand \U$11472 ( \12142 , \12050 , RIaa99480_65);
nand \U$11473 ( \12143 , \12141 , \12142 );
nor \U$11474 ( \12144 , \12138 , \12143 );
not \U$11475 ( \12145 , RIaa99390_63);
not \U$11476 ( \12146 , \11985 );
or \U$11477 ( \12147 , \12145 , \12146 );
nand \U$11478 ( \12148 , \11982 , RIaa99138_58);
nand \U$11479 ( \12149 , \12147 , \12148 );
not \U$11480 ( \12150 , RIaa98fd0_55);
not \U$11481 ( \12151 , \11994 );
or \U$11482 ( \12152 , \12150 , \12151 );
nand \U$11483 ( \12153 , \11998 , RIaa98e68_52);
nand \U$11484 ( \12154 , \12152 , \12153 );
nor \U$11485 ( \12155 , \12149 , \12154 );
not \U$11486 ( \12156 , RIaa99228_60);
not \U$11487 ( \12157 , \11951 );
or \U$11488 ( \12158 , \12156 , \12157 );
nand \U$11489 ( \12159 , \11990 , RIaa994f8_66);
nand \U$11490 ( \12160 , \12158 , \12159 );
not \U$11491 ( \12161 , RIaa992a0_61);
not \U$11492 ( \12162 , \11955 );
or \U$11493 ( \12163 , \12161 , \12162 );
nand \U$11494 ( \12164 , \12001 , RIaa99318_62);
nand \U$11495 ( \12165 , \12163 , \12164 );
nor \U$11496 ( \12166 , \12160 , \12165 );
nand \U$11497 ( \12167 , \12134 , \12144 , \12155 , \12166 );
buf \U$11498 ( \12168 , \12167 );
nand \U$11499 ( \12169 , \12123 , \12168 );
and \U$11500 ( \12170 , \12015 , \12067 , \12119 , \12169 );
and \U$11501 ( \12171 , \11946 , \12170 );
not \U$11502 ( \12172 , \12122 );
nor \U$11503 ( \12173 , \12172 , \12167 );
not \U$11504 ( \12174 , \12173 );
not \U$11505 ( \12175 , \12118 );
or \U$11506 ( \12176 , \12174 , \12175 );
not \U$11507 ( \12177 , \12113 );
not \U$11508 ( \12178 , \12117 );
nand \U$11509 ( \12179 , \12177 , \12178 );
nand \U$11510 ( \12180 , \12176 , \12179 );
and \U$11511 ( \12181 , \12180 , \12015 );
nor \U$11512 ( \12182 , \12005 , \12014 );
nor \U$11513 ( \12183 , \12181 , \12182 );
not \U$11514 ( \12184 , \12067 );
or \U$11515 ( \12185 , \12183 , \12184 );
not \U$11516 ( \12186 , \12019 );
nor \U$11517 ( \12187 , \12186 , \12066 );
not \U$11518 ( \12188 , \12187 );
nand \U$11519 ( \12189 , \12185 , \12188 );
nor \U$11520 ( \12190 , \12171 , \12189 );
not \U$11521 ( \12191 , RIaa98148_24);
not \U$11522 ( \12192 , \11960 );
or \U$11523 ( \12193 , \12191 , \12192 );
nand \U$11524 ( \12194 , RIaa97f68_20, RIaaa8a20_589);
nand \U$11525 ( \12195 , \12193 , \12194 );
not \U$11526 ( \12196 , \11969 );
nor \U$11527 ( \12197 , \12196 , \2016 );
nor \U$11528 ( \12198 , \12195 , \12197 );
and \U$11529 ( \12199 , RIaa983a0_29, \11948 );
buf \U$11530 ( \12200 , \11975 );
and \U$11531 ( \12201 , \12200 , RIaa98238_26);
nor \U$11532 ( \12202 , \12199 , \12201 );
nand \U$11533 ( \12203 , \12198 , \12202 );
and \U$11534 ( \12204 , \11985 , RIaa981c0_25);
not \U$11535 ( \12205 , RIaa98490_31);
not \U$11536 ( \12206 , \11966 );
nor \U$11537 ( \12207 , \12205 , \12206 );
nor \U$11538 ( \12208 , \12204 , \12207 );
buf \U$11539 ( \12209 , \11990 );
not \U$11540 ( \12210 , \12209 );
not \U$11541 ( \12211 , \12210 );
not \U$11542 ( \12212 , \2038 );
and \U$11543 ( \12213 , \12211 , \12212 );
not \U$11544 ( \12214 , \11982 );
not \U$11545 ( \12215 , \12214 );
and \U$11546 ( \12216 , \12215 , RIaa98580_33);
nor \U$11547 ( \12217 , \12213 , \12216 );
nand \U$11548 ( \12218 , \12208 , \12217 );
nor \U$11549 ( \12219 , \12203 , \12218 );
buf \U$11550 ( \12220 , \11993 );
not \U$11551 ( \12221 , \12220 );
nand \U$11552 ( \12222 , \12221 , RIaa980d0_23);
nand \U$11553 ( \12223 , \11953 , RIaa98328_28);
nand \U$11554 ( \12224 , \11951 , RIaa98418_30);
nand \U$11555 ( \12225 , \11473 , RIaa97e78_18);
nand \U$11556 ( \12226 , \12222 , \12223 , \12224 , \12225 );
not \U$11557 ( \12227 , \12106 );
and \U$11558 ( \12228 , \12227 , RIaa98058_22);
and \U$11559 ( \12229 , \12057 , RIaa97ef0_19);
nor \U$11560 ( \12230 , \12228 , \12229 );
buf \U$11561 ( \12231 , \12050 );
nand \U$11562 ( \12232 , \12231 , RIaa982b0_27);
buf \U$11563 ( \12233 , \12001 );
nand \U$11564 ( \12234 , \12233 , RIaa97fe0_21);
nand \U$11565 ( \12235 , \12230 , \12232 , \12234 );
nor \U$11566 ( \12236 , \12226 , \12235 );
nand \U$11567 ( \12237 , \12219 , \12236 );
not \U$11568 ( \12238 , \12237 );
xor \U$11569 ( \12239 , RIaaa95d8_614, \11369 );
nand \U$11570 ( \12240 , \12238 , \12239 );
and \U$11571 ( \12241 , \12190 , \12240 );
nor \U$11572 ( \12242 , \12238 , \12239 );
nor \U$11573 ( \12243 , \12241 , \12242 );
xor \U$11574 ( \12244 , \11370 , \12243 );
xnor \U$11575 ( \12245 , \12239 , \12238 );
and \U$11576 ( \12246 , \12190 , \12245 );
not \U$11577 ( \12247 , \12190 );
not \U$11578 ( \12248 , \12245 );
and \U$11579 ( \12249 , \12247 , \12248 );
nor \U$11580 ( \12250 , \12246 , \12249 );
not \U$11581 ( \12251 , \12250 );
xor \U$11582 ( \12252 , \12244 , \12251 );
not \U$11583 ( \12253 , \12250 );
not \U$11584 ( \12254 , \12253 );
and \U$11585 ( \12255 , \12015 , \12119 , \12169 );
not \U$11586 ( \12256 , \12255 );
not \U$11587 ( \12257 , \11946 );
or \U$11588 ( \12258 , \12256 , \12257 );
buf \U$11589 ( \12259 , \12183 );
nand \U$11590 ( \12260 , \12258 , \12259 );
not \U$11591 ( \12261 , \12260 );
not \U$11592 ( \12262 , \12187 );
nand \U$11593 ( \12263 , \12262 , \12067 );
not \U$11594 ( \12264 , \12263 );
and \U$11595 ( \12265 , \12261 , \12264 );
and \U$11596 ( \12266 , \12260 , \12263 );
nor \U$11597 ( \12267 , \12265 , \12266 );
not \U$11598 ( \12268 , \12267 );
not \U$11599 ( \12269 , \12268 );
or \U$11600 ( \12270 , \12254 , \12269 );
nand \U$11601 ( \12271 , \12267 , \12250 );
nand \U$11602 ( \12272 , \12270 , \12271 );
not \U$11603 ( \12273 , \12272 );
nand \U$11604 ( \12274 , \12252 , \12273 );
not \U$11605 ( \12275 , \12274 );
buf \U$11606 ( \12276 , \12244 );
not \U$11607 ( \12277 , \12276 );
nand \U$11608 ( \12278 , \12275 , \12277 );
not \U$11609 ( \12279 , \12278 );
buf \U$11610 ( \12280 , \12279 );
not \U$11611 ( \12281 , \12280 );
not \U$11612 ( \12282 , \12281 );
not \U$11613 ( \12283 , \11430 );
not \U$11614 ( \12284 , \12283 );
not \U$11615 ( \12285 , \11447 );
not \U$11616 ( \12286 , \12285 );
or \U$11617 ( \12287 , \12284 , \12286 );
not \U$11618 ( \12288 , \11417 );
or \U$11619 ( \12289 , \12284 , \12288 );
nand \U$11620 ( \12290 , \12287 , \12289 );
not \U$11621 ( \12291 , \12290 );
nand \U$11622 ( \12292 , \12284 , \12286 , \12288 );
nand \U$11623 ( \12293 , \12291 , \12292 );
buf \U$11624 ( \12294 , \12293 );
not \U$11625 ( \12295 , \12294 );
buf \U$11626 ( \12296 , \11454 );
not \U$11627 ( \12297 , \12296 );
not \U$11628 ( \12298 , \12297 );
buf \U$11629 ( \12299 , \11445 );
not \U$11630 ( \12300 , \12285 );
nand \U$11631 ( \12301 , \12299 , \12300 , \12288 );
not \U$11632 ( \12302 , \12301 );
or \U$11633 ( \12303 , \12298 , \12302 );
nand \U$11634 ( \12304 , \12299 , \12296 , \12286 , \12288 );
nand \U$11635 ( \12305 , \12303 , \12304 );
not \U$11636 ( \12306 , \12305 );
nor \U$11637 ( \12307 , \12295 , \12306 );
buf \U$11638 ( \12308 , \11502 );
not \U$11639 ( \12309 , \12308 );
not \U$11640 ( \12310 , \12309 );
not \U$11641 ( \12311 , \12301 );
or \U$11642 ( \12312 , \12310 , \12311 );
and \U$11643 ( \12313 , \12299 , \12300 , \12288 );
nor \U$11644 ( \12314 , \12297 , \12309 );
and \U$11645 ( \12315 , \12313 , \12314 );
nor \U$11646 ( \12316 , \12315 , \11483 );
nand \U$11647 ( \12317 , \12312 , \12316 );
not \U$11648 ( \12318 , \12317 );
not \U$11649 ( \12319 , \12318 );
not \U$11650 ( \12320 , \11421 );
not \U$11651 ( \12321 , \12288 );
and \U$11652 ( \12322 , \12320 , \12321 );
not \U$11653 ( \12323 , \11412 );
nor \U$11654 ( \12324 , \12322 , \12323 );
buf \U$11655 ( \12325 , \12324 );
and \U$11656 ( \12326 , \12307 , \12319 , \12325 );
buf \U$11657 ( \12327 , \12326 );
nand \U$11658 ( \12328 , \12327 , RIaa9ff60_293);
not \U$11659 ( \12329 , \12305 );
nand \U$11660 ( \12330 , \12329 , \12294 );
not \U$11661 ( \12331 , \12330 );
buf \U$11662 ( \12332 , \12317 );
buf \U$11663 ( \12333 , \12324 );
and \U$11664 ( \12334 , \12331 , \12332 , \12333 );
buf \U$11665 ( \12335 , \12334 );
nand \U$11666 ( \12336 , \12335 , RIaa9fd80_289);
nor \U$11667 ( \12337 , \12306 , \12294 );
nand \U$11668 ( \12338 , \12332 , \12337 , \12325 );
not \U$11669 ( \12339 , \12338 );
nand \U$11670 ( \12340 , \12339 , RIaa9fe70_291);
not \U$11671 ( \12341 , \12332 );
and \U$11672 ( \12342 , \12305 , \12294 );
nand \U$11673 ( \12343 , \12341 , \12342 , \12333 );
not \U$11674 ( \12344 , \12343 );
buf \U$11675 ( \12345 , \12344 );
nand \U$11676 ( \12346 , \12345 , RIaaa0140_297);
nand \U$11677 ( \12347 , \12328 , \12336 , \12340 , \12346 );
not \U$11678 ( \12348 , \12333 );
nor \U$11679 ( \12349 , \12348 , \12332 );
nand \U$11680 ( \12350 , \12349 , \12331 );
not \U$11681 ( \12351 , \12350 );
nand \U$11682 ( \12352 , \12351 , RIaa9fd08_288);
not \U$11683 ( \12353 , \12324 );
nand \U$11684 ( \12354 , \12318 , \12353 );
nor \U$11685 ( \12355 , \12330 , \12354 );
buf \U$11686 ( \12356 , \12355 );
nand \U$11687 ( \12357 , \12356 , RIaaa01b8_298);
not \U$11688 ( \12358 , \12354 );
nand \U$11689 ( \12359 , \12358 , \12307 );
not \U$11690 ( \12360 , \12359 );
nand \U$11691 ( \12361 , \12360 , RIaa9fdf8_290);
not \U$11692 ( \12362 , \12332 );
nor \U$11693 ( \12363 , \12362 , \12325 );
nand \U$11694 ( \12364 , \12363 , \12331 );
not \U$11695 ( \12365 , \12364 );
nand \U$11696 ( \12366 , \12365 , RIaa9fc90_287);
nand \U$11697 ( \12367 , \12352 , \12357 , \12361 , \12366 );
nor \U$11698 ( \12368 , \12347 , \12367 );
not \U$11699 ( \12369 , RIaa9fee8_292);
not \U$11700 ( \12370 , \12294 );
nand \U$11701 ( \12371 , \12370 , \12329 );
not \U$11702 ( \12372 , \12371 );
nand \U$11703 ( \12373 , \12372 , \12319 , \12325 );
buf \U$11704 ( \12374 , \12373 );
not \U$11705 ( \12375 , \12374 );
not \U$11706 ( \12376 , \12375 );
or \U$11707 ( \12377 , \12369 , \12376 );
not \U$11708 ( \12378 , \12332 );
and \U$11709 ( \12379 , \12378 , \12306 , \12295 , \12333 );
buf \U$11710 ( \12380 , \12379 );
nand \U$11711 ( \12381 , \12380 , RIaa9fa38_282);
nand \U$11712 ( \12382 , \12377 , \12381 );
nand \U$11713 ( \12383 , \12363 , \12342 );
not \U$11714 ( \12384 , \12383 );
nand \U$11715 ( \12385 , \12384 , RIaa9ffd8_294);
nor \U$11716 ( \12386 , \12293 , \12324 );
nand \U$11717 ( \12387 , \12305 , \12386 );
or \U$11718 ( \12388 , \12318 , \12387 );
not \U$11719 ( \12389 , \12388 );
not \U$11720 ( \12390 , \12389 );
not \U$11721 ( \12391 , \12390 );
and \U$11722 ( \12392 , \12391 , RIaaa0050_295);
not \U$11723 ( \12393 , RIaa9fba0_285);
or \U$11724 ( \12394 , \12332 , \12387 );
not \U$11725 ( \12395 , \12394 );
not \U$11726 ( \12396 , \12395 );
nor \U$11727 ( \12397 , \12393 , \12396 );
nor \U$11728 ( \12398 , \12392 , \12397 );
not \U$11729 ( \12399 , \12305 );
buf \U$11730 ( \12400 , \12386 );
and \U$11731 ( \12401 , \12332 , \12399 , \12400 );
buf \U$11732 ( \12402 , \12401 );
and \U$11733 ( \12403 , \12402 , RIaa9fab0_283);
not \U$11734 ( \12404 , RIaa9fc18_286);
nor \U$11735 ( \12405 , \12308 , \12297 );
not \U$11736 ( \12406 , \12405 );
not \U$11737 ( \12407 , \12313 );
or \U$11738 ( \12408 , \12406 , \12407 );
not \U$11739 ( \12409 , RIaaa8a20_589);
nand \U$11740 ( \12410 , \12408 , \12409 );
not \U$11741 ( \12411 , \12410 );
or \U$11742 ( \12412 , \12404 , \12411 );
nand \U$11743 ( \12413 , \11473 , RIaa9fb28_284);
nand \U$11744 ( \12414 , \12412 , \12413 );
nor \U$11745 ( \12415 , \12403 , \12414 );
nand \U$11746 ( \12416 , \12318 , \12306 , \12400 );
buf \U$11747 ( \12417 , \12416 );
not \U$11748 ( \12418 , \12417 );
nand \U$11749 ( \12419 , \12418 , RIaaa00c8_296);
nand \U$11750 ( \12420 , \12385 , \12398 , \12415 , \12419 );
nor \U$11751 ( \12421 , \12382 , \12420 );
nand \U$11752 ( \12422 , \12368 , \12421 );
buf \U$11753 ( \12423 , \12422 );
not \U$11754 ( \12424 , \12423 );
buf \U$11755 ( \12425 , \12424 );
not \U$11756 ( \12426 , \12425 );
not \U$11757 ( \12427 , \12426 );
and \U$11758 ( \12428 , \12282 , \12427 );
buf \U$11759 ( \12429 , \12244 );
buf \U$11760 ( \12430 , \12429 );
nand \U$11761 ( \12431 , \12275 , \12430 );
not \U$11762 ( \12432 , \12431 );
not \U$11763 ( \12433 , \12432 );
or \U$11764 ( \12434 , \12433 , \12425 );
nand \U$11765 ( \12435 , \12272 , \12277 );
buf \U$11766 ( \12436 , \12435 );
buf \U$11767 ( \12437 , \12436 );
not \U$11768 ( \12438 , \12437 );
not \U$11769 ( \12439 , \12327 );
not \U$11770 ( \12440 , \12439 );
not \U$11771 ( \12441 , \6961 );
and \U$11772 ( \12442 , \12440 , \12441 );
not \U$11773 ( \12443 , RIaa9f7e0_277);
nor \U$11774 ( \12444 , \12374 , \12443 );
nor \U$11775 ( \12445 , \12442 , \12444 );
not \U$11776 ( \12446 , \12350 );
and \U$11777 ( \12447 , \12446 , RIaa9f948_280);
not \U$11778 ( \12448 , \12334 );
not \U$11779 ( \12449 , \12448 );
and \U$11780 ( \12450 , \12449 , RIaa9f9c0_281);
nor \U$11781 ( \12451 , \12447 , \12450 );
buf \U$11782 ( \12452 , \12343 );
not \U$11783 ( \12453 , \12452 );
and \U$11784 ( \12454 , \12453 , RIaa9f330_267);
not \U$11785 ( \12455 , \12383 );
and \U$11786 ( \12456 , \12455 , RIaa9f6f0_275);
nor \U$11787 ( \12457 , \12454 , \12456 );
and \U$11788 ( \12458 , \12356 , RIaa9f2b8_266);
and \U$11789 ( \12459 , \12360 , RIaa9f420_269);
nor \U$11790 ( \12460 , \12458 , \12459 );
nand \U$11791 ( \12461 , \12445 , \12451 , \12457 , \12460 );
not \U$11792 ( \12462 , \12365 );
not \U$11793 ( \12463 , \12462 );
not \U$11794 ( \12464 , \6948 );
and \U$11795 ( \12465 , \12463 , \12464 );
not \U$11796 ( \12466 , RIaa9f8d0_279);
not \U$11797 ( \12467 , \12402 );
or \U$11798 ( \12468 , \12466 , \12467 );
not \U$11799 ( \12469 , \12417 );
nand \U$11800 ( \12470 , \12469 , RIaa9f498_270);
nand \U$11801 ( \12471 , \12468 , \12470 );
nor \U$11802 ( \12472 , \12465 , \12471 );
nand \U$11803 ( \12473 , \12339 , RIaa9f768_276);
nand \U$11804 ( \12474 , \12380 , RIaa9f858_278);
not \U$11805 ( \12475 , RIaa9f3a8_268);
not \U$11806 ( \12476 , \12388 );
not \U$11807 ( \12477 , \12476 );
or \U$11808 ( \12478 , \12475 , \12477 );
and \U$11809 ( \12479 , \12410 , RIaa9f588_272);
nand \U$11810 ( \12480 , \11473 , RIaa9f240_265);
not \U$11811 ( \12481 , \12480 );
nor \U$11812 ( \12482 , \12479 , \12481 );
nand \U$11813 ( \12483 , \12478 , \12482 );
not \U$11814 ( \12484 , RIaa9f510_271);
nor \U$11815 ( \12485 , \12484 , \12396 );
nor \U$11816 ( \12486 , \12483 , \12485 );
nand \U$11817 ( \12487 , \12472 , \12473 , \12474 , \12486 );
nor \U$11818 ( \12488 , \12461 , \12487 );
buf \U$11819 ( \12489 , \12488 );
not \U$11820 ( \12490 , \12489 );
not \U$11821 ( \12491 , \12490 );
and \U$11822 ( \12492 , \12438 , \12491 );
not \U$11823 ( \12493 , \12429 );
not \U$11824 ( \12494 , \12493 );
nand \U$11825 ( \12495 , \12494 , \12272 );
not \U$11826 ( \12496 , \12495 );
not \U$11827 ( \12497 , \12491 );
and \U$11828 ( \12498 , \12496 , \12497 );
nor \U$11829 ( \12499 , \12492 , \12498 );
nand \U$11830 ( \12500 , \12434 , \12499 );
nor \U$11831 ( \12501 , \12428 , \12500 );
not \U$11832 ( \12502 , \12439 );
nand \U$11833 ( \12503 , \12502 , RIaa9ee80_257);
nand \U$11834 ( \12504 , \12339 , RIaa9f0d8_262);
not \U$11835 ( \12505 , \12379 );
not \U$11836 ( \12506 , \12505 );
nand \U$11837 ( \12507 , \12506 , RIaa9f150_263);
nand \U$11838 ( \12508 , \12446 , RIaa9ef70_259);
nand \U$11839 ( \12509 , \12503 , \12504 , \12507 , \12508 );
not \U$11840 ( \12510 , RIaa9f060_261);
not \U$11841 ( \12511 , \12375 );
or \U$11842 ( \12512 , \12510 , \12511 );
buf \U$11843 ( \12513 , \12402 );
and \U$11844 ( \12514 , \12513 , RIaa9f1c8_264);
and \U$11845 ( \12515 , \12391 , RIaa9ed18_254);
not \U$11846 ( \12516 , RIaa9ebb0_251);
not \U$11847 ( \12517 , \12410 );
or \U$11848 ( \12518 , \12516 , \12517 );
nand \U$11849 ( \12519 , \11473 , RIaa9ea48_248);
nand \U$11850 ( \12520 , \12518 , \12519 );
nor \U$11851 ( \12521 , \12514 , \12515 , \12520 );
nand \U$11852 ( \12522 , \12512 , \12521 );
nor \U$11853 ( \12523 , \12509 , \12522 );
nand \U$11854 ( \12524 , \12453 , RIaa9eca0_253);
nand \U$11855 ( \12525 , \12356 , RIaa9ec28_252);
nand \U$11856 ( \12526 , \12365 , RIaa9eb38_250);
nand \U$11857 ( \12527 , \12384 , RIaa9eef8_258);
nand \U$11858 ( \12528 , \12524 , \12525 , \12526 , \12527 );
not \U$11859 ( \12529 , RIaa9efe8_260);
not \U$11860 ( \12530 , \12335 );
or \U$11861 ( \12531 , \12529 , \12530 );
not \U$11862 ( \12532 , \12359 );
buf \U$11863 ( \12533 , \12532 );
and \U$11864 ( \12534 , \12533 , RIaa9ee08_256);
not \U$11865 ( \12535 , RIaa9ed90_255);
not \U$11866 ( \12536 , \12469 );
or \U$11867 ( \12537 , \12535 , \12536 );
nand \U$11868 ( \12538 , \12395 , RIaa9eac0_249);
nand \U$11869 ( \12539 , \12537 , \12538 );
nor \U$11870 ( \12540 , \12534 , \12539 );
nand \U$11871 ( \12541 , \12531 , \12540 );
nor \U$11872 ( \12542 , \12528 , \12541 );
nand \U$11873 ( \12543 , \12523 , \12542 );
not \U$11874 ( \12544 , \12543 );
not \U$11875 ( \12545 , \12544 );
not \U$11876 ( \12546 , \12267 );
not \U$11877 ( \12547 , \12546 );
not \U$11878 ( \12548 , \12119 );
nand \U$11879 ( \12549 , \11945 , \12169 );
or \U$11880 ( \12550 , \12548 , \12549 );
not \U$11881 ( \12551 , \12180 );
nand \U$11882 ( \12552 , \12550 , \12551 );
not \U$11883 ( \12553 , \12182 );
nand \U$11884 ( \12554 , \12553 , \12015 );
not \U$11885 ( \12555 , \12554 );
and \U$11886 ( \12556 , \12552 , \12555 );
not \U$11887 ( \12557 , \12552 );
and \U$11888 ( \12558 , \12557 , \12554 );
nor \U$11889 ( \12559 , \12556 , \12558 );
not \U$11890 ( \12560 , \12559 );
or \U$11891 ( \12561 , \12547 , \12560 );
buf \U$11892 ( \12562 , \12559 );
buf \U$11893 ( \12563 , \12267 );
not \U$11894 ( \12564 , \12563 );
or \U$11895 ( \12565 , \12562 , \12564 );
nand \U$11896 ( \12566 , \12561 , \12565 );
buf \U$11897 ( \12567 , \12179 );
nand \U$11898 ( \12568 , \12567 , \12119 );
not \U$11899 ( \12569 , \12568 );
not \U$11900 ( \12570 , \12569 );
not \U$11901 ( \12571 , \12173 );
nand \U$11902 ( \12572 , \12549 , \12571 );
not \U$11903 ( \12573 , \12572 );
not \U$11904 ( \12574 , \12573 );
or \U$11905 ( \12575 , \12570 , \12574 );
not \U$11906 ( \12576 , \12571 );
not \U$11907 ( \12577 , \12549 );
or \U$11908 ( \12578 , \12576 , \12577 );
nand \U$11909 ( \12579 , \12578 , \12568 );
nand \U$11910 ( \12580 , \12575 , \12579 );
xor \U$11911 ( \12581 , \12580 , \12559 );
nor \U$11912 ( \12582 , \12566 , \12581 );
not \U$11913 ( \12583 , \12564 );
nand \U$11914 ( \12584 , \12582 , \12583 );
not \U$11915 ( \12585 , \12584 );
and \U$11916 ( \12586 , \12545 , \12585 );
not \U$11917 ( \12587 , \12562 );
not \U$11918 ( \12588 , \12546 );
not \U$11919 ( \12589 , \12588 );
buf \U$11920 ( \12590 , \12572 );
not \U$11921 ( \12591 , \12590 );
not \U$11922 ( \12592 , \12568 );
and \U$11923 ( \12593 , \12591 , \12592 );
and \U$11924 ( \12594 , \12590 , \12568 );
nor \U$11925 ( \12595 , \12593 , \12594 );
nand \U$11926 ( \12596 , \12587 , \12589 , \12595 );
buf \U$11927 ( \12597 , \12596 );
buf \U$11928 ( \12598 , \12597 );
or \U$11929 ( \12599 , \12598 , \12545 );
and \U$11930 ( \12600 , \12581 , \12589 );
buf \U$11931 ( \12601 , \12600 );
not \U$11932 ( \12602 , \12601 );
nand \U$11933 ( \12603 , \12599 , \12602 );
nor \U$11934 ( \12604 , \12586 , \12603 );
and \U$11935 ( \12605 , \11370 , \12243 );
buf \U$11936 ( \12606 , \12605 );
not \U$11937 ( \12607 , \12455 );
nor \U$11938 ( \12608 , \12607 , \7221 );
nor \U$11939 ( \12609 , \12462 , \7240 );
nor \U$11940 ( \12610 , \12608 , \12609 );
and \U$11941 ( \12611 , \12533 , RIaaa0410_303);
not \U$11942 ( \12612 , \12476 );
not \U$11943 ( \12613 , \12612 );
and \U$11944 ( \12614 , \12613 , RIaaa0488_304);
nor \U$11945 ( \12615 , \12611 , \12614 );
nand \U$11946 ( \12616 , \12610 , \12615 );
not \U$11947 ( \12617 , RIaaa0230_299);
not \U$11948 ( \12618 , \12339 );
or \U$11949 ( \12619 , \12617 , \12618 );
nand \U$11950 ( \12620 , \12345 , RIaaa0668_308);
nand \U$11951 ( \12621 , \12619 , \12620 );
nor \U$11952 ( \12622 , \12616 , \12621 );
not \U$11953 ( \12623 , RIaaa0578_306);
not \U$11954 ( \12624 , \12502 );
or \U$11955 ( \12625 , \12623 , \12624 );
nand \U$11956 ( \12626 , \12449 , RIaaa0398_302);
nand \U$11957 ( \12627 , \12625 , \12626 );
not \U$11958 ( \12628 , RIaaa02a8_300);
not \U$11959 ( \12629 , \12375 );
or \U$11960 ( \12630 , \12628 , \12629 );
nand \U$11961 ( \12631 , \12506 , RIaaa0938_314);
nand \U$11962 ( \12632 , \12630 , \12631 );
nor \U$11963 ( \12633 , \12627 , \12632 );
not \U$11964 ( \12634 , RIaaa0320_301);
not \U$11965 ( \12635 , \12351 );
or \U$11966 ( \12636 , \12634 , \12635 );
nand \U$11967 ( \12637 , \12356 , RIaaa06e0_309);
nand \U$11968 ( \12638 , \12636 , \12637 );
not \U$11969 ( \12639 , \12396 );
not \U$11970 ( \12640 , \7248 );
and \U$11971 ( \12641 , \12639 , \12640 );
and \U$11972 ( \12642 , \12513 , RIaaa08c0_313);
nor \U$11973 ( \12643 , \12641 , \12642 );
and \U$11974 ( \12644 , \12469 , RIaaa0500_305);
not \U$11975 ( \12645 , RIaaa07d0_311);
not \U$11976 ( \12646 , \12410 );
or \U$11977 ( \12647 , \12645 , \12646 );
nand \U$11978 ( \12648 , \11473 , RIaaa09b0_315);
nand \U$11979 ( \12649 , \12647 , \12648 );
nor \U$11980 ( \12650 , \12644 , \12649 );
nand \U$11981 ( \12651 , \12643 , \12650 );
nor \U$11982 ( \12652 , \12638 , \12651 );
nand \U$11983 ( \12653 , \12622 , \12633 , \12652 );
not \U$11984 ( \12654 , \12653 );
not \U$11985 ( \12655 , \12654 );
not \U$11986 ( \12656 , \12655 );
not \U$11987 ( \12657 , \12656 );
not \U$11988 ( \12658 , \12657 );
not \U$11989 ( \12659 , \12658 );
nand \U$11990 ( \12660 , \12606 , \12659 );
and \U$11991 ( \12661 , \12604 , \12660 );
and \U$11992 ( \12662 , \12501 , \12661 );
not \U$11993 ( \12663 , \12562 );
not \U$11994 ( \12664 , \12580 );
not \U$11995 ( \12665 , \12664 );
not \U$11996 ( \12666 , \12665 );
or \U$11997 ( \12667 , \12663 , \12666 );
buf \U$11998 ( \12668 , \12588 );
not \U$11999 ( \12669 , \12668 );
nand \U$12000 ( \12670 , \12667 , \12669 );
not \U$12001 ( \12671 , \12670 );
not \U$12002 ( \12672 , \12671 );
nand \U$12003 ( \12673 , \12606 , \12426 );
nand \U$12004 ( \12674 , \12672 , \12673 );
not \U$12005 ( \12675 , \12674 );
not \U$12006 ( \12676 , \12272 );
not \U$12007 ( \12677 , \12676 );
not \U$12008 ( \12678 , \12677 );
not \U$12009 ( \12679 , \12678 );
and \U$12010 ( \12680 , \12497 , \12430 );
not \U$12011 ( \12681 , \12497 );
not \U$12012 ( \12682 , \12430 );
and \U$12013 ( \12683 , \12681 , \12682 );
nor \U$12014 ( \12684 , \12680 , \12683 );
not \U$12015 ( \12685 , \12684 );
or \U$12016 ( \12686 , \12679 , \12685 );
not \U$12017 ( \12687 , \12275 );
or \U$12018 ( \12688 , \12430 , \12544 );
and \U$12019 ( \12689 , \12430 , \12544 );
nor \U$12020 ( \12690 , \12689 , \12678 );
nand \U$12021 ( \12691 , \12688 , \12690 );
nand \U$12022 ( \12692 , \12687 , \12691 );
nand \U$12023 ( \12693 , \12686 , \12692 );
not \U$12024 ( \12694 , \12693 );
or \U$12025 ( \12695 , \12675 , \12694 );
or \U$12026 ( \12696 , \12693 , \12674 );
nand \U$12027 ( \12697 , \12695 , \12696 );
nor \U$12028 ( \12698 , \12662 , \12697 );
or \U$12029 ( \12699 , \12281 , \12545 );
nand \U$12030 ( \12700 , \12432 , \12545 );
nand \U$12031 ( \12701 , \12699 , \12700 , \12437 );
not \U$12032 ( \12702 , \12701 );
nand \U$12033 ( \12703 , \12606 , \12497 );
nand \U$12034 ( \12704 , \12702 , \12703 );
not \U$12035 ( \12705 , \12687 );
or \U$12036 ( \12706 , \12705 , \12677 );
not \U$12037 ( \12707 , \12606 );
or \U$12038 ( \12708 , \12544 , \12707 );
nand \U$12039 ( \12709 , \12706 , \12708 , \12682 );
or \U$12040 ( \12710 , \12709 , \12703 );
nand \U$12041 ( \12711 , \12704 , \12710 );
and \U$12042 ( \12712 , \12693 , \12673 );
nor \U$12043 ( \12713 , \12712 , \12671 );
xor \U$12044 ( \12714 , \12711 , \12713 );
or \U$12045 ( \12715 , \12698 , \12714 );
not \U$12046 ( \12716 , \12715 );
not \U$12047 ( \12717 , \12665 );
buf \U$12048 ( \12718 , \11924 );
not \U$12049 ( \12719 , \11940 );
nor \U$12050 ( \12720 , \12719 , \11942 );
nor \U$12051 ( \12721 , \12718 , \12720 );
not \U$12052 ( \12722 , \12721 );
buf \U$12053 ( \12723 , \11726 );
not \U$12054 ( \12724 , \12723 );
nor \U$12055 ( \12725 , \11546 , \11918 );
not \U$12056 ( \12726 , \12725 );
nand \U$12057 ( \12727 , \11913 , \11862 );
not \U$12058 ( \12728 , \12727 );
or \U$12059 ( \12729 , \12726 , \12728 );
buf \U$12060 ( \12730 , \11538 );
nand \U$12061 ( \12731 , \12730 , \11545 );
nand \U$12062 ( \12732 , \12729 , \12731 );
not \U$12063 ( \12733 , \12732 );
or \U$12064 ( \12734 , \12724 , \12733 );
not \U$12065 ( \12735 , \11933 );
not \U$12066 ( \12736 , \11930 );
or \U$12067 ( \12737 , \12735 , \12736 );
buf \U$12068 ( \12738 , \11725 );
nand \U$12069 ( \12739 , \12737 , \12738 );
nand \U$12070 ( \12740 , \12734 , \12739 );
not \U$12071 ( \12741 , \12740 );
or \U$12072 ( \12742 , \12722 , \12741 );
not \U$12073 ( \12743 , \12732 );
not \U$12074 ( \12744 , \12743 );
nand \U$12075 ( \12745 , \12744 , \12723 );
buf \U$12076 ( \12746 , \11937 );
and \U$12077 ( \12747 , \12739 , \12720 , \12746 );
and \U$12078 ( \12748 , \12745 , \12747 );
not \U$12079 ( \12749 , \12718 );
not \U$12080 ( \12750 , \12720 );
or \U$12081 ( \12751 , \12749 , \12750 );
or \U$12082 ( \12752 , \12720 , \12746 );
nand \U$12083 ( \12753 , \12751 , \12752 );
nor \U$12084 ( \12754 , \12748 , \12753 );
nand \U$12085 ( \12755 , \12742 , \12754 );
not \U$12086 ( \12756 , \12755 );
not \U$12087 ( \12757 , \11946 );
buf \U$12088 ( \12758 , \12169 );
nand \U$12089 ( \12759 , \12571 , \12758 );
not \U$12090 ( \12760 , \12759 );
and \U$12091 ( \12761 , \12757 , \12760 );
and \U$12092 ( \12762 , \12759 , \11946 );
nor \U$12093 ( \12763 , \12761 , \12762 );
not \U$12094 ( \12764 , \12763 );
and \U$12095 ( \12765 , \12756 , \12764 );
not \U$12096 ( \12766 , \12756 );
and \U$12097 ( \12767 , \12766 , \12763 );
nor \U$12098 ( \12768 , \12765 , \12767 );
buf \U$12099 ( \12769 , \12768 );
nor \U$12100 ( \12770 , \12717 , \12769 );
not \U$12101 ( \12771 , \12770 );
not \U$12102 ( \12772 , \12424 );
or \U$12103 ( \12773 , \12771 , \12772 );
not \U$12104 ( \12774 , \12763 );
nor \U$12105 ( \12775 , \12580 , \12774 );
not \U$12106 ( \12776 , \12775 );
nand \U$12107 ( \12777 , \12580 , \12774 );
nand \U$12108 ( \12778 , \12776 , \12777 , \12768 );
buf \U$12109 ( \12779 , \12778 );
not \U$12110 ( \12780 , \12779 );
not \U$12111 ( \12781 , \12780 );
buf \U$12112 ( \12782 , \12580 );
not \U$12113 ( \12783 , \12782 );
and \U$12114 ( \12784 , \12783 , \12655 );
not \U$12115 ( \12785 , \12783 );
and \U$12116 ( \12786 , \12785 , \12656 );
or \U$12117 ( \12787 , \12784 , \12786 );
not \U$12118 ( \12788 , \12787 );
or \U$12119 ( \12789 , \12781 , \12788 );
nand \U$12120 ( \12790 , \12773 , \12789 );
not \U$12121 ( \12791 , \12374 );
not \U$12122 ( \12792 , RIaaa2378_370);
not \U$12123 ( \12793 , \12792 );
and \U$12124 ( \12794 , \12791 , \12793 );
nor \U$12125 ( \12795 , \12505 , \2453 );
nor \U$12126 ( \12796 , \12794 , \12795 );
not \U$12127 ( \12797 , \12384 );
not \U$12128 ( \12798 , \12797 );
not \U$12129 ( \12799 , \7989 );
and \U$12130 ( \12800 , \12798 , \12799 );
not \U$12131 ( \12801 , RIaaa25d0_375);
not \U$12132 ( \12802 , \12469 );
or \U$12133 ( \12803 , \12801 , \12802 );
nand \U$12134 ( \12804 , \12402 , RIaaa27b0_379);
nand \U$12135 ( \12805 , \12803 , \12804 );
nor \U$12136 ( \12806 , \12800 , \12805 );
and \U$12137 ( \12807 , \12613 , RIaaa2558_374);
not \U$12138 ( \12808 , RIaaa28a0_381);
not \U$12139 ( \12809 , \12410 );
or \U$12140 ( \12810 , \12808 , \12809 );
and \U$12141 ( \12811 , \11473 , RIaaa2990_383);
not \U$12142 ( \12812 , \12811 );
nand \U$12143 ( \12813 , \12810 , \12812 );
nor \U$12144 ( \12814 , \12807 , \12813 );
nand \U$12145 ( \12815 , \12395 , RIaaa2828_380);
and \U$12146 ( \12816 , \12814 , \12815 );
nand \U$12147 ( \12817 , \12796 , \12806 , \12816 );
and \U$12148 ( \12818 , \12342 , \12332 , \12333 );
and \U$12149 ( \12819 , \12818 , RIaaa2468_372);
and \U$12150 ( \12820 , \12344 , RIaaa2648_376);
nor \U$12151 ( \12821 , \12819 , \12820 );
and \U$12152 ( \12822 , \12449 , RIaaa2210_367);
and \U$12153 ( \12823 , \12339 , RIaaa2300_369);
nor \U$12154 ( \12824 , \12822 , \12823 );
and \U$12155 ( \12825 , \12356 , RIaaa26c0_377);
and \U$12156 ( \12826 , \12532 , RIaaa23f0_371);
nor \U$12157 ( \12827 , \12825 , \12826 );
nand \U$12158 ( \12828 , \12331 , \12341 , \12333 );
not \U$12159 ( \12829 , \12828 );
and \U$12160 ( \12830 , \12829 , RIaaa2288_368);
nor \U$12161 ( \12831 , \12378 , \12325 );
nand \U$12162 ( \12832 , \12831 , \12331 );
not \U$12163 ( \12833 , \12832 );
and \U$12164 ( \12834 , \12833 , RIaaa2918_382);
nor \U$12165 ( \12835 , \12830 , \12834 );
nand \U$12166 ( \12836 , \12821 , \12824 , \12827 , \12835 );
nor \U$12167 ( \12837 , \12817 , \12836 );
buf \U$12168 ( \12838 , \12837 );
not \U$12169 ( \12839 , \12838 );
not \U$12170 ( \12840 , \12839 );
buf \U$12171 ( \12841 , \12605 );
not \U$12172 ( \12842 , \12841 );
or \U$12173 ( \12843 , \12840 , \12842 );
not \U$12174 ( \12844 , \12580 );
not \U$12175 ( \12845 , \12768 );
nand \U$12176 ( \12846 , \12844 , \12845 );
or \U$12177 ( \12847 , \12846 , \12424 );
nand \U$12178 ( \12848 , \12843 , \12847 );
nor \U$12179 ( \12849 , \12790 , \12848 );
not \U$12180 ( \12850 , \12545 );
buf \U$12181 ( \12851 , \11675 );
nand \U$12182 ( \12852 , \11930 , \12851 );
not \U$12183 ( \12853 , \12852 );
not \U$12184 ( \12854 , \12743 );
not \U$12185 ( \12855 , \12854 );
or \U$12186 ( \12856 , \12853 , \12855 );
not \U$12187 ( \12857 , \12852 );
nand \U$12188 ( \12858 , \12743 , \12857 );
nand \U$12189 ( \12859 , \12856 , \12858 );
not \U$12190 ( \12860 , \12859 );
not \U$12191 ( \12861 , \12860 );
not \U$12192 ( \12862 , \12861 );
not \U$12193 ( \12863 , \12851 );
not \U$12194 ( \12864 , \12732 );
or \U$12195 ( \12865 , \12863 , \12864 );
nand \U$12196 ( \12866 , \12865 , \11930 );
and \U$12197 ( \12867 , \11933 , \12738 );
and \U$12198 ( \12868 , \12866 , \12867 );
not \U$12199 ( \12869 , \12866 );
not \U$12200 ( \12870 , \12867 );
and \U$12201 ( \12871 , \12869 , \12870 );
nor \U$12202 ( \12872 , \12868 , \12871 );
not \U$12203 ( \12873 , \12872 );
not \U$12204 ( \12874 , \12873 );
not \U$12205 ( \12875 , \12874 );
or \U$12206 ( \12876 , \12862 , \12875 );
not \U$12207 ( \12877 , \12872 );
and \U$12208 ( \12878 , \12877 , \12860 );
buf \U$12209 ( \12879 , \11920 );
not \U$12210 ( \12880 , \11546 );
nand \U$12211 ( \12881 , \12880 , \12731 );
xnor \U$12212 ( \12882 , \12879 , \12881 );
not \U$12213 ( \12883 , \12882 );
not \U$12214 ( \12884 , \12859 );
or \U$12215 ( \12885 , \12883 , \12884 );
not \U$12216 ( \12886 , \12881 );
and \U$12217 ( \12887 , \12879 , \12886 );
not \U$12218 ( \12888 , \12879 );
and \U$12219 ( \12889 , \12888 , \12881 );
nor \U$12220 ( \12890 , \12887 , \12889 );
or \U$12221 ( \12891 , \12859 , \12890 );
nand \U$12222 ( \12892 , \12885 , \12891 );
nor \U$12223 ( \12893 , \12878 , \12892 );
nand \U$12224 ( \12894 , \12876 , \12893 );
buf \U$12225 ( \12895 , \12874 );
nor \U$12226 ( \12896 , \12894 , \12895 );
buf \U$12227 ( \12897 , \12896 );
buf \U$12228 ( \12898 , \12897 );
not \U$12229 ( \12899 , \12898 );
or \U$12230 ( \12900 , \12850 , \12899 );
not \U$12231 ( \12901 , \12872 );
buf \U$12232 ( \12902 , \12901 );
or \U$12233 ( \12903 , \12894 , \12902 );
not \U$12234 ( \12904 , \12903 );
and \U$12235 ( \12905 , \12904 , \12544 );
not \U$12236 ( \12906 , \12901 );
not \U$12237 ( \12907 , \12892 );
not \U$12238 ( \12908 , \12907 );
nand \U$12239 ( \12909 , \12906 , \12908 );
not \U$12240 ( \12910 , \12909 );
buf \U$12241 ( \12911 , \12910 );
not \U$12242 ( \12912 , \12911 );
not \U$12243 ( \12913 , \12912 );
nor \U$12244 ( \12914 , \12905 , \12913 );
nand \U$12245 ( \12915 , \12900 , \12914 );
not \U$12246 ( \12916 , \12915 );
and \U$12247 ( \12917 , \12849 , \12916 );
not \U$12248 ( \12918 , \12849 );
and \U$12249 ( \12919 , \12918 , \12915 );
or \U$12250 ( \12920 , \12917 , \12919 );
not \U$12251 ( \12921 , \12920 );
not \U$12252 ( \12922 , \12916 );
not \U$12253 ( \12923 , \12839 );
not \U$12254 ( \12924 , \12430 );
or \U$12255 ( \12925 , \12923 , \12924 );
or \U$12256 ( \12926 , \12430 , \12839 );
nand \U$12257 ( \12927 , \12925 , \12926 );
not \U$12258 ( \12928 , \12927 );
not \U$12259 ( \12929 , \12275 );
or \U$12260 ( \12930 , \12928 , \12929 );
not \U$12261 ( \12931 , \12373 );
and \U$12262 ( \12932 , \12931 , RIaaa2cd8_390);
and \U$12263 ( \12933 , \12327 , RIaaa2a80_385);
nor \U$12264 ( \12934 , \12932 , \12933 );
and \U$12265 ( \12935 , \12335 , RIaaa2dc8_392);
and \U$12266 ( \12936 , \12339 , RIaaa2d50_391);
nor \U$12267 ( \12937 , \12935 , \12936 );
nand \U$12268 ( \12938 , \12934 , \12937 );
not \U$12269 ( \12939 , \12390 );
not \U$12270 ( \12940 , RIaaa2b70_387);
not \U$12271 ( \12941 , \12940 );
and \U$12272 ( \12942 , \12939 , \12941 );
and \U$12273 ( \12943 , \12365 , RIaaa3098_398);
nor \U$12274 ( \12944 , \12942 , \12943 );
nand \U$12275 ( \12945 , \12345 , RIaaa2c60_389);
nand \U$12276 ( \12946 , \12351 , RIaaa2e40_393);
nand \U$12277 ( \12947 , \12944 , \12945 , \12946 );
nor \U$12278 ( \12948 , \12938 , \12947 );
nand \U$12279 ( \12949 , \12356 , RIaaa2be8_388);
and \U$12280 ( \12950 , \12469 , RIaaa2af8_386);
not \U$12281 ( \12951 , \12394 );
buf \U$12282 ( \12952 , \12951 );
and \U$12283 ( \12953 , \12952 , RIaaa3020_397);
nor \U$12284 ( \12954 , \12950 , \12953 );
nand \U$12285 ( \12955 , \12455 , RIaaa2a08_384);
and \U$12286 ( \12956 , \12402 , RIaaa2f30_395);
not \U$12287 ( \12957 , RIaaa3110_399);
not \U$12288 ( \12958 , \12410 );
or \U$12289 ( \12959 , \12957 , \12958 );
nand \U$12290 ( \12960 , \11473 , RIaaa3188_400);
nand \U$12291 ( \12961 , \12959 , \12960 );
nor \U$12292 ( \12962 , \12956 , \12961 );
nand \U$12293 ( \12963 , \12949 , \12954 , \12955 , \12962 );
not \U$12294 ( \12964 , RIaaa2fa8_396);
not \U$12295 ( \12965 , \12506 );
or \U$12296 ( \12966 , \12964 , \12965 );
nand \U$12297 ( \12967 , \12360 , RIaaa2eb8_394);
nand \U$12298 ( \12968 , \12966 , \12967 );
nor \U$12299 ( \12969 , \12963 , \12968 );
nand \U$12300 ( \12970 , \12948 , \12969 );
buf \U$12301 ( \12971 , \12970 );
and \U$12302 ( \12972 , \12971 , \12495 );
not \U$12303 ( \12973 , \12971 );
and \U$12304 ( \12974 , \12973 , \12436 );
or \U$12305 ( \12975 , \12972 , \12974 );
nand \U$12306 ( \12976 , \12930 , \12975 );
not \U$12307 ( \12977 , \12976 );
or \U$12308 ( \12978 , \12922 , \12977 );
and \U$12309 ( \12979 , \12345 , RIaaa3f20_429);
and \U$12310 ( \12980 , \12327 , RIaaa39f8_418);
nor \U$12311 ( \12981 , \12979 , \12980 );
and \U$12312 ( \12982 , \12335 , RIaaa3d40_425);
and \U$12313 ( \12983 , \12339 , RIaaa3ae8_420);
nor \U$12314 ( \12984 , \12982 , \12983 );
nand \U$12315 ( \12985 , \12981 , \12984 );
and \U$12316 ( \12986 , \12446 , RIaaa3cc8_424);
and \U$12317 ( \12987 , \12365 , RIaaa4178_434);
nor \U$12318 ( \12988 , \12986 , \12987 );
and \U$12319 ( \12989 , \12356 , RIaaa3e30_427);
and \U$12320 ( \12990 , \12360 , RIaaa3f98_430);
nor \U$12321 ( \12991 , \12989 , \12990 );
nand \U$12322 ( \12992 , \12988 , \12991 );
nor \U$12323 ( \12993 , \12985 , \12992 );
not \U$12324 ( \12994 , RIaaa3b60_421);
not \U$12325 ( \12995 , \12931 );
or \U$12326 ( \12996 , \12994 , \12995 );
nand \U$12327 ( \12997 , \12506 , RIaaa3bd8_422);
nand \U$12328 ( \12998 , \12996 , \12997 );
not \U$12329 ( \12999 , \12612 );
not \U$12330 ( \13000 , RIaaa3ea8_428);
not \U$12331 ( \13001 , \13000 );
and \U$12332 ( \13002 , \12999 , \13001 );
and \U$12333 ( \13003 , \12418 , RIaaa4010_431);
nor \U$12334 ( \13004 , \13002 , \13003 );
nand \U$12335 ( \13005 , \12455 , RIaaa3a70_419);
not \U$12336 ( \13006 , \12401 );
not \U$12337 ( \13007 , \13006 );
and \U$12338 ( \13008 , \13007 , RIaaa3c50_423);
not \U$12339 ( \13009 , RIaaa4100_433);
not \U$12340 ( \13010 , \12410 );
or \U$12341 ( \13011 , \13009 , \13010 );
nand \U$12342 ( \13012 , \11473 , RIaaa3db8_426);
nand \U$12343 ( \13013 , \13011 , \13012 );
nor \U$12344 ( \13014 , \13008 , \13013 );
nand \U$12345 ( \13015 , \12952 , RIaaa4088_432);
nand \U$12346 ( \13016 , \13004 , \13005 , \13014 , \13015 );
nor \U$12347 ( \13017 , \12998 , \13016 );
nand \U$12348 ( \13018 , \12993 , \13017 );
buf \U$12349 ( \13019 , \13018 );
not \U$12350 ( \13020 , \13019 );
not \U$12351 ( \13021 , \13020 );
nand \U$12352 ( \13022 , \12606 , \13021 );
nand \U$12353 ( \13023 , \12978 , \13022 );
nand \U$12354 ( \13024 , \12921 , \13023 );
not \U$12355 ( \13025 , \13024 );
not \U$12356 ( \13026 , \12971 );
and \U$12357 ( \13027 , \12280 , \13026 );
or \U$12358 ( \13028 , \12433 , \13026 );
not \U$12359 ( \13029 , RIaaa1838_346);
not \U$12360 ( \13030 , \12339 );
or \U$12361 ( \13031 , \13029 , \13030 );
and \U$12362 ( \13032 , \12341 , \12306 , \12295 , \12325 );
nand \U$12363 ( \13033 , \13032 , RIaaa1928_348);
nand \U$12364 ( \13034 , \13031 , \13033 );
nand \U$12365 ( \13035 , \12365 , RIaaa1388_336);
nand \U$12366 ( \13036 , \12318 , \12305 , \12400 );
not \U$12367 ( \13037 , \13036 );
not \U$12368 ( \13038 , \7428 );
and \U$12369 ( \13039 , \13037 , \13038 );
and \U$12370 ( \13040 , \12402 , RIaaa19a0_349);
nor \U$12371 ( \13041 , \13039 , \13040 );
and \U$12372 ( \13042 , \12389 , RIaaa14f0_339);
not \U$12373 ( \13043 , RIaaa1310_335);
not \U$12374 ( \13044 , \12410 );
or \U$12375 ( \13045 , \13043 , \13044 );
nand \U$12376 ( \13046 , \11473 , RIaaa1220_333);
nand \U$12377 ( \13047 , \13045 , \13046 );
nor \U$12378 ( \13048 , \13042 , \13047 );
nand \U$12379 ( \13049 , \12418 , RIaaa15e0_341);
nand \U$12380 ( \13050 , \13035 , \13041 , \13048 , \13049 );
nor \U$12381 ( \13051 , \13034 , \13050 );
not \U$12382 ( \13052 , RIaaa1478_338);
not \U$12383 ( \13053 , \12453 );
or \U$12384 ( \13054 , \13052 , \13053 );
nand \U$12385 ( \13055 , \12455 , RIaaa16d0_343);
nand \U$12386 ( \13056 , \13054 , \13055 );
not \U$12387 ( \13057 , RIaaa1400_337);
not \U$12388 ( \13058 , \12356 );
or \U$12389 ( \13059 , \13057 , \13058 );
nand \U$12390 ( \13060 , \12532 , RIaaa1568_340);
nand \U$12391 ( \13061 , \13059 , \13060 );
nor \U$12392 ( \13062 , \13056 , \13061 );
and \U$12393 ( \13063 , \12931 , RIaaa18b0_347);
and \U$12394 ( \13064 , \12335 , RIaaa17c0_345);
nor \U$12395 ( \13065 , \13063 , \13064 );
and \U$12396 ( \13066 , \12446 , RIaaa1748_344);
and \U$12397 ( \13067 , \12327 , RIaaa1658_342);
nor \U$12398 ( \13068 , \13066 , \13067 );
nand \U$12399 ( \13069 , \13051 , \13062 , \13065 , \13068 );
buf \U$12400 ( \13070 , \13069 );
not \U$12401 ( \13071 , \13070 );
not \U$12402 ( \13072 , \13071 );
and \U$12403 ( \13073 , \13072 , \12495 );
not \U$12404 ( \13074 , \13072 );
and \U$12405 ( \13075 , \13074 , \12436 );
or \U$12406 ( \13076 , \13073 , \13075 );
nand \U$12407 ( \13077 , \13028 , \13076 );
nor \U$12408 ( \13078 , \13027 , \13077 );
not \U$12409 ( \13079 , \12581 );
not \U$12410 ( \13080 , \12589 );
nor \U$12411 ( \13081 , \13079 , \13080 );
not \U$12412 ( \13082 , \13081 );
not \U$12413 ( \13083 , RIaaa1ec8_360);
nor \U$12414 ( \13084 , \13083 , \12797 );
not \U$12415 ( \13085 , RIaaa1a90_351);
not \U$12416 ( \13086 , \12952 );
or \U$12417 ( \13087 , \13085 , \13086 );
nand \U$12418 ( \13088 , \12402 , RIaaa2198_366);
nand \U$12419 ( \13089 , \13087 , \13088 );
nor \U$12420 ( \13090 , \13084 , \13089 );
nand \U$12421 ( \13091 , \12339 , RIaaa2030_363);
nand \U$12422 ( \13092 , \12380 , RIaaa2120_365);
nand \U$12423 ( \13093 , \12418 , RIaaa1dd8_358);
nand \U$12424 ( \13094 , \12613 , RIaaa1ce8_356);
and \U$12425 ( \13095 , \12410 , RIaaa1b08_352);
nand \U$12426 ( \13096 , \11473 , RIaaa1a18_350);
not \U$12427 ( \13097 , \13096 );
nor \U$12428 ( \13098 , \13095 , \13097 );
and \U$12429 ( \13099 , \13093 , \13094 , \13098 );
nand \U$12430 ( \13100 , \13090 , \13091 , \13092 , \13099 );
not \U$12431 ( \13101 , \12448 );
not \U$12432 ( \13102 , RIaaa1fb8_362);
not \U$12433 ( \13103 , \13102 );
and \U$12434 ( \13104 , \13101 , \13103 );
not \U$12435 ( \13105 , RIaaa20a8_364);
nor \U$12436 ( \13106 , \12374 , \13105 );
nor \U$12437 ( \13107 , \13104 , \13106 );
not \U$12438 ( \13108 , \12439 );
not \U$12439 ( \13109 , \7181 );
and \U$12440 ( \13110 , \13108 , \13109 );
and \U$12441 ( \13111 , \12351 , RIaaa1f40_361);
nor \U$12442 ( \13112 , \13110 , \13111 );
and \U$12443 ( \13113 , \12453 , RIaaa1c70_355);
and \U$12444 ( \13114 , \12365 , RIaaa1b80_353);
nor \U$12445 ( \13115 , \13113 , \13114 );
and \U$12446 ( \13116 , \12356 , RIaaa1bf8_354);
and \U$12447 ( \13117 , \12360 , RIaaa1d60_357);
nor \U$12448 ( \13118 , \13116 , \13117 );
nand \U$12449 ( \13119 , \13107 , \13112 , \13115 , \13118 );
nor \U$12450 ( \13120 , \13100 , \13119 );
buf \U$12451 ( \13121 , \13120 );
buf \U$12452 ( \13122 , \13121 );
not \U$12453 ( \13123 , \13122 );
or \U$12454 ( \13124 , \13082 , \13123 );
nand \U$12455 ( \13125 , \12581 , \12583 );
buf \U$12456 ( \13126 , \13125 );
or \U$12457 ( \13127 , \13126 , \13122 );
nand \U$12458 ( \13128 , \13124 , \13127 );
nor \U$12459 ( \13129 , \12597 , \13072 );
nor \U$12460 ( \13130 , \13128 , \13129 );
nand \U$12461 ( \13131 , \12585 , \13072 );
nand \U$12462 ( \13132 , \13130 , \13131 );
not \U$12463 ( \13133 , \13132 );
not \U$12464 ( \13134 , \12423 );
buf \U$12465 ( \13135 , \12755 );
not \U$12466 ( \13136 , \13135 );
not \U$12467 ( \13137 , \12740 );
not \U$12468 ( \13138 , \12718 );
nand \U$12469 ( \13139 , \13138 , \12746 );
not \U$12470 ( \13140 , \13139 );
and \U$12471 ( \13141 , \13137 , \13140 );
and \U$12472 ( \13142 , \12740 , \13139 );
nor \U$12473 ( \13143 , \13141 , \13142 );
not \U$12474 ( \13144 , \13143 );
not \U$12475 ( \13145 , \13144 );
and \U$12476 ( \13146 , \13136 , \13145 );
not \U$12477 ( \13147 , \13143 );
and \U$12478 ( \13148 , \13135 , \13147 );
nor \U$12479 ( \13149 , \13146 , \13148 );
not \U$12480 ( \13150 , \13143 );
not \U$12481 ( \13151 , \12873 );
or \U$12482 ( \13152 , \13150 , \13151 );
not \U$12483 ( \13153 , \13143 );
nand \U$12484 ( \13154 , \13153 , \12872 );
nand \U$12485 ( \13155 , \13152 , \13154 );
nand \U$12486 ( \13156 , \13149 , \13155 );
buf \U$12487 ( \13157 , \12756 );
not \U$12488 ( \13158 , \13157 );
nor \U$12489 ( \13159 , \13156 , \13158 );
buf \U$12490 ( \13160 , \13159 );
not \U$12491 ( \13161 , \13160 );
or \U$12492 ( \13162 , \13134 , \13161 );
buf \U$12493 ( \13163 , \13157 );
nor \U$12494 ( \13164 , \13156 , \13163 );
not \U$12495 ( \13165 , \13164 );
not \U$12496 ( \13166 , \13165 );
and \U$12497 ( \13167 , \13166 , \12424 );
nor \U$12498 ( \13168 , \13155 , \13157 );
buf \U$12499 ( \13169 , \13168 );
and \U$12500 ( \13170 , \12491 , \13169 );
not \U$12501 ( \13171 , \12491 );
nor \U$12502 ( \13172 , \13155 , \13158 );
buf \U$12503 ( \13173 , \13172 );
and \U$12504 ( \13174 , \13171 , \13173 );
or \U$12505 ( \13175 , \13170 , \13174 );
nor \U$12506 ( \13176 , \13167 , \13175 );
nand \U$12507 ( \13177 , \13162 , \13176 );
not \U$12508 ( \13178 , \13177 );
nand \U$12509 ( \13179 , \13133 , \13178 );
not \U$12510 ( \13180 , \12797 );
not \U$12511 ( \13181 , RIaaa0b90_319);
not \U$12512 ( \13182 , \13181 );
and \U$12513 ( \13183 , \13180 , \13182 );
and \U$12514 ( \13184 , \12356 , RIaaa0c80_321);
nor \U$12515 ( \13185 , \13183 , \13184 );
and \U$12516 ( \13186 , \12365 , RIaaa1040_329);
and \U$12517 ( \13187 , \12476 , RIaaa0a28_316);
nor \U$12518 ( \13188 , \13186 , \13187 );
nand \U$12519 ( \13189 , \13185 , \13188 );
not \U$12520 ( \13190 , RIaaa0cf8_322);
not \U$12521 ( \13191 , \12339 );
or \U$12522 ( \13192 , \13190 , \13191 );
nand \U$12523 ( \13193 , \12351 , RIaaa0de8_324);
nand \U$12524 ( \13194 , \13192 , \13193 );
nor \U$12525 ( \13195 , \13189 , \13194 );
not \U$12526 ( \13196 , RIaaa0e60_325);
not \U$12527 ( \13197 , \12449 );
or \U$12528 ( \13198 , \13196 , \13197 );
nand \U$12529 ( \13199 , \12931 , RIaaa0d70_323);
nand \U$12530 ( \13200 , \13198 , \13199 );
not \U$12531 ( \13201 , RIaaa0b18_318);
not \U$12532 ( \13202 , \12327 );
or \U$12533 ( \13203 , \13201 , \13202 );
nand \U$12534 ( \13204 , \12379 , RIaaa1130_331);
nand \U$12535 ( \13205 , \13203 , \13204 );
nor \U$12536 ( \13206 , \13200 , \13205 );
not \U$12537 ( \13207 , RIaaa0c08_320);
not \U$12538 ( \13208 , \12453 );
or \U$12539 ( \13209 , \13207 , \13208 );
nand \U$12540 ( \13210 , \12360 , RIaaa0ed8_326);
nand \U$12541 ( \13211 , \13209 , \13210 );
and \U$12542 ( \13212 , \12513 , RIaaa10b8_330);
not \U$12543 ( \13213 , RIaaa0f50_327);
nor \U$12544 ( \13214 , \13213 , \12396 );
nor \U$12545 ( \13215 , \13212 , \13214 );
and \U$12546 ( \13216 , \12418 , RIaaa0aa0_317);
not \U$12547 ( \13217 , RIaaa0fc8_328);
not \U$12548 ( \13218 , \12410 );
or \U$12549 ( \13219 , \13217 , \13218 );
nand \U$12550 ( \13220 , \11473 , RIaaa11a8_332);
nand \U$12551 ( \13221 , \13219 , \13220 );
nor \U$12552 ( \13222 , \13216 , \13221 );
nand \U$12553 ( \13223 , \13215 , \13222 );
nor \U$12554 ( \13224 , \13211 , \13223 );
nand \U$12555 ( \13225 , \13195 , \13206 , \13224 );
not \U$12556 ( \13226 , \13225 );
buf \U$12557 ( \13227 , \13226 );
not \U$12558 ( \13228 , \13227 );
not \U$12559 ( \13229 , \13228 );
not \U$12560 ( \13230 , \12778 );
not \U$12561 ( \13231 , \12665 );
and \U$12562 ( \13232 , \13230 , \13231 );
not \U$12563 ( \13233 , \13232 );
or \U$12564 ( \13234 , \13229 , \13233 );
buf \U$12565 ( \13235 , \12664 );
not \U$12566 ( \13236 , \13235 );
not \U$12567 ( \13237 , \12774 );
and \U$12568 ( \13238 , \13163 , \13237 );
nand \U$12569 ( \13239 , \13236 , \13238 );
not \U$12570 ( \13240 , \13239 );
not \U$12571 ( \13241 , \13227 );
not \U$12572 ( \13242 , \13241 );
and \U$12573 ( \13243 , \13240 , \13242 );
not \U$12574 ( \13244 , \12845 );
not \U$12575 ( \13245 , \13244 );
and \U$12576 ( \13246 , \12787 , \13245 );
nor \U$12577 ( \13247 , \13243 , \13246 );
nand \U$12578 ( \13248 , \13234 , \13247 );
buf \U$12579 ( \13249 , \13248 );
and \U$12580 ( \13250 , \13179 , \13249 );
nor \U$12581 ( \13251 , \13133 , \13178 );
nor \U$12582 ( \13252 , \13250 , \13251 );
xor \U$12583 ( \13253 , \13078 , \13252 );
not \U$12584 ( \13254 , \12907 );
buf \U$12585 ( \13255 , \13254 );
not \U$12586 ( \13256 , \13255 );
not \U$12587 ( \13257 , \13256 );
not \U$12588 ( \13258 , \12894 );
or \U$12589 ( \13259 , \13257 , \13258 );
not \U$12590 ( \13260 , \12902 );
nand \U$12591 ( \13261 , \13259 , \13260 );
not \U$12592 ( \13262 , \12490 );
not \U$12593 ( \13263 , \13160 );
or \U$12594 ( \13264 , \13262 , \13263 );
nor \U$12595 ( \13265 , \13156 , \13163 );
not \U$12596 ( \13266 , \13265 );
not \U$12597 ( \13267 , \13266 );
and \U$12598 ( \13268 , \13267 , \12491 );
buf \U$12599 ( \13269 , \13172 );
and \U$12600 ( \13270 , \12545 , \13269 );
not \U$12601 ( \13271 , \12545 );
not \U$12602 ( \13272 , \13169 );
not \U$12603 ( \13273 , \13272 );
and \U$12604 ( \13274 , \13271 , \13273 );
or \U$12605 ( \13275 , \13270 , \13274 );
nor \U$12606 ( \13276 , \13268 , \13275 );
nand \U$12607 ( \13277 , \13264 , \13276 );
xor \U$12608 ( \13278 , \13261 , \13277 );
not \U$12609 ( \13279 , \13122 );
nor \U$12610 ( \13280 , \12598 , \13279 );
not \U$12611 ( \13281 , \13280 );
nand \U$12612 ( \13282 , \12585 , \13279 );
not \U$12613 ( \13283 , \13241 );
and \U$12614 ( \13284 , \13283 , \12601 );
not \U$12615 ( \13285 , \13283 );
not \U$12616 ( \13286 , \13125 );
and \U$12617 ( \13287 , \13285 , \13286 );
nor \U$12618 ( \13288 , \13284 , \13287 );
nand \U$12619 ( \13289 , \13281 , \13282 , \13288 );
xnor \U$12620 ( \13290 , \13278 , \13289 );
xor \U$12621 ( \13291 , \13253 , \13290 );
not \U$12622 ( \13292 , \13291 );
or \U$12623 ( \13293 , \13025 , \13292 );
not \U$12624 ( \13294 , \13023 );
nand \U$12625 ( \13295 , \13294 , \12920 );
nand \U$12626 ( \13296 , \13293 , \13295 );
not \U$12627 ( \13297 , \13296 );
not \U$12628 ( \13298 , \13169 );
buf \U$12629 ( \13299 , \13156 );
nand \U$12630 ( \13300 , \13298 , \13299 );
buf \U$12631 ( \13301 , \13155 );
not \U$12632 ( \13302 , \13163 );
and \U$12633 ( \13303 , \13301 , \13302 , \12545 );
and \U$12634 ( \13304 , \13163 , \12544 );
nor \U$12635 ( \13305 , \13303 , \13304 );
nand \U$12636 ( \13306 , \13300 , \13305 );
nand \U$12637 ( \13307 , \12606 , \12971 );
and \U$12638 ( \13308 , \13306 , \13307 );
or \U$12639 ( \13309 , \13277 , \13261 );
not \U$12640 ( \13310 , \13309 );
not \U$12641 ( \13311 , \13289 );
or \U$12642 ( \13312 , \13310 , \13311 );
nand \U$12643 ( \13313 , \13277 , \13261 );
nand \U$12644 ( \13314 , \13312 , \13313 );
xnor \U$12645 ( \13315 , \13308 , \13314 );
not \U$12646 ( \13316 , \13315 );
and \U$12647 ( \13317 , \12432 , \13072 );
and \U$12648 ( \13318 , \13122 , \12436 );
not \U$12649 ( \13319 , \13122 );
and \U$12650 ( \13320 , \13319 , \12495 );
nor \U$12651 ( \13321 , \13318 , \13320 );
nor \U$12652 ( \13322 , \13317 , \13321 );
nand \U$12653 ( \13323 , \12279 , \13071 );
nand \U$12654 ( \13324 , \13322 , \13323 );
not \U$12655 ( \13325 , \12849 );
nand \U$12656 ( \13326 , \13325 , \12915 );
xor \U$12657 ( \13327 , \13324 , \13326 );
buf \U$12658 ( \13328 , \13286 );
not \U$12659 ( \13329 , \13328 );
or \U$12660 ( \13330 , \13329 , \12658 );
nand \U$12661 ( \13331 , \12600 , \12658 );
nand \U$12662 ( \13332 , \13330 , \13331 );
nor \U$12663 ( \13333 , \12598 , \13241 );
nor \U$12664 ( \13334 , \13332 , \13333 );
nand \U$12665 ( \13335 , \12585 , \13241 );
nand \U$12666 ( \13336 , \13334 , \13335 );
not \U$12667 ( \13337 , \13336 );
not \U$12668 ( \13338 , \12779 );
and \U$12669 ( \13339 , \13338 , \12844 );
not \U$12670 ( \13340 , \13339 );
not \U$12671 ( \13341 , \13340 );
not \U$12672 ( \13342 , \12425 );
and \U$12673 ( \13343 , \13341 , \13342 );
not \U$12674 ( \13344 , \12425 );
nand \U$12675 ( \13345 , \13236 , \13238 );
not \U$12676 ( \13346 , \13345 );
not \U$12677 ( \13347 , \13346 );
or \U$12678 ( \13348 , \13344 , \13347 );
and \U$12679 ( \13349 , \12491 , \12770 );
not \U$12680 ( \13350 , \12491 );
not \U$12681 ( \13351 , \12846 );
and \U$12682 ( \13352 , \13350 , \13351 );
nor \U$12683 ( \13353 , \13349 , \13352 );
nand \U$12684 ( \13354 , \13348 , \13353 );
nor \U$12685 ( \13355 , \13343 , \13354 );
not \U$12686 ( \13356 , \13355 );
and \U$12687 ( \13357 , \13337 , \13356 );
and \U$12688 ( \13358 , \13336 , \13355 );
nor \U$12689 ( \13359 , \13357 , \13358 );
xnor \U$12690 ( \13360 , \13327 , \13359 );
not \U$12691 ( \13361 , \13360 );
xor \U$12692 ( \13362 , \13078 , \13252 );
and \U$12693 ( \13363 , \13362 , \13290 );
and \U$12694 ( \13364 , \13078 , \13252 );
or \U$12695 ( \13365 , \13363 , \13364 );
not \U$12696 ( \13366 , \13365 );
and \U$12697 ( \13367 , \13361 , \13366 );
and \U$12698 ( \13368 , \13360 , \13365 );
nor \U$12699 ( \13369 , \13367 , \13368 );
not \U$12700 ( \13370 , \13369 );
or \U$12701 ( \13371 , \13316 , \13370 );
or \U$12702 ( \13372 , \13315 , \13369 );
nand \U$12703 ( \13373 , \13371 , \13372 );
not \U$12704 ( \13374 , \13373 );
or \U$12705 ( \13375 , \13297 , \13374 );
not \U$12706 ( \13376 , \13369 );
nand \U$12707 ( \13377 , \13376 , \13315 );
nand \U$12708 ( \13378 , \13375 , \13377 );
not \U$12709 ( \13379 , \13365 );
not \U$12710 ( \13380 , \13326 );
not \U$12711 ( \13381 , \13355 );
buf \U$12712 ( \13382 , \13324 );
xor \U$12713 ( \13383 , \13381 , \13382 );
xor \U$12714 ( \13384 , \13383 , \13336 );
nand \U$12715 ( \13385 , \13380 , \13384 );
not \U$12716 ( \13386 , \13385 );
or \U$12717 ( \13387 , \13379 , \13386 );
not \U$12718 ( \13388 , \13384 );
nand \U$12719 ( \13389 , \13388 , \13326 );
nand \U$12720 ( \13390 , \13387 , \13389 );
not \U$12721 ( \13391 , \13390 );
not \U$12722 ( \13392 , \12433 );
not \U$12723 ( \13393 , \13122 );
and \U$12724 ( \13394 , \13392 , \13393 );
not \U$12725 ( \13395 , \12496 );
or \U$12726 ( \13396 , \13395 , \13283 );
or \U$12727 ( \13397 , \12437 , \13241 );
nand \U$12728 ( \13398 , \13396 , \13397 );
nor \U$12729 ( \13399 , \13394 , \13398 );
nand \U$12730 ( \13400 , \12280 , \13122 );
nand \U$12731 ( \13401 , \13399 , \13400 );
not \U$12732 ( \13402 , \13072 );
not \U$12733 ( \13403 , \12606 );
or \U$12734 ( \13404 , \13402 , \13403 );
nand \U$12735 ( \13405 , \13404 , \13306 );
nor \U$12736 ( \13406 , \13401 , \13405 );
not \U$12737 ( \13407 , \13406 );
nand \U$12738 ( \13408 , \13401 , \13405 );
nand \U$12739 ( \13409 , \13407 , \13408 );
not \U$12740 ( \13410 , \13306 );
not \U$12741 ( \13411 , \13314 );
or \U$12742 ( \13412 , \13410 , \13411 );
nand \U$12743 ( \13413 , \13412 , \13307 );
not \U$12744 ( \13414 , \13413 );
xor \U$12745 ( \13415 , \13409 , \13414 );
not \U$12746 ( \13416 , \13301 );
not \U$12747 ( \13417 , \13299 );
or \U$12748 ( \13418 , \13416 , \13417 );
nand \U$12749 ( \13419 , \13418 , \13302 );
not \U$12750 ( \13420 , \12497 );
not \U$12751 ( \13421 , \13340 );
not \U$12752 ( \13422 , \13421 );
or \U$12753 ( \13423 , \13420 , \13422 );
not \U$12754 ( \13424 , \13345 );
not \U$12755 ( \13425 , \12497 );
and \U$12756 ( \13426 , \13424 , \13425 );
and \U$12757 ( \13427 , \12545 , \12846 );
not \U$12758 ( \13428 , \12545 );
not \U$12759 ( \13429 , \12844 );
nand \U$12760 ( \13430 , \13429 , \12845 );
buf \U$12761 ( \13431 , \13430 );
and \U$12762 ( \13432 , \13428 , \13431 );
nor \U$12763 ( \13433 , \13427 , \13432 );
nor \U$12764 ( \13434 , \13426 , \13433 );
nand \U$12765 ( \13435 , \13423 , \13434 );
xor \U$12766 ( \13436 , \13419 , \13435 );
not \U$12767 ( \13437 , \13436 );
not \U$12768 ( \13438 , \12659 );
not \U$12769 ( \13439 , \12585 );
or \U$12770 ( \13440 , \13438 , \13439 );
not \U$12771 ( \13441 , \12598 );
not \U$12772 ( \13442 , \12659 );
and \U$12773 ( \13443 , \13441 , \13442 );
and \U$12774 ( \13444 , \12425 , \12601 );
not \U$12775 ( \13445 , \12425 );
and \U$12776 ( \13446 , \13445 , \13286 );
or \U$12777 ( \13447 , \13444 , \13446 );
nor \U$12778 ( \13448 , \13443 , \13447 );
nand \U$12779 ( \13449 , \13440 , \13448 );
not \U$12780 ( \13450 , \13449 );
not \U$12781 ( \13451 , \13450 );
or \U$12782 ( \13452 , \13437 , \13451 );
or \U$12783 ( \13453 , \13450 , \13436 );
nand \U$12784 ( \13454 , \13452 , \13453 );
not \U$12785 ( \13455 , \13336 );
not \U$12786 ( \13456 , \13381 );
or \U$12787 ( \13457 , \13455 , \13456 );
not \U$12788 ( \13458 , \13359 );
nand \U$12789 ( \13459 , \13458 , \13382 );
nand \U$12790 ( \13460 , \13457 , \13459 );
xor \U$12791 ( \13461 , \13454 , \13460 );
xnor \U$12792 ( \13462 , \13415 , \13461 );
not \U$12793 ( \13463 , \13462 );
or \U$12794 ( \13464 , \13391 , \13463 );
or \U$12795 ( \13465 , \13390 , \13462 );
nand \U$12796 ( \13466 , \13464 , \13465 );
or \U$12797 ( \13467 , \13378 , \13466 );
not \U$12798 ( \13468 , \13467 );
not \U$12799 ( \13469 , \11808 );
buf \U$12800 ( \13470 , \11806 );
not \U$12801 ( \13471 , \13470 );
not \U$12802 ( \13472 , \13471 );
or \U$12803 ( \13473 , \13469 , \13472 );
not \U$12804 ( \13474 , \13470 );
or \U$12805 ( \13475 , \13474 , \11808 );
nand \U$12806 ( \13476 , \13473 , \13475 );
buf \U$12807 ( \13477 , \11912 );
not \U$12808 ( \13478 , \13477 );
and \U$12809 ( \13479 , \13476 , \13478 );
not \U$12810 ( \13480 , \13476 );
and \U$12811 ( \13481 , \13480 , \13477 );
nor \U$12812 ( \13482 , \13479 , \13481 );
not \U$12813 ( \13483 , \13482 );
not \U$12814 ( \13484 , \13483 );
not \U$12815 ( \13485 , \13471 );
not \U$12816 ( \13486 , \11808 );
or \U$12817 ( \13487 , \13485 , \13486 );
nand \U$12818 ( \13488 , \13487 , \11913 );
not \U$12819 ( \13489 , \11916 );
and \U$12820 ( \13490 , \13489 , \11917 );
not \U$12821 ( \13491 , \13489 );
and \U$12822 ( \13492 , \13491 , \11814 );
nor \U$12823 ( \13493 , \13490 , \13492 );
not \U$12824 ( \13494 , \13493 );
and \U$12825 ( \13495 , \13488 , \13494 );
not \U$12826 ( \13496 , \13488 );
and \U$12827 ( \13497 , \13496 , \13493 );
nor \U$12828 ( \13498 , \13495 , \13497 );
not \U$12829 ( \13499 , \13498 );
not \U$12830 ( \13500 , \13499 );
or \U$12831 ( \13501 , \13484 , \13500 );
nand \U$12832 ( \13502 , \13498 , \13482 );
nand \U$12833 ( \13503 , \13501 , \13502 );
buf \U$12834 ( \13504 , \13503 );
not \U$12835 ( \13505 , \12882 );
not \U$12836 ( \13506 , \13498 );
not \U$12837 ( \13507 , \13506 );
and \U$12838 ( \13508 , \13505 , \13507 );
and \U$12839 ( \13509 , \12890 , \13506 );
nor \U$12840 ( \13510 , \13508 , \13509 );
nand \U$12841 ( \13511 , \13504 , \13510 );
buf \U$12842 ( \13512 , \13511 );
buf \U$12843 ( \13513 , \13504 );
nand \U$12844 ( \13514 , \13512 , \13513 );
buf \U$12845 ( \13515 , \12890 );
not \U$12846 ( \13516 , \13515 );
nand \U$12847 ( \13517 , \13514 , \13516 );
and \U$12848 ( \13518 , \12904 , \12491 );
nand \U$12849 ( \13519 , \13254 , \12902 );
buf \U$12850 ( \13520 , \13519 );
or \U$12851 ( \13521 , \13520 , \12544 );
nand \U$12852 ( \13522 , \12911 , \12544 );
nand \U$12853 ( \13523 , \13521 , \13522 );
nor \U$12854 ( \13524 , \13518 , \13523 );
buf \U$12855 ( \13525 , \12896 );
nand \U$12856 ( \13526 , \13525 , \12490 );
nand \U$12857 ( \13527 , \13524 , \13526 );
xor \U$12858 ( \13528 , \13517 , \13527 );
not \U$12859 ( \13529 , \12657 );
not \U$12860 ( \13530 , \13160 );
or \U$12861 ( \13531 , \13529 , \13530 );
buf \U$12862 ( \13532 , \13266 );
not \U$12863 ( \13533 , \13532 );
and \U$12864 ( \13534 , \13533 , \12658 );
and \U$12865 ( \13535 , \12423 , \13269 );
not \U$12866 ( \13536 , \12423 );
and \U$12867 ( \13537 , \13536 , \13169 );
or \U$12868 ( \13538 , \13535 , \13537 );
nor \U$12869 ( \13539 , \13534 , \13538 );
nand \U$12870 ( \13540 , \13531 , \13539 );
not \U$12871 ( \13541 , \13540 );
and \U$12872 ( \13542 , \13528 , \13541 );
not \U$12873 ( \13543 , \13528 );
and \U$12874 ( \13544 , \13543 , \13540 );
nor \U$12875 ( \13545 , \13542 , \13544 );
not \U$12876 ( \13546 , \13545 );
not \U$12877 ( \13547 , \12839 );
not \U$12878 ( \13548 , \12585 );
or \U$12879 ( \13549 , \13547 , \13548 );
not \U$12880 ( \13550 , \13081 );
not \U$12881 ( \13551 , \13026 );
or \U$12882 ( \13552 , \13550 , \13551 );
or \U$12883 ( \13553 , \13126 , \13026 );
nand \U$12884 ( \13554 , \13552 , \13553 );
nor \U$12885 ( \13555 , \12597 , \12839 );
nor \U$12886 ( \13556 , \13554 , \13555 );
nand \U$12887 ( \13557 , \13549 , \13556 );
nor \U$12888 ( \13558 , \13511 , \13515 );
buf \U$12889 ( \13559 , \13558 );
buf \U$12890 ( \13560 , \12488 );
and \U$12891 ( \13561 , \13559 , \13560 );
not \U$12892 ( \13562 , \12890 );
not \U$12893 ( \13563 , \13562 );
not \U$12894 ( \13564 , \13503 );
nand \U$12895 ( \13565 , \13563 , \13564 );
buf \U$12896 ( \13566 , \13565 );
not \U$12897 ( \13567 , \12543 );
or \U$12898 ( \13568 , \13566 , \13567 );
not \U$12899 ( \13569 , \12890 );
not \U$12900 ( \13570 , \13503 );
nand \U$12901 ( \13571 , \13569 , \13570 );
buf \U$12902 ( \13572 , \13571 );
not \U$12903 ( \13573 , \13572 );
nand \U$12904 ( \13574 , \13573 , \13567 );
nand \U$12905 ( \13575 , \13568 , \13574 );
nor \U$12906 ( \13576 , \13561 , \13575 );
nor \U$12907 ( \13577 , \13511 , \13516 );
buf \U$12908 ( \13578 , \13577 );
nand \U$12909 ( \13579 , \13578 , \12490 );
nand \U$12910 ( \13580 , \13576 , \13579 );
buf \U$12911 ( \13581 , \13483 );
not \U$12912 ( \13582 , \13581 );
buf \U$12913 ( \13583 , \13582 );
not \U$12914 ( \13584 , \13583 );
nor \U$12915 ( \13585 , \13580 , \13584 );
not \U$12916 ( \13586 , \13585 );
or \U$12917 ( \13587 , \13557 , \13586 );
not \U$12918 ( \13588 , \13072 );
not \U$12919 ( \13589 , \13339 );
or \U$12920 ( \13590 , \13588 , \13589 );
and \U$12921 ( \13591 , \13346 , \13071 );
or \U$12922 ( \13592 , \12846 , \13122 );
nand \U$12923 ( \13593 , \12770 , \13122 );
nand \U$12924 ( \13594 , \13592 , \13593 );
nor \U$12925 ( \13595 , \13591 , \13594 );
nand \U$12926 ( \13596 , \13590 , \13595 );
nand \U$12927 ( \13597 , \13587 , \13596 );
nand \U$12928 ( \13598 , \13557 , \13586 );
nand \U$12929 ( \13599 , \13597 , \13598 );
not \U$12930 ( \13600 , \13599 );
not \U$12931 ( \13601 , \13600 );
or \U$12932 ( \13602 , \13546 , \13601 );
not \U$12933 ( \13603 , \13279 );
not \U$12934 ( \13604 , \13339 );
or \U$12935 ( \13605 , \13603 , \13604 );
not \U$12936 ( \13606 , \13345 );
not \U$12937 ( \13607 , \13279 );
and \U$12938 ( \13608 , \13606 , \13607 );
and \U$12939 ( \13609 , \13283 , \13431 );
not \U$12940 ( \13610 , \13283 );
and \U$12941 ( \13611 , \13610 , \12846 );
nor \U$12942 ( \13612 , \13609 , \13611 );
nor \U$12943 ( \13613 , \13608 , \13612 );
nand \U$12944 ( \13614 , \13605 , \13613 );
nand \U$12945 ( \13615 , \13512 , \13572 );
nand \U$12946 ( \13616 , \13516 , \12545 , \13513 );
nand \U$12947 ( \13617 , \13515 , \12544 );
and \U$12948 ( \13618 , \13615 , \13616 , \13617 );
nor \U$12949 ( \13619 , \13614 , \13618 );
not \U$12950 ( \13620 , \13619 );
nand \U$12951 ( \13621 , \13614 , \13618 );
nand \U$12952 ( \13622 , \13620 , \13621 );
not \U$12953 ( \13623 , \13622 );
not \U$12954 ( \13624 , \12971 );
not \U$12955 ( \13625 , \12585 );
or \U$12956 ( \13626 , \13624 , \13625 );
not \U$12957 ( \13627 , \13286 );
or \U$12958 ( \13628 , \13627 , \13071 );
nand \U$12959 ( \13629 , \12601 , \13071 );
nand \U$12960 ( \13630 , \13628 , \13629 );
nor \U$12961 ( \13631 , \12598 , \12971 );
nor \U$12962 ( \13632 , \13630 , \13631 );
nand \U$12963 ( \13633 , \13626 , \13632 );
not \U$12964 ( \13634 , \13633 );
and \U$12965 ( \13635 , \13623 , \13634 );
and \U$12966 ( \13636 , \13622 , \13633 );
nor \U$12967 ( \13637 , \13635 , \13636 );
not \U$12968 ( \13638 , \13637 );
nand \U$12969 ( \13639 , \13602 , \13638 );
not \U$12970 ( \13640 , \13545 );
nand \U$12971 ( \13641 , \13599 , \13640 );
nand \U$12972 ( \13642 , \13639 , \13641 );
nand \U$12973 ( \13643 , \12327 , RIaaa3818_414);
nand \U$12974 ( \13644 , \12449 , RIaaa3980_417);
nand \U$12975 ( \13645 , \12931 , RIaaa37a0_413);
nand \U$12976 ( \13646 , \12446 , RIaaa3908_416);
nand \U$12977 ( \13647 , \13643 , \13644 , \13645 , \13646 );
nand \U$12978 ( \13648 , \12344 , RIaaa3368_404);
nand \U$12979 ( \13649 , \12356 , RIaaa3278_402);
nand \U$12980 ( \13650 , \12365 , RIaaa35c0_409);
nand \U$12981 ( \13651 , \12360 , RIaaa33e0_405);
nand \U$12982 ( \13652 , \13648 , \13649 , \13650 , \13651 );
nor \U$12983 ( \13653 , \13647 , \13652 );
not \U$12984 ( \13654 , RIaaa3728_412);
not \U$12985 ( \13655 , \12339 );
or \U$12986 ( \13656 , \13654 , \13655 );
nand \U$12987 ( \13657 , \12379 , RIaaa3638_410);
nand \U$12988 ( \13658 , \13656 , \13657 );
and \U$12989 ( \13659 , \12418 , RIaaa3458_406);
and \U$12990 ( \13660 , \12402 , RIaaa36b0_411);
nor \U$12991 ( \13661 , \13659 , \13660 );
nand \U$12992 ( \13662 , \12384 , RIaaa3890_415);
and \U$12993 ( \13663 , \12476 , RIaaa32f0_403);
not \U$12994 ( \13664 , RIaaa3548_408);
not \U$12995 ( \13665 , \12410 );
or \U$12996 ( \13666 , \13664 , \13665 );
nand \U$12997 ( \13667 , \11473 , RIaaa3200_401);
nand \U$12998 ( \13668 , \13666 , \13667 );
nor \U$12999 ( \13669 , \13663 , \13668 );
nand \U$13000 ( \13670 , \12395 , RIaaa34d0_407);
nand \U$13001 ( \13671 , \13661 , \13662 , \13669 , \13670 );
nor \U$13002 ( \13672 , \13658 , \13671 );
nand \U$13003 ( \13673 , \13653 , \13672 );
not \U$13004 ( \13674 , \13673 );
buf \U$13005 ( \13675 , \13674 );
not \U$13006 ( \13676 , \13675 );
nand \U$13007 ( \13677 , \12605 , \13676 );
not \U$13008 ( \13678 , \13677 );
not \U$13009 ( \13679 , \12274 );
not \U$13010 ( \13680 , \13679 );
not \U$13011 ( \13681 , \13021 );
not \U$13012 ( \13682 , \12493 );
not \U$13013 ( \13683 , \13682 );
or \U$13014 ( \13684 , \13681 , \13683 );
or \U$13015 ( \13685 , \12494 , \13021 );
nand \U$13016 ( \13686 , \13684 , \13685 );
not \U$13017 ( \13687 , \13686 );
or \U$13018 ( \13688 , \13680 , \13687 );
nand \U$13019 ( \13689 , \12927 , \12677 );
nand \U$13020 ( \13690 , \13688 , \13689 );
not \U$13021 ( \13691 , \13690 );
not \U$13022 ( \13692 , \13691 );
or \U$13023 ( \13693 , \13678 , \13692 );
not \U$13024 ( \13694 , \13677 );
nand \U$13025 ( \13695 , \13694 , \13690 );
nand \U$13026 ( \13696 , \13693 , \13695 );
not \U$13027 ( \13697 , \13241 );
not \U$13028 ( \13698 , \13160 );
or \U$13029 ( \13699 , \13697 , \13698 );
and \U$13030 ( \13700 , \13267 , \13283 );
not \U$13031 ( \13701 , \13169 );
or \U$13032 ( \13702 , \13701 , \12657 );
not \U$13033 ( \13703 , \12656 );
buf \U$13034 ( \13704 , \13173 );
nand \U$13035 ( \13705 , \13703 , \13704 );
nand \U$13036 ( \13706 , \13702 , \13705 );
nor \U$13037 ( \13707 , \13700 , \13706 );
nand \U$13038 ( \13708 , \13699 , \13707 );
not \U$13039 ( \13709 , \13708 );
not \U$13040 ( \13710 , \13618 );
not \U$13041 ( \13711 , \12423 );
not \U$13042 ( \13712 , \13525 );
or \U$13043 ( \13713 , \13711 , \13712 );
not \U$13044 ( \13714 , \12903 );
and \U$13045 ( \13715 , \13714 , \12424 );
or \U$13046 ( \13716 , \13520 , \13560 );
buf \U$13047 ( \13717 , \12909 );
not \U$13048 ( \13718 , \13717 );
nand \U$13049 ( \13719 , \13718 , \13560 );
nand \U$13050 ( \13720 , \13716 , \13719 );
nor \U$13051 ( \13721 , \13715 , \13720 );
nand \U$13052 ( \13722 , \13713 , \13721 );
not \U$13053 ( \13723 , \13722 );
or \U$13054 ( \13724 , \13710 , \13723 );
or \U$13055 ( \13725 , \13722 , \13618 );
nand \U$13056 ( \13726 , \13724 , \13725 );
not \U$13057 ( \13727 , \13726 );
or \U$13058 ( \13728 , \13709 , \13727 );
not \U$13059 ( \13729 , \13618 );
nand \U$13060 ( \13730 , \13729 , \13722 );
nand \U$13061 ( \13731 , \13728 , \13730 );
not \U$13062 ( \13732 , \13731 );
xor \U$13063 ( \13733 , \13696 , \13732 );
not \U$13064 ( \13734 , \12841 );
nand \U$13065 ( \13735 , \12449 , RIaaa4790_447);
nand \U$13066 ( \13736 , \12327 , RIaaa4628_444);
nand \U$13067 ( \13737 , \12931 , RIaaa4880_449);
nand \U$13068 ( \13738 , \12446 , RIaaa4718_446);
nand \U$13069 ( \13739 , \13735 , \13736 , \13737 , \13738 );
nand \U$13070 ( \13740 , \12344 , RIaaa4448_440);
nand \U$13071 ( \13741 , \12356 , RIaaa43d0_439);
nand \U$13072 ( \13742 , \12360 , RIaaa4538_442);
nand \U$13073 ( \13743 , \12365 , RIaaa4358_438);
nand \U$13074 ( \13744 , \13740 , \13741 , \13742 , \13743 );
nor \U$13075 ( \13745 , \13739 , \13744 );
not \U$13076 ( \13746 , RIaaa4808_448);
not \U$13077 ( \13747 , \12339 );
or \U$13078 ( \13748 , \13746 , \13747 );
nand \U$13079 ( \13749 , \12379 , RIaaa48f8_450);
nand \U$13080 ( \13750 , \13748 , \13749 );
and \U$13081 ( \13751 , \12613 , RIaaa44c0_441);
not \U$13082 ( \13752 , RIaaa42e0_437);
not \U$13083 ( \13753 , \12410 );
or \U$13084 ( \13754 , \13752 , \13753 );
nand \U$13085 ( \13755 , \11473 , RIaaa41f0_435);
nand \U$13086 ( \13756 , \13754 , \13755 );
nor \U$13087 ( \13757 , \13751 , \13756 );
not \U$13088 ( \13758 , \12951 );
not \U$13089 ( \13759 , \13758 );
not \U$13090 ( \13760 , RIaaa4268_436);
not \U$13091 ( \13761 , \13760 );
and \U$13092 ( \13762 , \13759 , \13761 );
and \U$13093 ( \13763 , \13007 , RIaaa4970_451);
nor \U$13094 ( \13764 , \13762 , \13763 );
nand \U$13095 ( \13765 , \12384 , RIaaa46a0_445);
nand \U$13096 ( \13766 , \12469 , RIaaa45b0_443);
nand \U$13097 ( \13767 , \13757 , \13764 , \13765 , \13766 );
nor \U$13098 ( \13768 , \13750 , \13767 );
nand \U$13099 ( \13769 , \13745 , \13768 );
buf \U$13100 ( \13770 , \13769 );
not \U$13101 ( \13771 , \13770 );
nor \U$13102 ( \13772 , \13734 , \13771 );
not \U$13103 ( \13773 , \13772 );
not \U$13104 ( \13774 , \13773 );
not \U$13105 ( \13775 , \12422 );
not \U$13106 ( \13776 , \13775 );
not \U$13107 ( \13777 , \13776 );
not \U$13108 ( \13778 , \13578 );
or \U$13109 ( \13779 , \13777 , \13778 );
and \U$13110 ( \13780 , \13559 , \12424 );
not \U$13111 ( \13781 , \13571 );
not \U$13112 ( \13782 , \13781 );
not \U$13113 ( \13783 , \12488 );
or \U$13114 ( \13784 , \13782 , \13783 );
or \U$13115 ( \13785 , \13566 , \12489 );
nand \U$13116 ( \13786 , \13784 , \13785 );
nor \U$13117 ( \13787 , \13780 , \13786 );
nand \U$13118 ( \13788 , \13779 , \13787 );
not \U$13119 ( \13789 , \13581 );
not \U$13120 ( \13790 , RIaaa9560_613);
not \U$13121 ( \13791 , \11910 );
not \U$13122 ( \13792 , \13791 );
or \U$13123 ( \13793 , \13790 , \13792 );
nand \U$13124 ( \13794 , \13793 , \13477 );
not \U$13125 ( \13795 , \13794 );
nand \U$13126 ( \13796 , \13789 , \13795 );
not \U$13127 ( \13797 , \13796 );
not \U$13128 ( \13798 , \13797 );
not \U$13129 ( \13799 , \13798 );
not \U$13130 ( \13800 , \13799 );
not \U$13131 ( \13801 , \13567 );
or \U$13132 ( \13802 , \13800 , \13801 );
nand \U$13133 ( \13803 , \13582 , \13794 );
buf \U$13134 ( \13804 , \13803 );
nand \U$13135 ( \13805 , \13802 , \13804 );
nand \U$13136 ( \13806 , \13788 , \13805 );
not \U$13137 ( \13807 , \12656 );
not \U$13138 ( \13808 , \13714 );
or \U$13139 ( \13809 , \13807 , \13808 );
and \U$13140 ( \13810 , \12424 , \12911 );
not \U$13141 ( \13811 , \12424 );
not \U$13142 ( \13812 , \12877 );
not \U$13143 ( \13813 , \13812 );
nand \U$13144 ( \13814 , \13813 , \13254 );
not \U$13145 ( \13815 , \13814 );
and \U$13146 ( \13816 , \13811 , \13815 );
nor \U$13147 ( \13817 , \13810 , \13816 );
nand \U$13148 ( \13818 , \13809 , \13817 );
not \U$13149 ( \13819 , \13525 );
nor \U$13150 ( \13820 , \13819 , \12656 );
nor \U$13151 ( \13821 , \13818 , \13820 );
xor \U$13152 ( \13822 , \13806 , \13821 );
not \U$13153 ( \13823 , \13122 );
not \U$13154 ( \13824 , \13267 );
or \U$13155 ( \13825 , \13823 , \13824 );
and \U$13156 ( \13826 , \13273 , \13283 );
and \U$13157 ( \13827 , \13173 , \13241 );
nor \U$13158 ( \13828 , \13826 , \13827 );
nand \U$13159 ( \13829 , \13825 , \13828 );
not \U$13160 ( \13830 , \13160 );
nor \U$13161 ( \13831 , \13830 , \13122 );
nor \U$13162 ( \13832 , \13829 , \13831 );
and \U$13163 ( \13833 , \13822 , \13832 );
and \U$13164 ( \13834 , \13806 , \13821 );
or \U$13165 ( \13835 , \13833 , \13834 );
not \U$13166 ( \13836 , \13835 );
or \U$13167 ( \13837 , \13774 , \13836 );
not \U$13168 ( \13838 , \13676 );
not \U$13169 ( \13839 , \12430 );
or \U$13170 ( \13840 , \13838 , \13839 );
not \U$13171 ( \13841 , \13673 );
not \U$13172 ( \13842 , \13841 );
or \U$13173 ( \13843 , \12430 , \13842 );
nand \U$13174 ( \13844 , \13840 , \13843 );
not \U$13175 ( \13845 , \13844 );
not \U$13176 ( \13846 , \12275 );
or \U$13177 ( \13847 , \13845 , \13846 );
nand \U$13178 ( \13848 , \13686 , \12677 );
nand \U$13179 ( \13849 , \13847 , \13848 );
nand \U$13180 ( \13850 , \13837 , \13849 );
xnor \U$13181 ( \13851 , \13733 , \13850 );
xor \U$13182 ( \13852 , \13586 , \13596 );
xnor \U$13183 ( \13853 , \13852 , \13557 );
not \U$13184 ( \13854 , \13853 );
not \U$13185 ( \13855 , \12971 );
not \U$13186 ( \13856 , \13235 );
or \U$13187 ( \13857 , \13855 , \13856 );
or \U$13188 ( \13858 , \13231 , \12971 );
nand \U$13189 ( \13859 , \13857 , \13858 );
not \U$13190 ( \13860 , \13859 );
not \U$13191 ( \13861 , \12779 );
not \U$13192 ( \13862 , \13861 );
or \U$13193 ( \13863 , \13860 , \13862 );
not \U$13194 ( \13864 , \13072 );
not \U$13195 ( \13865 , \12664 );
or \U$13196 ( \13866 , \13864 , \13865 );
or \U$13197 ( \13867 , \13235 , \13072 );
nand \U$13198 ( \13868 , \13866 , \13867 );
buf \U$13199 ( \13869 , \12845 );
nand \U$13200 ( \13870 , \13868 , \13869 );
nand \U$13201 ( \13871 , \13863 , \13870 );
not \U$13202 ( \13872 , \13871 );
and \U$13203 ( \13873 , \13580 , \13584 );
nor \U$13204 ( \13874 , \13873 , \13585 );
not \U$13205 ( \13875 , \13874 );
or \U$13206 ( \13876 , \13872 , \13875 );
or \U$13207 ( \13877 , \13871 , \13874 );
nand \U$13208 ( \13878 , \13876 , \13877 );
not \U$13209 ( \13879 , \13878 );
not \U$13210 ( \13880 , \12838 );
not \U$13211 ( \13881 , \12601 );
or \U$13212 ( \13882 , \13880 , \13881 );
and \U$13213 ( \13883 , \13328 , \12839 );
buf \U$13214 ( \13884 , \12582 );
not \U$13215 ( \13885 , \13018 );
not \U$13216 ( \13886 , \13885 );
not \U$13217 ( \13887 , \13886 );
not \U$13218 ( \13888 , \12668 );
or \U$13219 ( \13889 , \13887 , \13888 );
buf \U$13220 ( \13890 , \12564 );
not \U$13221 ( \13891 , \13890 );
or \U$13222 ( \13892 , \13891 , \13021 );
nand \U$13223 ( \13893 , \13889 , \13892 );
and \U$13224 ( \13894 , \13884 , \13893 );
nor \U$13225 ( \13895 , \13883 , \13894 );
nand \U$13226 ( \13896 , \13882 , \13895 );
not \U$13227 ( \13897 , \13896 );
or \U$13228 ( \13898 , \13879 , \13897 );
not \U$13229 ( \13899 , \13874 );
nand \U$13230 ( \13900 , \13899 , \13871 );
nand \U$13231 ( \13901 , \13898 , \13900 );
nand \U$13232 ( \13902 , \13851 , \13854 , \13901 );
not \U$13233 ( \13903 , \13901 );
nand \U$13234 ( \13904 , \13853 , \13903 );
not \U$13235 ( \13905 , \13708 );
and \U$13236 ( \13906 , \13726 , \13905 );
not \U$13237 ( \13907 , \13726 );
and \U$13238 ( \13908 , \13907 , \13708 );
nor \U$13239 ( \13909 , \13906 , \13908 );
not \U$13240 ( \13910 , \13909 );
nand \U$13241 ( \13911 , \13851 , \13904 , \13910 );
not \U$13242 ( \13912 , \13850 );
xor \U$13243 ( \13913 , \13732 , \13696 );
nand \U$13244 ( \13914 , \13912 , \13913 );
nand \U$13245 ( \13915 , \13902 , \13911 , \13914 );
xor \U$13246 ( \13916 , \13642 , \13915 );
not \U$13247 ( \13917 , \13619 );
not \U$13248 ( \13918 , \13917 );
not \U$13249 ( \13919 , \13633 );
or \U$13250 ( \13920 , \13918 , \13919 );
nand \U$13251 ( \13921 , \13920 , \13621 );
not \U$13252 ( \13922 , \13921 );
not \U$13253 ( \13923 , \13922 );
and \U$13254 ( \13924 , \13528 , \13540 );
and \U$13255 ( \13925 , \13517 , \13527 );
nor \U$13256 ( \13926 , \13924 , \13925 );
and \U$13257 ( \13927 , \13248 , \13177 );
not \U$13258 ( \13928 , \13248 );
and \U$13259 ( \13929 , \13928 , \13178 );
nor \U$13260 ( \13930 , \13927 , \13929 );
and \U$13261 ( \13931 , \13930 , \13132 );
not \U$13262 ( \13932 , \13930 );
and \U$13263 ( \13933 , \13932 , \13133 );
nor \U$13264 ( \13934 , \13931 , \13933 );
xnor \U$13265 ( \13935 , \13926 , \13934 );
buf \U$13266 ( \13936 , \13935 );
not \U$13267 ( \13937 , \13936 );
or \U$13268 ( \13938 , \13923 , \13937 );
or \U$13269 ( \13939 , \13936 , \13922 );
nand \U$13270 ( \13940 , \13938 , \13939 );
not \U$13271 ( \13941 , \13940 );
nand \U$13272 ( \13942 , \12916 , \13022 );
xor \U$13273 ( \13943 , \13942 , \12976 );
not \U$13274 ( \13944 , \13677 );
not \U$13275 ( \13945 , \13732 );
or \U$13276 ( \13946 , \13944 , \13945 );
nand \U$13277 ( \13947 , \13946 , \13690 );
xnor \U$13278 ( \13948 , \13943 , \13947 );
not \U$13279 ( \13949 , \13948 );
and \U$13280 ( \13950 , \13941 , \13949 );
and \U$13281 ( \13951 , \13940 , \13948 );
nor \U$13282 ( \13952 , \13950 , \13951 );
not \U$13283 ( \13953 , \13952 );
and \U$13284 ( \13954 , \13916 , \13953 );
and \U$13285 ( \13955 , \13642 , \13915 );
nor \U$13286 ( \13956 , \13954 , \13955 );
not \U$13287 ( \13957 , \13956 );
nand \U$13288 ( \13958 , \13947 , \13943 );
and \U$13289 ( \13959 , \13940 , \13958 );
nor \U$13290 ( \13960 , \13947 , \13943 );
nor \U$13291 ( \13961 , \13959 , \13960 );
not \U$13292 ( \13962 , \13961 );
xnor \U$13293 ( \13963 , \13023 , \12920 );
not \U$13294 ( \13964 , \13921 );
not \U$13295 ( \13965 , \13935 );
or \U$13296 ( \13966 , \13964 , \13965 );
not \U$13297 ( \13967 , \13926 );
nand \U$13298 ( \13968 , \13967 , \13934 );
nand \U$13299 ( \13969 , \13966 , \13968 );
xor \U$13300 ( \13970 , \13963 , \13969 );
xnor \U$13301 ( \13971 , \13970 , \13291 );
not \U$13302 ( \13972 , \13971 );
or \U$13303 ( \13973 , \13962 , \13972 );
or \U$13304 ( \13974 , \13971 , \13961 );
nand \U$13305 ( \13975 , \13973 , \13974 );
nand \U$13306 ( \13976 , \13957 , \13975 );
not \U$13307 ( \13977 , \13976 );
not \U$13308 ( \13978 , \13640 );
not \U$13309 ( \13979 , \13600 );
or \U$13310 ( \13980 , \13978 , \13979 );
nand \U$13311 ( \13981 , \13599 , \13545 );
nand \U$13312 ( \13982 , \13980 , \13981 );
and \U$13313 ( \13983 , \13982 , \13637 );
not \U$13314 ( \13984 , \13982 );
and \U$13315 ( \13985 , \13984 , \13638 );
nor \U$13316 ( \13986 , \13983 , \13985 );
not \U$13317 ( \13987 , \13835 );
not \U$13318 ( \13988 , \13772 );
not \U$13319 ( \13989 , \13849 );
or \U$13320 ( \13990 , \13988 , \13989 );
or \U$13321 ( \13991 , \13849 , \13772 );
nand \U$13322 ( \13992 , \13990 , \13991 );
not \U$13323 ( \13993 , \13992 );
or \U$13324 ( \13994 , \13987 , \13993 );
or \U$13325 ( \13995 , \13992 , \13835 );
nand \U$13326 ( \13996 , \13994 , \13995 );
not \U$13327 ( \13997 , \12605 );
not \U$13328 ( \13998 , \12341 );
and \U$13329 ( \13999 , \12331 , \13998 , \12333 );
nand \U$13330 ( \14000 , \13999 , RIaaa6950_519);
nand \U$13331 ( \14001 , \12818 , RIaaa6860_517);
nand \U$13332 ( \14002 , \12339 , RIaaa6680_513);
nand \U$13333 ( \14003 , \12831 , \12307 );
not \U$13334 ( \14004 , \14003 );
nand \U$13335 ( \14005 , \14004 , RIaaa67e8_516);
nand \U$13336 ( \14006 , \14000 , \14001 , \14002 , \14005 );
not \U$13337 ( \14007 , RIaaa6608_512);
not \U$13338 ( \14008 , \12373 );
not \U$13339 ( \14009 , \14008 );
or \U$13340 ( \14010 , \14007 , \14009 );
not \U$13341 ( \14011 , \12832 );
not \U$13342 ( \14012 , \8537 );
and \U$13343 ( \14013 , \14011 , \14012 );
not \U$13344 ( \14014 , RIaaa6770_515);
not \U$13345 ( \14015 , \12401 );
or \U$13346 ( \14016 , \14014 , \14015 );
nand \U$13347 ( \14017 , \12476 , RIaaa64a0_509);
nand \U$13348 ( \14018 , \14016 , \14017 );
nor \U$13349 ( \14019 , \14013 , \14018 );
nand \U$13350 ( \14020 , \14010 , \14019 );
nor \U$13351 ( \14021 , \14006 , \14020 );
nand \U$13352 ( \14022 , \12344 , RIaaa6428_508);
nand \U$13353 ( \14023 , \12829 , RIaaa68d8_518);
nand \U$13354 ( \14024 , \12356 , RIaaa63b0_507);
nand \U$13355 ( \14025 , \12532 , RIaaa6590_511);
nand \U$13356 ( \14026 , \14022 , \14023 , \14024 , \14025 );
not \U$13357 ( \14027 , RIaaa66f8_514);
not \U$13358 ( \14028 , \12379 );
or \U$13359 ( \14029 , \14027 , \14028 );
not \U$13360 ( \14030 , RIaaa6518_510);
nor \U$13361 ( \14031 , \14030 , \12417 );
not \U$13362 ( \14032 , RIaaa6248_504);
not \U$13363 ( \14033 , \12951 );
or \U$13364 ( \14034 , \14032 , \14033 );
and \U$13365 ( \14035 , \12410 , RIaaa62c0_505);
nand \U$13366 ( \14036 , \11473 , RIaaa61d0_503);
not \U$13367 ( \14037 , \14036 );
nor \U$13368 ( \14038 , \14035 , \14037 );
nand \U$13369 ( \14039 , \14034 , \14038 );
nor \U$13370 ( \14040 , \14031 , \14039 );
nand \U$13371 ( \14041 , \14029 , \14040 );
nor \U$13372 ( \14042 , \14026 , \14041 );
nand \U$13373 ( \14043 , \14021 , \14042 );
not \U$13374 ( \14044 , \14043 );
buf \U$13375 ( \14045 , \14044 );
nor \U$13376 ( \14046 , \13997 , \14045 );
not \U$13377 ( \14047 , \14046 );
not \U$13378 ( \14048 , \14047 );
not \U$13379 ( \14049 , \12655 );
not \U$13380 ( \14050 , \13578 );
or \U$13381 ( \14051 , \14049 , \14050 );
and \U$13382 ( \14052 , \13559 , \12654 );
or \U$13383 ( \14053 , \13566 , \13775 );
not \U$13384 ( \14054 , \13571 );
nand \U$13385 ( \14055 , \14054 , \13775 );
nand \U$13386 ( \14056 , \14053 , \14055 );
nor \U$13387 ( \14057 , \14052 , \14056 );
nand \U$13388 ( \14058 , \14051 , \14057 );
and \U$13389 ( \14059 , \13789 , \13794 );
buf \U$13390 ( \14060 , \14059 );
not \U$13391 ( \14061 , \14060 );
not \U$13392 ( \14062 , \13567 );
or \U$13393 ( \14063 , \14061 , \14062 );
nor \U$13394 ( \14064 , \13789 , \13795 );
buf \U$13395 ( \14065 , \14064 );
not \U$13396 ( \14066 , \14065 );
buf \U$13397 ( \14067 , \14066 );
or \U$13398 ( \14068 , \12544 , \14067 );
nand \U$13399 ( \14069 , \14063 , \14068 );
nor \U$13400 ( \14070 , \13798 , \12490 );
nor \U$13401 ( \14071 , \14069 , \14070 );
not \U$13402 ( \14072 , \14071 );
and \U$13403 ( \14073 , \14058 , \14072 );
and \U$13404 ( \14074 , \13714 , \13283 );
or \U$13405 ( \14075 , \13520 , \12656 );
nand \U$13406 ( \14076 , \12911 , \12656 );
nand \U$13407 ( \14077 , \14075 , \14076 );
nor \U$13408 ( \14078 , \14074 , \14077 );
nand \U$13409 ( \14079 , \12898 , \13228 );
nand \U$13410 ( \14080 , \14078 , \14079 );
xor \U$13411 ( \14081 , \14073 , \14080 );
not \U$13412 ( \14082 , \13072 );
not \U$13413 ( \14083 , \13160 );
or \U$13414 ( \14084 , \14082 , \14083 );
not \U$13415 ( \14085 , \13532 );
and \U$13416 ( \14086 , \14085 , \13071 );
or \U$13417 ( \14087 , \13272 , \13279 );
not \U$13418 ( \14088 , \13122 );
nand \U$13419 ( \14089 , \14088 , \13704 );
nand \U$13420 ( \14090 , \14087 , \14089 );
nor \U$13421 ( \14091 , \14086 , \14090 );
nand \U$13422 ( \14092 , \14084 , \14091 );
and \U$13423 ( \14093 , \14081 , \14092 );
and \U$13424 ( \14094 , \14073 , \14080 );
nor \U$13425 ( \14095 , \14093 , \14094 );
not \U$13426 ( \14096 , \14095 );
or \U$13427 ( \14097 , \14048 , \14096 );
not \U$13428 ( \14098 , \13770 );
not \U$13429 ( \14099 , \12430 );
or \U$13430 ( \14100 , \14098 , \14099 );
not \U$13431 ( \14101 , \13769 );
buf \U$13432 ( \14102 , \14101 );
not \U$13433 ( \14103 , \14102 );
or \U$13434 ( \14104 , \12276 , \14103 );
nand \U$13435 ( \14105 , \14100 , \14104 );
not \U$13436 ( \14106 , \14105 );
not \U$13437 ( \14107 , \12274 );
not \U$13438 ( \14108 , \14107 );
or \U$13439 ( \14109 , \14106 , \14108 );
nand \U$13440 ( \14110 , \13844 , \12677 );
nand \U$13441 ( \14111 , \14109 , \14110 );
nand \U$13442 ( \14112 , \14097 , \14111 );
xor \U$13443 ( \14113 , \13996 , \14112 );
not \U$13444 ( \14114 , \13676 );
not \U$13445 ( \14115 , \12585 );
or \U$13446 ( \14116 , \14114 , \14115 );
not \U$13447 ( \14117 , \12597 );
not \U$13448 ( \14118 , \13676 );
and \U$13449 ( \14119 , \14117 , \14118 );
not \U$13450 ( \14120 , \13079 );
and \U$13451 ( \14121 , \14120 , \13893 );
nor \U$13452 ( \14122 , \14119 , \14121 );
nand \U$13453 ( \14123 , \14116 , \14122 );
not \U$13454 ( \14124 , \14123 );
not \U$13455 ( \14125 , \13788 );
not \U$13456 ( \14126 , \13805 );
not \U$13457 ( \14127 , \14126 );
and \U$13458 ( \14128 , \14125 , \14127 );
and \U$13459 ( \14129 , \13788 , \14126 );
nor \U$13460 ( \14130 , \14128 , \14129 );
not \U$13461 ( \14131 , \14130 );
not \U$13462 ( \14132 , \12780 );
and \U$13463 ( \14133 , \12783 , \12838 );
not \U$13464 ( \14134 , \12783 );
and \U$13465 ( \14135 , \14134 , \12839 );
nor \U$13466 ( \14136 , \14133 , \14135 );
not \U$13467 ( \14137 , \14136 );
or \U$13468 ( \14138 , \14132 , \14137 );
not \U$13469 ( \14139 , \12769 );
nand \U$13470 ( \14140 , \14139 , \13859 );
nand \U$13471 ( \14141 , \14138 , \14140 );
not \U$13472 ( \14142 , \14141 );
or \U$13473 ( \14143 , \14131 , \14142 );
or \U$13474 ( \14144 , \14141 , \14130 );
nand \U$13475 ( \14145 , \14143 , \14144 );
not \U$13476 ( \14146 , \14145 );
or \U$13477 ( \14147 , \14124 , \14146 );
not \U$13478 ( \14148 , \14130 );
nand \U$13479 ( \14149 , \14148 , \14141 );
nand \U$13480 ( \14150 , \14147 , \14149 );
not \U$13481 ( \14151 , \14150 );
not \U$13482 ( \14152 , \13878 );
not \U$13483 ( \14153 , \13896 );
not \U$13484 ( \14154 , \14153 );
or \U$13485 ( \14155 , \14152 , \14154 );
not \U$13486 ( \14156 , \13878 );
nand \U$13487 ( \14157 , \14156 , \13896 );
nand \U$13488 ( \14158 , \14155 , \14157 );
not \U$13489 ( \14159 , \14158 );
nand \U$13490 ( \14160 , \14151 , \14159 );
xor \U$13491 ( \14161 , \13806 , \13821 );
xor \U$13492 ( \14162 , \14161 , \13832 );
not \U$13493 ( \14163 , \14162 );
and \U$13494 ( \14164 , \14160 , \14163 );
and \U$13495 ( \14165 , \14150 , \14158 );
nor \U$13496 ( \14166 , \14164 , \14165 );
and \U$13497 ( \14167 , \14113 , \14166 );
and \U$13498 ( \14168 , \13996 , \14112 );
or \U$13499 ( \14169 , \14167 , \14168 );
xor \U$13500 ( \14170 , \13986 , \14169 );
not \U$13501 ( \14171 , \13901 );
not \U$13502 ( \14172 , \13854 );
or \U$13503 ( \14173 , \14171 , \14172 );
nand \U$13504 ( \14174 , \13904 , \13910 );
nand \U$13505 ( \14175 , \14173 , \14174 );
not \U$13506 ( \14176 , \14175 );
not \U$13507 ( \14177 , \13851 );
not \U$13508 ( \14178 , \14177 );
and \U$13509 ( \14179 , \14176 , \14178 );
not \U$13510 ( \14180 , \13851 );
and \U$13511 ( \14181 , \14175 , \14180 );
nor \U$13512 ( \14182 , \14179 , \14181 );
and \U$13513 ( \14183 , \14170 , \14182 );
and \U$13514 ( \14184 , \13986 , \14169 );
or \U$13515 ( \14185 , \14183 , \14184 );
not \U$13516 ( \14186 , \14185 );
not \U$13517 ( \14187 , \13916 );
not \U$13518 ( \14188 , \13952 );
and \U$13519 ( \14189 , \14187 , \14188 );
and \U$13520 ( \14190 , \13952 , \13916 );
nor \U$13521 ( \14191 , \14189 , \14190 );
not \U$13522 ( \14192 , \14191 );
nand \U$13523 ( \14193 , \14186 , \14192 );
not \U$13524 ( \14194 , \14193 );
or \U$13525 ( \14195 , \13977 , \14194 );
not \U$13526 ( \14196 , \13975 );
nand \U$13527 ( \14197 , \14196 , \13956 );
nand \U$13528 ( \14198 , \14195 , \14197 );
not \U$13529 ( \14199 , \13296 );
not \U$13530 ( \14200 , \14199 );
not \U$13531 ( \14201 , \13373 );
or \U$13532 ( \14202 , \14200 , \14201 );
or \U$13533 ( \14203 , \13373 , \14199 );
nand \U$13534 ( \14204 , \14202 , \14203 );
not \U$13535 ( \14205 , \13969 );
buf \U$13536 ( \14206 , \13963 );
not \U$13537 ( \14207 , \14206 );
not \U$13538 ( \14208 , \13291 );
or \U$13539 ( \14209 , \14207 , \14208 );
or \U$13540 ( \14210 , \13291 , \14206 );
nand \U$13541 ( \14211 , \14209 , \14210 );
not \U$13542 ( \14212 , \14211 );
or \U$13543 ( \14213 , \14205 , \14212 );
nand \U$13544 ( \14214 , \14213 , \13961 );
or \U$13545 ( \14215 , \14211 , \13969 );
nand \U$13546 ( \14216 , \14214 , \14215 );
nand \U$13547 ( \14217 , \14204 , \14216 );
buf \U$13548 ( \14218 , \14217 );
not \U$13549 ( \14219 , \14218 );
or \U$13550 ( \14220 , \14198 , \14219 );
or \U$13551 ( \14221 , \14204 , \14216 );
nand \U$13552 ( \14222 , \14220 , \14221 );
nand \U$13553 ( \14223 , \13466 , \13378 );
buf \U$13554 ( \14224 , \14223 );
nand \U$13555 ( \14225 , \14222 , \14224 );
not \U$13556 ( \14226 , \14225 );
or \U$13557 ( \14227 , \13468 , \14226 );
not \U$13558 ( \14228 , \13390 );
not \U$13559 ( \14229 , \13462 );
not \U$13560 ( \14230 , \14229 );
or \U$13561 ( \14231 , \14228 , \14230 );
buf \U$13562 ( \14232 , \13454 );
xor \U$13563 ( \14233 , \13409 , \14232 );
not \U$13564 ( \14234 , \13460 );
xnor \U$13565 ( \14235 , \14233 , \14234 );
nand \U$13566 ( \14236 , \14235 , \13414 );
nand \U$13567 ( \14237 , \14231 , \14236 );
buf \U$13568 ( \14238 , \13283 );
not \U$13569 ( \14239 , \14238 );
not \U$13570 ( \14240 , \12280 );
or \U$13571 ( \14241 , \14239 , \14240 );
not \U$13572 ( \14242 , \14238 );
and \U$13573 ( \14243 , \12432 , \14242 );
and \U$13574 ( \14244 , \12659 , \13395 );
not \U$13575 ( \14245 , \12659 );
and \U$13576 ( \14246 , \14245 , \12437 );
nor \U$13577 ( \14247 , \14244 , \14246 );
nor \U$13578 ( \14248 , \14243 , \14247 );
nand \U$13579 ( \14249 , \14241 , \14248 );
not \U$13580 ( \14250 , \12545 );
not \U$13581 ( \14251 , \13421 );
or \U$13582 ( \14252 , \14250 , \14251 );
and \U$13583 ( \14253 , \13346 , \12544 );
or \U$13584 ( \14254 , \12707 , \13122 );
nand \U$13585 ( \14255 , \14254 , \13431 );
nor \U$13586 ( \14256 , \14253 , \14255 );
nand \U$13587 ( \14257 , \14252 , \14256 );
xnor \U$13588 ( \14258 , \14249 , \14257 );
and \U$13589 ( \14259 , \12585 , \12426 );
not \U$13590 ( \14260 , \12425 );
not \U$13591 ( \14261 , \12598 );
not \U$13592 ( \14262 , \14261 );
or \U$13593 ( \14263 , \14260 , \14262 );
and \U$13594 ( \14264 , \12497 , \13286 );
not \U$13595 ( \14265 , \12497 );
and \U$13596 ( \14266 , \14265 , \12601 );
nor \U$13597 ( \14267 , \14264 , \14266 );
nand \U$13598 ( \14268 , \14263 , \14267 );
nor \U$13599 ( \14269 , \14259 , \14268 );
not \U$13600 ( \14270 , \14269 );
xor \U$13601 ( \14271 , \13408 , \14270 );
not \U$13602 ( \14272 , \13436 );
not \U$13603 ( \14273 , \13449 );
or \U$13604 ( \14274 , \14272 , \14273 );
nand \U$13605 ( \14275 , \13435 , \13419 );
nand \U$13606 ( \14276 , \14274 , \14275 );
xnor \U$13607 ( \14277 , \14271 , \14276 );
xor \U$13608 ( \14278 , \14258 , \14277 );
not \U$13609 ( \14279 , \14232 );
and \U$13610 ( \14280 , \14234 , \14279 );
nor \U$13611 ( \14281 , \14280 , \13409 );
and \U$13612 ( \14282 , \13454 , \13460 );
nor \U$13613 ( \14283 , \14281 , \14282 );
xor \U$13614 ( \14284 , \14278 , \14283 );
nand \U$13615 ( \14285 , \14237 , \14284 );
not \U$13616 ( \14286 , \12490 );
not \U$13617 ( \14287 , \13891 );
not \U$13618 ( \14288 , \14287 );
or \U$13619 ( \14289 , \14286 , \14288 );
or \U$13620 ( \14290 , \14287 , \12497 );
nand \U$13621 ( \14291 , \14289 , \14290 );
not \U$13622 ( \14292 , \14291 );
not \U$13623 ( \14293 , \13079 );
or \U$13624 ( \14294 , \14292 , \14293 );
xor \U$13625 ( \14295 , \12544 , \13891 );
not \U$13626 ( \14296 , \14295 );
not \U$13627 ( \14297 , \14120 );
or \U$13628 ( \14298 , \14296 , \14297 );
not \U$13629 ( \14299 , \13884 );
nand \U$13630 ( \14300 , \14298 , \14299 );
nand \U$13631 ( \14301 , \14294 , \14300 );
not \U$13632 ( \14302 , \13869 );
and \U$13633 ( \14303 , \12781 , \14302 );
nor \U$13634 ( \14304 , \14303 , \12844 );
xor \U$13635 ( \14305 , \14301 , \14304 );
not \U$13636 ( \14306 , \12281 );
not \U$13637 ( \14307 , \12659 );
and \U$13638 ( \14308 , \14306 , \14307 );
or \U$13639 ( \14309 , \12433 , \12658 );
and \U$13640 ( \14310 , \12496 , \12426 );
nor \U$13641 ( \14311 , \12437 , \12426 );
nor \U$13642 ( \14312 , \14310 , \14311 );
nand \U$13643 ( \14313 , \14309 , \14312 );
nor \U$13644 ( \14314 , \14308 , \14313 );
and \U$13645 ( \14315 , \14305 , \14314 );
and \U$13646 ( \14316 , \14301 , \14304 );
or \U$13647 ( \14317 , \14315 , \14316 );
xor \U$13648 ( \14318 , \12501 , \12661 );
xor \U$13649 ( \14319 , \14317 , \14318 );
not \U$13650 ( \14320 , \14242 );
not \U$13651 ( \14321 , \12606 );
or \U$13652 ( \14322 , \14320 , \14321 );
nand \U$13653 ( \14323 , \14322 , \14269 );
xor \U$13654 ( \14324 , \14301 , \14304 );
xor \U$13655 ( \14325 , \14324 , \14314 );
not \U$13656 ( \14326 , \14325 );
nand \U$13657 ( \14327 , \14323 , \14326 );
xor \U$13658 ( \14328 , \14319 , \14327 );
and \U$13659 ( \14329 , \14249 , \14257 );
not \U$13660 ( \14330 , \13408 );
not \U$13661 ( \14331 , \14330 );
xnor \U$13662 ( \14332 , \14270 , \14276 );
not \U$13663 ( \14333 , \14332 );
or \U$13664 ( \14334 , \14331 , \14333 );
not \U$13665 ( \14335 , \14270 );
nand \U$13666 ( \14336 , \14335 , \14276 );
nand \U$13667 ( \14337 , \14334 , \14336 );
xor \U$13668 ( \14338 , \14329 , \14337 );
not \U$13669 ( \14339 , \14326 );
not \U$13670 ( \14340 , \14323 );
not \U$13671 ( \14341 , \14340 );
or \U$13672 ( \14342 , \14339 , \14341 );
nand \U$13673 ( \14343 , \14325 , \14323 );
nand \U$13674 ( \14344 , \14342 , \14343 );
and \U$13675 ( \14345 , \14338 , \14344 );
and \U$13676 ( \14346 , \14329 , \14337 );
nor \U$13677 ( \14347 , \14345 , \14346 );
nand \U$13678 ( \14348 , \14328 , \14347 );
xor \U$13679 ( \14349 , \14329 , \14344 );
xnor \U$13680 ( \14350 , \14349 , \14337 );
xor \U$13681 ( \14351 , \14258 , \14277 );
and \U$13682 ( \14352 , \14351 , \14283 );
and \U$13683 ( \14353 , \14258 , \14277 );
or \U$13684 ( \14354 , \14352 , \14353 );
nand \U$13685 ( \14355 , \14350 , \14354 );
xor \U$13686 ( \14356 , \14317 , \14318 );
and \U$13687 ( \14357 , \14356 , \14327 );
and \U$13688 ( \14358 , \14317 , \14318 );
or \U$13689 ( \14359 , \14357 , \14358 );
xor \U$13690 ( \14360 , \12604 , \12697 );
not \U$13691 ( \14361 , \14360 );
not \U$13692 ( \14362 , \12501 );
nand \U$13693 ( \14363 , \14362 , \12661 );
nand \U$13694 ( \14364 , \14363 , \12660 );
not \U$13695 ( \14365 , \14364 );
or \U$13696 ( \14366 , \14361 , \14365 );
or \U$13697 ( \14367 , \14364 , \14360 );
nand \U$13698 ( \14368 , \14366 , \14367 );
nand \U$13699 ( \14369 , \14359 , \14368 );
and \U$13700 ( \14370 , \14285 , \14348 , \14355 , \14369 );
nand \U$13701 ( \14371 , \14227 , \14370 );
xor \U$13702 ( \14372 , \14150 , \14162 );
xor \U$13703 ( \14373 , \14372 , \14159 );
not \U$13704 ( \14374 , \12971 );
not \U$13705 ( \14375 , \13160 );
or \U$13706 ( \14376 , \14374 , \14375 );
and \U$13707 ( \14377 , \14085 , \13026 );
or \U$13708 ( \14378 , \13272 , \13072 );
nand \U$13709 ( \14379 , \13269 , \13072 );
nand \U$13710 ( \14380 , \14378 , \14379 );
nor \U$13711 ( \14381 , \14377 , \14380 );
nand \U$13712 ( \14382 , \14376 , \14381 );
not \U$13713 ( \14383 , \14382 );
not \U$13714 ( \14384 , \13122 );
not \U$13715 ( \14385 , \12904 );
or \U$13716 ( \14386 , \14384 , \14385 );
and \U$13717 ( \14387 , \12913 , \13227 );
nor \U$13718 ( \14388 , \13520 , \13227 );
nor \U$13719 ( \14389 , \14387 , \14388 );
nand \U$13720 ( \14390 , \14386 , \14389 );
not \U$13721 ( \14391 , \14390 );
nand \U$13722 ( \14392 , \13578 , \13228 );
not \U$13723 ( \14393 , \14392 );
and \U$13724 ( \14394 , \13559 , \13227 );
or \U$13725 ( \14395 , \13572 , \12655 );
or \U$13726 ( \14396 , \13566 , \12654 );
nand \U$13727 ( \14397 , \14395 , \14396 );
nor \U$13728 ( \14398 , \14394 , \14397 );
not \U$13729 ( \14399 , \14398 );
or \U$13730 ( \14400 , \14393 , \14399 );
not \U$13731 ( \14401 , \14067 );
nand \U$13732 ( \14402 , \14401 , \12490 );
nand \U$13733 ( \14403 , \14060 , \13560 );
buf \U$13734 ( \14404 , \13796 );
not \U$13735 ( \14405 , \14404 );
nand \U$13736 ( \14406 , \14405 , \12424 );
and \U$13737 ( \14407 , \14402 , \14403 , \14406 );
not \U$13738 ( \14408 , \14407 );
nand \U$13739 ( \14409 , \14400 , \14408 );
nand \U$13740 ( \14410 , \12898 , \13279 );
nand \U$13741 ( \14411 , \14391 , \14409 , \14410 );
not \U$13742 ( \14412 , \14411 );
or \U$13743 ( \14413 , \14383 , \14412 );
not \U$13744 ( \14414 , \14410 );
or \U$13745 ( \14415 , \14390 , \14414 );
not \U$13746 ( \14416 , \14409 );
nand \U$13747 ( \14417 , \14415 , \14416 );
nand \U$13748 ( \14418 , \14413 , \14417 );
nand \U$13749 ( \14419 , \12327 , RIaaa5618_478);
nand \U$13750 ( \14420 , \13999 , RIaaa58e8_484);
nand \U$13751 ( \14421 , RIaaa5708_480, \12339 );
nand \U$13752 ( \14422 , \12829 , RIaaa5960_485);
nand \U$13753 ( \14423 , \14419 , \14420 , \14421 , \14422 );
not \U$13754 ( \14424 , \12452 );
nand \U$13755 ( \14425 , \14424 , RIaaa5348_472);
nand \U$13756 ( \14426 , \12356 , RIaaa5258_470);
nand \U$13757 ( \14427 , \12833 , RIaaa5528_476);
nand \U$13758 ( \14428 , \12532 , RIaaa53c0_473);
nand \U$13759 ( \14429 , \14425 , \14426 , \14427 , \14428 );
nor \U$13760 ( \14430 , \14423 , \14429 );
not \U$13761 ( \14431 , RIaaa5780_481);
not \U$13762 ( \14432 , \14008 );
or \U$13763 ( \14433 , \14431 , \14432 );
nand \U$13764 ( \14434 , \13032 , RIaaa57f8_482);
nand \U$13765 ( \14435 , \14433 , \14434 );
not \U$13766 ( \14436 , \13006 );
not \U$13767 ( \14437 , RIaaa5870_483);
not \U$13768 ( \14438 , \14437 );
and \U$13769 ( \14439 , \14436 , \14438 );
nor \U$13770 ( \14440 , \12417 , \8953 );
nor \U$13771 ( \14441 , \14439 , \14440 );
nand \U$13772 ( \14442 , \14004 , RIaaa5690_479);
and \U$13773 ( \14443 , \12476 , RIaaa52d0_471);
not \U$13774 ( \14444 , RIaaa55a0_477);
not \U$13775 ( \14445 , \12410 );
or \U$13776 ( \14446 , \14444 , \14445 );
nand \U$13777 ( \14447 , \11473 , RIaaa51e0_469);
nand \U$13778 ( \14448 , \14446 , \14447 );
nor \U$13779 ( \14449 , \14443 , \14448 );
nand \U$13780 ( \14450 , \12395 , RIaaa54b0_475);
nand \U$13781 ( \14451 , \14441 , \14442 , \14449 , \14450 );
nor \U$13782 ( \14452 , \14435 , \14451 );
and \U$13783 ( \14453 , \14430 , \14452 );
buf \U$13784 ( \14454 , \14453 );
not \U$13785 ( \14455 , \14454 );
and \U$13786 ( \14456 , \12605 , \14455 );
not \U$13787 ( \14457 , \14045 );
not \U$13788 ( \14458 , \12277 );
or \U$13789 ( \14459 , \14457 , \14458 );
or \U$13790 ( \14460 , \12682 , \14045 );
nand \U$13791 ( \14461 , \14459 , \14460 );
not \U$13792 ( \14462 , \14461 );
not \U$13793 ( \14463 , \12275 );
or \U$13794 ( \14464 , \14462 , \14463 );
nand \U$13795 ( \14465 , \14105 , \12677 );
nand \U$13796 ( \14466 , \14464 , \14465 );
xor \U$13797 ( \14467 , \14456 , \14466 );
and \U$13798 ( \14468 , \14418 , \14467 );
not \U$13799 ( \14469 , \14418 );
not \U$13800 ( \14470 , \14467 );
and \U$13801 ( \14471 , \14469 , \14470 );
nor \U$13802 ( \14472 , \14468 , \14471 );
nand \U$13803 ( \14473 , \13032 , RIaaa49e8_452);
nand \U$13804 ( \14474 , \12829 , RIaaa4d30_459);
nand \U$13805 ( \14475 , \12356 , RIaaa5000_465);
nand \U$13806 ( \14476 , \12532 , RIaaa4da8_460);
nand \U$13807 ( \14477 , \14473 , \14474 , \14475 , \14476 );
not \U$13808 ( \14478 , RIaaa5078_466);
not \U$13809 ( \14479 , \12453 );
or \U$13810 ( \14480 , \14478 , \14479 );
not \U$13811 ( \14481 , \13758 );
not \U$13812 ( \14482 , \8768 );
and \U$13813 ( \14483 , \14481 , \14482 );
not \U$13814 ( \14484 , RIaaa4f10_463);
nand \U$13815 ( \14485 , \12399 , \12400 );
not \U$13816 ( \14486 , \14485 );
not \U$13817 ( \14487 , \12319 );
nand \U$13818 ( \14488 , \14486 , \14487 );
not \U$13819 ( \14489 , \14488 );
not \U$13820 ( \14490 , \14489 );
or \U$13821 ( \14491 , \14484 , \14490 );
and \U$13822 ( \14492 , \12410 , RIaaa4bc8_456);
nand \U$13823 ( \14493 , \11473 , RIaaa4ad8_454);
not \U$13824 ( \14494 , \14493 );
nor \U$13825 ( \14495 , \14492 , \14494 );
nand \U$13826 ( \14496 , \14491 , \14495 );
nor \U$13827 ( \14497 , \14483 , \14496 );
nand \U$13828 ( \14498 , \14480 , \14497 );
nor \U$13829 ( \14499 , \14477 , \14498 );
nand \U$13830 ( \14500 , \14008 , RIaaa5168_468);
and \U$13831 ( \14501 , \12402 , RIaaa4a60_453);
and \U$13832 ( \14502 , \12476 , RIaaa4f88_464);
nor \U$13833 ( \14503 , \14501 , \14502 );
nand \U$13834 ( \14504 , \12833 , RIaaa4c40_457);
nand \U$13835 ( \14505 , \14500 , \14503 , \14504 );
nand \U$13836 ( \14506 , \12339 , RIaaa50f0_467);
nand \U$13837 ( \14507 , \12818 , RIaaa4e98_462);
nand \U$13838 ( \14508 , \13999 , RIaaa4cb8_458);
nand \U$13839 ( \14509 , \14004 , RIaaa4e20_461);
nand \U$13840 ( \14510 , \14506 , \14507 , \14508 , \14509 );
nor \U$13841 ( \14511 , \14505 , \14510 );
and \U$13842 ( \14512 , \14499 , \14511 );
buf \U$13843 ( \14513 , \14512 );
not \U$13844 ( \14514 , \14513 );
nand \U$13845 ( \14515 , \12605 , \14514 );
not \U$13846 ( \14516 , \14515 );
not \U$13847 ( \14517 , \14454 );
not \U$13848 ( \14518 , \14517 );
not \U$13849 ( \14519 , \12276 );
or \U$13850 ( \14520 , \14518 , \14519 );
or \U$13851 ( \14521 , \13682 , \14517 );
nand \U$13852 ( \14522 , \14520 , \14521 );
not \U$13853 ( \14523 , \14522 );
not \U$13854 ( \14524 , \12275 );
or \U$13855 ( \14525 , \14523 , \14524 );
nand \U$13856 ( \14526 , \14461 , \12677 );
nand \U$13857 ( \14527 , \14525 , \14526 );
not \U$13858 ( \14528 , \14527 );
or \U$13859 ( \14529 , \14516 , \14528 );
or \U$13860 ( \14530 , \14527 , \14515 );
nand \U$13861 ( \14531 , \14529 , \14530 );
not \U$13862 ( \14532 , \14531 );
not \U$13863 ( \14533 , \12838 );
not \U$13864 ( \14534 , \13267 );
or \U$13865 ( \14535 , \14533 , \14534 );
and \U$13866 ( \14536 , \13026 , \13169 );
not \U$13867 ( \14537 , \13026 );
and \U$13868 ( \14538 , \14537 , \13704 );
nor \U$13869 ( \14539 , \14536 , \14538 );
nand \U$13870 ( \14540 , \14535 , \14539 );
not \U$13871 ( \14541 , \13160 );
nor \U$13872 ( \14542 , \14541 , \12838 );
nor \U$13873 ( \14543 , \14540 , \14542 );
not \U$13874 ( \14544 , \14543 );
not \U$13875 ( \14545 , \14544 );
not \U$13876 ( \14546 , \13121 );
not \U$13877 ( \14547 , \14546 );
not \U$13878 ( \14548 , \13578 );
or \U$13879 ( \14549 , \14547 , \14548 );
and \U$13880 ( \14550 , \13559 , \13121 );
and \U$13881 ( \14551 , \13226 , \13572 );
not \U$13882 ( \14552 , \13226 );
and \U$13883 ( \14553 , \14552 , \13566 );
nor \U$13884 ( \14554 , \14551 , \14553 );
nor \U$13885 ( \14555 , \14550 , \14554 );
nand \U$13886 ( \14556 , \14549 , \14555 );
not \U$13887 ( \14557 , \12656 );
not \U$13888 ( \14558 , \13799 );
or \U$13889 ( \14559 , \14557 , \14558 );
not \U$13890 ( \14560 , \12423 );
not \U$13891 ( \14561 , \13804 );
and \U$13892 ( \14562 , \14560 , \14561 );
and \U$13893 ( \14563 , \14401 , \13776 );
nor \U$13894 ( \14564 , \14562 , \14563 );
nand \U$13895 ( \14565 , \14559 , \14564 );
nand \U$13896 ( \14566 , \14556 , \14565 );
not \U$13897 ( \14567 , \14566 );
and \U$13898 ( \14568 , \12904 , \13071 );
not \U$13899 ( \14569 , \13121 );
not \U$13900 ( \14570 , \13718 );
or \U$13901 ( \14571 , \14569 , \14570 );
or \U$13902 ( \14572 , \13520 , \13122 );
nand \U$13903 ( \14573 , \14571 , \14572 );
nor \U$13904 ( \14574 , \14568 , \14573 );
nand \U$13905 ( \14575 , \12898 , \13072 );
nand \U$13906 ( \14576 , \14574 , \14575 );
not \U$13907 ( \14577 , \14576 );
or \U$13908 ( \14578 , \14567 , \14577 );
nand \U$13909 ( \14579 , \14574 , \14575 , \14556 , \14565 );
nand \U$13910 ( \14580 , \14578 , \14579 );
not \U$13911 ( \14581 , \14580 );
or \U$13912 ( \14582 , \14545 , \14581 );
not \U$13913 ( \14583 , \14575 );
not \U$13914 ( \14584 , \14574 );
or \U$13915 ( \14585 , \14583 , \14584 );
not \U$13916 ( \14586 , \14566 );
nand \U$13917 ( \14587 , \14585 , \14586 );
nand \U$13918 ( \14588 , \14582 , \14587 );
not \U$13919 ( \14589 , \14588 );
or \U$13920 ( \14590 , \14532 , \14589 );
not \U$13921 ( \14591 , \14515 );
nand \U$13922 ( \14592 , \14591 , \14527 );
nand \U$13923 ( \14593 , \14590 , \14592 );
xor \U$13924 ( \14594 , \14472 , \14593 );
not \U$13925 ( \14595 , \13770 );
not \U$13926 ( \14596 , \12585 );
or \U$13927 ( \14597 , \14595 , \14596 );
or \U$13928 ( \14598 , \13627 , \14118 );
nand \U$13929 ( \14599 , \13081 , \14118 );
nand \U$13930 ( \14600 , \14598 , \14599 );
nor \U$13931 ( \14601 , \12597 , \13770 );
nor \U$13932 ( \14602 , \14600 , \14601 );
nand \U$13933 ( \14603 , \14597 , \14602 );
not \U$13934 ( \14604 , \13886 );
not \U$13935 ( \14605 , \12844 );
or \U$13936 ( \14606 , \14604 , \14605 );
or \U$13937 ( \14607 , \12844 , \13021 );
nand \U$13938 ( \14608 , \14606 , \14607 );
not \U$13939 ( \14609 , \14608 );
not \U$13940 ( \14610 , \13861 );
or \U$13941 ( \14611 , \14609 , \14610 );
nand \U$13942 ( \14612 , \14136 , \13245 );
nand \U$13943 ( \14613 , \14611 , \14612 );
not \U$13944 ( \14614 , \14613 );
not \U$13945 ( \14615 , \14058 );
not \U$13946 ( \14616 , \14071 );
and \U$13947 ( \14617 , \14615 , \14616 );
and \U$13948 ( \14618 , \14058 , \14071 );
nor \U$13949 ( \14619 , \14617 , \14618 );
not \U$13950 ( \14620 , \14619 );
or \U$13951 ( \14621 , \14614 , \14620 );
or \U$13952 ( \14622 , \14613 , \14619 );
nand \U$13953 ( \14623 , \14621 , \14622 );
xor \U$13954 ( \14624 , \14603 , \14623 );
not \U$13955 ( \14625 , \14624 );
not \U$13956 ( \14626 , \13771 );
not \U$13957 ( \14627 , \12601 );
or \U$13958 ( \14628 , \14626 , \14627 );
and \U$13959 ( \14629 , \13328 , \13770 );
not \U$13960 ( \14630 , \14044 );
not \U$13961 ( \14631 , \12564 );
or \U$13962 ( \14632 , \14630 , \14631 );
or \U$13963 ( \14633 , \12669 , \14045 );
nand \U$13964 ( \14634 , \14632 , \14633 );
and \U$13965 ( \14635 , \13884 , \14634 );
nor \U$13966 ( \14636 , \14629 , \14635 );
nand \U$13967 ( \14637 , \14628 , \14636 );
not \U$13968 ( \14638 , \14637 );
nand \U$13969 ( \14639 , \14398 , \14392 );
not \U$13970 ( \14640 , \14639 );
not \U$13971 ( \14641 , \14407 );
and \U$13972 ( \14642 , \14640 , \14641 );
and \U$13973 ( \14643 , \14639 , \14407 );
nor \U$13974 ( \14644 , \14642 , \14643 );
not \U$13975 ( \14645 , \14644 );
not \U$13976 ( \14646 , \14645 );
not \U$13977 ( \14647 , \13842 );
not \U$13978 ( \14648 , \12844 );
not \U$13979 ( \14649 , \14648 );
not \U$13980 ( \14650 , \14649 );
or \U$13981 ( \14651 , \14647 , \14650 );
or \U$13982 ( \14652 , \13231 , \13676 );
nand \U$13983 ( \14653 , \14651 , \14652 );
not \U$13984 ( \14654 , \14653 );
not \U$13985 ( \14655 , \13861 );
or \U$13986 ( \14656 , \14654 , \14655 );
not \U$13987 ( \14657 , \13430 );
not \U$13988 ( \14658 , \13021 );
and \U$13989 ( \14659 , \14657 , \14658 );
and \U$13990 ( \14660 , \12783 , \12845 );
not \U$13991 ( \14661 , \13886 );
not \U$13992 ( \14662 , \14661 );
and \U$13993 ( \14663 , \14660 , \14662 );
nor \U$13994 ( \14664 , \14659 , \14663 );
nand \U$13995 ( \14665 , \14656 , \14664 );
not \U$13996 ( \14666 , \14665 );
not \U$13997 ( \14667 , \14666 );
or \U$13998 ( \14668 , \14646 , \14667 );
nand \U$13999 ( \14669 , \14665 , \14644 );
nand \U$14000 ( \14670 , \14668 , \14669 );
not \U$14001 ( \14671 , \14670 );
or \U$14002 ( \14672 , \14638 , \14671 );
nand \U$14003 ( \14673 , \14665 , \14645 );
nand \U$14004 ( \14674 , \14672 , \14673 );
not \U$14005 ( \14675 , \14674 );
or \U$14006 ( \14676 , \14625 , \14675 );
or \U$14007 ( \14677 , \14674 , \14624 );
nand \U$14008 ( \14678 , \14411 , \14417 );
not \U$14009 ( \14679 , \14678 );
not \U$14010 ( \14680 , \14382 );
and \U$14011 ( \14681 , \14679 , \14680 );
and \U$14012 ( \14682 , \14678 , \14382 );
nor \U$14013 ( \14683 , \14681 , \14682 );
not \U$14014 ( \14684 , \14683 );
nand \U$14015 ( \14685 , \14677 , \14684 );
nand \U$14016 ( \14686 , \14676 , \14685 );
and \U$14017 ( \14687 , \14594 , \14686 );
and \U$14018 ( \14688 , \14472 , \14593 );
or \U$14019 ( \14689 , \14687 , \14688 );
xor \U$14020 ( \14690 , \14373 , \14689 );
and \U$14021 ( \14691 , \14418 , \14467 );
and \U$14022 ( \14692 , \14456 , \14466 );
nor \U$14023 ( \14693 , \14691 , \14692 );
not \U$14024 ( \14694 , \14693 );
not \U$14025 ( \14695 , \14111 );
not \U$14026 ( \14696 , \14046 );
and \U$14027 ( \14697 , \14695 , \14696 );
and \U$14028 ( \14698 , \14111 , \14046 );
nor \U$14029 ( \14699 , \14697 , \14698 );
not \U$14030 ( \14700 , \14699 );
not \U$14031 ( \14701 , \14095 );
or \U$14032 ( \14702 , \14700 , \14701 );
or \U$14033 ( \14703 , \14095 , \14699 );
nand \U$14034 ( \14704 , \14702 , \14703 );
nand \U$14035 ( \14705 , \14694 , \14704 );
not \U$14036 ( \14706 , \14704 );
nand \U$14037 ( \14707 , \14706 , \14693 );
nand \U$14038 ( \14708 , \14705 , \14707 );
xnor \U$14039 ( \14709 , \14123 , \14145 );
not \U$14040 ( \14710 , \14613 );
not \U$14041 ( \14711 , \14710 );
not \U$14042 ( \14712 , \14619 );
and \U$14043 ( \14713 , \14711 , \14712 );
and \U$14044 ( \14714 , \14603 , \14623 );
nor \U$14045 ( \14715 , \14713 , \14714 );
nand \U$14046 ( \14716 , \14709 , \14715 );
xor \U$14047 ( \14717 , \14092 , \14081 );
and \U$14048 ( \14718 , \14716 , \14717 );
nor \U$14049 ( \14719 , \14709 , \14715 );
nor \U$14050 ( \14720 , \14718 , \14719 );
and \U$14051 ( \14721 , \14708 , \14720 );
not \U$14052 ( \14722 , \14708 );
not \U$14053 ( \14723 , \14720 );
and \U$14054 ( \14724 , \14722 , \14723 );
nor \U$14055 ( \14725 , \14721 , \14724 );
xor \U$14056 ( \14726 , \14690 , \14725 );
not \U$14057 ( \14727 , \14726 );
not \U$14058 ( \14728 , \14709 );
not \U$14059 ( \14729 , \14728 );
not \U$14060 ( \14730 , \14715 );
not \U$14061 ( \14731 , \14717 );
and \U$14062 ( \14732 , \14730 , \14731 );
and \U$14063 ( \14733 , \14717 , \14715 );
nor \U$14064 ( \14734 , \14732 , \14733 );
not \U$14065 ( \14735 , \14734 );
not \U$14066 ( \14736 , \14735 );
or \U$14067 ( \14737 , \14729 , \14736 );
not \U$14068 ( \14738 , \14728 );
nand \U$14069 ( \14739 , \14738 , \14734 );
nand \U$14070 ( \14740 , \14737 , \14739 );
and \U$14071 ( \14741 , \14513 , \12493 );
not \U$14072 ( \14742 , \14513 );
and \U$14073 ( \14743 , \14742 , \12276 );
or \U$14074 ( \14744 , \14741 , \14743 );
not \U$14075 ( \14745 , \14744 );
not \U$14076 ( \14746 , \12274 );
not \U$14077 ( \14747 , \14746 );
or \U$14078 ( \14748 , \14745 , \14747 );
nand \U$14079 ( \14749 , \14522 , \12677 );
nand \U$14080 ( \14750 , \14748 , \14749 );
not \U$14081 ( \14751 , \14750 );
not \U$14082 ( \14752 , \14751 );
and \U$14083 ( \14753 , \12418 , RIaaa5ac8_488);
and \U$14084 ( \14754 , \12951 , RIaaa5e10_495);
nor \U$14085 ( \14755 , \14753 , \14754 );
nand \U$14086 ( \14756 , \12356 , RIaaa5bb8_490);
nand \U$14087 ( \14757 , \14004 , RIaaa5a50_487);
and \U$14088 ( \14758 , \12402 , RIaaa5d20_493);
not \U$14089 ( \14759 , RIaaa5e88_496);
not \U$14090 ( \14760 , \12410 );
or \U$14091 ( \14761 , \14759 , \14760 );
nand \U$14092 ( \14762 , \11473 , RIaaa5d98_494);
nand \U$14093 ( \14763 , \14761 , \14762 );
nor \U$14094 ( \14764 , \14758 , \14763 );
nand \U$14095 ( \14765 , \14755 , \14756 , \14757 , \14764 );
not \U$14096 ( \14766 , RIaaa5ca8_492);
not \U$14097 ( \14767 , \12379 );
or \U$14098 ( \14768 , \14766 , \14767 );
nand \U$14099 ( \14769 , \12360 , RIaaa6068_500);
nand \U$14100 ( \14770 , \14768 , \14769 );
nor \U$14101 ( \14771 , \14765 , \14770 );
not \U$14102 ( \14772 , RIaaa59d8_486);
not \U$14103 ( \14773 , \12327 );
or \U$14104 ( \14774 , \14772 , \14773 );
not \U$14105 ( \14775 , \12612 );
not \U$14106 ( \14776 , \4153 );
and \U$14107 ( \14777 , \14775 , \14776 );
and \U$14108 ( \14778 , \12365 , RIaaa5f00_497);
nor \U$14109 ( \14779 , \14777 , \14778 );
nand \U$14110 ( \14780 , \14774 , \14779 );
not \U$14111 ( \14781 , RIaaa5f78_498);
not \U$14112 ( \14782 , \12449 );
or \U$14113 ( \14783 , \14781 , \14782 );
nand \U$14114 ( \14784 , \14008 , RIaaa6158_502);
nand \U$14115 ( \14785 , \14783 , \14784 );
nor \U$14116 ( \14786 , \14780 , \14785 );
and \U$14117 ( \14787 , \12339 , RIaaa60e0_501);
not \U$14118 ( \14788 , RIaaa5c30_491);
not \U$14119 ( \14789 , \12453 );
or \U$14120 ( \14790 , \14788 , \14789 );
not \U$14121 ( \14791 , \12350 );
nand \U$14122 ( \14792 , \14791 , RIaaa5ff0_499);
nand \U$14123 ( \14793 , \14790 , \14792 );
nor \U$14124 ( \14794 , \14787 , \14793 );
and \U$14125 ( \14795 , \14771 , \14786 , \14794 );
buf \U$14126 ( \14796 , \14795 );
not \U$14127 ( \14797 , \14796 );
nand \U$14128 ( \14798 , \12841 , \14797 );
not \U$14129 ( \14799 , \14798 );
and \U$14130 ( \14800 , \14752 , \14799 );
not \U$14131 ( \14801 , \13070 );
not \U$14132 ( \14802 , \13578 );
or \U$14133 ( \14803 , \14801 , \14802 );
not \U$14134 ( \14804 , \13570 );
nand \U$14135 ( \14805 , \14804 , \13510 );
nor \U$14136 ( \14806 , \14805 , \13515 );
buf \U$14137 ( \14807 , \14806 );
and \U$14138 ( \14808 , \14807 , \13071 );
not \U$14139 ( \14809 , \13781 );
not \U$14140 ( \14810 , \13120 );
or \U$14141 ( \14811 , \14809 , \14810 );
not \U$14142 ( \14812 , \13562 );
and \U$14143 ( \14813 , \14812 , \13564 );
not \U$14144 ( \14814 , \14813 );
or \U$14145 ( \14815 , \14814 , \13120 );
nand \U$14146 ( \14816 , \14811 , \14815 );
nor \U$14147 ( \14817 , \14808 , \14816 );
nand \U$14148 ( \14818 , \14803 , \14817 );
not \U$14149 ( \14819 , \14065 );
or \U$14150 ( \14820 , \12654 , \14819 );
nand \U$14151 ( \14821 , \14405 , \13226 );
nand \U$14152 ( \14822 , \14060 , \12654 );
nand \U$14153 ( \14823 , \14820 , \14821 , \14822 );
and \U$14154 ( \14824 , \14818 , \14823 );
not \U$14155 ( \14825 , \14824 );
not \U$14156 ( \14826 , \12971 );
not \U$14157 ( \14827 , \13525 );
or \U$14158 ( \14828 , \14826 , \14827 );
not \U$14159 ( \14829 , \12894 );
nand \U$14160 ( \14830 , \14829 , \13812 );
not \U$14161 ( \14831 , \14830 );
and \U$14162 ( \14832 , \14831 , \13026 );
not \U$14163 ( \14833 , \13070 );
or \U$14164 ( \14834 , \13814 , \14833 );
or \U$14165 ( \14835 , \13717 , \13070 );
nand \U$14166 ( \14836 , \14834 , \14835 );
nor \U$14167 ( \14837 , \14832 , \14836 );
nand \U$14168 ( \14838 , \14828 , \14837 );
not \U$14169 ( \14839 , \14838 );
nand \U$14170 ( \14840 , \14825 , \14839 );
not \U$14171 ( \14841 , \14840 );
not \U$14172 ( \14842 , \13021 );
not \U$14173 ( \14843 , \13160 );
or \U$14174 ( \14844 , \14842 , \14843 );
and \U$14175 ( \14845 , \13267 , \13020 );
and \U$14176 ( \14846 , \12838 , \13169 );
not \U$14177 ( \14847 , \12838 );
and \U$14178 ( \14848 , \14847 , \13269 );
or \U$14179 ( \14849 , \14846 , \14848 );
nor \U$14180 ( \14850 , \14845 , \14849 );
nand \U$14181 ( \14851 , \14844 , \14850 );
not \U$14182 ( \14852 , \14851 );
or \U$14183 ( \14853 , \14841 , \14852 );
nand \U$14184 ( \14854 , \14838 , \14824 );
nand \U$14185 ( \14855 , \14853 , \14854 );
not \U$14186 ( \14856 , \14750 );
not \U$14187 ( \14857 , \14798 );
and \U$14188 ( \14858 , \14856 , \14857 );
and \U$14189 ( \14859 , \14750 , \14798 );
nor \U$14190 ( \14860 , \14858 , \14859 );
not \U$14191 ( \14861 , \14860 );
and \U$14192 ( \14862 , \14855 , \14861 );
nor \U$14193 ( \14863 , \14800 , \14862 );
xnor \U$14194 ( \14864 , \14588 , \14531 );
xor \U$14195 ( \14865 , \14863 , \14864 );
not \U$14196 ( \14866 , \14543 );
not \U$14197 ( \14867 , \14580 );
or \U$14198 ( \14868 , \14866 , \14867 );
or \U$14199 ( \14869 , \14580 , \14543 );
nand \U$14200 ( \14870 , \14868 , \14869 );
not \U$14201 ( \14871 , \14870 );
xnor \U$14202 ( \14872 , \14637 , \14670 );
nand \U$14203 ( \14873 , \14871 , \14872 );
not \U$14204 ( \14874 , \13770 );
not \U$14205 ( \14875 , \13232 );
or \U$14206 ( \14876 , \14874 , \14875 );
not \U$14207 ( \14877 , \13239 );
not \U$14208 ( \14878 , \14103 );
and \U$14209 ( \14879 , \14877 , \14878 );
and \U$14210 ( \14880 , \14653 , \13869 );
nor \U$14211 ( \14881 , \14879 , \14880 );
nand \U$14212 ( \14882 , \14876 , \14881 );
not \U$14213 ( \14883 , \14565 );
not \U$14214 ( \14884 , \14883 );
not \U$14215 ( \14885 , \14556 );
or \U$14216 ( \14886 , \14884 , \14885 );
or \U$14217 ( \14887 , \14556 , \14883 );
nand \U$14218 ( \14888 , \14886 , \14887 );
nand \U$14219 ( \14889 , \14882 , \14888 );
not \U$14220 ( \14890 , \14889 );
and \U$14221 ( \14891 , \12585 , \14455 );
not \U$14222 ( \14892 , \14634 );
not \U$14223 ( \14893 , \12581 );
or \U$14224 ( \14894 , \14892 , \14893 );
or \U$14225 ( \14895 , \12597 , \14517 );
nand \U$14226 ( \14896 , \14894 , \14895 );
nor \U$14227 ( \14897 , \14891 , \14896 );
not \U$14228 ( \14898 , \14897 );
or \U$14229 ( \14899 , \14890 , \14898 );
not \U$14230 ( \14900 , \14882 );
not \U$14231 ( \14901 , \14888 );
nand \U$14232 ( \14902 , \14900 , \14901 );
nand \U$14233 ( \14903 , \14899 , \14902 );
not \U$14234 ( \14904 , \14903 );
and \U$14235 ( \14905 , \14873 , \14904 );
nor \U$14236 ( \14906 , \14871 , \14872 );
nor \U$14237 ( \14907 , \14905 , \14906 );
and \U$14238 ( \14908 , \14865 , \14907 );
and \U$14239 ( \14909 , \14863 , \14864 );
or \U$14240 ( \14910 , \14908 , \14909 );
xor \U$14241 ( \14911 , \14740 , \14910 );
xor \U$14242 ( \14912 , \14472 , \14593 );
xor \U$14243 ( \14913 , \14912 , \14686 );
not \U$14244 ( \14914 , \14913 );
and \U$14245 ( \14915 , \14911 , \14914 );
and \U$14246 ( \14916 , \14740 , \14910 );
nor \U$14247 ( \14917 , \14915 , \14916 );
not \U$14248 ( \14918 , \14917 );
nand \U$14249 ( \14919 , \14727 , \14918 );
not \U$14250 ( \14920 , \14913 );
not \U$14251 ( \14921 , \14911 );
or \U$14252 ( \14922 , \14920 , \14921 );
or \U$14253 ( \14923 , \14911 , \14913 );
nand \U$14254 ( \14924 , \14922 , \14923 );
xor \U$14255 ( \14925 , \14863 , \14864 );
xor \U$14256 ( \14926 , \14925 , \14907 );
not \U$14257 ( \14927 , \14926 );
not \U$14258 ( \14928 , \14855 );
not \U$14259 ( \14929 , \14860 );
and \U$14260 ( \14930 , \14928 , \14929 );
and \U$14261 ( \14931 , \14855 , \14860 );
nor \U$14262 ( \14932 , \14930 , \14931 );
and \U$14263 ( \14933 , \14831 , \12838 );
not \U$14264 ( \14934 , \12910 );
not \U$14265 ( \14935 , \12970 );
not \U$14266 ( \14936 , \14935 );
or \U$14267 ( \14937 , \14934 , \14936 );
not \U$14268 ( \14938 , \12971 );
or \U$14269 ( \14939 , \13814 , \14938 );
nand \U$14270 ( \14940 , \14937 , \14939 );
nor \U$14271 ( \14941 , \14933 , \14940 );
nand \U$14272 ( \14942 , \12897 , \12839 );
nand \U$14273 ( \14943 , \14941 , \14942 );
not \U$14274 ( \14944 , \14943 );
or \U$14275 ( \14945 , \14805 , \13516 );
not \U$14276 ( \14946 , \14945 );
nand \U$14277 ( \14947 , \14946 , \12971 );
not \U$14278 ( \14948 , \14947 );
buf \U$14279 ( \14949 , \14806 );
and \U$14280 ( \14950 , \14949 , \14935 );
or \U$14281 ( \14951 , \14814 , \14833 );
not \U$14282 ( \14952 , \13069 );
nand \U$14283 ( \14953 , \14952 , \13781 );
nand \U$14284 ( \14954 , \14951 , \14953 );
nor \U$14285 ( \14955 , \14950 , \14954 );
not \U$14286 ( \14956 , \14955 );
or \U$14287 ( \14957 , \14948 , \14956 );
not \U$14288 ( \14958 , \14810 );
not \U$14289 ( \14959 , \14405 );
or \U$14290 ( \14960 , \14958 , \14959 );
nand \U$14291 ( \14961 , \13584 , \13226 );
nand \U$14292 ( \14962 , \14960 , \14961 );
not \U$14293 ( \14963 , \14404 );
and \U$14294 ( \14964 , \13225 , \13583 );
nor \U$14295 ( \14965 , \14964 , \13795 );
nor \U$14296 ( \14966 , \14963 , \14965 );
nor \U$14297 ( \14967 , \14962 , \14966 );
nand \U$14298 ( \14968 , \14957 , \14967 );
not \U$14299 ( \14969 , \14968 );
and \U$14300 ( \14970 , \14944 , \14969 );
and \U$14301 ( \14971 , \14943 , \14968 );
nor \U$14302 ( \14972 , \14970 , \14971 );
not \U$14303 ( \14973 , \14972 );
not \U$14304 ( \14974 , \13676 );
not \U$14305 ( \14975 , \13160 );
or \U$14306 ( \14976 , \14974 , \14975 );
not \U$14307 ( \14977 , \13842 );
and \U$14308 ( \14978 , \13267 , \14977 );
or \U$14309 ( \14979 , \13272 , \13021 );
nand \U$14310 ( \14980 , \13269 , \13021 );
nand \U$14311 ( \14981 , \14979 , \14980 );
nor \U$14312 ( \14982 , \14978 , \14981 );
nand \U$14313 ( \14983 , \14976 , \14982 );
nand \U$14314 ( \14984 , \14973 , \14983 );
not \U$14315 ( \14985 , \14941 );
not \U$14316 ( \14986 , \14942 );
or \U$14317 ( \14987 , \14985 , \14986 );
not \U$14318 ( \14988 , \14968 );
nand \U$14319 ( \14989 , \14987 , \14988 );
nand \U$14320 ( \14990 , \14984 , \14989 );
not \U$14321 ( \14991 , \14990 );
not \U$14322 ( \14992 , \14991 );
and \U$14323 ( \14993 , \12335 , RIaaa6d10_527);
and \U$14324 ( \14994 , \12339 , RIaaa6d88_528);
nor \U$14325 ( \14995 , \14993 , \14994 );
not \U$14326 ( \14996 , RIaaa6e00_529);
not \U$14327 ( \14997 , \14008 );
or \U$14328 ( \14998 , \14996 , \14997 );
not \U$14329 ( \14999 , RIaaa6a40_521);
not \U$14330 ( \15000 , \14488 );
not \U$14331 ( \15001 , \15000 );
or \U$14332 ( \15002 , \14999 , \15001 );
nor \U$14333 ( \15003 , \14485 , \14487 );
nand \U$14334 ( \15004 , \15003 , RIaaa6f68_532);
nand \U$14335 ( \15005 , \15002 , \15004 );
not \U$14336 ( \15006 , RIaaa69c8_520);
not \U$14337 ( \15007 , \12389 );
or \U$14338 ( \15008 , \15006 , \15007 );
and \U$14339 ( \15009 , \12410 , RIaaa7058_534);
nand \U$14340 ( \15010 , \11473 , RIaaa7148_536);
not \U$14341 ( \15011 , \15010 );
nor \U$14342 ( \15012 , \15009 , \15011 );
nand \U$14343 ( \15013 , \15008 , \15012 );
nor \U$14344 ( \15014 , \15005 , \15013 );
nand \U$14345 ( \15015 , \14998 , \15014 );
not \U$14346 ( \15016 , RIaaa6ef0_531);
not \U$14347 ( \15017 , \13032 );
or \U$14348 ( \15018 , \15016 , \15017 );
not \U$14349 ( \15019 , \13036 );
not \U$14350 ( \15020 , \8889 );
and \U$14351 ( \15021 , \15019 , \15020 );
and \U$14352 ( \15022 , \12833 , RIaaa70d0_535);
nor \U$14353 ( \15023 , \15021 , \15022 );
nand \U$14354 ( \15024 , \15018 , \15023 );
nor \U$14355 ( \15025 , \15015 , \15024 );
not \U$14356 ( \15026 , \12828 );
not \U$14357 ( \15027 , \4324 );
and \U$14358 ( \15028 , \15026 , \15027 );
and \U$14359 ( \15029 , \12327 , RIaaa6b30_523);
nor \U$14360 ( \15030 , \15028 , \15029 );
not \U$14361 ( \15031 , RIaaa6ba8_524);
not \U$14362 ( \15032 , \12344 );
or \U$14363 ( \15033 , \15031 , \15032 );
nand \U$14364 ( \15034 , \12532 , RIaaa6e78_530);
nand \U$14365 ( \15035 , \15033 , \15034 );
not \U$14366 ( \15036 , RIaaa6c20_525);
not \U$14367 ( \15037 , \12356 );
or \U$14368 ( \15038 , \15036 , \15037 );
nand \U$14369 ( \15039 , \14004 , RIaaa6ab8_522);
nand \U$14370 ( \15040 , \15038 , \15039 );
nor \U$14371 ( \15041 , \15035 , \15040 );
and \U$14372 ( \15042 , \14995 , \15025 , \15030 , \15041 );
buf \U$14373 ( \15043 , \15042 );
buf \U$14374 ( \15044 , \15043 );
not \U$14375 ( \15045 , \15044 );
and \U$14376 ( \15046 , \12841 , \15045 );
not \U$14377 ( \15047 , \15046 );
and \U$14378 ( \15048 , \14744 , \12677 );
not \U$14379 ( \15049 , \12251 );
not \U$14380 ( \15050 , \15049 );
nand \U$14381 ( \15051 , \15050 , \12668 , \14796 );
and \U$14382 ( \15052 , \12493 , \15051 );
not \U$14383 ( \15053 , \12493 );
not \U$14384 ( \15054 , \14796 );
nand \U$14385 ( \15055 , \15049 , \15054 );
or \U$14386 ( \15056 , \12668 , \15055 );
and \U$14387 ( \15057 , \15053 , \15056 );
nor \U$14388 ( \15058 , \15052 , \15057 );
nor \U$14389 ( \15059 , \15048 , \15058 );
not \U$14390 ( \15060 , \15059 );
or \U$14391 ( \15061 , \15047 , \15060 );
or \U$14392 ( \15062 , \15059 , \15046 );
nand \U$14393 ( \15063 , \15061 , \15062 );
not \U$14394 ( \15064 , \15063 );
not \U$14395 ( \15065 , \15064 );
and \U$14396 ( \15066 , \14992 , \15065 );
not \U$14397 ( \15067 , \15059 );
and \U$14398 ( \15068 , \15067 , \15046 );
nor \U$14399 ( \15069 , \15066 , \15068 );
xor \U$14400 ( \15070 , \14932 , \15069 );
not \U$14401 ( \15071 , \14818 );
not \U$14402 ( \15072 , \14823 );
not \U$14403 ( \15073 , \15072 );
and \U$14404 ( \15074 , \15071 , \15073 );
and \U$14405 ( \15075 , \14818 , \15072 );
nor \U$14406 ( \15076 , \15074 , \15075 );
not \U$14407 ( \15077 , \14044 );
not \U$14408 ( \15078 , \15077 );
not \U$14409 ( \15079 , \13235 );
or \U$14410 ( \15080 , \15078 , \15079 );
or \U$14411 ( \15081 , \13235 , \15077 );
nand \U$14412 ( \15082 , \15080 , \15081 );
not \U$14413 ( \15083 , \15082 );
not \U$14414 ( \15084 , \12780 );
or \U$14415 ( \15085 , \15083 , \15084 );
and \U$14416 ( \15086 , \14660 , \14103 );
nor \U$14417 ( \15087 , \13430 , \14103 );
nor \U$14418 ( \15088 , \15086 , \15087 );
nand \U$14419 ( \15089 , \15085 , \15088 );
not \U$14420 ( \15090 , \15089 );
xor \U$14421 ( \15091 , \15076 , \15090 );
not \U$14422 ( \15092 , \14517 );
not \U$14423 ( \15093 , \13286 );
or \U$14424 ( \15094 , \15092 , \15093 );
not \U$14425 ( \15095 , \14513 );
not \U$14426 ( \15096 , \15095 );
not \U$14427 ( \15097 , \15096 );
not \U$14428 ( \15098 , \13890 );
or \U$14429 ( \15099 , \15097 , \15098 );
not \U$14430 ( \15100 , \14513 );
not \U$14431 ( \15101 , \15100 );
or \U$14432 ( \15102 , \12669 , \15101 );
nand \U$14433 ( \15103 , \15099 , \15102 );
nand \U$14434 ( \15104 , \13884 , \15103 );
nand \U$14435 ( \15105 , \15094 , \15104 );
not \U$14436 ( \15106 , \12600 );
nor \U$14437 ( \15107 , \15106 , \14455 );
nor \U$14438 ( \15108 , \15105 , \15107 );
and \U$14439 ( \15109 , \15091 , \15108 );
and \U$14440 ( \15110 , \15076 , \15090 );
or \U$14441 ( \15111 , \15109 , \15110 );
xor \U$14442 ( \15112 , \14824 , \14838 );
xnor \U$14443 ( \15113 , \15112 , \14851 );
nand \U$14444 ( \15114 , \15111 , \15113 );
not \U$14445 ( \15115 , \14897 );
xor \U$14446 ( \15116 , \14882 , \14888 );
not \U$14447 ( \15117 , \15116 );
or \U$14448 ( \15118 , \15115 , \15117 );
buf \U$14449 ( \15119 , \14897 );
or \U$14450 ( \15120 , \15119 , \15116 );
nand \U$14451 ( \15121 , \15118 , \15120 );
and \U$14452 ( \15122 , \15114 , \15121 );
nor \U$14453 ( \15123 , \15111 , \15113 );
nor \U$14454 ( \15124 , \15122 , \15123 );
and \U$14455 ( \15125 , \15070 , \15124 );
and \U$14456 ( \15126 , \14932 , \15069 );
or \U$14457 ( \15127 , \15125 , \15126 );
not \U$14458 ( \15128 , \15127 );
xnor \U$14459 ( \15129 , \14683 , \14674 );
buf \U$14460 ( \15130 , \14624 );
and \U$14461 ( \15131 , \15129 , \15130 );
not \U$14462 ( \15132 , \15129 );
not \U$14463 ( \15133 , \15130 );
and \U$14464 ( \15134 , \15132 , \15133 );
nor \U$14465 ( \15135 , \15131 , \15134 );
not \U$14466 ( \15136 , \15135 );
and \U$14467 ( \15137 , \15128 , \15136 );
and \U$14468 ( \15138 , \15127 , \15135 );
nor \U$14469 ( \15139 , \15137 , \15138 );
not \U$14470 ( \15140 , \15139 );
not \U$14471 ( \15141 , \15140 );
or \U$14472 ( \15142 , \14927 , \15141 );
not \U$14473 ( \15143 , \15135 );
nand \U$14474 ( \15144 , \15143 , \15127 );
nand \U$14475 ( \15145 , \15142 , \15144 );
nand \U$14476 ( \15146 , \14924 , \15145 );
nand \U$14477 ( \15147 , \14919 , \15146 );
xor \U$14478 ( \15148 , \14373 , \14689 );
and \U$14479 ( \15149 , \15148 , \14725 );
and \U$14480 ( \15150 , \14373 , \14689 );
or \U$14481 ( \15151 , \15149 , \15150 );
not \U$14482 ( \15152 , \15151 );
not \U$14483 ( \15153 , \13910 );
not \U$14484 ( \15154 , \13903 );
or \U$14485 ( \15155 , \15153 , \15154 );
nand \U$14486 ( \15156 , \13901 , \13909 );
nand \U$14487 ( \15157 , \15155 , \15156 );
and \U$14488 ( \15158 , \15157 , \13854 );
not \U$14489 ( \15159 , \15157 );
and \U$14490 ( \15160 , \15159 , \13853 );
nor \U$14491 ( \15161 , \15158 , \15160 );
not \U$14492 ( \15162 , \14705 );
not \U$14493 ( \15163 , \14720 );
or \U$14494 ( \15164 , \15162 , \15163 );
nand \U$14495 ( \15165 , \15164 , \14707 );
nor \U$14496 ( \15166 , \15161 , \15165 );
not \U$14497 ( \15167 , \15166 );
nand \U$14498 ( \15168 , \15165 , \15161 );
xor \U$14499 ( \15169 , \13996 , \14112 );
xor \U$14500 ( \15170 , \15169 , \14166 );
nand \U$14501 ( \15171 , \15167 , \15168 , \15170 );
not \U$14502 ( \15172 , \15170 );
not \U$14503 ( \15173 , \15166 );
nand \U$14504 ( \15174 , \15173 , \15168 );
nand \U$14505 ( \15175 , \15172 , \15174 );
nand \U$14506 ( \15176 , \15171 , \15175 );
nand \U$14507 ( \15177 , \15152 , \15176 );
not \U$14508 ( \15178 , \15170 );
not \U$14509 ( \15179 , \15174 );
or \U$14510 ( \15180 , \15178 , \15179 );
not \U$14511 ( \15181 , \15161 );
nand \U$14512 ( \15182 , \15181 , \15165 );
nand \U$14513 ( \15183 , \15180 , \15182 );
xor \U$14514 ( \15184 , \13986 , \14169 );
xor \U$14515 ( \15185 , \15184 , \14182 );
nand \U$14516 ( \15186 , \15183 , \15185 );
nand \U$14517 ( \15187 , \15177 , \15186 );
nor \U$14518 ( \15188 , \15147 , \15187 );
not \U$14519 ( \15189 , \15188 );
xor \U$14520 ( \15190 , \15113 , \15111 );
xnor \U$14521 ( \15191 , \15190 , \15121 );
not \U$14522 ( \15192 , \15044 );
not \U$14523 ( \15193 , \12279 );
or \U$14524 ( \15194 , \15192 , \15193 );
and \U$14525 ( \15195 , \14796 , \12277 );
not \U$14526 ( \15196 , \14796 );
and \U$14527 ( \15197 , \15196 , \12276 );
nor \U$14528 ( \15198 , \15195 , \15197 );
not \U$14529 ( \15199 , \15198 );
not \U$14530 ( \15200 , \12678 );
and \U$14531 ( \15201 , \15199 , \15200 );
not \U$14532 ( \15202 , \12431 );
and \U$14533 ( \15203 , \15202 , \15045 );
nor \U$14534 ( \15204 , \15201 , \15203 );
nand \U$14535 ( \15205 , \15194 , \15204 );
and \U$14536 ( \15206 , \12904 , \14661 );
and \U$14537 ( \15207 , \12838 , \12912 );
not \U$14538 ( \15208 , \12838 );
and \U$14539 ( \15209 , \15208 , \13520 );
nor \U$14540 ( \15210 , \15207 , \15209 );
nor \U$14541 ( \15211 , \15206 , \15210 );
nand \U$14542 ( \15212 , \12898 , \13021 );
nand \U$14543 ( \15213 , \15211 , \15212 );
not \U$14544 ( \15214 , \15213 );
not \U$14545 ( \15215 , \13770 );
not \U$14546 ( \15216 , \13160 );
or \U$14547 ( \15217 , \15215 , \15216 );
and \U$14548 ( \15218 , \14085 , \13771 );
and \U$14549 ( \15219 , \13676 , \13704 );
not \U$14550 ( \15220 , \13676 );
and \U$14551 ( \15221 , \15220 , \13169 );
or \U$14552 ( \15222 , \15219 , \15221 );
nor \U$14553 ( \15223 , \15218 , \15222 );
nand \U$14554 ( \15224 , \15217 , \15223 );
not \U$14555 ( \15225 , \15224 );
or \U$14556 ( \15226 , \15214 , \15225 );
and \U$14557 ( \15227 , \13999 , RIaaa7760_549);
and \U$14558 ( \15228 , \12818 , RIaaa75f8_546);
nor \U$14559 ( \15229 , \15227 , \15228 );
and \U$14560 ( \15230 , \13032 , RIaaa78c8_552);
not \U$14561 ( \15231 , RIaaa7580_545);
not \U$14562 ( \15232 , \14489 );
or \U$14563 ( \15233 , \15231 , \15232 );
nand \U$14564 ( \15234 , RIaaa7490_543, \12476 );
nand \U$14565 ( \15235 , \15233 , \15234 );
nor \U$14566 ( \15236 , \15230 , \15235 );
and \U$14567 ( \15237 , \14008 , RIaaa7850_551);
not \U$14568 ( \15238 , \13036 );
nand \U$14569 ( \15239 , \15238 , RIaaa7238_538);
nand \U$14570 ( \15240 , \15003 , RIaaa7940_553);
and \U$14571 ( \15241 , \12410 , RIaaa72b0_539);
nand \U$14572 ( \15242 , \11473 , RIaaa71c0_537);
not \U$14573 ( \15243 , \15242 );
nor \U$14574 ( \15244 , \15241 , \15243 );
nand \U$14575 ( \15245 , \15239 , \15240 , \15244 );
nor \U$14576 ( \15246 , \15237 , \15245 );
nand \U$14577 ( \15247 , \15229 , \15236 , \15246 );
not \U$14578 ( \15248 , \15247 );
nand \U$14579 ( \15249 , \12339 , RIaaa77d8_550);
nand \U$14580 ( \15250 , \12344 , RIaaa7418_542);
nand \U$14581 ( \15251 , \12829 , RIaaa76e8_548);
nand \U$14582 ( \15252 , \15249 , \15250 , \15251 );
nand \U$14583 ( \15253 , \12356 , RIaaa73a0_541);
nand \U$14584 ( \15254 , \12532 , RIaaa7508_544);
nand \U$14585 ( \15255 , \12833 , RIaaa7328_540);
nand \U$14586 ( \15256 , \14004 , RIaaa7670_547);
nand \U$14587 ( \15257 , \15253 , \15254 , \15255 , \15256 );
nor \U$14588 ( \15258 , \15252 , \15257 );
nand \U$14589 ( \15259 , \15248 , \15258 );
not \U$14590 ( \15260 , \15259 );
buf \U$14591 ( \15261 , \15260 );
not \U$14592 ( \15262 , \15261 );
nand \U$14593 ( \15263 , \12606 , \15262 );
nand \U$14594 ( \15264 , \15226 , \15263 );
xor \U$14595 ( \15265 , \15205 , \15264 );
not \U$14596 ( \15266 , \15265 );
not \U$14597 ( \15267 , \15266 );
xor \U$14598 ( \15268 , \15076 , \15090 );
xor \U$14599 ( \15269 , \15268 , \15108 );
not \U$14600 ( \15270 , \15269 );
not \U$14601 ( \15271 , \15270 );
or \U$14602 ( \15272 , \15267 , \15271 );
nand \U$14603 ( \15273 , \15269 , \15265 );
nand \U$14604 ( \15274 , \15272 , \15273 );
not \U$14605 ( \15275 , \15274 );
not \U$14606 ( \15276 , \15261 );
not \U$14607 ( \15277 , \12279 );
or \U$14608 ( \15278 , \15276 , \15277 );
and \U$14609 ( \15279 , \12430 , \15262 );
and \U$14610 ( \15280 , \12275 , \15279 );
and \U$14611 ( \15281 , \15044 , \12435 );
not \U$14612 ( \15282 , \15044 );
and \U$14613 ( \15283 , \15282 , \12495 );
nor \U$14614 ( \15284 , \15281 , \15283 );
nor \U$14615 ( \15285 , \15280 , \15284 );
nand \U$14616 ( \15286 , \15278 , \15285 );
and \U$14617 ( \15287 , \13559 , \12838 );
or \U$14618 ( \15288 , \13572 , \12970 );
or \U$14619 ( \15289 , \14935 , \13566 );
nand \U$14620 ( \15290 , \15288 , \15289 );
nor \U$14621 ( \15291 , \15287 , \15290 );
nand \U$14622 ( \15292 , \12839 , \13578 );
nand \U$14623 ( \15293 , \14060 , \13121 );
not \U$14624 ( \15294 , \13121 );
nand \U$14625 ( \15295 , \15294 , \14401 );
nand \U$14626 ( \15296 , \14405 , \13071 );
and \U$14627 ( \15297 , \15293 , \15295 , \15296 );
nand \U$14628 ( \15298 , \15291 , \15292 , \15297 );
not \U$14629 ( \15299 , \15298 );
and \U$14630 ( \15300 , \14977 , \12904 );
not \U$14631 ( \15301 , \12911 );
not \U$14632 ( \15302 , \13020 );
or \U$14633 ( \15303 , \15301 , \15302 );
or \U$14634 ( \15304 , \14661 , \13520 );
nand \U$14635 ( \15305 , \15303 , \15304 );
nor \U$14636 ( \15306 , \15300 , \15305 );
nand \U$14637 ( \15307 , \12898 , \13676 );
nand \U$14638 ( \15308 , \15306 , \15307 );
not \U$14639 ( \15309 , \15308 );
or \U$14640 ( \15310 , \15299 , \15309 );
not \U$14641 ( \15311 , \13997 );
nand \U$14642 ( \15312 , \12335 , RIaaa8750_583);
nand \U$14643 ( \15313 , \12502 , RIaaa85e8_580);
nand \U$14644 ( \15314 , \12339 , RIaaa87c8_584);
nand \U$14645 ( \15315 , \12351 , RIaaa86d8_582);
nand \U$14646 ( \15316 , \15312 , \15313 , \15314 , \15315 );
and \U$14647 ( \15317 , \12453 , RIaaa8480_577);
and \U$14648 ( \15318 , \12455 , RIaaa8660_581);
nor \U$14649 ( \15319 , \15317 , \15318 );
and \U$14650 ( \15320 , \12356 , RIaaa8390_575);
and \U$14651 ( \15321 , \12360 , RIaaa84f8_578);
nor \U$14652 ( \15322 , \15320 , \15321 );
nand \U$14653 ( \15323 , \15319 , \15322 );
nor \U$14654 ( \15324 , \15316 , \15323 );
not \U$14655 ( \15325 , RIaaa8840_585);
not \U$14656 ( \15326 , \12375 );
or \U$14657 ( \15327 , \15325 , \15326 );
nand \U$14658 ( \15328 , \12380 , RIaaa88b8_586);
nand \U$14659 ( \15329 , \15327 , \15328 );
and \U$14660 ( \15330 , \12513 , RIaaa8930_587);
not \U$14661 ( \15331 , RIaaa8228_572);
nor \U$14662 ( \15332 , \15331 , \12396 );
nor \U$14663 ( \15333 , \15330 , \15332 );
nand \U$14664 ( \15334 , \12365 , RIaaa8318_574);
and \U$14665 ( \15335 , \12476 , RIaaa8408_576);
not \U$14666 ( \15336 , RIaaa82a0_573);
not \U$14667 ( \15337 , \12410 );
or \U$14668 ( \15338 , \15336 , \15337 );
nand \U$14669 ( \15339 , \11473 , RIaaa81b0_571);
nand \U$14670 ( \15340 , \15338 , \15339 );
nor \U$14671 ( \15341 , \15335 , \15340 );
nand \U$14672 ( \15342 , \12418 , RIaaa8570_579);
nand \U$14673 ( \15343 , \15333 , \15334 , \15341 , \15342 );
nor \U$14674 ( \15344 , \15329 , \15343 );
nand \U$14675 ( \15345 , \15324 , \15344 );
buf \U$14676 ( \15346 , \15345 );
not \U$14677 ( \15347 , \15346 );
not \U$14678 ( \15348 , \15347 );
and \U$14679 ( \15349 , \15311 , \15348 );
nand \U$14680 ( \15350 , \15291 , \15292 );
not \U$14681 ( \15351 , \15297 );
and \U$14682 ( \15352 , \15350 , \15351 );
nor \U$14683 ( \15353 , \15349 , \15352 );
nand \U$14684 ( \15354 , \15310 , \15353 );
nand \U$14685 ( \15355 , \15286 , \15354 );
not \U$14686 ( \15356 , \15355 );
not \U$14687 ( \15357 , \14983 );
and \U$14688 ( \15358 , \14972 , \15357 );
not \U$14689 ( \15359 , \14972 );
and \U$14690 ( \15360 , \15359 , \14983 );
nor \U$14691 ( \15361 , \15358 , \15360 );
not \U$14692 ( \15362 , \15361 );
not \U$14693 ( \15363 , \15362 );
not \U$14694 ( \15364 , \14797 );
not \U$14695 ( \15365 , \12585 );
or \U$14696 ( \15366 , \15364 , \15365 );
not \U$14697 ( \15367 , \12597 );
not \U$14698 ( \15368 , \14797 );
and \U$14699 ( \15369 , \15367 , \15368 );
and \U$14700 ( \15370 , \14120 , \15103 );
nor \U$14701 ( \15371 , \15369 , \15370 );
nand \U$14702 ( \15372 , \15366 , \15371 );
and \U$14703 ( \15373 , \14955 , \14947 );
not \U$14704 ( \15374 , \14967 );
and \U$14705 ( \15375 , \15373 , \15374 );
not \U$14706 ( \15376 , \15373 );
and \U$14707 ( \15377 , \15376 , \14967 );
nor \U$14708 ( \15378 , \15375 , \15377 );
not \U$14709 ( \15379 , \14517 );
not \U$14710 ( \15380 , \13235 );
or \U$14711 ( \15381 , \15379 , \15380 );
or \U$14712 ( \15382 , \12783 , \14517 );
nand \U$14713 ( \15383 , \15381 , \15382 );
not \U$14714 ( \15384 , \15383 );
not \U$14715 ( \15385 , \12780 );
or \U$14716 ( \15386 , \15384 , \15385 );
not \U$14717 ( \15387 , \12769 );
nand \U$14718 ( \15388 , \15387 , \15082 );
nand \U$14719 ( \15389 , \15386 , \15388 );
xor \U$14720 ( \15390 , \15378 , \15389 );
and \U$14721 ( \15391 , \15372 , \15390 );
and \U$14722 ( \15392 , \15378 , \15389 );
nor \U$14723 ( \15393 , \15391 , \15392 );
not \U$14724 ( \15394 , \15393 );
not \U$14725 ( \15395 , \15394 );
or \U$14726 ( \15396 , \15363 , \15395 );
nand \U$14727 ( \15397 , \15393 , \15361 );
nand \U$14728 ( \15398 , \15396 , \15397 );
not \U$14729 ( \15399 , \15398 );
or \U$14730 ( \15400 , \15356 , \15399 );
or \U$14731 ( \15401 , \15355 , \15398 );
nand \U$14732 ( \15402 , \15400 , \15401 );
not \U$14733 ( \15403 , \15402 );
or \U$14734 ( \15404 , \15275 , \15403 );
nand \U$14735 ( \15405 , \15270 , \15265 );
nand \U$14736 ( \15406 , \15404 , \15405 );
not \U$14737 ( \15407 , \15406 );
xor \U$14738 ( \15408 , \15191 , \15407 );
and \U$14739 ( \15409 , \15205 , \15264 );
and \U$14740 ( \15410 , \14984 , \14989 );
nor \U$14741 ( \15411 , \15410 , \15063 );
not \U$14742 ( \15412 , \15411 );
or \U$14743 ( \15413 , \14972 , \15357 );
nand \U$14744 ( \15414 , \15413 , \15063 , \14989 );
nand \U$14745 ( \15415 , \15412 , \15414 );
xor \U$14746 ( \15416 , \15409 , \15415 );
not \U$14747 ( \15417 , \15355 );
or \U$14748 ( \15418 , \15361 , \15417 );
nand \U$14749 ( \15419 , \15418 , \15394 );
nand \U$14750 ( \15420 , \15417 , \15361 );
nand \U$14751 ( \15421 , \15419 , \15420 );
xnor \U$14752 ( \15422 , \15416 , \15421 );
xor \U$14753 ( \15423 , \15408 , \15422 );
xor \U$14754 ( \15424 , \15372 , \15390 );
not \U$14755 ( \15425 , \15424 );
nor \U$14756 ( \15426 , \15286 , \15354 );
not \U$14757 ( \15427 , \15426 );
nand \U$14758 ( \15428 , \15427 , \15355 );
nand \U$14759 ( \15429 , \15425 , \15428 );
not \U$14760 ( \15430 , \15429 );
xor \U$14761 ( \15431 , \15350 , \15297 );
xnor \U$14762 ( \15432 , \15308 , \15431 );
not \U$14763 ( \15433 , \15262 );
not \U$14764 ( \15434 , \12585 );
or \U$14765 ( \15435 , \15433 , \15434 );
not \U$14766 ( \15436 , \12597 );
not \U$14767 ( \15437 , \15262 );
and \U$14768 ( \15438 , \15436 , \15437 );
not \U$14769 ( \15439 , \15045 );
not \U$14770 ( \15440 , \12583 );
or \U$14771 ( \15441 , \15439 , \15440 );
not \U$14772 ( \15442 , \15044 );
or \U$14773 ( \15443 , \13080 , \15442 );
nand \U$14774 ( \15444 , \15441 , \15443 );
and \U$14775 ( \15445 , \14120 , \15444 );
nor \U$14776 ( \15446 , \15438 , \15445 );
nand \U$14777 ( \15447 , \15435 , \15446 );
not \U$14778 ( \15448 , \15447 );
not \U$14779 ( \15449 , \13019 );
not \U$14780 ( \15450 , \13578 );
or \U$14781 ( \15451 , \15449 , \15450 );
and \U$14782 ( \15452 , \14949 , \13885 );
not \U$14783 ( \15453 , \14054 );
not \U$14784 ( \15454 , \12837 );
or \U$14785 ( \15455 , \15453 , \15454 );
or \U$14786 ( \15456 , \13566 , \12838 );
nand \U$14787 ( \15457 , \15455 , \15456 );
nor \U$14788 ( \15458 , \15452 , \15457 );
nand \U$14789 ( \15459 , \15451 , \15458 );
not \U$14790 ( \15460 , \15459 );
not \U$14791 ( \15461 , \14404 );
not \U$14792 ( \15462 , \12971 );
and \U$14793 ( \15463 , \15461 , \15462 );
and \U$14794 ( \15464 , \14833 , \13804 );
not \U$14795 ( \15465 , \14833 );
and \U$14796 ( \15466 , \15465 , \14067 );
nor \U$14797 ( \15467 , \15464 , \15466 );
nor \U$14798 ( \15468 , \15463 , \15467 );
not \U$14799 ( \15469 , \15468 );
and \U$14800 ( \15470 , \15460 , \15469 );
and \U$14801 ( \15471 , \15459 , \15468 );
nor \U$14802 ( \15472 , \15470 , \15471 );
not \U$14803 ( \15473 , \15472 );
not \U$14804 ( \15474 , \15054 );
not \U$14805 ( \15475 , \12844 );
or \U$14806 ( \15476 , \15474 , \15475 );
or \U$14807 ( \15477 , \13235 , \15054 );
nand \U$14808 ( \15478 , \15476 , \15477 );
not \U$14809 ( \15479 , \15478 );
not \U$14810 ( \15480 , \12780 );
or \U$14811 ( \15481 , \15479 , \15480 );
not \U$14812 ( \15482 , \15095 );
not \U$14813 ( \15483 , \13235 );
or \U$14814 ( \15484 , \15482 , \15483 );
or \U$14815 ( \15485 , \12783 , \14514 );
nand \U$14816 ( \15486 , \15484 , \15485 );
nand \U$14817 ( \15487 , \15486 , \13245 );
nand \U$14818 ( \15488 , \15481 , \15487 );
not \U$14819 ( \15489 , \15488 );
or \U$14820 ( \15490 , \15473 , \15489 );
or \U$14821 ( \15491 , \15488 , \15472 );
nand \U$14822 ( \15492 , \15490 , \15491 );
not \U$14823 ( \15493 , \15492 );
or \U$14824 ( \15494 , \15448 , \15493 );
not \U$14825 ( \15495 , \15472 );
nand \U$14826 ( \15496 , \15495 , \15488 );
nand \U$14827 ( \15497 , \15494 , \15496 );
xor \U$14828 ( \15498 , \15432 , \15497 );
not \U$14829 ( \15499 , \14455 );
not \U$14830 ( \15500 , \13160 );
or \U$14831 ( \15501 , \15499 , \15500 );
and \U$14832 ( \15502 , \13533 , \14454 );
not \U$14833 ( \15503 , \14045 );
or \U$14834 ( \15504 , \13701 , \15503 );
nand \U$14835 ( \15505 , \13269 , \15503 );
nand \U$14836 ( \15506 , \15504 , \15505 );
nor \U$14837 ( \15507 , \15502 , \15506 );
nand \U$14838 ( \15508 , \15501 , \15507 );
not \U$14839 ( \15509 , \15508 );
not \U$14840 ( \15510 , \14103 );
not \U$14841 ( \15511 , \13525 );
or \U$14842 ( \15512 , \15510 , \15511 );
and \U$14843 ( \15513 , \13714 , \14102 );
or \U$14844 ( \15514 , \13520 , \13841 );
nand \U$14845 ( \15515 , \13718 , \13841 );
nand \U$14846 ( \15516 , \15514 , \15515 );
nor \U$14847 ( \15517 , \15513 , \15516 );
nand \U$14848 ( \15518 , \15512 , \15517 );
not \U$14849 ( \15519 , \15518 );
not \U$14850 ( \15520 , \15049 );
nand \U$14851 ( \15521 , \15520 , \12668 );
nand \U$14852 ( \15522 , \12339 , RIaaa80c0_569);
not \U$14853 ( \15523 , \12832 );
nand \U$14854 ( \15524 , \15523 , RIaaa7df0_563);
nand \U$14855 ( \15525 , \14004 , RIaaa7a30_555);
nand \U$14856 ( \15526 , \15522 , \15524 , \15525 );
and \U$14857 ( \15527 , \13999 , RIaaa7fd0_567);
not \U$14858 ( \15528 , RIaaa8138_570);
nor \U$14859 ( \15529 , \12373 , \15528 );
nor \U$14860 ( \15530 , \15527 , \15529 );
and \U$14861 ( \15531 , \12818 , RIaaa79b8_554);
not \U$14862 ( \15532 , RIaaa7c88_560);
not \U$14863 ( \15533 , \15003 );
or \U$14864 ( \15534 , \15532 , \15533 );
nand \U$14865 ( \15535 , \12389 , RIaaa7aa8_556);
nand \U$14866 ( \15536 , \15534 , \15535 );
nor \U$14867 ( \15537 , \15531 , \15536 );
nand \U$14868 ( \15538 , \15530 , \15537 );
nor \U$14869 ( \15539 , \15526 , \15538 );
and \U$14870 ( \15540 , \12532 , RIaaa8048_568);
not \U$14871 ( \15541 , RIaaa7d78_562);
not \U$14872 ( \15542 , \15238 );
or \U$14873 ( \15543 , \15541 , \15542 );
and \U$14874 ( \15544 , \12410 , RIaaa7e68_564);
nand \U$14875 ( \15545 , \11473 , RIaaa7ee0_565);
not \U$14876 ( \15546 , \15545 );
nor \U$14877 ( \15547 , \15544 , \15546 );
nand \U$14878 ( \15548 , \15543 , \15547 );
nor \U$14879 ( \15549 , \15540 , \15548 );
nand \U$14880 ( \15550 , \13032 , RIaaa7d00_561);
nand \U$14881 ( \15551 , \12344 , RIaaa7c10_559);
nand \U$14882 ( \15552 , \15549 , \15550 , \15551 );
not \U$14883 ( \15553 , RIaaa7f58_566);
not \U$14884 ( \15554 , \12829 );
or \U$14885 ( \15555 , \15553 , \15554 );
not \U$14886 ( \15556 , \14488 );
not \U$14887 ( \15557 , \4774 );
and \U$14888 ( \15558 , \15556 , \15557 );
and \U$14889 ( \15559 , \12356 , RIaaa7b98_558);
nor \U$14890 ( \15560 , \15558 , \15559 );
nand \U$14891 ( \15561 , \15555 , \15560 );
nor \U$14892 ( \15562 , \15552 , \15561 );
nand \U$14893 ( \15563 , \15539 , \15562 );
not \U$14894 ( \15564 , \15563 );
not \U$14895 ( \15565 , \15564 );
buf \U$14896 ( \15566 , \15565 );
not \U$14897 ( \15567 , \15566 );
not \U$14898 ( \15568 , \15567 );
and \U$14899 ( \15569 , \15521 , \15568 );
not \U$14900 ( \15570 , \15049 );
nor \U$14901 ( \15571 , \12583 , \15570 );
nor \U$14902 ( \15572 , \15569 , \15571 );
nand \U$14903 ( \15573 , \12682 , \15572 );
not \U$14904 ( \15574 , \15573 );
and \U$14905 ( \15575 , \15519 , \15574 );
and \U$14906 ( \15576 , \15573 , \15518 );
nor \U$14907 ( \15577 , \15575 , \15576 );
or \U$14908 ( \15578 , \15509 , \15577 );
not \U$14909 ( \15579 , \15573 );
nand \U$14910 ( \15580 , \15579 , \15518 );
nand \U$14911 ( \15581 , \15578 , \15580 );
and \U$14912 ( \15582 , \15498 , \15581 );
and \U$14913 ( \15583 , \15432 , \15497 );
or \U$14914 ( \15584 , \15582 , \15583 );
not \U$14915 ( \15585 , \15584 );
or \U$14916 ( \15586 , \15430 , \15585 );
not \U$14917 ( \15587 , \15417 );
not \U$14918 ( \15588 , \15426 );
nand \U$14919 ( \15589 , \15587 , \15424 , \15588 );
nand \U$14920 ( \15590 , \15586 , \15589 );
not \U$14921 ( \15591 , \15590 );
not \U$14922 ( \15592 , \15345 );
and \U$14923 ( \15593 , \12279 , \15592 );
not \U$14924 ( \15594 , \15279 );
or \U$14925 ( \15595 , \15594 , \12678 );
nand \U$14926 ( \15596 , \12682 , \12677 , \15261 );
nor \U$14927 ( \15597 , \15570 , \15592 );
nand \U$14928 ( \15598 , \12430 , \12678 , \15597 );
nand \U$14929 ( \15599 , \15595 , \15596 , \15598 );
nor \U$14930 ( \15600 , \15593 , \15599 );
not \U$14931 ( \15601 , \15600 );
not \U$14932 ( \15602 , \15601 );
not \U$14933 ( \15603 , \15486 );
not \U$14934 ( \15604 , \12780 );
or \U$14935 ( \15605 , \15603 , \15604 );
nand \U$14936 ( \15606 , \15383 , \13869 );
nand \U$14937 ( \15607 , \15605 , \15606 );
not \U$14938 ( \15608 , \15607 );
not \U$14939 ( \15609 , \15106 );
not \U$14940 ( \15610 , \15054 );
and \U$14941 ( \15611 , \15609 , \15610 );
not \U$14942 ( \15612 , \15054 );
not \U$14943 ( \15613 , \13286 );
or \U$14944 ( \15614 , \15612 , \15613 );
nand \U$14945 ( \15615 , \13884 , \15444 );
nand \U$14946 ( \15616 , \15614 , \15615 );
nor \U$14947 ( \15617 , \15611 , \15616 );
not \U$14948 ( \15618 , \15617 );
or \U$14949 ( \15619 , \15608 , \15618 );
or \U$14950 ( \15620 , \15617 , \15607 );
nand \U$14951 ( \15621 , \15619 , \15620 );
not \U$14952 ( \15622 , \15621 );
or \U$14953 ( \15623 , \15602 , \15622 );
not \U$14954 ( \15624 , \15617 );
nand \U$14955 ( \15625 , \15624 , \15607 );
nand \U$14956 ( \15626 , \15623 , \15625 );
not \U$14957 ( \15627 , \15626 );
not \U$14958 ( \15628 , \15503 );
not \U$14959 ( \15629 , \13160 );
or \U$14960 ( \15630 , \15628 , \15629 );
and \U$14961 ( \15631 , \14085 , \14045 );
and \U$14962 ( \15632 , \14102 , \13169 );
not \U$14963 ( \15633 , \14102 );
and \U$14964 ( \15634 , \15633 , \13704 );
or \U$14965 ( \15635 , \15632 , \15634 );
nor \U$14966 ( \15636 , \15631 , \15635 );
nand \U$14967 ( \15637 , \15630 , \15636 );
not \U$14968 ( \15638 , \15565 );
buf \U$14969 ( \15639 , \15638 );
not \U$14970 ( \15640 , \15639 );
and \U$14971 ( \15641 , \12841 , \15640 );
or \U$14972 ( \15642 , \15637 , \15641 );
not \U$14973 ( \15643 , \15459 );
nor \U$14974 ( \15644 , \15643 , \15468 );
nand \U$14975 ( \15645 , \15642 , \15644 );
not \U$14976 ( \15646 , \15213 );
not \U$14977 ( \15647 , \15224 );
not \U$14978 ( \15648 , \15647 );
or \U$14979 ( \15649 , \15646 , \15648 );
not \U$14980 ( \15650 , \15213 );
nand \U$14981 ( \15651 , \15650 , \15224 );
nand \U$14982 ( \15652 , \15649 , \15651 );
xor \U$14983 ( \15653 , \15645 , \15652 );
not \U$14984 ( \15654 , \15653 );
not \U$14985 ( \15655 , \15654 );
or \U$14986 ( \15656 , \15627 , \15655 );
not \U$14987 ( \15657 , \15645 );
nand \U$14988 ( \15658 , \15657 , \15652 );
nand \U$14989 ( \15659 , \15656 , \15658 );
not \U$14990 ( \15660 , \15659 );
nand \U$14991 ( \15661 , \15591 , \15660 );
not \U$14992 ( \15662 , \15661 );
xnor \U$14993 ( \15663 , \15274 , \15402 );
not \U$14994 ( \15664 , \15663 );
not \U$14995 ( \15665 , \15664 );
or \U$14996 ( \15666 , \15662 , \15665 );
or \U$14997 ( \15667 , \15591 , \15660 );
nand \U$14998 ( \15668 , \15666 , \15667 );
not \U$14999 ( \15669 , \15668 );
nand \U$15000 ( \15670 , \15423 , \15669 );
or \U$15001 ( \15671 , \15423 , \15669 );
not \U$15002 ( \15672 , \15584 );
not \U$15003 ( \15673 , \15428 );
not \U$15004 ( \15674 , \15424 );
and \U$15005 ( \15675 , \15673 , \15674 );
and \U$15006 ( \15676 , \15428 , \15424 );
nor \U$15007 ( \15677 , \15675 , \15676 );
not \U$15008 ( \15678 , \15677 );
and \U$15009 ( \15679 , \15672 , \15678 );
and \U$15010 ( \15680 , \15584 , \15677 );
nor \U$15011 ( \15681 , \15679 , \15680 );
not \U$15012 ( \15682 , \15681 );
not \U$15013 ( \15683 , \15682 );
or \U$15014 ( \15684 , \15644 , \15641 );
xor \U$15015 ( \15685 , \15684 , \15637 );
and \U$15016 ( \15686 , \14405 , \12838 );
and \U$15017 ( \15687 , \14935 , \13804 );
not \U$15018 ( \15688 , \14935 );
not \U$15019 ( \15689 , \14065 );
and \U$15020 ( \15690 , \15688 , \15689 );
nor \U$15021 ( \15691 , \15687 , \15690 );
nor \U$15022 ( \15692 , \15686 , \15691 );
not \U$15023 ( \15693 , \13674 );
nand \U$15024 ( \15694 , \15693 , \14946 );
not \U$15025 ( \15695 , \15694 );
not \U$15026 ( \15696 , \13674 );
not \U$15027 ( \15697 , \13558 );
or \U$15028 ( \15698 , \15696 , \15697 );
and \U$15029 ( \15699 , \13885 , \13781 );
not \U$15030 ( \15700 , \13885 );
not \U$15031 ( \15701 , \13566 );
and \U$15032 ( \15702 , \15700 , \15701 );
nor \U$15033 ( \15703 , \15699 , \15702 );
nand \U$15034 ( \15704 , \15698 , \15703 );
nor \U$15035 ( \15705 , \15695 , \15704 );
xor \U$15036 ( \15706 , \15692 , \15705 );
nand \U$15037 ( \15707 , \12272 , \15568 );
and \U$15038 ( \15708 , \15706 , \15707 );
and \U$15039 ( \15709 , \15692 , \15705 );
or \U$15040 ( \15710 , \15708 , \15709 );
not \U$15041 ( \15711 , \15710 );
not \U$15042 ( \15712 , \15639 );
not \U$15043 ( \15713 , \15712 );
not \U$15044 ( \15714 , \12276 );
or \U$15045 ( \15715 , \15713 , \15714 );
or \U$15046 ( \15716 , \12276 , \15712 );
nand \U$15047 ( \15717 , \15715 , \15716 );
not \U$15048 ( \15718 , \15717 );
not \U$15049 ( \15719 , \14107 );
or \U$15050 ( \15720 , \15718 , \15719 );
not \U$15051 ( \15721 , \12495 );
not \U$15052 ( \15722 , \15347 );
and \U$15053 ( \15723 , \15721 , \15722 );
nor \U$15054 ( \15724 , \12435 , \15346 );
nor \U$15055 ( \15725 , \15723 , \15724 );
nand \U$15056 ( \15726 , \15720 , \15725 );
not \U$15057 ( \15727 , \15726 );
or \U$15058 ( \15728 , \15711 , \15727 );
or \U$15059 ( \15729 , \15726 , \15710 );
nand \U$15060 ( \15730 , \15728 , \15729 );
not \U$15061 ( \15731 , \15730 );
not \U$15062 ( \15732 , \13830 );
not \U$15063 ( \15733 , \14514 );
not \U$15064 ( \15734 , \15733 );
and \U$15065 ( \15735 , \15732 , \15734 );
not \U$15066 ( \15736 , \15733 );
not \U$15067 ( \15737 , \13267 );
or \U$15068 ( \15738 , \15736 , \15737 );
and \U$15069 ( \15739 , \14517 , \13269 );
not \U$15070 ( \15740 , \14517 );
and \U$15071 ( \15741 , \15740 , \13169 );
nor \U$15072 ( \15742 , \15739 , \15741 );
nand \U$15073 ( \15743 , \15738 , \15742 );
nor \U$15074 ( \15744 , \15735 , \15743 );
not \U$15075 ( \15745 , \15744 );
not \U$15076 ( \15746 , \15745 );
not \U$15077 ( \15747 , \13798 );
not \U$15078 ( \15748 , \13019 );
and \U$15079 ( \15749 , \15747 , \15748 );
and \U$15080 ( \15750 , \12838 , \14060 );
not \U$15081 ( \15751 , \12838 );
buf \U$15082 ( \15752 , \14065 );
and \U$15083 ( \15753 , \15751 , \15752 );
or \U$15084 ( \15754 , \15750 , \15753 );
nor \U$15085 ( \15755 , \15749 , \15754 );
not \U$15086 ( \15756 , \15755 );
not \U$15087 ( \15757 , \13770 );
not \U$15088 ( \15758 , \13578 );
or \U$15089 ( \15759 , \15757 , \15758 );
and \U$15090 ( \15760 , \13559 , \13771 );
or \U$15091 ( \15761 , \13566 , \13841 );
not \U$15092 ( \15762 , \13572 );
nand \U$15093 ( \15763 , \15762 , \13674 );
nand \U$15094 ( \15764 , \15761 , \15763 );
nor \U$15095 ( \15765 , \15760 , \15764 );
nand \U$15096 ( \15766 , \15759 , \15765 );
nand \U$15097 ( \15767 , \15756 , \15766 );
not \U$15098 ( \15768 , \15767 );
not \U$15099 ( \15769 , \14830 );
and \U$15100 ( \15770 , \15769 , \14045 );
not \U$15101 ( \15771 , \12910 );
not \U$15102 ( \15772 , \14101 );
or \U$15103 ( \15773 , \15771 , \15772 );
not \U$15104 ( \15774 , \13815 );
or \U$15105 ( \15775 , \15774 , \13771 );
nand \U$15106 ( \15776 , \15773 , \15775 );
nor \U$15107 ( \15777 , \15770 , \15776 );
not \U$15108 ( \15778 , \14045 );
nand \U$15109 ( \15779 , \15778 , \13525 );
nand \U$15110 ( \15780 , \15777 , \15779 );
not \U$15111 ( \15781 , \15780 );
or \U$15112 ( \15782 , \15768 , \15781 );
or \U$15113 ( \15783 , \15780 , \15767 );
nand \U$15114 ( \15784 , \15782 , \15783 );
not \U$15115 ( \15785 , \15784 );
or \U$15116 ( \15786 , \15746 , \15785 );
not \U$15117 ( \15787 , \15767 );
nand \U$15118 ( \15788 , \15787 , \15780 );
nand \U$15119 ( \15789 , \15786 , \15788 );
not \U$15120 ( \15790 , \15789 );
or \U$15121 ( \15791 , \15731 , \15790 );
not \U$15122 ( \15792 , \15710 );
nand \U$15123 ( \15793 , \15792 , \15726 );
nand \U$15124 ( \15794 , \15791 , \15793 );
xor \U$15125 ( \15795 , \15685 , \15794 );
not \U$15126 ( \15796 , \15600 );
not \U$15127 ( \15797 , \15621 );
or \U$15128 ( \15798 , \15796 , \15797 );
or \U$15129 ( \15799 , \15621 , \15600 );
nand \U$15130 ( \15800 , \15798 , \15799 );
and \U$15131 ( \15801 , \15795 , \15800 );
and \U$15132 ( \15802 , \15685 , \15794 );
or \U$15133 ( \15803 , \15801 , \15802 );
not \U$15134 ( \15804 , \15626 );
not \U$15135 ( \15805 , \15804 );
not \U$15136 ( \15806 , \15654 );
or \U$15137 ( \15807 , \15805 , \15806 );
nand \U$15138 ( \15808 , \15653 , \15626 );
nand \U$15139 ( \15809 , \15807 , \15808 );
and \U$15140 ( \15810 , \15803 , \15809 );
not \U$15141 ( \15811 , \15803 );
not \U$15142 ( \15812 , \15809 );
and \U$15143 ( \15813 , \15811 , \15812 );
nor \U$15144 ( \15814 , \15810 , \15813 );
not \U$15145 ( \15815 , \15814 );
or \U$15146 ( \15816 , \15683 , \15815 );
not \U$15147 ( \15817 , \15812 );
nand \U$15148 ( \15818 , \15817 , \15803 );
nand \U$15149 ( \15819 , \15816 , \15818 );
xor \U$15150 ( \15820 , \15659 , \15590 );
xnor \U$15151 ( \15821 , \15820 , \15663 );
nand \U$15152 ( \15822 , \15819 , \15821 );
nand \U$15153 ( \15823 , \15671 , \15822 );
nand \U$15154 ( \15824 , \15670 , \15823 );
not \U$15155 ( \15825 , \15824 );
not \U$15156 ( \15826 , \14904 );
not \U$15157 ( \15827 , \14871 );
or \U$15158 ( \15828 , \15826 , \15827 );
or \U$15159 ( \15829 , \14904 , \14871 );
nand \U$15160 ( \15830 , \15828 , \15829 );
not \U$15161 ( \15831 , \15830 );
not \U$15162 ( \15832 , \14872 );
not \U$15163 ( \15833 , \15832 );
and \U$15164 ( \15834 , \15831 , \15833 );
and \U$15165 ( \15835 , \15830 , \15832 );
nor \U$15166 ( \15836 , \15834 , \15835 );
xor \U$15167 ( \15837 , \14932 , \15069 );
xor \U$15168 ( \15838 , \15837 , \15124 );
xor \U$15169 ( \15839 , \15836 , \15838 );
not \U$15170 ( \15840 , \15421 );
not \U$15171 ( \15841 , \15409 );
not \U$15172 ( \15842 , \15841 );
not \U$15173 ( \15843 , \15415 );
or \U$15174 ( \15844 , \15842 , \15843 );
or \U$15175 ( \15845 , \15415 , \15841 );
nand \U$15176 ( \15846 , \15844 , \15845 );
not \U$15177 ( \15847 , \15846 );
or \U$15178 ( \15848 , \15840 , \15847 );
not \U$15179 ( \15849 , \15841 );
nand \U$15180 ( \15850 , \15849 , \15415 );
nand \U$15181 ( \15851 , \15848 , \15850 );
xor \U$15182 ( \15852 , \15839 , \15851 );
xor \U$15183 ( \15853 , \15191 , \15407 );
and \U$15184 ( \15854 , \15853 , \15422 );
and \U$15185 ( \15855 , \15191 , \15407 );
or \U$15186 ( \15856 , \15854 , \15855 );
nand \U$15187 ( \15857 , \15852 , \15856 );
not \U$15188 ( \15858 , \15836 );
nand \U$15189 ( \15859 , \15851 , \15858 );
not \U$15190 ( \15860 , \15859 );
not \U$15191 ( \15861 , \15851 );
nand \U$15192 ( \15862 , \15861 , \15836 );
not \U$15193 ( \15863 , \15862 );
or \U$15194 ( \15864 , \15860 , \15863 );
nand \U$15195 ( \15865 , \15864 , \15838 );
nand \U$15196 ( \15866 , \15861 , \15858 );
nand \U$15197 ( \15867 , \15865 , \15866 );
not \U$15198 ( \15868 , \14926 );
not \U$15199 ( \15869 , \15139 );
or \U$15200 ( \15870 , \15868 , \15869 );
or \U$15201 ( \15871 , \15139 , \14926 );
nand \U$15202 ( \15872 , \15870 , \15871 );
nand \U$15203 ( \15873 , \15867 , \15872 );
nand \U$15204 ( \15874 , \15857 , \15873 );
not \U$15205 ( \15875 , \15874 );
nand \U$15206 ( \15876 , \15825 , \15875 );
not \U$15207 ( \15877 , \15873 );
not \U$15208 ( \15878 , \15856 );
not \U$15209 ( \15879 , \15852 );
nand \U$15210 ( \15880 , \15878 , \15879 );
or \U$15211 ( \15881 , \15877 , \15880 );
not \U$15212 ( \15882 , \15872 );
nand \U$15213 ( \15883 , \15882 , \15865 , \15866 );
nand \U$15214 ( \15884 , \15881 , \15883 );
not \U$15215 ( \15885 , \15884 );
nand \U$15216 ( \15886 , \15876 , \15885 );
not \U$15217 ( \15887 , \15886 );
or \U$15218 ( \15888 , \15189 , \15887 );
not \U$15219 ( \15889 , \15681 );
not \U$15220 ( \15890 , \15814 );
or \U$15221 ( \15891 , \15889 , \15890 );
or \U$15222 ( \15892 , \15681 , \15814 );
nand \U$15223 ( \15893 , \15891 , \15892 );
not \U$15224 ( \15894 , \15577 );
not \U$15225 ( \15895 , \15508 );
and \U$15226 ( \15896 , \15894 , \15895 );
and \U$15227 ( \15897 , \15577 , \15508 );
nor \U$15228 ( \15898 , \15896 , \15897 );
not \U$15229 ( \15899 , \15898 );
xor \U$15230 ( \15900 , \15447 , \15492 );
nand \U$15231 ( \15901 , \15899 , \15900 );
not \U$15232 ( \15902 , \15043 );
not \U$15233 ( \15903 , \15902 );
not \U$15234 ( \15904 , \13235 );
or \U$15235 ( \15905 , \15903 , \15904 );
or \U$15236 ( \15906 , \12844 , \15902 );
nand \U$15237 ( \15907 , \15905 , \15906 );
not \U$15238 ( \15908 , \15907 );
not \U$15239 ( \15909 , \12780 );
or \U$15240 ( \15910 , \15908 , \15909 );
nand \U$15241 ( \15911 , \15478 , \13869 );
nand \U$15242 ( \15912 , \15910 , \15911 );
not \U$15243 ( \15913 , \15912 );
xor \U$15244 ( \15914 , \15692 , \15705 );
xor \U$15245 ( \15915 , \15914 , \15707 );
not \U$15246 ( \15916 , \15915 );
or \U$15247 ( \15917 , \15913 , \15916 );
or \U$15248 ( \15918 , \15915 , \15912 );
nand \U$15249 ( \15919 , \15917 , \15918 );
not \U$15250 ( \15920 , \15919 );
not \U$15251 ( \15921 , \15592 );
not \U$15252 ( \15922 , \15921 );
not \U$15253 ( \15923 , \12585 );
or \U$15254 ( \15924 , \15922 , \15923 );
not \U$15255 ( \15925 , \12600 );
not \U$15256 ( \15926 , \15261 );
or \U$15257 ( \15927 , \15925 , \15926 );
or \U$15258 ( \15928 , \13627 , \15261 );
nand \U$15259 ( \15929 , \15927 , \15928 );
nor \U$15260 ( \15930 , \12598 , \15921 );
nor \U$15261 ( \15931 , \15929 , \15930 );
nand \U$15262 ( \15932 , \15924 , \15931 );
not \U$15263 ( \15933 , \15932 );
or \U$15264 ( \15934 , \15920 , \15933 );
not \U$15265 ( \15935 , \15915 );
nand \U$15266 ( \15936 , \15935 , \15912 );
nand \U$15267 ( \15937 , \15934 , \15936 );
nand \U$15268 ( \15938 , \15937 , \15900 );
nand \U$15269 ( \15939 , \15937 , \15899 );
nand \U$15270 ( \15940 , \15901 , \15938 , \15939 );
not \U$15271 ( \15941 , \15940 );
xor \U$15272 ( \15942 , \15432 , \15497 );
xor \U$15273 ( \15943 , \15942 , \15581 );
not \U$15274 ( \15944 , \15943 );
nand \U$15275 ( \15945 , \15941 , \15944 );
not \U$15276 ( \15946 , \15945 );
xor \U$15277 ( \15947 , \15685 , \15794 );
xor \U$15278 ( \15948 , \15947 , \15800 );
not \U$15279 ( \15949 , \15948 );
or \U$15280 ( \15950 , \15946 , \15949 );
nand \U$15281 ( \15951 , \15943 , \15940 );
nand \U$15282 ( \15952 , \15950 , \15951 );
nor \U$15283 ( \15953 , \15893 , \15952 );
not \U$15284 ( \15954 , \15953 );
not \U$15285 ( \15955 , \15954 );
xor \U$15286 ( \15956 , \15730 , \15789 );
not \U$15287 ( \15957 , \15755 );
not \U$15288 ( \15958 , \15766 );
or \U$15289 ( \15959 , \15957 , \15958 );
or \U$15290 ( \15960 , \15766 , \15755 );
nand \U$15291 ( \15961 , \15959 , \15960 );
and \U$15292 ( \15962 , \15261 , \13235 );
not \U$15293 ( \15963 , \15261 );
and \U$15294 ( \15964 , \15963 , \14648 );
nor \U$15295 ( \15965 , \15962 , \15964 );
not \U$15296 ( \15966 , \15965 );
not \U$15297 ( \15967 , \13861 );
or \U$15298 ( \15968 , \15966 , \15967 );
nand \U$15299 ( \15969 , \15907 , \13869 );
nand \U$15300 ( \15970 , \15968 , \15969 );
not \U$15301 ( \15971 , \15970 );
and \U$15302 ( \15972 , \15961 , \15971 );
not \U$15303 ( \15973 , \15961 );
and \U$15304 ( \15974 , \15973 , \15970 );
or \U$15305 ( \15975 , \15972 , \15974 );
not \U$15306 ( \15976 , \15975 );
not \U$15307 ( \15977 , \15640 );
not \U$15308 ( \15978 , \12585 );
or \U$15309 ( \15979 , \15977 , \15978 );
not \U$15310 ( \15980 , \12600 );
not \U$15311 ( \15981 , \15592 );
or \U$15312 ( \15982 , \15980 , \15981 );
or \U$15313 ( \15983 , \13627 , \15592 );
nand \U$15314 ( \15984 , \15982 , \15983 );
and \U$15315 ( \15985 , \14117 , \15639 );
nor \U$15316 ( \15986 , \15984 , \15985 );
nand \U$15317 ( \15987 , \15979 , \15986 );
not \U$15318 ( \15988 , \15987 );
or \U$15319 ( \15989 , \15976 , \15988 );
nand \U$15320 ( \15990 , \15970 , \15961 );
nand \U$15321 ( \15991 , \15989 , \15990 );
not \U$15322 ( \15992 , \15991 );
not \U$15323 ( \15993 , \13159 );
not \U$15324 ( \15994 , \15993 );
not \U$15325 ( \15995 , \14796 );
and \U$15326 ( \15996 , \15994 , \15995 );
not \U$15327 ( \15997 , \14796 );
not \U$15328 ( \15998 , \13164 );
or \U$15329 ( \15999 , \15997 , \15998 );
and \U$15330 ( \16000 , \15100 , \13269 );
not \U$15331 ( \16001 , \15100 );
and \U$15332 ( \16002 , \16001 , \13169 );
nor \U$15333 ( \16003 , \16000 , \16002 );
nand \U$15334 ( \16004 , \15999 , \16003 );
nor \U$15335 ( \16005 , \15996 , \16004 );
not \U$15336 ( \16006 , \16005 );
not \U$15337 ( \16007 , \16006 );
and \U$15338 ( \16008 , \13235 , \12587 );
nor \U$15339 ( \16009 , \16008 , \15567 );
nor \U$15340 ( \16010 , \12670 , \16009 );
not \U$15341 ( \16011 , \16010 );
not \U$15342 ( \16012 , \14454 );
not \U$15343 ( \16013 , \14831 );
or \U$15344 ( \16014 , \16012 , \16013 );
and \U$15345 ( \16015 , \15077 , \13815 );
not \U$15346 ( \16016 , \15077 );
not \U$15347 ( \16017 , \13717 );
and \U$15348 ( \16018 , \16016 , \16017 );
nor \U$15349 ( \16019 , \16015 , \16018 );
nand \U$15350 ( \16020 , \16014 , \16019 );
and \U$15351 ( \16021 , \12897 , \14517 );
nor \U$15352 ( \16022 , \16020 , \16021 );
not \U$15353 ( \16023 , \16022 );
or \U$15354 ( \16024 , \16011 , \16023 );
not \U$15355 ( \16025 , \16021 );
not \U$15356 ( \16026 , \16025 );
not \U$15357 ( \16027 , \16020 );
not \U$15358 ( \16028 , \16027 );
or \U$15359 ( \16029 , \16026 , \16028 );
not \U$15360 ( \16030 , \16010 );
nand \U$15361 ( \16031 , \16029 , \16030 );
nand \U$15362 ( \16032 , \16024 , \16031 );
not \U$15363 ( \16033 , \16032 );
or \U$15364 ( \16034 , \16007 , \16033 );
not \U$15365 ( \16035 , \16025 );
not \U$15366 ( \16036 , \16027 );
or \U$15367 ( \16037 , \16035 , \16036 );
nand \U$15368 ( \16038 , \16037 , \16010 );
nand \U$15369 ( \16039 , \16034 , \16038 );
not \U$15370 ( \16040 , \16039 );
not \U$15371 ( \16041 , \15744 );
not \U$15372 ( \16042 , \15784 );
or \U$15373 ( \16043 , \16041 , \16042 );
or \U$15374 ( \16044 , \15784 , \15744 );
nand \U$15375 ( \16045 , \16043 , \16044 );
not \U$15376 ( \16046 , \16045 );
not \U$15377 ( \16047 , \16046 );
or \U$15378 ( \16048 , \16040 , \16047 );
not \U$15379 ( \16049 , \16039 );
nand \U$15380 ( \16050 , \16049 , \16045 );
nand \U$15381 ( \16051 , \16048 , \16050 );
not \U$15382 ( \16052 , \16051 );
or \U$15383 ( \16053 , \15992 , \16052 );
nand \U$15384 ( \16054 , \16045 , \16039 );
nand \U$15385 ( \16055 , \16053 , \16054 );
not \U$15386 ( \16056 , \16055 );
xor \U$15387 ( \16057 , \15956 , \16056 );
not \U$15388 ( \16058 , \15899 );
not \U$15389 ( \16059 , \15900 );
not \U$15390 ( \16060 , \16059 );
or \U$15391 ( \16061 , \16058 , \16060 );
nand \U$15392 ( \16062 , \15898 , \15900 );
nand \U$15393 ( \16063 , \16061 , \16062 );
and \U$15394 ( \16064 , \16063 , \15937 );
not \U$15395 ( \16065 , \16063 );
not \U$15396 ( \16066 , \15937 );
and \U$15397 ( \16067 , \16065 , \16066 );
nor \U$15398 ( \16068 , \16064 , \16067 );
xnor \U$15399 ( \16069 , \16057 , \16068 );
not \U$15400 ( \16070 , \16069 );
buf \U$15401 ( \16071 , \15932 );
buf \U$15402 ( \16072 , \15919 );
and \U$15403 ( \16073 , \16071 , \16072 );
not \U$15404 ( \16074 , \16071 );
not \U$15405 ( \16075 , \16072 );
and \U$15406 ( \16076 , \16074 , \16075 );
nor \U$15407 ( \16077 , \16073 , \16076 );
and \U$15408 ( \16078 , \16051 , \15991 );
not \U$15409 ( \16079 , \16051 );
not \U$15410 ( \16080 , \15991 );
and \U$15411 ( \16081 , \16079 , \16080 );
nor \U$15412 ( \16082 , \16078 , \16081 );
xor \U$15413 ( \16083 , \16077 , \16082 );
not \U$15414 ( \16084 , \15045 );
not \U$15415 ( \16085 , \13160 );
or \U$15416 ( \16086 , \16084 , \16085 );
and \U$15417 ( \16087 , \13267 , \15044 );
not \U$15418 ( \16088 , \13169 );
or \U$15419 ( \16089 , \16088 , \14797 );
not \U$15420 ( \16090 , \14796 );
nand \U$15421 ( \16091 , \16090 , \13173 );
nand \U$15422 ( \16092 , \16089 , \16091 );
nor \U$15423 ( \16093 , \16087 , \16092 );
nand \U$15424 ( \16094 , \16086 , \16093 );
not \U$15425 ( \16095 , \16094 );
nand \U$15426 ( \16096 , \13578 , \14517 );
not \U$15427 ( \16097 , \16096 );
and \U$15428 ( \16098 , \14807 , \14454 );
or \U$15429 ( \16099 , \13566 , \14044 );
not \U$15430 ( \16100 , \14043 );
nand \U$15431 ( \16101 , \16100 , \13781 );
nand \U$15432 ( \16102 , \16099 , \16101 );
nor \U$15433 ( \16103 , \16098 , \16102 );
not \U$15434 ( \16104 , \16103 );
or \U$15435 ( \16105 , \16097 , \16104 );
and \U$15436 ( \16106 , \15752 , \13673 );
nor \U$15437 ( \16107 , \13804 , \13673 );
nor \U$15438 ( \16108 , \16106 , \16107 );
nand \U$15439 ( \16109 , \14405 , \14101 );
nand \U$15440 ( \16110 , \16108 , \16109 );
nand \U$15441 ( \16111 , \16105 , \16110 );
not \U$15442 ( \16112 , \16111 );
not \U$15443 ( \16113 , \12903 );
not \U$15444 ( \16114 , \15100 );
and \U$15445 ( \16115 , \16113 , \16114 );
or \U$15446 ( \16116 , \13520 , \14454 );
not \U$15447 ( \16117 , \13717 );
nand \U$15448 ( \16118 , \16117 , \14454 );
nand \U$15449 ( \16119 , \16116 , \16118 );
nor \U$15450 ( \16120 , \16115 , \16119 );
nand \U$15451 ( \16121 , \13525 , \14514 );
nand \U$15452 ( \16122 , \16120 , \16121 );
not \U$15453 ( \16123 , \16122 );
or \U$15454 ( \16124 , \16112 , \16123 );
or \U$15455 ( \16125 , \16122 , \16111 );
nand \U$15456 ( \16126 , \16124 , \16125 );
not \U$15457 ( \16127 , \16126 );
or \U$15458 ( \16128 , \16095 , \16127 );
not \U$15459 ( \16129 , \16111 );
nand \U$15460 ( \16130 , \16129 , \16122 );
nand \U$15461 ( \16131 , \16128 , \16130 );
not \U$15462 ( \16132 , \16131 );
xor \U$15463 ( \16133 , \16005 , \16032 );
not \U$15464 ( \16134 , \13019 );
not \U$15465 ( \16135 , \13804 );
and \U$15466 ( \16136 , \16134 , \16135 );
and \U$15467 ( \16137 , \14401 , \13886 );
nor \U$15468 ( \16138 , \16136 , \16137 );
not \U$15469 ( \16139 , \14404 );
nand \U$15470 ( \16140 , \16139 , \13675 );
nand \U$15471 ( \16141 , \16138 , \16140 );
and \U$15472 ( \16142 , \13559 , \14044 );
or \U$15473 ( \16143 , \14809 , \13769 );
or \U$15474 ( \16144 , \13566 , \14101 );
nand \U$15475 ( \16145 , \16143 , \16144 );
nor \U$15476 ( \16146 , \16142 , \16145 );
nand \U$15477 ( \16147 , \13578 , \15077 );
nand \U$15478 ( \16148 , \16146 , \16147 );
xor \U$15479 ( \16149 , \16141 , \16148 );
not \U$15480 ( \16150 , \13079 );
nand \U$15481 ( \16151 , \16150 , \15712 );
not \U$15482 ( \16152 , \16151 );
and \U$15483 ( \16153 , \16149 , \16152 );
and \U$15484 ( \16154 , \16141 , \16148 );
nor \U$15485 ( \16155 , \16153 , \16154 );
xor \U$15486 ( \16156 , \16133 , \16155 );
not \U$15487 ( \16157 , \16156 );
or \U$15488 ( \16158 , \16132 , \16157 );
buf \U$15489 ( \16159 , \16032 );
nand \U$15490 ( \16160 , \16159 , \16005 );
not \U$15491 ( \16161 , \16160 );
not \U$15492 ( \16162 , \16159 );
nand \U$15493 ( \16163 , \16162 , \16006 );
not \U$15494 ( \16164 , \16163 );
or \U$15495 ( \16165 , \16161 , \16164 );
not \U$15496 ( \16166 , \16155 );
nand \U$15497 ( \16167 , \16165 , \16166 );
nand \U$15498 ( \16168 , \16158 , \16167 );
and \U$15499 ( \16169 , \16083 , \16168 );
and \U$15500 ( \16170 , \16077 , \16082 );
or \U$15501 ( \16171 , \16169 , \16170 );
not \U$15502 ( \16172 , \16171 );
nand \U$15503 ( \16173 , \16070 , \16172 );
not \U$15504 ( \16174 , \16171 );
not \U$15505 ( \16175 , \16069 );
or \U$15506 ( \16176 , \16174 , \16175 );
xor \U$15507 ( \16177 , \16077 , \16082 );
xor \U$15508 ( \16178 , \16177 , \16168 );
and \U$15509 ( \16179 , \16156 , \16131 );
not \U$15510 ( \16180 , \16156 );
not \U$15511 ( \16181 , \16131 );
and \U$15512 ( \16182 , \16180 , \16181 );
nor \U$15513 ( \16183 , \16179 , \16182 );
not \U$15514 ( \16184 , \16183 );
xor \U$15515 ( \16185 , \15987 , \15975 );
not \U$15516 ( \16186 , \16151 );
and \U$15517 ( \16187 , \16149 , \16186 );
not \U$15518 ( \16188 , \16149 );
and \U$15519 ( \16189 , \16188 , \16151 );
nor \U$15520 ( \16190 , \16187 , \16189 );
not \U$15521 ( \16191 , \16190 );
not \U$15522 ( \16192 , \15346 );
not \U$15523 ( \16193 , \13339 );
or \U$15524 ( \16194 , \16192 , \16193 );
not \U$15525 ( \16195 , \13345 );
not \U$15526 ( \16196 , \15346 );
and \U$15527 ( \16197 , \16195 , \16196 );
and \U$15528 ( \16198 , \15261 , \13430 );
not \U$15529 ( \16199 , \15261 );
not \U$15530 ( \16200 , \14660 );
and \U$15531 ( \16201 , \16199 , \16200 );
nor \U$15532 ( \16202 , \16198 , \16201 );
nor \U$15533 ( \16203 , \16197 , \16202 );
nand \U$15534 ( \16204 , \16194 , \16203 );
not \U$15535 ( \16205 , \16204 );
not \U$15536 ( \16206 , \16205 );
not \U$15537 ( \16207 , \13235 );
not \U$15538 ( \16208 , \15639 );
not \U$15539 ( \16209 , \13163 );
or \U$15540 ( \16210 , \16208 , \16209 );
not \U$15541 ( \16211 , \13237 );
nand \U$15542 ( \16212 , \16210 , \16211 );
nand \U$15543 ( \16213 , \13302 , \15640 );
and \U$15544 ( \16214 , \16207 , \16212 , \16213 );
not \U$15545 ( \16215 , \16110 );
not \U$15546 ( \16216 , \16215 );
nand \U$15547 ( \16217 , \16103 , \16096 );
not \U$15548 ( \16218 , \16217 );
or \U$15549 ( \16219 , \16216 , \16218 );
nand \U$15550 ( \16220 , \16103 , \16096 , \16110 );
nand \U$15551 ( \16221 , \16219 , \16220 );
xor \U$15552 ( \16222 , \16214 , \16221 );
and \U$15553 ( \16223 , \15769 , \14796 );
not \U$15554 ( \16224 , \13718 );
not \U$15555 ( \16225 , \14513 );
or \U$15556 ( \16226 , \16224 , \16225 );
or \U$15557 ( \16227 , \13520 , \15096 );
nand \U$15558 ( \16228 , \16226 , \16227 );
nor \U$15559 ( \16229 , \16223 , \16228 );
nand \U$15560 ( \16230 , \13525 , \15054 );
nand \U$15561 ( \16231 , \16229 , \16230 );
and \U$15562 ( \16232 , \16222 , \16231 );
and \U$15563 ( \16233 , \16214 , \16221 );
or \U$15564 ( \16234 , \16232 , \16233 );
not \U$15565 ( \16235 , \16234 );
or \U$15566 ( \16236 , \16206 , \16235 );
or \U$15567 ( \16237 , \16234 , \16205 );
nand \U$15568 ( \16238 , \16236 , \16237 );
not \U$15569 ( \16239 , \16238 );
or \U$15570 ( \16240 , \16191 , \16239 );
not \U$15571 ( \16241 , \16205 );
buf \U$15572 ( \16242 , \16234 );
nand \U$15573 ( \16243 , \16241 , \16242 );
nand \U$15574 ( \16244 , \16240 , \16243 );
and \U$15575 ( \16245 , \16185 , \16244 );
not \U$15576 ( \16246 , \16185 );
not \U$15577 ( \16247 , \16244 );
and \U$15578 ( \16248 , \16246 , \16247 );
nor \U$15579 ( \16249 , \16245 , \16248 );
not \U$15580 ( \16250 , \16249 );
or \U$15581 ( \16251 , \16184 , \16250 );
nand \U$15582 ( \16252 , \16244 , \16185 );
nand \U$15583 ( \16253 , \16251 , \16252 );
nand \U$15584 ( \16254 , \16178 , \16253 );
nand \U$15585 ( \16255 , \16176 , \16254 );
nand \U$15586 ( \16256 , \16173 , \16255 );
nand \U$15587 ( \16257 , \15945 , \15951 );
and \U$15588 ( \16258 , \16257 , \15948 );
not \U$15589 ( \16259 , \16257 );
not \U$15590 ( \16260 , \15948 );
and \U$15591 ( \16261 , \16259 , \16260 );
nor \U$15592 ( \16262 , \16258 , \16261 );
buf \U$15593 ( \16263 , \15956 );
not \U$15594 ( \16264 , \16056 );
xor \U$15595 ( \16265 , \16263 , \16264 );
buf \U$15596 ( \16266 , \16068 );
and \U$15597 ( \16267 , \16265 , \16266 );
and \U$15598 ( \16268 , \16263 , \16264 );
nor \U$15599 ( \16269 , \16267 , \16268 );
nand \U$15600 ( \16270 , \16262 , \16269 );
not \U$15601 ( \16271 , \16270 );
or \U$15602 ( \16272 , \16256 , \16271 );
and \U$15603 ( \16273 , \15893 , \15952 );
nor \U$15604 ( \16274 , \16269 , \16262 );
nor \U$15605 ( \16275 , \16273 , \16274 );
nand \U$15606 ( \16276 , \16272 , \16275 );
not \U$15607 ( \16277 , \16276 );
or \U$15608 ( \16278 , \15955 , \16277 );
not \U$15609 ( \16279 , \16178 );
not \U$15610 ( \16280 , \16253 );
nand \U$15611 ( \16281 , \16279 , \16280 );
and \U$15612 ( \16282 , \16173 , \16281 );
xor \U$15613 ( \16283 , \16185 , \16247 );
xnor \U$15614 ( \16284 , \16283 , \16183 );
not \U$15615 ( \16285 , \16284 );
xor \U$15616 ( \16286 , \16126 , \16094 );
not \U$15617 ( \16287 , \16286 );
not \U$15618 ( \16288 , \15262 );
not \U$15619 ( \16289 , \13160 );
or \U$15620 ( \16290 , \16288 , \16289 );
and \U$15621 ( \16291 , \13166 , \15261 );
not \U$15622 ( \16292 , \15902 );
not \U$15623 ( \16293 , \13269 );
or \U$15624 ( \16294 , \16292 , \16293 );
not \U$15625 ( \16295 , \13169 );
or \U$15626 ( \16296 , \16295 , \15442 );
nand \U$15627 ( \16297 , \16294 , \16296 );
nor \U$15628 ( \16298 , \16291 , \16297 );
nand \U$15629 ( \16299 , \16290 , \16298 );
not \U$15630 ( \16300 , \16299 );
not \U$15631 ( \16301 , \14945 );
not \U$15632 ( \16302 , \14513 );
and \U$15633 ( \16303 , \16301 , \16302 );
not \U$15634 ( \16304 , \14513 );
not \U$15635 ( \16305 , \14806 );
or \U$15636 ( \16306 , \16304 , \16305 );
and \U$15637 ( \16307 , \14453 , \13781 );
not \U$15638 ( \16308 , \14453 );
and \U$15639 ( \16309 , \16308 , \14813 );
nor \U$15640 ( \16310 , \16307 , \16309 );
nand \U$15641 ( \16311 , \16306 , \16310 );
nor \U$15642 ( \16312 , \16303 , \16311 );
not \U$15643 ( \16313 , \14044 );
not \U$15644 ( \16314 , \13797 );
or \U$15645 ( \16315 , \16313 , \16314 );
not \U$15646 ( \16316 , \14819 );
not \U$15647 ( \16317 , \14101 );
and \U$15648 ( \16318 , \16316 , \16317 );
and \U$15649 ( \16319 , \14060 , \14101 );
nor \U$15650 ( \16320 , \16318 , \16319 );
nand \U$15651 ( \16321 , \16315 , \16320 );
not \U$15652 ( \16322 , \16321 );
and \U$15653 ( \16323 , \16312 , \16322 );
not \U$15654 ( \16324 , \16312 );
and \U$15655 ( \16325 , \16324 , \16321 );
nor \U$15656 ( \16326 , \16323 , \16325 );
not \U$15657 ( \16327 , \16326 );
and \U$15658 ( \16328 , \12845 , \15712 );
not \U$15659 ( \16329 , \16328 );
or \U$15660 ( \16330 , \16327 , \16329 );
not \U$15661 ( \16331 , \16312 );
nand \U$15662 ( \16332 , \16331 , \16321 );
nand \U$15663 ( \16333 , \16330 , \16332 );
not \U$15664 ( \16334 , \16333 );
and \U$15665 ( \16335 , \16300 , \16334 );
not \U$15666 ( \16336 , \15640 );
not \U$15667 ( \16337 , \13339 );
or \U$15668 ( \16338 , \16336 , \16337 );
not \U$15669 ( \16339 , \13345 );
not \U$15670 ( \16340 , \15640 );
and \U$15671 ( \16341 , \16339 , \16340 );
or \U$15672 ( \16342 , \12846 , \15347 );
nand \U$15673 ( \16343 , \12770 , \15347 );
nand \U$15674 ( \16344 , \16342 , \16343 );
nor \U$15675 ( \16345 , \16341 , \16344 );
nand \U$15676 ( \16346 , \16338 , \16345 );
not \U$15677 ( \16347 , \16346 );
nor \U$15678 ( \16348 , \16335 , \16347 );
and \U$15679 ( \16349 , \16333 , \16299 );
nor \U$15680 ( \16350 , \16348 , \16349 );
not \U$15681 ( \16351 , \16350 );
or \U$15682 ( \16352 , \16287 , \16351 );
or \U$15683 ( \16353 , \16350 , \16286 );
nand \U$15684 ( \16354 , \16352 , \16353 );
not \U$15685 ( \16355 , \16354 );
xor \U$15686 ( \16356 , \16190 , \16205 );
xor \U$15687 ( \16357 , \16356 , \16242 );
not \U$15688 ( \16358 , \16357 );
not \U$15689 ( \16359 , \16358 );
or \U$15690 ( \16360 , \16355 , \16359 );
not \U$15691 ( \16361 , \16350 );
nand \U$15692 ( \16362 , \16361 , \16286 );
nand \U$15693 ( \16363 , \16360 , \16362 );
not \U$15694 ( \16364 , \16363 );
nand \U$15695 ( \16365 , \16285 , \16364 );
and \U$15696 ( \16366 , \16270 , \16365 );
not \U$15697 ( \16367 , \16354 );
not \U$15698 ( \16368 , \16357 );
or \U$15699 ( \16369 , \16367 , \16368 );
or \U$15700 ( \16370 , \16354 , \16357 );
nand \U$15701 ( \16371 , \16369 , \16370 );
not \U$15702 ( \16372 , \16371 );
xor \U$15703 ( \16373 , \16333 , \16299 );
and \U$15704 ( \16374 , \16373 , \16346 );
not \U$15705 ( \16375 , \16373 );
and \U$15706 ( \16376 , \16375 , \16347 );
nor \U$15707 ( \16377 , \16374 , \16376 );
xor \U$15708 ( \16378 , \16214 , \16221 );
xor \U$15709 ( \16379 , \16378 , \16231 );
not \U$15710 ( \16380 , \16379 );
not \U$15711 ( \16381 , \15902 );
and \U$15712 ( \16382 , \14831 , \16381 );
not \U$15713 ( \16383 , \13815 );
or \U$15714 ( \16384 , \16383 , \14796 );
nand \U$15715 ( \16385 , \12910 , \14796 );
nand \U$15716 ( \16386 , \16384 , \16385 );
nor \U$15717 ( \16387 , \16382 , \16386 );
nand \U$15718 ( \16388 , \15902 , \13525 );
not \U$15719 ( \16389 , \13147 );
not \U$15720 ( \16390 , \16389 );
not \U$15721 ( \16391 , \15638 );
or \U$15722 ( \16392 , \16390 , \16391 );
nand \U$15723 ( \16393 , \16392 , \13812 );
not \U$15724 ( \16394 , \16389 );
nand \U$15725 ( \16395 , \16394 , \15566 );
and \U$15726 ( \16396 , \14043 , \14065 );
nor \U$15727 ( \16397 , \13803 , \14043 );
nor \U$15728 ( \16398 , \16396 , \16397 );
nand \U$15729 ( \16399 , \13797 , \14453 );
nand \U$15730 ( \16400 , \16398 , \16399 );
nand \U$15731 ( \16401 , \16393 , \13302 , \16395 , \16400 );
buf \U$15732 ( \16402 , \16401 );
nand \U$15733 ( \16403 , \16387 , \16388 , \16402 );
nor \U$15734 ( \16404 , \13165 , \15346 );
not \U$15735 ( \16405 , \16404 );
not \U$15736 ( \16406 , \15993 );
nand \U$15737 ( \16407 , \16406 , \15921 );
and \U$15738 ( \16408 , \15262 , \13269 );
not \U$15739 ( \16409 , \15262 );
and \U$15740 ( \16410 , \16409 , \13169 );
nor \U$15741 ( \16411 , \16408 , \16410 );
nand \U$15742 ( \16412 , \16405 , \16407 , \16411 );
and \U$15743 ( \16413 , \16403 , \16412 );
not \U$15744 ( \16414 , \16402 );
nand \U$15745 ( \16415 , \16387 , \16388 );
nand \U$15746 ( \16416 , \16414 , \16415 );
not \U$15747 ( \16417 , \16416 );
nor \U$15748 ( \16418 , \16413 , \16417 );
nand \U$15749 ( \16419 , \16380 , \16418 );
nand \U$15750 ( \16420 , \16377 , \16419 );
not \U$15751 ( \16421 , \16418 );
nand \U$15752 ( \16422 , \16421 , \16379 );
nand \U$15753 ( \16423 , \16420 , \16422 );
not \U$15754 ( \16424 , \16423 );
nand \U$15755 ( \16425 , \16372 , \16424 );
xor \U$15756 ( \16426 , \16326 , \16328 );
not \U$15757 ( \16427 , \15262 );
not \U$15758 ( \16428 , \12898 );
or \U$15759 ( \16429 , \16427 , \16428 );
and \U$15760 ( \16430 , \12904 , \15261 );
or \U$15761 ( \16431 , \13520 , \15044 );
not \U$15762 ( \16432 , \16017 );
or \U$15763 ( \16433 , \16432 , \15902 );
nand \U$15764 ( \16434 , \16431 , \16433 );
nor \U$15765 ( \16435 , \16430 , \16434 );
nand \U$15766 ( \16436 , \16429 , \16435 );
not \U$15767 ( \16437 , \16436 );
not \U$15768 ( \16438 , \16400 );
not \U$15769 ( \16439 , \16438 );
nand \U$15770 ( \16440 , \16393 , \13158 , \16395 );
not \U$15771 ( \16441 , \16440 );
or \U$15772 ( \16442 , \16439 , \16441 );
nand \U$15773 ( \16443 , \16442 , \16401 );
not \U$15774 ( \16444 , \14796 );
not \U$15775 ( \16445 , \13558 );
or \U$15776 ( \16446 , \16444 , \16445 );
and \U$15777 ( \16447 , \14513 , \13781 );
not \U$15778 ( \16448 , \14513 );
and \U$15779 ( \16449 , \16448 , \14813 );
nor \U$15780 ( \16450 , \16447 , \16449 );
nand \U$15781 ( \16451 , \16446 , \16450 );
not \U$15782 ( \16452 , \13578 );
nor \U$15783 ( \16453 , \16452 , \14796 );
nor \U$15784 ( \16454 , \16451 , \16453 );
nor \U$15785 ( \16455 , \16443 , \16454 );
not \U$15786 ( \16456 , \16455 );
and \U$15787 ( \16457 , \16437 , \16456 );
nand \U$15788 ( \16458 , \16443 , \16454 );
not \U$15789 ( \16459 , \16458 );
nor \U$15790 ( \16460 , \16457 , \16459 );
xor \U$15791 ( \16461 , \16426 , \16460 );
nand \U$15792 ( \16462 , \16416 , \16403 );
not \U$15793 ( \16463 , \16412 );
and \U$15794 ( \16464 , \16462 , \16463 );
not \U$15795 ( \16465 , \16462 );
and \U$15796 ( \16466 , \16465 , \16412 );
nor \U$15797 ( \16467 , \16464 , \16466 );
not \U$15798 ( \16468 , \16467 );
and \U$15799 ( \16469 , \16461 , \16468 );
not \U$15800 ( \16470 , \16461 );
and \U$15801 ( \16471 , \16470 , \16467 );
nor \U$15802 ( \16472 , \16469 , \16471 );
not \U$15803 ( \16473 , \16455 );
nand \U$15804 ( \16474 , \16473 , \16458 );
not \U$15805 ( \16475 , \16474 );
not \U$15806 ( \16476 , \16436 );
and \U$15807 ( \16477 , \16475 , \16476 );
and \U$15808 ( \16478 , \16436 , \16474 );
nor \U$15809 ( \16479 , \16477 , \16478 );
not \U$15810 ( \16480 , \16479 );
not \U$15811 ( \16481 , \15993 );
not \U$15812 ( \16482 , \15639 );
and \U$15813 ( \16483 , \16481 , \16482 );
not \U$15814 ( \16484 , \15639 );
not \U$15815 ( \16485 , \13164 );
or \U$15816 ( \16486 , \16484 , \16485 );
and \U$15817 ( \16487 , \15921 , \13173 );
not \U$15818 ( \16488 , \15921 );
and \U$15819 ( \16489 , \16488 , \13169 );
nor \U$15820 ( \16490 , \16487 , \16489 );
nand \U$15821 ( \16491 , \16486 , \16490 );
nor \U$15822 ( \16492 , \16483 , \16491 );
or \U$15823 ( \16493 , \15689 , \14453 );
nand \U$15824 ( \16494 , \14059 , \14453 );
nand \U$15825 ( \16495 , \16493 , \16494 );
nor \U$15826 ( \16496 , \13798 , \15095 );
nor \U$15827 ( \16497 , \16495 , \16496 );
not \U$15828 ( \16498 , \13301 );
nand \U$15829 ( \16499 , \16498 , \15640 );
xor \U$15830 ( \16500 , \16497 , \16499 );
not \U$15831 ( \16501 , \14949 );
not \U$15832 ( \16502 , \15043 );
or \U$15833 ( \16503 , \16501 , \16502 );
and \U$15834 ( \16504 , \14795 , \14054 );
not \U$15835 ( \16505 , \14795 );
and \U$15836 ( \16506 , \16505 , \14813 );
nor \U$15837 ( \16507 , \16504 , \16506 );
nand \U$15838 ( \16508 , \16503 , \16507 );
nor \U$15839 ( \16509 , \14945 , \15043 );
nor \U$15840 ( \16510 , \16508 , \16509 );
and \U$15841 ( \16511 , \16500 , \16510 );
and \U$15842 ( \16512 , \16497 , \16499 );
or \U$15843 ( \16513 , \16511 , \16512 );
nand \U$15844 ( \16514 , \16492 , \16513 );
and \U$15845 ( \16515 , \16480 , \16514 );
nor \U$15846 ( \16516 , \16492 , \16513 );
buf \U$15847 ( \16517 , \16516 );
nor \U$15848 ( \16518 , \16515 , \16517 );
nand \U$15849 ( \16519 , \16472 , \16518 );
not \U$15850 ( \16520 , \16519 );
not \U$15851 ( \16521 , \16516 );
nand \U$15852 ( \16522 , \16521 , \16514 );
not \U$15853 ( \16523 , \16522 );
not \U$15854 ( \16524 , \16479 );
or \U$15855 ( \16525 , \16523 , \16524 );
or \U$15856 ( \16526 , \16479 , \16522 );
nand \U$15857 ( \16527 , \16525 , \16526 );
not \U$15858 ( \16528 , \16527 );
not \U$15859 ( \16529 , \16528 );
not \U$15860 ( \16530 , \15564 );
not \U$15861 ( \16531 , \13515 );
or \U$15862 ( \16532 , \16530 , \16531 );
nand \U$15863 ( \16533 , \16532 , \12861 );
not \U$15864 ( \16534 , \13515 );
nand \U$15865 ( \16535 , \16534 , \15565 );
and \U$15866 ( \16536 , \16533 , \16535 , \12895 );
not \U$15867 ( \16537 , \13797 );
not \U$15868 ( \16538 , \14795 );
or \U$15869 ( \16539 , \16537 , \16538 );
and \U$15870 ( \16540 , \14512 , \14059 );
not \U$15871 ( \16541 , \14512 );
and \U$15872 ( \16542 , \16541 , \14065 );
nor \U$15873 ( \16543 , \16540 , \16542 );
nand \U$15874 ( \16544 , \16539 , \16543 );
nand \U$15875 ( \16545 , \16536 , \16544 );
not \U$15876 ( \16546 , \13525 );
not \U$15877 ( \16547 , \16546 );
not \U$15878 ( \16548 , \15592 );
and \U$15879 ( \16549 , \16547 , \16548 );
not \U$15880 ( \16550 , \15347 );
not \U$15881 ( \16551 , \14831 );
or \U$15882 ( \16552 , \16550 , \16551 );
and \U$15883 ( \16553 , \15261 , \16017 );
not \U$15884 ( \16554 , \15261 );
and \U$15885 ( \16555 , \16554 , \13815 );
nor \U$15886 ( \16556 , \16553 , \16555 );
nand \U$15887 ( \16557 , \16552 , \16556 );
nor \U$15888 ( \16558 , \16549 , \16557 );
xor \U$15889 ( \16559 , \16545 , \16558 );
xor \U$15890 ( \16560 , \16497 , \16499 );
xor \U$15891 ( \16561 , \16560 , \16510 );
and \U$15892 ( \16562 , \16559 , \16561 );
and \U$15893 ( \16563 , \16545 , \16558 );
or \U$15894 ( \16564 , \16562 , \16563 );
not \U$15895 ( \16565 , \16564 );
not \U$15896 ( \16566 , \16565 );
or \U$15897 ( \16567 , \16529 , \16566 );
not \U$15898 ( \16568 , \16564 );
not \U$15899 ( \16569 , \16527 );
or \U$15900 ( \16570 , \16568 , \16569 );
not \U$15901 ( \16571 , \15640 );
not \U$15902 ( \16572 , \13525 );
or \U$15903 ( \16573 , \16571 , \16572 );
not \U$15904 ( \16574 , \12903 );
and \U$15905 ( \16575 , \16574 , \15639 );
or \U$15906 ( \16576 , \13520 , \15592 );
nand \U$15907 ( \16577 , \16117 , \15592 );
nand \U$15908 ( \16578 , \16576 , \16577 );
nor \U$15909 ( \16579 , \16575 , \16578 );
nand \U$15910 ( \16580 , \16573 , \16579 );
xor \U$15911 ( \16581 , \15259 , \13515 );
nand \U$15912 ( \16582 , \16581 , \13513 );
not \U$15913 ( \16583 , \15042 );
not \U$15914 ( \16584 , \13515 );
or \U$15915 ( \16585 , \16583 , \16584 );
or \U$15916 ( \16586 , \13515 , \15042 );
nand \U$15917 ( \16587 , \16585 , \16586 );
nand \U$15918 ( \16588 , \16587 , \13512 );
and \U$15919 ( \16589 , \16582 , \13514 , \16588 );
not \U$15920 ( \16590 , \16589 );
nor \U$15921 ( \16591 , \16536 , \16544 );
not \U$15922 ( \16592 , \16591 );
nand \U$15923 ( \16593 , \16592 , \16545 );
not \U$15924 ( \16594 , \16593 );
or \U$15925 ( \16595 , \16590 , \16594 );
or \U$15926 ( \16596 , \16593 , \16589 );
nand \U$15927 ( \16597 , \16595 , \16596 );
or \U$15928 ( \16598 , \16580 , \16597 );
nand \U$15929 ( \16599 , \16580 , \16597 );
nand \U$15930 ( \16600 , \16598 , \16599 );
nand \U$15931 ( \16601 , \16581 , \13512 );
xor \U$15932 ( \16602 , \13515 , \15345 );
nand \U$15933 ( \16603 , \16602 , \13513 );
nand \U$15934 ( \16604 , \16601 , \16603 , \13514 );
not \U$15935 ( \16605 , \16604 );
nand \U$15936 ( \16606 , \13255 , \15566 );
and \U$15937 ( \16607 , \14795 , \14059 );
not \U$15938 ( \16608 , \14795 );
not \U$15939 ( \16609 , \15689 );
and \U$15940 ( \16610 , \16608 , \16609 );
nor \U$15941 ( \16611 , \16607 , \16610 );
nand \U$15942 ( \16612 , \14405 , \15043 );
nand \U$15943 ( \16613 , \16611 , \16612 );
not \U$15944 ( \16614 , \16613 );
nand \U$15945 ( \16615 , \16606 , \16614 );
and \U$15946 ( \16616 , \16605 , \16615 );
nor \U$15947 ( \16617 , \16606 , \16614 );
nor \U$15948 ( \16618 , \16616 , \16617 );
and \U$15949 ( \16619 , \16600 , \16618 );
not \U$15950 ( \16620 , \13506 );
not \U$15951 ( \16621 , \13583 );
nand \U$15952 ( \16622 , \16621 , \15564 );
nand \U$15953 ( \16623 , \16620 , \16622 );
nand \U$15954 ( \16624 , \15566 , \13583 );
nand \U$15955 ( \16625 , \16623 , \13516 , \16624 );
not \U$15956 ( \16626 , \16625 );
not \U$15957 ( \16627 , \14405 );
and \U$15958 ( \16628 , \13583 , \15259 );
not \U$15959 ( \16629 , \13583 );
and \U$15960 ( \16630 , \16629 , \15260 );
nor \U$15961 ( \16631 , \16628 , \16630 );
not \U$15962 ( \16632 , \16631 );
or \U$15963 ( \16633 , \16627 , \16632 );
and \U$15964 ( \16634 , \15042 , \14059 );
not \U$15965 ( \16635 , \15042 );
not \U$15966 ( \16636 , \14066 );
and \U$15967 ( \16637 , \16635 , \16636 );
nor \U$15968 ( \16638 , \16634 , \16637 );
nand \U$15969 ( \16639 , \16633 , \16638 );
not \U$15970 ( \16640 , \16639 );
and \U$15971 ( \16641 , \16626 , \16640 );
and \U$15972 ( \16642 , \16625 , \16639 );
nor \U$15973 ( \16643 , \16641 , \16642 );
not \U$15974 ( \16644 , \16643 );
not \U$15975 ( \16645 , \15762 );
not \U$15976 ( \16646 , \15592 );
or \U$15977 ( \16647 , \16645 , \16646 );
or \U$15978 ( \16648 , \13566 , \15347 );
nand \U$15979 ( \16649 , \16647 , \16648 );
and \U$15980 ( \16650 , \13515 , \15639 );
not \U$15981 ( \16651 , \13515 );
and \U$15982 ( \16652 , \16651 , \15566 );
or \U$15983 ( \16653 , \16650 , \16652 );
nor \U$15984 ( \16654 , \16653 , \13512 );
nor \U$15985 ( \16655 , \16649 , \16654 );
not \U$15986 ( \16656 , \16655 );
or \U$15987 ( \16657 , \16644 , \16656 );
not \U$15988 ( \16658 , \15639 );
nand \U$15989 ( \16659 , \16658 , \16631 , \13794 );
nand \U$15990 ( \16660 , \16659 , \15921 );
not \U$15991 ( \16661 , \16631 );
or \U$15992 ( \16662 , \16661 , \13795 );
nand \U$15993 ( \16663 , \16662 , \14404 );
and \U$15994 ( \16664 , \13513 , \15712 );
not \U$15995 ( \16665 , \16622 );
nor \U$15996 ( \16666 , \16664 , \16665 );
and \U$15997 ( \16667 , \16660 , \16663 , \16666 );
nand \U$15998 ( \16668 , \16657 , \16667 );
not \U$15999 ( \16669 , \16643 );
not \U$16000 ( \16670 , \16655 );
nand \U$16001 ( \16671 , \16669 , \16670 );
and \U$16002 ( \16672 , \16668 , \16671 );
not \U$16003 ( \16673 , \16625 );
nand \U$16004 ( \16674 , \16673 , \16639 );
nor \U$16005 ( \16675 , \16672 , \16674 );
xor \U$16006 ( \16676 , \16613 , \16606 );
xor \U$16007 ( \16677 , \16676 , \16604 );
or \U$16008 ( \16678 , \16675 , \16677 );
nand \U$16009 ( \16679 , \16668 , \16671 , \16674 );
nand \U$16010 ( \16680 , \16678 , \16679 );
nor \U$16011 ( \16681 , \16619 , \16680 );
nor \U$16012 ( \16682 , \16600 , \16618 );
or \U$16013 ( \16683 , \16681 , \16682 );
xor \U$16014 ( \16684 , \16545 , \16558 );
xor \U$16015 ( \16685 , \16684 , \16561 );
not \U$16016 ( \16686 , \16597 );
not \U$16017 ( \16687 , \16580 );
not \U$16018 ( \16688 , \16687 );
or \U$16019 ( \16689 , \16686 , \16688 );
not \U$16020 ( \16690 , \16589 );
nand \U$16021 ( \16691 , \16690 , \16593 );
nand \U$16022 ( \16692 , \16689 , \16691 );
nand \U$16023 ( \16693 , \16685 , \16692 );
nand \U$16024 ( \16694 , \16683 , \16693 );
not \U$16025 ( \16695 , \16685 );
not \U$16026 ( \16696 , \16692 );
nand \U$16027 ( \16697 , \16695 , \16696 );
nand \U$16028 ( \16698 , \16694 , \16697 );
nand \U$16029 ( \16699 , \16570 , \16698 );
nand \U$16030 ( \16700 , \16567 , \16699 );
not \U$16031 ( \16701 , \16700 );
or \U$16032 ( \16702 , \16520 , \16701 );
not \U$16033 ( \16703 , \16472 );
not \U$16034 ( \16704 , \16518 );
nand \U$16035 ( \16705 , \16703 , \16704 );
nand \U$16036 ( \16706 , \16702 , \16705 );
not \U$16037 ( \16707 , \16706 );
or \U$16038 ( \16708 , \16426 , \16460 );
and \U$16039 ( \16709 , \16467 , \16708 );
and \U$16040 ( \16710 , \16426 , \16460 );
nor \U$16041 ( \16711 , \16709 , \16710 );
not \U$16042 ( \16712 , \16711 );
not \U$16043 ( \16713 , \16418 );
not \U$16044 ( \16714 , \16379 );
or \U$16045 ( \16715 , \16713 , \16714 );
or \U$16046 ( \16716 , \16379 , \16418 );
nand \U$16047 ( \16717 , \16715 , \16716 );
and \U$16048 ( \16718 , \16717 , \16377 );
not \U$16049 ( \16719 , \16717 );
not \U$16050 ( \16720 , \16377 );
and \U$16051 ( \16721 , \16719 , \16720 );
nor \U$16052 ( \16722 , \16718 , \16721 );
not \U$16053 ( \16723 , \16722 );
or \U$16054 ( \16724 , \16712 , \16723 );
or \U$16055 ( \16725 , \16722 , \16711 );
nand \U$16056 ( \16726 , \16724 , \16725 );
not \U$16057 ( \16727 , \16726 );
or \U$16058 ( \16728 , \16707 , \16727 );
not \U$16059 ( \16729 , \16711 );
nand \U$16060 ( \16730 , \16729 , \16722 );
nand \U$16061 ( \16731 , \16728 , \16730 );
nand \U$16062 ( \16732 , \16425 , \16731 );
nand \U$16063 ( \16733 , \16284 , \16363 );
nand \U$16064 ( \16734 , \16371 , \16423 );
nand \U$16065 ( \16735 , \16732 , \16733 , \16734 );
nand \U$16066 ( \16736 , \16282 , \16366 , \15954 , \16735 );
nand \U$16067 ( \16737 , \16278 , \16736 );
nor \U$16068 ( \16738 , \15819 , \15821 );
not \U$16069 ( \16739 , \16738 );
nand \U$16070 ( \16740 , \15670 , \16739 );
nor \U$16071 ( \16741 , \16740 , \15874 );
and \U$16072 ( \16742 , \16737 , \16741 , \15188 );
nand \U$16073 ( \16743 , \15171 , \15175 , \15151 );
nand \U$16074 ( \16744 , \14726 , \14917 );
not \U$16075 ( \16745 , \15185 );
not \U$16076 ( \16746 , \15183 );
nand \U$16077 ( \16747 , \16745 , \16746 );
and \U$16078 ( \16748 , \16743 , \16744 , \16747 );
nor \U$16079 ( \16749 , \14924 , \15145 );
nand \U$16080 ( \16750 , \16749 , \14919 );
and \U$16081 ( \16751 , \16748 , \16750 );
buf \U$16082 ( \16752 , \16747 );
and \U$16083 ( \16753 , \16752 , \15187 );
nor \U$16084 ( \16754 , \16751 , \16753 );
nor \U$16085 ( \16755 , \16742 , \16754 );
nand \U$16086 ( \16756 , \15888 , \16755 );
nand \U$16087 ( \16757 , \14217 , \14223 );
nand \U$16088 ( \16758 , \14191 , \14185 );
nand \U$16089 ( \16759 , \14197 , \16758 );
nor \U$16090 ( \16760 , \16757 , \16759 );
and \U$16091 ( \16761 , \14285 , \14348 , \14355 );
and \U$16092 ( \16762 , \16760 , \16761 , \14369 );
nand \U$16093 ( \16763 , \16756 , \16762 );
not \U$16094 ( \16764 , \14369 );
not \U$16095 ( \16765 , \14348 );
not \U$16096 ( \16766 , \14355 );
nor \U$16097 ( \16767 , \14237 , \14284 );
not \U$16098 ( \16768 , \16767 );
or \U$16099 ( \16769 , \16766 , \16768 );
or \U$16100 ( \16770 , \14350 , \14354 );
nand \U$16101 ( \16771 , \16769 , \16770 );
not \U$16102 ( \16772 , \16771 );
or \U$16103 ( \16773 , \16765 , \16772 );
or \U$16104 ( \16774 , \14347 , \14328 );
nand \U$16105 ( \16775 , \16773 , \16774 );
not \U$16106 ( \16776 , \16775 );
or \U$16107 ( \16777 , \16764 , \16776 );
or \U$16108 ( \16778 , \14359 , \14368 );
nand \U$16109 ( \16779 , \16777 , \16778 );
not \U$16110 ( \16780 , \16779 );
nand \U$16111 ( \16781 , \14371 , \16763 , \16780 );
not \U$16112 ( \16782 , \16781 );
or \U$16113 ( \16783 , \12716 , \16782 );
nand \U$16114 ( \16784 , \12698 , \12714 );
not \U$16115 ( \16785 , \12703 );
not \U$16116 ( \16786 , \12709 );
or \U$16117 ( \16787 , \16785 , \16786 );
nand \U$16118 ( \16788 , \16787 , \12710 );
not \U$16119 ( \16789 , \16788 );
and \U$16120 ( \16790 , \12711 , \12713 );
and \U$16121 ( \16791 , \12701 , \12703 );
nor \U$16122 ( \16792 , \16790 , \16791 );
not \U$16123 ( \16793 , \16792 );
or \U$16124 ( \16794 , \16789 , \16793 );
or \U$16125 ( \16795 , \16792 , \16788 );
nand \U$16126 ( \16796 , \16794 , \16795 );
not \U$16127 ( \16797 , RIaaa89a8_588);
nand \U$16128 ( \16798 , \16797 , RIaaa91a0_605);
nor \U$16129 ( \16799 , \16798 , \11810 );
nand \U$16130 ( \16800 , \16799 , RIaaa90b0_603);
not \U$16131 ( \16801 , \16800 );
nand \U$16132 ( \16802 , \16801 , RIaaa9218_606);
not \U$16133 ( \16803 , \16802 );
nand \U$16134 ( \16804 , \16803 , RIaaa9290_607);
nor \U$16135 ( \16805 , \16804 , \11757 );
and \U$16136 ( \16806 , \16805 , RIaaa9380_609);
nand \U$16137 ( \16807 , \16806 , RIaaa93f8_610);
not \U$16138 ( \16808 , RIaaa9038_602);
and \U$16139 ( \16809 , \16807 , \16808 );
buf \U$16140 ( \16810 , \12005 );
nor \U$16141 ( \16811 , \16807 , \16808 );
or \U$16142 ( \16812 , \16811 , RIaaa9470_611);
nand \U$16143 ( \16813 , \16811 , RIaaa9470_611);
nand \U$16144 ( \16814 , \16812 , \16813 );
and \U$16145 ( \16815 , \16810 , \16814 );
not \U$16146 ( \16816 , \16813 );
or \U$16147 ( \16817 , \16816 , RIaaa94e8_612);
not \U$16148 ( \16818 , \16806 );
or \U$16149 ( \16819 , \16818 , \11368 );
nand \U$16150 ( \16820 , \16817 , \16819 );
and \U$16151 ( \16821 , \12066 , \16820 );
nor \U$16152 ( \16822 , \16815 , \16821 );
not \U$16153 ( \16823 , \16822 );
nor \U$16154 ( \16824 , \16809 , \16823 , \16811 );
buf \U$16155 ( \16825 , \12113 );
not \U$16156 ( \16826 , \16825 );
and \U$16157 ( \16827 , \16824 , \16826 );
buf \U$16158 ( \16828 , \13474 );
and \U$16159 ( \16829 , \11808 , RIaaa89a8_588);
not \U$16160 ( \16830 , \16798 );
nor \U$16161 ( \16831 , \16829 , \16830 );
nand \U$16162 ( \16832 , \16828 , \16831 );
and \U$16163 ( \16833 , \13478 , \16832 );
not \U$16164 ( \16834 , RIaaa9128_604);
not \U$16165 ( \16835 , \16798 );
or \U$16166 ( \16836 , \16834 , \16835 );
or \U$16167 ( \16837 , \16798 , RIaaa9128_604);
nand \U$16168 ( \16838 , \16836 , \16837 );
not \U$16169 ( \16839 , \13489 );
or \U$16170 ( \16840 , \16838 , \16839 );
or \U$16171 ( \16841 , \16799 , RIaaa90b0_603);
nand \U$16172 ( \16842 , \16841 , \16800 );
not \U$16173 ( \16843 , \16842 );
or \U$16174 ( \16844 , \12730 , \16843 );
or \U$16175 ( \16845 , \16831 , \16828 );
nand \U$16176 ( \16846 , \16840 , \16844 , \16845 );
nor \U$16177 ( \16847 , \16833 , \16846 );
nand \U$16178 ( \16848 , \16839 , \16838 );
and \U$16179 ( \16849 , \16848 , \16842 );
not \U$16180 ( \16850 , \16848 );
not \U$16181 ( \16851 , \16842 );
and \U$16182 ( \16852 , \16850 , \16851 );
nor \U$16183 ( \16853 , \16852 , \12730 );
nor \U$16184 ( \16854 , \16849 , \16853 );
or \U$16185 ( \16855 , \16847 , \16854 );
buf \U$16186 ( \16856 , \11669 );
not \U$16187 ( \16857 , \16856 );
not \U$16188 ( \16858 , RIaaa9218_606);
not \U$16189 ( \16859 , \16800 );
or \U$16190 ( \16860 , \16858 , \16859 );
or \U$16191 ( \16861 , \16800 , RIaaa9218_606);
nand \U$16192 ( \16862 , \16860 , \16861 );
or \U$16193 ( \16863 , \16857 , \16862 );
nand \U$16194 ( \16864 , \16855 , \16863 );
buf \U$16195 ( \16865 , \11721 );
not \U$16196 ( \16866 , \16865 );
not \U$16197 ( \16867 , \16802 );
not \U$16198 ( \16868 , RIaaa9290_607);
and \U$16199 ( \16869 , \16867 , \16868 );
and \U$16200 ( \16870 , \16802 , RIaaa9290_607);
nor \U$16201 ( \16871 , \16869 , \16870 );
not \U$16202 ( \16872 , \16871 );
and \U$16203 ( \16873 , \16866 , \16872 );
and \U$16204 ( \16874 , \16857 , \16862 );
nor \U$16205 ( \16875 , \16873 , \16874 );
and \U$16206 ( \16876 , \16864 , \16875 );
and \U$16207 ( \16877 , \16865 , \16871 );
buf \U$16208 ( \16878 , \11754 );
not \U$16209 ( \16879 , \16804 );
not \U$16210 ( \16880 , RIaaa9308_608);
and \U$16211 ( \16881 , \16879 , \16880 );
and \U$16212 ( \16882 , \16804 , RIaaa9308_608);
nor \U$16213 ( \16883 , \16881 , \16882 );
and \U$16214 ( \16884 , \16878 , \16883 );
buf \U$16215 ( \16885 , \11939 );
not \U$16216 ( \16886 , \16885 );
or \U$16217 ( \16887 , \16805 , RIaaa9380_609);
nand \U$16218 ( \16888 , \16887 , \16818 );
and \U$16219 ( \16889 , \16886 , \16888 );
nor \U$16220 ( \16890 , \16877 , \16884 , \16889 );
not \U$16221 ( \16891 , \16890 );
nor \U$16222 ( \16892 , \16876 , \16891 );
or \U$16223 ( \16893 , \16889 , \16878 , \16883 );
or \U$16224 ( \16894 , \16886 , \16888 );
nand \U$16225 ( \16895 , \16893 , \16894 );
or \U$16226 ( \16896 , \16892 , \16895 );
not \U$16227 ( \16897 , RIaaa93f8_610);
not \U$16228 ( \16898 , \16818 );
or \U$16229 ( \16899 , \16897 , \16898 );
or \U$16230 ( \16900 , \16818 , RIaaa93f8_610);
nand \U$16231 ( \16901 , \16899 , \16900 );
nand \U$16232 ( \16902 , \16896 , \16901 );
or \U$16233 ( \16903 , \16892 , \16895 , \16901 );
not \U$16234 ( \16904 , \12168 );
nand \U$16235 ( \16905 , \16903 , \16904 );
and \U$16236 ( \16906 , \16902 , \16905 );
and \U$16237 ( \16907 , \16822 , \16826 );
nor \U$16238 ( \16908 , \16907 , \16824 );
nor \U$16239 ( \16909 , \16906 , \16908 );
or \U$16240 ( \16910 , \16821 , \16810 , \16814 );
or \U$16241 ( \16911 , \12066 , \16820 );
nand \U$16242 ( \16912 , \16910 , \16911 );
nor \U$16243 ( \16913 , \16827 , \16909 , \16912 );
not \U$16244 ( \16914 , RIaaa95d8_614);
not \U$16245 ( \16915 , \16819 );
or \U$16246 ( \16916 , \16914 , \16915 );
or \U$16247 ( \16917 , \16819 , RIaaa95d8_614);
nand \U$16248 ( \16918 , \16916 , \16917 );
nor \U$16249 ( \16919 , RIaaa8e58_598, RIaaa8fc0_601);
nor \U$16250 ( \16920 , RIaaa8ed0_599, RIaaa8f48_600);
and \U$16251 ( \16921 , \16919 , \16920 , \11374 );
not \U$16252 ( \16922 , \16921 );
not \U$16253 ( \16923 , \16922 );
and \U$16254 ( \16924 , \16923 , RIaa97e78_18);
not \U$16255 ( \16925 , RIaa981c0_25);
not \U$16256 ( \16926 , RIaaa8e58_598);
nor \U$16257 ( \16927 , \16926 , RIaaa8fc0_601);
nor \U$16258 ( \16928 , RIaaa8ed0_599, RIaaa8f48_600);
and \U$16259 ( \16929 , \16927 , \16928 );
not \U$16260 ( \16930 , \16929 );
not \U$16261 ( \16931 , \16930 );
not \U$16262 ( \16932 , \16931 );
or \U$16263 ( \16933 , \16925 , \16932 );
nand \U$16264 ( \16934 , \16933 , \12194 );
nor \U$16265 ( \16935 , \16924 , \16934 );
not \U$16266 ( \16936 , RIaaa8ed0_599);
not \U$16267 ( \16937 , RIaaa8fc0_601);
nand \U$16268 ( \16938 , \16936 , \16937 , RIaaa8f48_600, RIaaa8e58_598);
not \U$16269 ( \16939 , \16938 );
buf \U$16270 ( \16940 , \16939 );
buf \U$16271 ( \16941 , \16940 );
and \U$16272 ( \16942 , \16941 , RIaa983a0_29);
not \U$16273 ( \16943 , RIaaa8ed0_599);
nor \U$16274 ( \16944 , \16943 , RIaaa8f48_600);
nand \U$16275 ( \16945 , RIaaa8e58_598, RIaaa8fc0_601);
not \U$16276 ( \16946 , \16945 );
and \U$16277 ( \16947 , \16944 , \16946 );
buf \U$16278 ( \16948 , \16947 );
buf \U$16279 ( \16949 , \16948 );
and \U$16280 ( \16950 , \16949 , RIaa98328_28);
nor \U$16281 ( \16951 , \16942 , \16950 );
nand \U$16282 ( \16952 , \16944 , \16919 );
not \U$16283 ( \16953 , \16952 );
not \U$16284 ( \16954 , \16953 );
not \U$16285 ( \16955 , \16954 );
and \U$16286 ( \16956 , \16955 , RIaa98580_33);
not \U$16287 ( \16957 , RIaaa8ed0_599);
nor \U$16288 ( \16958 , \16957 , RIaaa8f48_600);
and \U$16289 ( \16959 , \16958 , \16927 );
buf \U$16290 ( \16960 , \16959 );
and \U$16291 ( \16961 , \16960 , RIaa982b0_27);
nor \U$16292 ( \16962 , \16956 , \16961 );
not \U$16293 ( \16963 , RIaaa8fc0_601);
nand \U$16294 ( \16964 , \16963 , RIaaa8ed0_599, RIaaa8f48_600, RIaaa8e58_598);
not \U$16295 ( \16965 , \16964 );
buf \U$16296 ( \16966 , \16965 );
and \U$16297 ( \16967 , \16966 , RIaa980d0_23);
nor \U$16298 ( \16968 , \11405 , \16945 );
buf \U$16299 ( \16969 , \16968 );
and \U$16300 ( \16970 , \16969 , RIaa98148_24);
nor \U$16301 ( \16971 , \16967 , \16970 );
nand \U$16302 ( \16972 , \16935 , \16951 , \16962 , \16971 );
not \U$16303 ( \16973 , \11409 );
nand \U$16304 ( \16974 , \16973 , \16920 );
not \U$16305 ( \16975 , \16974 );
not \U$16306 ( \16976 , \16975 );
not \U$16307 ( \16977 , \16976 );
and \U$16308 ( \16978 , \16977 , RIaa97ef0_19);
and \U$16309 ( \16979 , \16973 , \16958 );
not \U$16310 ( \16980 , \16979 );
not \U$16311 ( \16981 , \16980 );
buf \U$16312 ( \16982 , \16981 );
and \U$16313 ( \16983 , \16982 , RIaa98508_32);
nor \U$16314 ( \16984 , \16978 , \16983 );
not \U$16315 ( \16985 , RIaaa8f48_600);
nor \U$16316 ( \16986 , \16985 , RIaaa8ed0_599);
nor \U$16317 ( \16987 , RIaaa8e58_598, RIaaa8fc0_601);
and \U$16318 ( \16988 , \16986 , \16987 );
buf \U$16319 ( \16989 , \16988 );
not \U$16320 ( \16990 , \16989 );
not \U$16321 ( \16991 , \16990 );
and \U$16322 ( \16992 , \16991 , RIaa97fe0_21);
not \U$16323 ( \16993 , RIaaa8e58_598);
not \U$16324 ( \16994 , RIaaa8ed0_599);
nand \U$16325 ( \16995 , \16993 , \16994 , RIaaa8fc0_601, RIaaa8f48_600);
not \U$16326 ( \16996 , \16995 );
and \U$16327 ( \16997 , \16996 , RIaa98058_22);
nor \U$16328 ( \16998 , \16992 , \16997 );
not \U$16329 ( \16999 , \11405 );
and \U$16330 ( \17000 , \16999 , \16987 );
not \U$16331 ( \17001 , \17000 );
not \U$16332 ( \17002 , \17001 );
and \U$16333 ( \17003 , \17002 , RIaa98490_31);
and \U$16334 ( \17004 , \16973 , \16999 );
not \U$16335 ( \17005 , \17004 );
not \U$16336 ( \17006 , \17005 );
buf \U$16337 ( \17007 , \17006 );
and \U$16338 ( \17008 , \17007 , RIaa985f8_34);
nor \U$16339 ( \17009 , \17003 , \17008 );
and \U$16340 ( \17010 , \16946 , \16928 );
not \U$16341 ( \17011 , \17010 );
not \U$16342 ( \17012 , \17011 );
and \U$16343 ( \17013 , \17012 , RIaa98238_26);
not \U$16344 ( \17014 , RIaaa8ed0_599);
nand \U$16345 ( \17015 , \17014 , RIaaa8e58_598, RIaaa8fc0_601, RIaaa8f48_600);
not \U$16346 ( \17016 , \17015 );
and \U$16347 ( \17017 , \17016 , RIaa98418_30);
nor \U$16348 ( \17018 , \17013 , \17017 );
nand \U$16349 ( \17019 , \16984 , \16998 , \17009 , \17018 );
nor \U$16350 ( \17020 , \16972 , \17019 );
and \U$16351 ( \17021 , \12237 , \16918 , \17020 );
not \U$16352 ( \17022 , \12238 );
not \U$16353 ( \17023 , \16918 );
and \U$16354 ( \17024 , \17022 , \17023 );
not \U$16355 ( \17025 , \12730 );
and \U$16356 ( \17026 , \16965 , RIaa9afb0_123);
and \U$16357 ( \17027 , \16969 , RIaa9b028_124);
nor \U$16358 ( \17028 , \17026 , \17027 );
and \U$16359 ( \17029 , \16960 , RIaa9b280_129);
not \U$16360 ( \17030 , \11475 );
nor \U$16361 ( \17031 , \17029 , \17030 );
nand \U$16362 ( \17032 , \16923 , RIaa9aec0_121);
nand \U$16363 ( \17033 , \17028 , \17031 , \17032 );
nand \U$16364 ( \17034 , \16979 , RIaa9b190_127);
nand \U$16365 ( \17035 , \16996 , RIaa9b550_135);
nand \U$16366 ( \17036 , \17006 , RIaa9b3e8_132);
nand \U$16367 ( \17037 , \17000 , RIaa9b208_128);
nand \U$16368 ( \17038 , \17034 , \17035 , \17036 , \17037 );
nor \U$16369 ( \17039 , \17033 , \17038 );
nand \U$16370 ( \17040 , \16931 , RIaa9b460_133);
nand \U$16371 ( \17041 , \16940 , RIaa9b370_131);
nand \U$16372 ( \17042 , \17016 , RIaa9b2f8_130);
nand \U$16373 ( \17043 , \17012 , RIaa9b4d8_134);
nand \U$16374 ( \17044 , \17040 , \17041 , \17042 , \17043 );
nand \U$16375 ( \17045 , \16977 , RIaa9ae48_120);
nand \U$16376 ( \17046 , \16989 , RIaa9b5c8_136);
nand \U$16377 ( \17047 , \16955 , RIaa9b0a0_125);
nand \U$16378 ( \17048 , \16948 , RIaa9b118_126);
nand \U$16379 ( \17049 , \17045 , \17046 , \17047 , \17048 );
nor \U$16380 ( \17050 , \17044 , \17049 );
nand \U$16381 ( \17051 , \17039 , \17050 );
not \U$16382 ( \17052 , \17051 );
or \U$16383 ( \17053 , \17025 , \17052 );
nand \U$16384 ( \17054 , \16975 , RIaa9c018_158);
nand \U$16385 ( \17055 , \16996 , RIaa9bfa0_157);
and \U$16386 ( \17056 , \16973 , \16958 );
nand \U$16387 ( \17057 , \17056 , RIaa9c270_163);
nand \U$16388 ( \17058 , \16988 , RIaa9bf28_156);
nand \U$16389 ( \17059 , \17054 , \17055 , \17057 , \17058 );
nand \U$16390 ( \17060 , \16947 , RIaa9c5b8_170);
not \U$16391 ( \17061 , \17015 );
nand \U$16392 ( \17062 , \17061 , RIaa9c3d8_166);
nand \U$16393 ( \17063 , \16959 , RIaa9be38_154);
nand \U$16394 ( \17064 , \17010 , RIaa9c4c8_168);
nand \U$16395 ( \17065 , \17060 , \17062 , \17063 , \17064 );
nor \U$16396 ( \17066 , \17059 , \17065 );
nand \U$16397 ( \17067 , \16921 , RIaa9c090_159);
and \U$16398 ( \17068 , \16953 , RIaa9c2e8_164);
not \U$16399 ( \17069 , \11769 );
nor \U$16400 ( \17070 , \17068 , \17069 );
nand \U$16401 ( \17071 , \16939 , RIaa9c360_165);
nand \U$16402 ( \17072 , \16968 , RIaa9c180_161);
nand \U$16403 ( \17073 , \17067 , \17070 , \17071 , \17072 );
nand \U$16404 ( \17074 , \17004 , RIaa9beb0_155);
nand \U$16405 ( \17075 , \16965 , RIaa9c1f8_162);
nand \U$16406 ( \17076 , \17000 , RIaa9c540_169);
nand \U$16407 ( \17077 , \16929 , RIaa9c450_167);
nand \U$16408 ( \17078 , \17074 , \17075 , \17076 , \17077 );
nor \U$16409 ( \17079 , \17073 , \17078 );
nand \U$16410 ( \17080 , \17066 , \17079 );
buf \U$16411 ( \17081 , \17080 );
and \U$16412 ( \17082 , \16828 , \17081 );
nand \U$16413 ( \17083 , \16975 , RIaa9c6a8_172);
nand \U$16414 ( \17084 , \17004 , RIaa9cdb0_187);
nand \U$16415 ( \17085 , \16988 , RIaa9cae0_181);
nand \U$16416 ( \17086 , \17000 , RIaa9c900_177);
nand \U$16417 ( \17087 , \17083 , \17084 , \17085 , \17086 );
nand \U$16418 ( \17088 , \16939 , RIaa9c9f0_179);
nand \U$16419 ( \17089 , \16959 , RIaa9cd38_186);
nand \U$16420 ( \17090 , \17061 , RIaa9cbd0_183);
nand \U$16421 ( \17091 , \17010 , RIaa9cb58_182);
nand \U$16422 ( \17092 , \17088 , \17089 , \17090 , \17091 );
nor \U$16423 ( \17093 , \17087 , \17092 );
nand \U$16424 ( \17094 , \16921 , RIaa9c798_174);
and \U$16425 ( \17095 , \16929 , RIaa9ca68_180);
not \U$16426 ( \17096 , \11869 );
nor \U$16427 ( \17097 , \17095 , \17096 );
nand \U$16428 ( \17098 , \16965 , RIaa9c630_171);
nand \U$16429 ( \17099 , \16947 , RIaa9c888_176);
nand \U$16430 ( \17100 , \17094 , \17097 , \17098 , \17099 );
nand \U$16431 ( \17101 , RIaaa8ed0_599, RIaaa8f48_600, RIaaa8e58_598, RIaaa8fc0_601);
not \U$16432 ( \17102 , \17101 );
not \U$16433 ( \17103 , \6268 );
and \U$16434 ( \17104 , \17102 , \17103 );
and \U$16435 ( \17105 , \16953 , RIaa9ccc0_185);
nor \U$16436 ( \17106 , \17104 , \17105 );
nand \U$16437 ( \17107 , \17056 , RIaa9cc48_184);
nand \U$16438 ( \17108 , \16996 , RIaa9c978_178);
nand \U$16439 ( \17109 , \17106 , \17107 , \17108 );
nor \U$16440 ( \17110 , \17100 , \17109 );
nand \U$16441 ( \17111 , \17093 , \17110 );
not \U$16442 ( \17112 , \17111 );
not \U$16443 ( \17113 , \17112 );
nor \U$16444 ( \17114 , \17082 , \13791 , \17113 );
nor \U$16445 ( \17115 , \16828 , \17081 );
and \U$16446 ( \17116 , \16959 , RIaa9ba78_146);
not \U$16447 ( \17117 , \11817 );
nor \U$16448 ( \17118 , \17116 , \17117 );
and \U$16449 ( \17119 , \16965 , RIaa9b988_144);
nor \U$16450 ( \17120 , \17101 , \6363 );
nor \U$16451 ( \17121 , \17119 , \17120 );
nand \U$16452 ( \17122 , \16921 , RIaa9b898_142);
nand \U$16453 ( \17123 , \17118 , \17121 , \17122 );
nand \U$16454 ( \17124 , \17056 , RIaa9b730_139);
nand \U$16455 ( \17125 , \17004 , RIaa9bbe0_149);
nand \U$16456 ( \17126 , \16996 , RIaa9bc58_150);
nand \U$16457 ( \17127 , \17000 , RIaa9b7a8_140);
nand \U$16458 ( \17128 , \17124 , \17125 , \17126 , \17127 );
nor \U$16459 ( \17129 , \17123 , \17128 );
nand \U$16460 ( \17130 , \16975 , RIaa9b820_141);
nand \U$16461 ( \17131 , \16953 , RIaa9b6b8_138);
nand \U$16462 ( \17132 , \16947 , RIaa9b640_137);
nand \U$16463 ( \17133 , \17010 , RIaa9bdc0_153);
nand \U$16464 ( \17134 , \17130 , \17131 , \17132 , \17133 );
nand \U$16465 ( \17135 , \16929 , RIaa9bd48_152);
nand \U$16466 ( \17136 , \16939 , RIaa9bb68_148);
nand \U$16467 ( \17137 , \16988 , RIaa9bcd0_151);
nand \U$16468 ( \17138 , \17061 , RIaa9baf0_147);
nand \U$16469 ( \17139 , \17135 , \17136 , \17137 , \17138 );
nor \U$16470 ( \17140 , \17134 , \17139 );
nand \U$16471 ( \17141 , \17129 , \17140 );
buf \U$16472 ( \17142 , \17141 );
not \U$16473 ( \17143 , \17142 );
nor \U$16474 ( \17144 , \17114 , \17115 , \17143 );
or \U$16475 ( \17145 , \17144 , \16839 );
or \U$16476 ( \17146 , \17114 , \17115 );
nand \U$16477 ( \17147 , \17146 , \17143 );
nand \U$16478 ( \17148 , \17145 , \17147 );
nand \U$16479 ( \17149 , \17053 , \17148 );
not \U$16480 ( \17150 , \17011 );
not \U$16481 ( \17151 , RIaa9a218_94);
not \U$16482 ( \17152 , \17151 );
and \U$16483 ( \17153 , \17150 , \17152 );
nor \U$16484 ( \17154 , \17153 , \11732 );
and \U$16485 ( \17155 , \16965 , RIaa99f48_88);
and \U$16486 ( \17156 , \16969 , RIaa9a038_90);
nor \U$16487 ( \17157 , \17155 , \17156 );
nand \U$16488 ( \17158 , \16923 , RIaa99fc0_89);
nand \U$16489 ( \17159 , \17154 , \17157 , \17158 );
nand \U$16490 ( \17160 , \17002 , RIaa9a3f8_98);
nand \U$16491 ( \17161 , \16960 , RIaa9a470_99);
nand \U$16492 ( \17162 , \17006 , RIaa9a5d8_102);
nand \U$16493 ( \17163 , \17016 , RIaa9a560_101);
nand \U$16494 ( \17164 , \17160 , \17161 , \17162 , \17163 );
nor \U$16495 ( \17165 , \17159 , \17164 );
nand \U$16496 ( \17166 , \16977 , RIaa99e58_86);
nand \U$16497 ( \17167 , \16981 , RIaa9a380_97);
nand \U$16498 ( \17168 , \16996 , RIaa9a128_92);
nand \U$16499 ( \17169 , \16989 , RIaa9a1a0_93);
nand \U$16500 ( \17170 , \17166 , \17167 , \17168 , \17169 );
nand \U$16501 ( \17171 , \16940 , RIaa9a4e8_100);
nand \U$16502 ( \17172 , \16948 , RIaa9a308_96);
nand \U$16503 ( \17173 , \16955 , RIaa9a290_95);
nand \U$16504 ( \17174 , \16931 , RIaa9a0b0_91);
nand \U$16505 ( \17175 , \17171 , \17172 , \17173 , \17174 );
nor \U$16506 ( \17176 , \17170 , \17175 );
nand \U$16507 ( \17177 , \17165 , \17176 );
not \U$16508 ( \17178 , \17177 );
and \U$16509 ( \17179 , \16878 , \17178 );
not \U$16510 ( \17180 , \17015 );
not \U$16511 ( \17181 , \11677 );
and \U$16512 ( \17182 , \17180 , \17181 );
not \U$16513 ( \17183 , \16976 );
and \U$16514 ( \17184 , \17183 , RIaa9a650_103);
nor \U$16515 ( \17185 , \17182 , \17184 );
not \U$16516 ( \17186 , \16979 );
nor \U$16517 ( \17187 , \17186 , \11691 );
not \U$16518 ( \17188 , RIaa9ace0_117);
nor \U$16519 ( \17189 , \17188 , \16995 );
nor \U$16520 ( \17190 , \17187 , \17189 );
nand \U$16521 ( \17191 , \17185 , \17190 );
not \U$16522 ( \17192 , \16947 );
not \U$16523 ( \17193 , \17192 );
not \U$16524 ( \17194 , \11704 );
and \U$16525 ( \17195 , \17193 , \17194 );
and \U$16526 ( \17196 , \16955 , RIaa9a8a8_108);
nor \U$16527 ( \17197 , \17195 , \17196 );
and \U$16528 ( \17198 , \16929 , RIaa9ad58_118);
nor \U$16529 ( \17199 , \16938 , \11707 );
nor \U$16530 ( \17200 , \17198 , \17199 );
nand \U$16531 ( \17201 , \17197 , \17200 );
nor \U$16532 ( \17202 , \17191 , \17201 );
not \U$16533 ( \17203 , \17000 );
not \U$16534 ( \17204 , \17203 );
not \U$16535 ( \17205 , \11710 );
and \U$16536 ( \17206 , \17204 , \17205 );
and \U$16537 ( \17207 , \17004 , RIaa9abf0_115);
nor \U$16538 ( \17208 , \17206 , \17207 );
nand \U$16539 ( \17209 , \16960 , RIaa9aa88_112);
nand \U$16540 ( \17210 , \17010 , RIaa9add0_119);
nand \U$16541 ( \17211 , \17208 , \17209 , \17210 );
nand \U$16542 ( \17212 , \16921 , RIaa9a6c8_104);
and \U$16543 ( \17213 , \16965 , RIaa9a7b8_106);
not \U$16544 ( \17214 , RIaa9a830_107);
nor \U$16545 ( \17215 , \17214 , \17101 );
nor \U$16546 ( \17216 , \17213 , \17215 );
and \U$16547 ( \17217 , \16988 , RIaa9ac68_116);
nor \U$16548 ( \17218 , \17217 , \11683 );
nand \U$16549 ( \17219 , \17212 , \17216 , \17218 );
nor \U$16550 ( \17220 , \17211 , \17219 );
nand \U$16551 ( \17221 , \17202 , \17220 );
not \U$16552 ( \17222 , \17221 );
not \U$16553 ( \17223 , \17222 );
not \U$16554 ( \17224 , \16865 );
or \U$16555 ( \17225 , \17223 , \17224 );
and \U$16556 ( \17226 , \16996 , RIaa99a98_78);
not \U$16557 ( \17227 , RIaa99660_69);
nor \U$16558 ( \17228 , \17227 , \16980 );
nor \U$16559 ( \17229 , \17226 , \17228 );
and \U$16560 ( \17230 , \16977 , RIaa99840_73);
and \U$16561 ( \17231 , \17016 , RIaa997c8_72);
nor \U$16562 ( \17232 , \17230 , \17231 );
nand \U$16563 ( \17233 , \17229 , \17232 );
nand \U$16564 ( \17234 , \16940 , RIaa99750_71);
nand \U$16565 ( \17235 , \16948 , RIaa99c78_82);
nand \U$16566 ( \17236 , \16931 , RIaa99b88_80);
nand \U$16567 ( \17237 , \16955 , RIaa99d68_84);
nand \U$16568 ( \17238 , \17234 , \17235 , \17236 , \17237 );
nor \U$16569 ( \17239 , \17233 , \17238 );
nand \U$16570 ( \17240 , \16923 , RIaa998b8_74);
and \U$16571 ( \17241 , \16965 , RIaa999a8_76);
nor \U$16572 ( \17242 , \17101 , \11548 );
nor \U$16573 ( \17243 , \17241 , \17242 );
and \U$16574 ( \17244 , \16989 , RIaa99b10_79);
not \U$16575 ( \17245 , \11551 );
nor \U$16576 ( \17246 , \17244 , \17245 );
nand \U$16577 ( \17247 , \17240 , \17243 , \17246 );
nand \U$16578 ( \17248 , \17006 , RIaa99de0_85);
nand \U$16579 ( \17249 , \17012 , RIaa99c00_81);
nand \U$16580 ( \17250 , \17000 , RIaa996d8_70);
nand \U$16581 ( \17251 , \16960 , RIaa99cf0_83);
nand \U$16582 ( \17252 , \17248 , \17249 , \17250 , \17251 );
nor \U$16583 ( \17253 , \17247 , \17252 );
nand \U$16584 ( \17254 , \17239 , \17253 );
not \U$16585 ( \17255 , \17254 );
nand \U$16586 ( \17256 , \17255 , \16886 );
nand \U$16587 ( \17257 , \17225 , \17256 );
nor \U$16588 ( \17258 , \17179 , \17257 );
not \U$16589 ( \17259 , \17005 );
not \U$16590 ( \17260 , \11640 );
and \U$16591 ( \17261 , \17259 , \17260 );
nor \U$16592 ( \17262 , \17203 , \11637 );
nor \U$16593 ( \17263 , \17261 , \17262 );
not \U$16594 ( \17264 , \17011 );
not \U$16595 ( \17265 , RIaa9d620_205);
not \U$16596 ( \17266 , \17265 );
and \U$16597 ( \17267 , \17264 , \17266 );
and \U$16598 ( \17268 , \16960 , RIaa9d2d8_198);
nor \U$16599 ( \17269 , \17267 , \17268 );
nand \U$16600 ( \17270 , \17263 , \17269 );
nand \U$16601 ( \17271 , \16921 , RIaa9d080_193);
and \U$16602 ( \17272 , \17061 , RIaa9d350_199);
nor \U$16603 ( \17273 , \17272 , \11632 );
nand \U$16604 ( \17274 , \16965 , RIaa9cf18_190);
nand \U$16605 ( \17275 , \16969 , RIaa9cf90_191);
nand \U$16606 ( \17276 , \17271 , \17273 , \17274 , \17275 );
nor \U$16607 ( \17277 , \17270 , \17276 );
nand \U$16608 ( \17278 , \17183 , RIaa9d008_192);
nand \U$16609 ( \17279 , \16979 , RIaa9d1e8_196);
nand \U$16610 ( \17280 , \16996 , RIaa9d4b8_202);
nand \U$16611 ( \17281 , \16988 , RIaa9d530_203);
nand \U$16612 ( \17282 , \17278 , \17279 , \17280 , \17281 );
and \U$16613 ( \17283 , \16929 , RIaa9d5a8_204);
and \U$16614 ( \17284 , \16939 , RIaa9d3c8_200);
nor \U$16615 ( \17285 , \17283 , \17284 );
and \U$16616 ( \17286 , \16953 , RIaa9d170_195);
and \U$16617 ( \17287 , \16947 , RIaa9d0f8_194);
nor \U$16618 ( \17288 , \17286 , \17287 );
nand \U$16619 ( \17289 , \17285 , \17288 );
nor \U$16620 ( \17290 , \17282 , \17289 );
nand \U$16621 ( \17291 , \17277 , \17290 );
buf \U$16622 ( \17292 , \17291 );
not \U$16623 ( \17293 , \17292 );
and \U$16624 ( \17294 , \16856 , \17293 );
and \U$16625 ( \17295 , \17025 , \17052 );
nor \U$16626 ( \17296 , \17294 , \17295 );
and \U$16627 ( \17297 , \17149 , \17258 , \17296 );
or \U$16628 ( \17298 , \17179 , \16865 , \17222 );
or \U$16629 ( \17299 , \16878 , \17178 );
nand \U$16630 ( \17300 , \17298 , \17299 );
and \U$16631 ( \17301 , \17300 , \17256 );
and \U$16632 ( \17302 , \16885 , \17254 );
nor \U$16633 ( \17303 , \17301 , \17302 );
nand \U$16634 ( \17304 , \17258 , \16857 , \17292 );
nand \U$16635 ( \17305 , \17303 , \17304 );
nor \U$16636 ( \17306 , \17297 , \17305 );
not \U$16637 ( \17307 , RIaa992a0_61);
nor \U$16638 ( \17308 , \17307 , \16995 );
not \U$16639 ( \17309 , RIaa99570_67);
nor \U$16640 ( \17310 , \17309 , \16980 );
nor \U$16641 ( \17311 , \17308 , \17310 );
and \U$16642 ( \17312 , \17006 , RIaa994f8_66);
not \U$16643 ( \17313 , RIaa995e8_68);
nor \U$16644 ( \17314 , \17313 , \17001 );
nor \U$16645 ( \17315 , \17312 , \17314 );
nand \U$16646 ( \17316 , \17311 , \17315 );
nand \U$16647 ( \17317 , \16940 , RIaa991b0_59);
nand \U$16648 ( \17318 , \16948 , RIaa990c0_57);
nand \U$16649 ( \17319 , \16931 , RIaa99390_63);
nand \U$16650 ( \17320 , \16955 , RIaa99138_58);
nand \U$16651 ( \17321 , \17317 , \17318 , \17319 , \17320 );
nor \U$16652 ( \17322 , \17316 , \17321 );
and \U$16653 ( \17323 , \16965 , RIaa98fd0_55);
not \U$16654 ( \17324 , RIaa99048_56);
nor \U$16655 ( \17325 , \17324 , \17101 );
nor \U$16656 ( \17326 , \17323 , \17325 );
and \U$16657 ( \17327 , \17016 , RIaa99228_60);
not \U$16658 ( \17328 , \12137 );
nor \U$16659 ( \17329 , \17327 , \17328 );
nand \U$16660 ( \17330 , \16923 , RIaa98ee0_53);
nand \U$16661 ( \17331 , \17326 , \17329 , \17330 );
and \U$16662 ( \17332 , \16977 , RIaa98e68_52);
and \U$16663 ( \17333 , \16960 , RIaa99480_65);
nor \U$16664 ( \17334 , \17332 , \17333 );
not \U$16665 ( \17335 , \17011 );
not \U$16666 ( \17336 , RIaa99408_64);
not \U$16667 ( \17337 , \17336 );
and \U$16668 ( \17338 , \17335 , \17337 );
and \U$16669 ( \17339 , \16989 , RIaa99318_62);
nor \U$16670 ( \17340 , \17338 , \17339 );
nand \U$16671 ( \17341 , \17334 , \17340 );
nor \U$16672 ( \17342 , \17331 , \17341 );
nand \U$16673 ( \17343 , \17322 , \17342 );
not \U$16674 ( \17344 , \17343 );
and \U$16675 ( \17345 , \12168 , \17344 );
not \U$16676 ( \17346 , \16922 );
not \U$16677 ( \17347 , \1750 );
and \U$16678 ( \17348 , \17346 , \17347 );
not \U$16679 ( \17349 , RIaa9e1d8_230);
or \U$16680 ( \17350 , \16930 , \17349 );
nand \U$16681 ( \17351 , \17350 , \11963 );
nor \U$16682 ( \17352 , \17348 , \17351 );
and \U$16683 ( \17353 , \16941 , RIaa9e3b8_234);
and \U$16684 ( \17354 , \16949 , RIaa9e340_233);
nor \U$16685 ( \17355 , \17353 , \17354 );
and \U$16686 ( \17356 , \16955 , RIaa9e598_238);
and \U$16687 ( \17357 , \16960 , RIaa9e2c8_232);
nor \U$16688 ( \17358 , \17356 , \17357 );
and \U$16689 ( \17359 , \16966 , RIaa9e0e8_228);
and \U$16690 ( \17360 , \16969 , RIaa9e160_229);
nor \U$16691 ( \17361 , \17359 , \17360 );
nand \U$16692 ( \17362 , \17352 , \17355 , \17358 , \17361 );
and \U$16693 ( \17363 , \16982 , RIaa9e520_237);
and \U$16694 ( \17364 , \17007 , RIaa9e610_239);
nor \U$16695 ( \17365 , \17363 , \17364 );
not \U$16696 ( \17366 , \17001 );
not \U$16697 ( \17367 , RIaa9e4a8_236);
not \U$16698 ( \17368 , \17367 );
and \U$16699 ( \17369 , \17366 , \17368 );
and \U$16700 ( \17370 , \16996 , RIaa9e070_227);
nor \U$16701 ( \17371 , \17369 , \17370 );
and \U$16702 ( \17372 , \16977 , RIaa9de90_223);
not \U$16703 ( \17373 , RIaa9dff8_226);
nor \U$16704 ( \17374 , \17373 , \16990 );
nor \U$16705 ( \17375 , \17372 , \17374 );
and \U$16706 ( \17376 , \17012 , RIaa9e250_231);
and \U$16707 ( \17377 , \17016 , RIaa9e430_235);
nor \U$16708 ( \17378 , \17376 , \17377 );
nand \U$16709 ( \17379 , \17365 , \17371 , \17375 , \17378 );
nor \U$16710 ( \17380 , \17362 , \17379 );
not \U$16711 ( \17381 , \17380 );
not \U$16712 ( \17382 , \16810 );
or \U$16713 ( \17383 , \17381 , \17382 );
and \U$16714 ( \17384 , \16923 , RIaa986e8_36);
not \U$16715 ( \17385 , RIaa989b8_42);
not \U$16716 ( \17386 , \16931 );
or \U$16717 ( \17387 , \17385 , \17386 );
nand \U$16718 ( \17388 , \17387 , \12023 );
nor \U$16719 ( \17389 , \17384 , \17388 );
and \U$16720 ( \17390 , \16960 , RIaa98c88_48);
and \U$16721 ( \17391 , \16941 , RIaa98b98_46);
nor \U$16722 ( \17392 , \17390 , \17391 );
and \U$16723 ( \17393 , \16955 , RIaa98b20_45);
and \U$16724 ( \17394 , \16949 , RIaa98aa8_44);
nor \U$16725 ( \17395 , \17393 , \17394 );
and \U$16726 ( \17396 , \16966 , RIaa987d8_38);
and \U$16727 ( \17397 , \16969 , RIaa98850_39);
nor \U$16728 ( \17398 , \17396 , \17397 );
nand \U$16729 ( \17399 , \17389 , \17392 , \17395 , \17398 );
and \U$16730 ( \17400 , \16982 , RIaa98df0_51);
and \U$16731 ( \17401 , \16996 , RIaa98940_41);
nor \U$16732 ( \17402 , \17400 , \17401 );
and \U$16733 ( \17403 , \16977 , RIaa98670_35);
and \U$16734 ( \17404 , \17016 , RIaa98c10_47);
nor \U$16735 ( \17405 , \17403 , \17404 );
and \U$16736 ( \17406 , \17002 , RIaa98d78_50);
and \U$16737 ( \17407 , \17007 , RIaa98d00_49);
nor \U$16738 ( \17408 , \17406 , \17407 );
and \U$16739 ( \17409 , \16991 , RIaa988c8_40);
and \U$16740 ( \17410 , \17012 , RIaa98a30_43);
nor \U$16741 ( \17411 , \17409 , \17410 );
nand \U$16742 ( \17412 , \17402 , \17405 , \17408 , \17411 );
nor \U$16743 ( \17413 , \17399 , \17412 );
nand \U$16744 ( \17414 , \12066 , \17413 );
nand \U$16745 ( \17415 , \17383 , \17414 );
nand \U$16746 ( \17416 , \16923 , RIaa9dad0_215);
nand \U$16747 ( \17417 , \16960 , RIaa9d698_206);
and \U$16748 ( \17418 , \17416 , \17417 , \12070 );
and \U$16749 ( \17419 , \16955 , RIaa9d788_208);
and \U$16750 ( \17420 , \16941 , RIaa9d878_210);
nor \U$16751 ( \17421 , \17419 , \17420 );
and \U$16752 ( \17422 , \16931 , RIaa9dcb0_219);
and \U$16753 ( \17423 , \16949 , RIaa9d710_207);
nor \U$16754 ( \17424 , \17422 , \17423 );
and \U$16755 ( \17425 , \16966 , RIaa9dda0_221);
and \U$16756 ( \17426 , \16969 , RIaa9de18_222);
nor \U$16757 ( \17427 , \17425 , \17426 );
nand \U$16758 ( \17428 , \17418 , \17421 , \17424 , \17427 );
and \U$16759 ( \17429 , \16982 , RIaa9d9e0_213);
and \U$16760 ( \17430 , \16996 , RIaa9dc38_218);
nor \U$16761 ( \17431 , \17429 , \17430 );
and \U$16762 ( \17432 , \16991 , RIaa9dbc0_217);
and \U$16763 ( \17433 , \17016 , RIaa9d8f0_211);
nor \U$16764 ( \17434 , \17432 , \17433 );
and \U$16765 ( \17435 , \16977 , RIaa9da58_214);
and \U$16766 ( \17436 , \17010 , RIaa9dd28_220);
nor \U$16767 ( \17437 , \17435 , \17436 );
not \U$16768 ( \17438 , \17001 );
not \U$16769 ( \17439 , \1615 );
and \U$16770 ( \17440 , \17438 , \17439 );
and \U$16771 ( \17441 , \17007 , RIaa9d800_209);
nor \U$16772 ( \17442 , \17440 , \17441 );
nand \U$16773 ( \17443 , \17431 , \17434 , \17437 , \17442 );
nor \U$16774 ( \17444 , \17428 , \17443 );
and \U$16775 ( \17445 , \16825 , \17444 );
nor \U$16776 ( \17446 , \17345 , \17415 , \17445 );
not \U$16777 ( \17447 , \17446 );
or \U$16778 ( \17448 , \17306 , \17447 );
or \U$16779 ( \17449 , \17445 , \12168 , \17344 );
or \U$16780 ( \17450 , \16825 , \17444 );
nand \U$16781 ( \17451 , \17449 , \17450 );
not \U$16782 ( \17452 , \17451 );
or \U$16783 ( \17453 , \17452 , \17415 );
or \U$16784 ( \17454 , \12237 , \17020 );
or \U$16785 ( \17455 , \17413 , \12066 );
not \U$16786 ( \17456 , \17380 );
not \U$16787 ( \17457 , \16810 );
nand \U$16788 ( \17458 , \17456 , \17414 , \17457 );
nand \U$16789 ( \17459 , \17454 , \17455 , \17458 );
not \U$16790 ( \17460 , \17459 );
nand \U$16791 ( \17461 , \17448 , \17453 , \17460 );
nor \U$16792 ( \17462 , \17024 , \17461 );
nor \U$16793 ( \17463 , \17021 , \17462 );
or \U$16794 ( \17464 , \16913 , \17463 );
not \U$16795 ( \17465 , \17461 );
nand \U$16796 ( \17466 , \17465 , \12238 , \16918 );
nand \U$16797 ( \17467 , \17464 , \17466 );
not \U$16798 ( \17468 , \17467 );
not \U$16799 ( \17469 , \17468 );
not \U$16800 ( \17470 , \17469 );
not \U$16801 ( \17471 , \17470 );
and \U$16802 ( \17472 , \16784 , \16796 , \17471 );
nand \U$16803 ( \17473 , \16783 , \17472 );
buf \U$16804 ( \17474 , \11955 );
not \U$16805 ( \17475 , \17474 );
not \U$16806 ( \17476 , \17475 );
not \U$16807 ( \17477 , \6967 );
and \U$16808 ( \17478 , \17476 , \17477 );
not \U$16809 ( \17479 , RIaa9f2b8_266);
nor \U$16810 ( \17480 , \17479 , \12210 );
nor \U$16811 ( \17481 , \17478 , \17480 );
and \U$16812 ( \17482 , \12233 , RIaa9f330_267);
not \U$16813 ( \17483 , RIaa9f588_272);
not \U$16814 ( \17484 , \12288 );
not \U$16815 ( \17485 , \16969 );
or \U$16816 ( \17486 , \17484 , \17485 );
nand \U$16817 ( \17487 , \17486 , \12409 );
not \U$16818 ( \17488 , \17487 );
or \U$16819 ( \17489 , \17483 , \17488 );
and \U$16820 ( \17490 , \12288 , \16966 );
not \U$16821 ( \17491 , \12288 );
and \U$16822 ( \17492 , \17491 , \16969 );
or \U$16823 ( \17493 , \17490 , \17492 );
not \U$16824 ( \17494 , \17493 );
or \U$16825 ( \17495 , \17494 , \6948 );
nand \U$16826 ( \17496 , \17489 , \17495 );
nor \U$16827 ( \17497 , \17482 , \17496 );
nand \U$16828 ( \17498 , \17481 , \17497 );
not \U$16829 ( \17499 , \12231 );
or \U$16830 ( \17500 , \17499 , \12443 );
not \U$16831 ( \17501 , \12196 );
nand \U$16832 ( \17502 , \17501 , RIaa9f498_270);
nand \U$16833 ( \17503 , \17500 , \17502 , \12480 );
nor \U$16834 ( \17504 , \17498 , \17503 );
not \U$16835 ( \17505 , \11948 );
not \U$16836 ( \17506 , \17505 );
and \U$16837 ( \17507 , \17506 , RIaa9f678_274);
not \U$16838 ( \17508 , \11985 );
nor \U$16839 ( \17509 , \17508 , \1427 );
nor \U$16840 ( \17510 , \17507 , \17509 );
not \U$16841 ( \17511 , \11950 );
not \U$16842 ( \17512 , \1416 );
and \U$16843 ( \17513 , \17511 , \17512 );
and \U$16844 ( \17514 , \12057 , RIaa9f510_271);
nor \U$16845 ( \17515 , \17513 , \17514 );
nand \U$16846 ( \17516 , \12215 , RIaa9f858_278);
and \U$16847 ( \17517 , \17510 , \17515 , \17516 );
not \U$16848 ( \17518 , \12200 );
not \U$16849 ( \17519 , \17518 );
not \U$16850 ( \17520 , RIaa9f3a8_268);
not \U$16851 ( \17521 , \17520 );
and \U$16852 ( \17522 , \17519 , \17521 );
and \U$16853 ( \17523 , \12221 , RIaa9f9c0_281);
nor \U$16854 ( \17524 , \17522 , \17523 );
not \U$16855 ( \17525 , \12206 );
not \U$16856 ( \17526 , RIaa9f948_280);
not \U$16857 ( \17527 , \17526 );
and \U$16858 ( \17528 , \17525 , \17527 );
and \U$16859 ( \17529 , \11953 , RIaa9f8d0_279);
nor \U$16860 ( \17530 , \17528 , \17529 );
and \U$16861 ( \17531 , \17524 , \17530 );
and \U$16862 ( \17532 , \17504 , \17517 , \17531 );
buf \U$16863 ( \17533 , \17532 );
not \U$16864 ( \17534 , \17533 );
not \U$16865 ( \17535 , \17534 );
not \U$16866 ( \17536 , \11370 );
or \U$16867 ( \17537 , \12019 , \17413 );
not \U$16868 ( \17538 , \17537 );
not \U$16869 ( \17539 , \17380 );
nand \U$16870 ( \17540 , \17539 , \12013 );
not \U$16871 ( \17541 , \17540 );
not \U$16872 ( \17542 , \17444 );
nand \U$16873 ( \17543 , \17542 , \12116 );
not \U$16874 ( \17544 , \17543 );
nand \U$16875 ( \17545 , \17254 , \11618 );
nand \U$16876 ( \17546 , \17343 , \12121 );
nand \U$16877 ( \17547 , \17545 , \17546 );
nand \U$16878 ( \17548 , \17177 , \11759 );
nand \U$16879 ( \17549 , \17291 , \11674 );
nand \U$16880 ( \17550 , \17221 , \11724 );
nand \U$16881 ( \17551 , \17548 , \17549 , \17550 );
nor \U$16882 ( \17552 , \17547 , \17551 );
not \U$16883 ( \17553 , \17552 );
nand \U$16884 ( \17554 , \17111 , \11911 );
not \U$16885 ( \17555 , \17554 );
not \U$16886 ( \17556 , \17080 );
nand \U$16887 ( \17557 , \17556 , \11808 );
nand \U$16888 ( \17558 , \17555 , \17557 );
nand \U$16889 ( \17559 , \17080 , RIaaa91a0_605);
nand \U$16890 ( \17560 , \17141 , \11814 );
nand \U$16891 ( \17561 , \17559 , \17560 );
not \U$16892 ( \17562 , \17561 );
and \U$16893 ( \17563 , \17558 , \17562 );
nor \U$16894 ( \17564 , \17142 , \11814 );
nor \U$16895 ( \17565 , \17563 , \17564 );
nand \U$16896 ( \17566 , \17052 , \11545 );
and \U$16897 ( \17567 , \17565 , \17566 );
nor \U$16898 ( \17568 , \17052 , \11545 );
nor \U$16899 ( \17569 , \17567 , \17568 );
not \U$16900 ( \17570 , \17569 );
or \U$16901 ( \17571 , \17553 , \17570 );
not \U$16902 ( \17572 , \17548 );
not \U$16903 ( \17573 , \17550 );
nor \U$16904 ( \17574 , \17291 , \11674 );
not \U$16905 ( \17575 , \17574 );
or \U$16906 ( \17576 , \17573 , \17575 );
nand \U$16907 ( \17577 , \17222 , \11932 );
nand \U$16908 ( \17578 , \17576 , \17577 );
not \U$16909 ( \17579 , \17578 );
or \U$16910 ( \17580 , \17572 , \17579 );
nand \U$16911 ( \17581 , \17178 , \11923 );
nand \U$16912 ( \17582 , \17580 , \17581 );
not \U$16913 ( \17583 , \17547 );
and \U$16914 ( \17584 , \17582 , \17583 );
nor \U$16915 ( \17585 , \17254 , \11618 );
not \U$16916 ( \17586 , \17585 );
not \U$16917 ( \17587 , \17546 );
or \U$16918 ( \17588 , \17586 , \17587 );
nand \U$16919 ( \17589 , \17344 , \12122 );
nand \U$16920 ( \17590 , \17588 , \17589 );
nor \U$16921 ( \17591 , \17584 , \17590 );
nand \U$16922 ( \17592 , \17571 , \17591 );
not \U$16923 ( \17593 , \17592 );
or \U$16924 ( \17594 , \17544 , \17593 );
not \U$16925 ( \17595 , \12116 );
nand \U$16926 ( \17596 , \17595 , \17444 );
nand \U$16927 ( \17597 , \17594 , \17596 );
not \U$16928 ( \17598 , \17597 );
or \U$16929 ( \17599 , \17541 , \17598 );
not \U$16930 ( \17600 , \12013 );
nand \U$16931 ( \17601 , \17600 , \17380 );
nand \U$16932 ( \17602 , \17599 , \17601 );
not \U$16933 ( \17603 , \17602 );
or \U$16934 ( \17604 , \17538 , \17603 );
nand \U$16935 ( \17605 , \12019 , \17413 );
nand \U$16936 ( \17606 , \17604 , \17605 );
or \U$16937 ( \17607 , \17020 , \12239 );
nand \U$16938 ( \17608 , \17606 , \17607 );
nand \U$16939 ( \17609 , \17020 , \12239 );
nand \U$16940 ( \17610 , \17608 , \17609 );
not \U$16941 ( \17611 , \17610 );
or \U$16942 ( \17612 , \17536 , \17611 );
not \U$16943 ( \17613 , \11370 );
nand \U$16944 ( \17614 , \17613 , \17608 , \17609 );
nand \U$16945 ( \17615 , \17612 , \17614 );
not \U$16946 ( \17616 , \17615 );
nand \U$16947 ( \17617 , \17609 , \17607 );
not \U$16948 ( \17618 , \17617 );
not \U$16949 ( \17619 , \17606 );
or \U$16950 ( \17620 , \17618 , \17619 );
or \U$16951 ( \17621 , \17606 , \17617 );
nand \U$16952 ( \17622 , \17620 , \17621 );
not \U$16953 ( \17623 , \17622 );
nand \U$16954 ( \17624 , \17616 , \17623 );
nand \U$16955 ( \17625 , \17615 , \17622 );
not \U$16956 ( \17626 , \17602 );
nand \U$16957 ( \17627 , \17537 , \17605 );
not \U$16958 ( \17628 , \17627 );
and \U$16959 ( \17629 , \17626 , \17628 );
and \U$16960 ( \17630 , \17602 , \17627 );
nor \U$16961 ( \17631 , \17629 , \17630 );
not \U$16962 ( \17632 , \17631 );
not \U$16963 ( \17633 , \17632 );
not \U$16964 ( \17634 , \17633 );
not \U$16965 ( \17635 , \17634 );
not \U$16966 ( \17636 , \17622 );
or \U$16967 ( \17637 , \17635 , \17636 );
or \U$16968 ( \17638 , \17634 , \17622 );
nand \U$16969 ( \17639 , \17637 , \17638 );
nand \U$16970 ( \17640 , \17624 , \17625 , \17639 );
not \U$16971 ( \17641 , \17640 );
buf \U$16972 ( \17642 , \17615 );
not \U$16973 ( \17643 , \17642 );
nand \U$16974 ( \17644 , \17641 , \17643 );
not \U$16975 ( \17645 , \17644 );
not \U$16976 ( \17646 , \17645 );
or \U$16977 ( \17647 , \17535 , \17646 );
not \U$16978 ( \17648 , \17640 );
nand \U$16979 ( \17649 , \17648 , \17642 );
not \U$16980 ( \17650 , \17649 );
and \U$16981 ( \17651 , \17650 , \17533 );
not \U$16982 ( \17652 , \17639 );
buf \U$16983 ( \17653 , \17652 );
not \U$16984 ( \17654 , \17642 );
nand \U$16985 ( \17655 , \17653 , \17654 );
buf \U$16986 ( \17656 , \17655 );
not \U$16987 ( \17657 , \17656 );
not \U$16988 ( \17658 , RIaa9ed18_254);
nor \U$16989 ( \17659 , \17658 , \17518 );
not \U$16990 ( \17660 , RIaa9f0d8_262);
nor \U$16991 ( \17661 , \17660 , \17508 );
nor \U$16992 ( \17662 , \17659 , \17661 );
not \U$16993 ( \17663 , \12210 );
not \U$16994 ( \17664 , \6850 );
and \U$16995 ( \17665 , \17663 , \17664 );
and \U$16996 ( \17666 , \12057 , RIaa9eac0_249);
nor \U$16997 ( \17667 , \17665 , \17666 );
nand \U$16998 ( \17668 , \17662 , \17667 );
not \U$16999 ( \17669 , \12233 );
not \U$17000 ( \17670 , \17669 );
not \U$17001 ( \17671 , RIaa9eca0_253);
not \U$17002 ( \17672 , \17671 );
and \U$17003 ( \17673 , \17670 , \17672 );
and \U$17004 ( \17674 , \17493 , RIaa9eb38_250);
and \U$17005 ( \17675 , \17487 , RIaa9ebb0_251);
nor \U$17006 ( \17676 , \17674 , \17675 );
not \U$17007 ( \17677 , \17676 );
nor \U$17008 ( \17678 , \17673 , \17677 );
nand \U$17009 ( \17679 , \17506 , RIaa9ee80_257);
nand \U$17010 ( \17680 , \11978 , RIaa9f060_261);
nand \U$17011 ( \17681 , \12215 , RIaa9f150_263);
nand \U$17012 ( \17682 , \17678 , \17679 , \17680 , \17681 );
nor \U$17013 ( \17683 , \17668 , \17682 );
buf \U$17014 ( \17684 , \11966 );
and \U$17015 ( \17685 , \17684 , RIaa9ef70_259);
not \U$17016 ( \17686 , \11993 );
and \U$17017 ( \17687 , \17686 , RIaa9efe8_260);
nor \U$17018 ( \17688 , \17685 , \17687 );
not \U$17019 ( \17689 , RIaa9eef8_258);
not \U$17020 ( \17690 , \11951 );
nor \U$17021 ( \17691 , \17689 , \17690 );
not \U$17022 ( \17692 , RIaa9ee08_256);
nor \U$17023 ( \17693 , \17692 , \17475 );
nor \U$17024 ( \17694 , \17691 , \17693 );
nand \U$17025 ( \17695 , \17688 , \17694 );
nand \U$17026 ( \17696 , \11953 , RIaa9f1c8_264);
nand \U$17027 ( \17697 , \17501 , RIaa9ed90_255);
nand \U$17028 ( \17698 , \17696 , \17697 , \12519 );
nor \U$17029 ( \17699 , \17695 , \17698 );
and \U$17030 ( \17700 , \17683 , \17699 );
not \U$17031 ( \17701 , \17700 );
buf \U$17032 ( \17702 , \17701 );
and \U$17033 ( \17703 , \17657 , \17702 );
nand \U$17034 ( \17704 , \17642 , \17652 );
not \U$17035 ( \17705 , \17704 );
not \U$17036 ( \17706 , \17702 );
and \U$17037 ( \17707 , \17705 , \17706 );
nor \U$17038 ( \17708 , \17651 , \17703 , \17707 );
nand \U$17039 ( \17709 , \17647 , \17708 );
not \U$17040 ( \17710 , \17597 );
nand \U$17041 ( \17711 , \17601 , \17540 );
not \U$17042 ( \17712 , \17711 );
and \U$17043 ( \17713 , \17710 , \17712 );
and \U$17044 ( \17714 , \17597 , \17711 );
nor \U$17045 ( \17715 , \17713 , \17714 );
buf \U$17046 ( \17716 , \17715 );
not \U$17047 ( \17717 , \17716 );
not \U$17048 ( \17718 , \17717 );
not \U$17049 ( \17719 , \17632 );
or \U$17050 ( \17720 , \17718 , \17719 );
not \U$17051 ( \17721 , \17716 );
not \U$17052 ( \17722 , \17631 );
or \U$17053 ( \17723 , \17721 , \17722 );
buf \U$17054 ( \17724 , \17592 );
not \U$17055 ( \17725 , \17724 );
nand \U$17056 ( \17726 , \17596 , \17543 );
not \U$17057 ( \17727 , \17726 );
and \U$17058 ( \17728 , \17725 , \17727 );
and \U$17059 ( \17729 , \17724 , \17726 );
nor \U$17060 ( \17730 , \17728 , \17729 );
not \U$17061 ( \17731 , \17730 );
not \U$17062 ( \17732 , \17715 );
or \U$17063 ( \17733 , \17731 , \17732 );
or \U$17064 ( \17734 , \17715 , \17730 );
nand \U$17065 ( \17735 , \17733 , \17734 );
nand \U$17066 ( \17736 , \17723 , \17735 );
not \U$17067 ( \17737 , \17736 );
nand \U$17068 ( \17738 , \17720 , \17737 );
buf \U$17069 ( \17739 , \17738 );
buf \U$17070 ( \17740 , \17735 );
nand \U$17071 ( \17741 , \17739 , \17740 );
buf \U$17072 ( \17742 , \17633 );
not \U$17073 ( \17743 , \17742 );
and \U$17074 ( \17744 , \17741 , \17743 );
nand \U$17075 ( \17745 , \17610 , \11370 );
not \U$17076 ( \17746 , \17745 );
not \U$17077 ( \17747 , \17746 );
and \U$17078 ( \17748 , \11953 , RIaa9fab0_283);
not \U$17079 ( \17749 , RIaa9fd80_289);
nor \U$17080 ( \17750 , \17749 , \12220 );
nor \U$17081 ( \17751 , \17748 , \17750 );
and \U$17082 ( \17752 , \12057 , RIaa9fba0_285);
not \U$17083 ( \17753 , RIaaa0140_297);
nor \U$17084 ( \17754 , \17753 , \17669 );
nor \U$17085 ( \17755 , \17752 , \17754 );
nand \U$17086 ( \17756 , \11985 , RIaa9fe70_291);
nand \U$17087 ( \17757 , \17751 , \17755 , \17756 );
not \U$17088 ( \17758 , \12214 );
not \U$17089 ( \17759 , RIaa9fa38_282);
not \U$17090 ( \17760 , \17759 );
and \U$17091 ( \17761 , \17758 , \17760 );
and \U$17092 ( \17762 , \17506 , RIaa9ff60_293);
nor \U$17093 ( \17763 , \17761 , \17762 );
not \U$17094 ( \17764 , \12210 );
not \U$17095 ( \17765 , RIaaa01b8_298);
not \U$17096 ( \17766 , \17765 );
and \U$17097 ( \17767 , \17764 , \17766 );
and \U$17098 ( \17768 , \12200 , RIaaa0050_295);
nor \U$17099 ( \17769 , \17767 , \17768 );
nand \U$17100 ( \17770 , \17763 , \17769 );
nor \U$17101 ( \17771 , \17757 , \17770 );
not \U$17102 ( \17772 , \12206 );
not \U$17103 ( \17773 , \7005 );
and \U$17104 ( \17774 , \17772 , \17773 );
not \U$17105 ( \17775 , \17690 );
and \U$17106 ( \17776 , \17775 , RIaa9ffd8_294);
nor \U$17107 ( \17777 , \17774 , \17776 );
not \U$17108 ( \17778 , \17499 );
not \U$17109 ( \17779 , RIaa9fee8_292);
not \U$17110 ( \17780 , \17779 );
and \U$17111 ( \17781 , \17778 , \17780 );
and \U$17112 ( \17782 , \17501 , RIaaa00c8_296);
nor \U$17113 ( \17783 , \17781 , \17782 );
and \U$17114 ( \17784 , \12227 , RIaa9fdf8_290);
and \U$17115 ( \17785 , \17493 , RIaa9fc90_287);
and \U$17116 ( \17786 , \17487 , RIaa9fc18_286);
nor \U$17117 ( \17787 , \17784 , \17785 , \17786 );
and \U$17118 ( \17788 , \17777 , \17783 , \17787 , \12413 );
and \U$17119 ( \17789 , \17771 , \17788 );
buf \U$17120 ( \17790 , \17789 );
buf \U$17121 ( \17791 , \17790 );
buf \U$17122 ( \17792 , \17791 );
nor \U$17123 ( \17793 , \17747 , \17792 );
nor \U$17124 ( \17794 , \17744 , \17793 );
and \U$17125 ( \17795 , \17709 , \17794 );
nor \U$17126 ( \17796 , \17795 , \17793 );
and \U$17127 ( \17797 , \17645 , \17702 );
or \U$17128 ( \17798 , \17649 , \17702 );
not \U$17129 ( \17799 , \17705 );
nand \U$17130 ( \17800 , \17798 , \17799 );
nor \U$17131 ( \17801 , \17797 , \17800 );
nor \U$17132 ( \17802 , \17747 , \17533 );
not \U$17133 ( \17803 , \17802 );
and \U$17134 ( \17804 , \17801 , \17803 );
and \U$17135 ( \17805 , \17746 , \17702 );
buf \U$17136 ( \17806 , \17640 );
buf \U$17137 ( \17807 , \17806 );
buf \U$17138 ( \17808 , \17653 );
not \U$17139 ( \17809 , \17808 );
nand \U$17140 ( \17810 , \17807 , \17809 );
not \U$17141 ( \17811 , \17810 );
buf \U$17142 ( \17812 , \17642 );
not \U$17143 ( \17813 , \17812 );
nor \U$17144 ( \17814 , \17805 , \17811 , \17813 );
and \U$17145 ( \17815 , \17802 , \17814 );
nor \U$17146 ( \17816 , \17804 , \17815 );
or \U$17147 ( \17817 , \17796 , \17816 );
or \U$17148 ( \17818 , \17801 , \17802 );
nand \U$17149 ( \17819 , \17817 , \17818 );
not \U$17150 ( \17820 , \17819 );
xor \U$17151 ( \17821 , \17802 , \17814 );
not \U$17152 ( \17822 , \17821 );
and \U$17153 ( \17823 , \17820 , \17822 );
and \U$17154 ( \17824 , \17819 , \17821 );
nor \U$17155 ( \17825 , \17823 , \17824 );
not \U$17156 ( \17826 , \17825 );
xnor \U$17157 ( \17827 , \17709 , \17794 );
not \U$17158 ( \17828 , \17827 );
not \U$17159 ( \17829 , \17792 );
not \U$17160 ( \17830 , \17829 );
not \U$17161 ( \17831 , \17645 );
or \U$17162 ( \17832 , \17830 , \17831 );
not \U$17163 ( \17833 , \17649 );
not \U$17164 ( \17834 , \17829 );
and \U$17165 ( \17835 , \17833 , \17834 );
or \U$17166 ( \17836 , \17656 , \17533 );
or \U$17167 ( \17837 , \17799 , \17534 );
nand \U$17168 ( \17838 , \17836 , \17837 );
nor \U$17169 ( \17839 , \17835 , \17838 );
nand \U$17170 ( \17840 , \17832 , \17839 );
not \U$17171 ( \17841 , \17738 );
nand \U$17172 ( \17842 , \17841 , \17742 );
buf \U$17173 ( \17843 , \17842 );
not \U$17174 ( \17844 , \17843 );
not \U$17175 ( \17845 , \17844 );
or \U$17176 ( \17846 , \17845 , \17706 );
nor \U$17177 ( \17847 , \17738 , \17742 );
buf \U$17178 ( \17848 , \17847 );
buf \U$17179 ( \17849 , \17848 );
and \U$17180 ( \17850 , \17849 , \17706 );
nand \U$17181 ( \17851 , \11982 , RIaaa0938_314);
not \U$17182 ( \17852 , \12057 );
not \U$17183 ( \17853 , \17852 );
nand \U$17184 ( \17854 , \17853 , RIaaa0758_310);
nand \U$17185 ( \17855 , \12233 , RIaaa0668_308);
and \U$17186 ( \17856 , \12221 , RIaaa0398_302);
and \U$17187 ( \17857 , \11953 , RIaaa08c0_313);
nor \U$17188 ( \17858 , \17856 , \17857 );
nand \U$17189 ( \17859 , \17851 , \17854 , \17855 , \17858 );
buf \U$17190 ( \17860 , \11974 );
not \U$17191 ( \17861 , \17860 );
and \U$17192 ( \17862 , \17861 , RIaaa0488_304);
and \U$17193 ( \17863 , \11985 , RIaaa0230_299);
nor \U$17194 ( \17864 , \17862 , \17863 );
and \U$17195 ( \17865 , \12209 , RIaaa06e0_309);
and \U$17196 ( \17866 , \17506 , RIaaa0578_306);
nor \U$17197 ( \17867 , \17865 , \17866 );
nand \U$17198 ( \17868 , \17864 , \17867 );
nor \U$17199 ( \17869 , \17859 , \17868 );
not \U$17200 ( \17870 , \12206 );
and \U$17201 ( \17871 , \17870 , RIaaa0320_301);
and \U$17202 ( \17872 , \17501 , RIaaa0500_305);
nor \U$17203 ( \17873 , \17871 , \17872 );
and \U$17204 ( \17874 , \12227 , RIaaa0410_303);
not \U$17205 ( \17875 , RIaaa07d0_311);
not \U$17206 ( \17876 , \17487 );
or \U$17207 ( \17877 , \17875 , \17876 );
or \U$17208 ( \17878 , \17494 , \7240 );
nand \U$17209 ( \17879 , \17877 , \17878 );
nor \U$17210 ( \17880 , \17874 , \17879 );
nand \U$17211 ( \17881 , \17873 , \17880 );
or \U$17212 ( \17882 , \17690 , \7221 );
nand \U$17213 ( \17883 , \11978 , RIaaa02a8_300);
nand \U$17214 ( \17884 , \17882 , \17883 , \12648 );
nor \U$17215 ( \17885 , \17881 , \17884 );
nand \U$17216 ( \17886 , \17869 , \17885 );
buf \U$17217 ( \17887 , \17886 );
and \U$17218 ( \17888 , \17746 , \17887 );
not \U$17219 ( \17889 , \17632 );
nor \U$17220 ( \17890 , \17889 , \17740 );
not \U$17221 ( \17891 , \17890 );
not \U$17222 ( \17892 , \17891 );
nor \U$17223 ( \17893 , \17850 , \17888 , \17892 );
nand \U$17224 ( \17894 , \17846 , \17893 );
or \U$17225 ( \17895 , \17840 , \17894 );
nand \U$17226 ( \17896 , \17828 , \17895 );
not \U$17227 ( \17897 , \17896 );
xor \U$17228 ( \17898 , \17796 , \17816 );
not \U$17229 ( \17899 , \17898 );
or \U$17230 ( \17900 , \17897 , \17899 );
or \U$17231 ( \17901 , \17898 , \17896 );
nand \U$17232 ( \17902 , \17900 , \17901 );
not \U$17233 ( \17903 , \17902 );
nor \U$17234 ( \17904 , \17622 , \17743 );
and \U$17235 ( \17905 , \12209 , RIaaa7b98_558);
and \U$17236 ( \17906 , \11953 , RIaaa7c88_560);
nor \U$17237 ( \17907 , \17905 , \17906 );
and \U$17238 ( \17908 , \17870 , RIaaa7f58_566);
and \U$17239 ( \17909 , \17686 , RIaaa7fd0_567);
nor \U$17240 ( \17910 , \17908 , \17909 );
and \U$17241 ( \17911 , \12215 , RIaaa7d00_561);
and \U$17242 ( \17912 , \11985 , RIaaa80c0_569);
nor \U$17243 ( \17913 , \17911 , \17912 );
and \U$17244 ( \17914 , \17775 , RIaaa7a30_555);
and \U$17245 ( \17915 , \11948 , RIaaa79b8_554);
nor \U$17246 ( \17916 , \17914 , \17915 );
nand \U$17247 ( \17917 , \17907 , \17910 , \17913 , \17916 );
and \U$17248 ( \17918 , \11969 , RIaaa7b20_557);
not \U$17249 ( \17919 , \17860 );
and \U$17250 ( \17920 , \17919 , RIaaa7aa8_556);
nor \U$17251 ( \17921 , \17918 , \17920 );
not \U$17252 ( \17922 , \17499 );
not \U$17253 ( \17923 , \15528 );
and \U$17254 ( \17924 , \17922 , \17923 );
or \U$17255 ( \17925 , \17669 , \9632 );
and \U$17256 ( \17926 , \17493 , RIaaa7df0_563);
and \U$17257 ( \17927 , \17487 , RIaaa7e68_564);
nor \U$17258 ( \17928 , \17926 , \17927 );
nand \U$17259 ( \17929 , \17925 , \17928 );
nor \U$17260 ( \17930 , \17924 , \17929 );
and \U$17261 ( \17931 , \17474 , RIaaa8048_568);
and \U$17262 ( \17932 , \17853 , RIaaa7d78_562);
nor \U$17263 ( \17933 , \17931 , \17932 );
nand \U$17264 ( \17934 , \17921 , \17930 , \17933 , \15545 );
or \U$17265 ( \17935 , \17917 , \17934 );
not \U$17266 ( \17936 , \17935 );
or \U$17267 ( \17937 , \17904 , \17936 );
nand \U$17268 ( \17938 , \17622 , \17743 );
nand \U$17269 ( \17939 , \17937 , \17938 , \17642 );
not \U$17270 ( \17940 , \17939 );
not \U$17271 ( \17941 , \12196 );
not \U$17272 ( \17942 , \7454 );
and \U$17273 ( \17943 , \17941 , \17942 );
and \U$17274 ( \17944 , \17870 , RIaaa1748_344);
nor \U$17275 ( \17945 , \17943 , \17944 );
and \U$17276 ( \17946 , \12221 , RIaaa17c0_345);
and \U$17277 ( \17947 , \11978 , RIaaa18b0_347);
nor \U$17278 ( \17948 , \17946 , \17947 );
nand \U$17279 ( \17949 , \17945 , \17948 );
and \U$17280 ( \17950 , \12233 , RIaaa1478_338);
and \U$17281 ( \17951 , \17493 , RIaaa1388_336);
and \U$17282 ( \17952 , \17487 , RIaaa1310_335);
nor \U$17283 ( \17953 , \17951 , \17952 );
not \U$17284 ( \17954 , \17953 );
nor \U$17285 ( \17955 , \17950 , \17954 );
nand \U$17286 ( \17956 , \17775 , RIaaa16d0_343);
nand \U$17287 ( \17957 , \12209 , RIaaa1400_337);
nand \U$17288 ( \17958 , \11948 , RIaaa1658_342);
nand \U$17289 ( \17959 , \17955 , \17956 , \17957 , \17958 );
nor \U$17290 ( \17960 , \17949 , \17959 );
nand \U$17291 ( \17961 , \17919 , RIaaa14f0_339);
nand \U$17292 ( \17962 , \11985 , RIaaa1838_346);
nand \U$17293 ( \17963 , \12057 , RIaaa1298_334);
nand \U$17294 ( \17964 , \17474 , RIaaa1568_340);
nand \U$17295 ( \17965 , \17961 , \17962 , \17963 , \17964 );
nand \U$17296 ( \17966 , \11953 , RIaaa19a0_349);
nand \U$17297 ( \17967 , \11982 , RIaaa1928_348);
nand \U$17298 ( \17968 , \17966 , \17967 , \13046 );
nor \U$17299 ( \17969 , \17965 , \17968 );
nand \U$17300 ( \17970 , \17960 , \17969 );
not \U$17301 ( \17971 , \17558 );
buf \U$17302 ( \17972 , \17559 );
not \U$17303 ( \17973 , \17972 );
not \U$17304 ( \17974 , \17973 );
and \U$17305 ( \17975 , \17971 , \17974 );
buf \U$17306 ( \17976 , \17557 );
and \U$17307 ( \17977 , \17972 , \17976 );
buf \U$17308 ( \17978 , \17554 );
not \U$17309 ( \17979 , \17978 );
nor \U$17310 ( \17980 , \17977 , \17979 );
nor \U$17311 ( \17981 , \17975 , \17980 );
buf \U$17312 ( \17982 , \17981 );
not \U$17313 ( \17983 , \17982 );
and \U$17314 ( \17984 , \17970 , \17983 );
not \U$17315 ( \17985 , RIaaa9560_613);
not \U$17316 ( \17986 , \17112 );
or \U$17317 ( \17987 , \17985 , \17986 );
nand \U$17318 ( \17988 , \17987 , \17554 );
not \U$17319 ( \17989 , \17988 );
nor \U$17320 ( \17990 , \17984 , \17989 );
not \U$17321 ( \17991 , \17990 );
or \U$17322 ( \17992 , \17981 , \17988 );
not \U$17323 ( \17993 , \17992 );
not \U$17324 ( \17994 , \17993 );
and \U$17325 ( \17995 , \17991 , \17994 );
not \U$17326 ( \17996 , \17993 );
not \U$17327 ( \17997 , \12214 );
not \U$17328 ( \17998 , \2131 );
and \U$17329 ( \17999 , \17997 , \17998 );
not \U$17330 ( \18000 , RIaaa2cd8_390);
not \U$17331 ( \18001 , \11978 );
nor \U$17332 ( \18002 , \18000 , \18001 );
nor \U$17333 ( \18003 , \17999 , \18002 );
not \U$17334 ( \18004 , \12220 );
not \U$17335 ( \18005 , \7685 );
and \U$17336 ( \18006 , \18004 , \18005 );
not \U$17337 ( \18007 , RIaaa2f30_395);
not \U$17338 ( \18008 , \11953 );
nor \U$17339 ( \18009 , \18007 , \18008 );
nor \U$17340 ( \18010 , \18006 , \18009 );
nand \U$17341 ( \18011 , \18003 , \18010 );
not \U$17342 ( \18012 , \17860 );
not \U$17343 ( \18013 , \12940 );
and \U$17344 ( \18014 , \18012 , \18013 );
not \U$17345 ( \18015 , \11969 );
nor \U$17346 ( \18016 , \18015 , \7700 );
nor \U$17347 ( \18017 , \18014 , \18016 );
not \U$17348 ( \18018 , \12106 );
not \U$17349 ( \18019 , \7672 );
and \U$17350 ( \18020 , \18018 , \18019 );
and \U$17351 ( \18021 , \17506 , RIaaa2a80_385);
nor \U$17352 ( \18022 , \18020 , \18021 );
nand \U$17353 ( \18023 , \18017 , \18022 );
nor \U$17354 ( \18024 , \18011 , \18023 );
not \U$17355 ( \18025 , RIaaa2d50_391);
not \U$17356 ( \18026 , \11985 );
or \U$17357 ( \18027 , \18025 , \18026 );
and \U$17358 ( \18028 , \12233 , RIaaa2c60_389);
and \U$17359 ( \18029 , RIaaa3110_399, \17487 );
and \U$17360 ( \18030 , \17493 , RIaaa3098_398);
nor \U$17361 ( \18031 , \18028 , \18029 , \18030 );
nand \U$17362 ( \18032 , \18027 , \18031 );
not \U$17363 ( \18033 , RIaaa2be8_388);
not \U$17364 ( \18034 , \12209 );
or \U$17365 ( \18035 , \18033 , \18034 );
nand \U$17366 ( \18036 , \12057 , RIaaa3020_397);
nand \U$17367 ( \18037 , \18035 , \18036 );
nor \U$17368 ( \18038 , \18032 , \18037 );
nand \U$17369 ( \18039 , \17684 , RIaaa2e40_393);
nand \U$17370 ( \18040 , \11951 , RIaaa2a08_384);
and \U$17371 ( \18041 , \18039 , \18040 , \12960 );
nand \U$17372 ( \18042 , \18024 , \18038 , \18041 );
not \U$17373 ( \18043 , \18042 );
or \U$17374 ( \18044 , \17996 , \18043 );
not \U$17375 ( \18045 , \17988 );
not \U$17376 ( \18046 , \17970 );
or \U$17377 ( \18047 , \18045 , \18046 );
nand \U$17378 ( \18048 , \18047 , \17982 );
nand \U$17379 ( \18049 , \18044 , \18048 );
nor \U$17380 ( \18050 , \17995 , \18049 );
and \U$17381 ( \18051 , RIaaa3f98_430, \17474 );
and \U$17382 ( \18052 , \12233 , RIaaa3f20_429);
nor \U$17383 ( \18053 , \12196 , \7950 );
nor \U$17384 ( \18054 , \18051 , \18052 , \18053 );
and \U$17385 ( \18055 , \11953 , RIaaa3c50_423);
and \U$17386 ( \18056 , \11948 , RIaaa39f8_418);
nor \U$17387 ( \18057 , \18055 , \18056 );
nand \U$17388 ( \18058 , \18054 , \18057 );
not \U$17389 ( \18059 , \12057 );
not \U$17390 ( \18060 , \18059 );
not \U$17391 ( \18061 , \7953 );
and \U$17392 ( \18062 , \18060 , \18061 );
and \U$17393 ( \18063 , RIaaa3ae8_420, \11985 );
nor \U$17394 ( \18064 , \18062 , \18063 );
not \U$17395 ( \18065 , \12214 );
not \U$17396 ( \18066 , \2680 );
and \U$17397 ( \18067 , \18065 , \18066 );
and \U$17398 ( \18068 , \17919 , RIaaa3ea8_428);
nor \U$17399 ( \18069 , \18067 , \18068 );
nand \U$17400 ( \18070 , \18064 , \18069 );
nor \U$17401 ( \18071 , \18058 , \18070 );
nand \U$17402 ( \18072 , \17684 , RIaaa3cc8_424);
nand \U$17403 ( \18073 , \12221 , RIaaa3d40_425);
nand \U$17404 ( \18074 , \11951 , RIaaa3a70_419);
and \U$17405 ( \18075 , \17493 , RIaaa4178_434);
and \U$17406 ( \18076 , \17487 , RIaaa4100_433);
nor \U$17407 ( \18077 , \18075 , \18076 );
nand \U$17408 ( \18078 , \18072 , \18073 , \18074 , \18077 );
nand \U$17409 ( \18079 , \12209 , RIaaa3e30_427);
nand \U$17410 ( \18080 , \12231 , RIaaa3b60_421);
nand \U$17411 ( \18081 , \18079 , \18080 , \13012 );
nor \U$17412 ( \18082 , \18078 , \18081 );
nand \U$17413 ( \18083 , \18071 , \18082 );
not \U$17414 ( \18084 , \18083 );
not \U$17415 ( \18085 , \18084 );
not \U$17416 ( \18086 , \18085 );
not \U$17417 ( \18087 , \17972 );
not \U$17418 ( \18088 , \17978 );
or \U$17419 ( \18089 , \18087 , \18088 );
nand \U$17420 ( \18090 , \18089 , \17976 );
not \U$17421 ( \18091 , \18090 );
not \U$17422 ( \18092 , \17564 );
buf \U$17423 ( \18093 , \17560 );
nand \U$17424 ( \18094 , \18092 , \18093 );
not \U$17425 ( \18095 , \18094 );
and \U$17426 ( \18096 , \18091 , \18095 );
and \U$17427 ( \18097 , \18090 , \18094 );
nor \U$17428 ( \18098 , \18096 , \18097 );
not \U$17429 ( \18099 , \18098 );
not \U$17430 ( \18100 , \17981 );
and \U$17431 ( \18101 , \18099 , \18100 );
and \U$17432 ( \18102 , \18098 , \17981 );
nor \U$17433 ( \18103 , \18101 , \18102 );
not \U$17434 ( \18104 , \18098 );
buf \U$17435 ( \18105 , \17565 );
not \U$17436 ( \18106 , \18105 );
and \U$17437 ( \18107 , \17051 , \11544 );
not \U$17438 ( \18108 , \17051 );
and \U$17439 ( \18109 , \18108 , \11545 );
nor \U$17440 ( \18110 , \18107 , \18109 );
not \U$17441 ( \18111 , \18110 );
and \U$17442 ( \18112 , \18106 , \18111 );
and \U$17443 ( \18113 , \18105 , \18110 );
nor \U$17444 ( \18114 , \18112 , \18113 );
not \U$17445 ( \18115 , \18114 );
or \U$17446 ( \18116 , \18104 , \18115 );
or \U$17447 ( \18117 , \18114 , \18098 );
nand \U$17448 ( \18118 , \18116 , \18117 );
nor \U$17449 ( \18119 , \18103 , \18118 );
buf \U$17450 ( \18120 , \18114 );
buf \U$17451 ( \18121 , \18120 );
nand \U$17452 ( \18122 , \18119 , \18121 );
not \U$17453 ( \18123 , \18122 );
not \U$17454 ( \18124 , \18123 );
or \U$17455 ( \18125 , \18086 , \18124 );
not \U$17456 ( \18126 , \18120 );
nand \U$17457 ( \18127 , \18119 , \18126 );
not \U$17458 ( \18128 , \18127 );
and \U$17459 ( \18129 , \18128 , \18084 );
not \U$17460 ( \18130 , \18001 );
not \U$17461 ( \18131 , \12792 );
and \U$17462 ( \18132 , \18130 , \18131 );
and \U$17463 ( \18133 , \17919 , RIaaa2558_374);
nor \U$17464 ( \18134 , \18132 , \18133 );
and \U$17465 ( \18135 , \17474 , RIaaa23f0_371);
and \U$17466 ( \18136 , \17853 , RIaaa2828_380);
nor \U$17467 ( \18137 , \18135 , \18136 );
nand \U$17468 ( \18138 , \12209 , RIaaa26c0_377);
nand \U$17469 ( \18139 , \18134 , \18137 , \18138 );
and \U$17470 ( \18140 , \11969 , RIaaa25d0_375);
and \U$17471 ( \18141 , \11953 , RIaaa27b0_379);
nor \U$17472 ( \18142 , \18140 , \18141 );
and \U$17473 ( \18143 , \12221 , RIaaa2210_367);
and \U$17474 ( \18144 , \11948 , RIaaa2468_372);
nor \U$17475 ( \18145 , \18143 , \18144 );
nand \U$17476 ( \18146 , \18142 , \18145 );
nor \U$17477 ( \18147 , \18139 , \18146 );
and \U$17478 ( \18148 , \12215 , RIaaa2738_378);
nor \U$17479 ( \18149 , \17690 , \7989 );
nor \U$17480 ( \18150 , \18148 , \18149 , \12811 );
and \U$17481 ( \18151 , \11966 , RIaaa2288_368);
and \U$17482 ( \18152 , \11985 , RIaaa2300_369);
nor \U$17483 ( \18153 , \18151 , \18152 );
and \U$17484 ( \18154 , \12233 , RIaaa2648_376);
and \U$17485 ( \18155 , \17493 , RIaaa2918_382);
and \U$17486 ( \18156 , \17487 , RIaaa28a0_381);
nor \U$17487 ( \18157 , \18154 , \18155 , \18156 );
and \U$17488 ( \18158 , \18150 , \18153 , \18157 );
nand \U$17489 ( \18159 , \18147 , \18158 );
and \U$17490 ( \18160 , \18103 , \18120 );
not \U$17491 ( \18161 , \18160 );
and \U$17492 ( \18162 , \18159 , \18161 );
not \U$17493 ( \18163 , \18159 );
not \U$17494 ( \18164 , \18103 );
not \U$17495 ( \18165 , \18164 );
nand \U$17496 ( \18166 , \18165 , \18126 );
and \U$17497 ( \18167 , \18163 , \18166 );
nor \U$17498 ( \18168 , \18162 , \18167 );
nor \U$17499 ( \18169 , \18129 , \18168 );
nand \U$17500 ( \18170 , \18125 , \18169 );
xor \U$17501 ( \18171 , \18050 , \18170 );
not \U$17502 ( \18172 , \17574 );
nand \U$17503 ( \18173 , \18172 , \17549 );
xor \U$17504 ( \18174 , \17569 , \18173 );
not \U$17505 ( \18175 , \17549 );
not \U$17506 ( \18176 , \17569 );
or \U$17507 ( \18177 , \18175 , \18176 );
nand \U$17508 ( \18178 , \18177 , \18172 );
nand \U$17509 ( \18179 , \17577 , \17550 );
not \U$17510 ( \18180 , \18179 );
and \U$17511 ( \18181 , \18178 , \18180 );
not \U$17512 ( \18182 , \18178 );
and \U$17513 ( \18183 , \18182 , \18179 );
nor \U$17514 ( \18184 , \18181 , \18183 );
not \U$17515 ( \18185 , \18184 );
xor \U$17516 ( \18186 , \18174 , \18185 );
not \U$17517 ( \18187 , \18120 );
not \U$17518 ( \18188 , \18174 );
nand \U$17519 ( \18189 , \18187 , \18188 );
nand \U$17520 ( \18190 , \18120 , \18174 );
nand \U$17521 ( \18191 , \18189 , \18190 );
nand \U$17522 ( \18192 , \18186 , \18191 );
not \U$17523 ( \18193 , \18184 );
not \U$17524 ( \18194 , \18193 );
nor \U$17525 ( \18195 , \18192 , \18194 );
buf \U$17526 ( \18196 , \18195 );
not \U$17527 ( \18197 , \18196 );
not \U$17528 ( \18198 , \12214 );
not \U$17529 ( \18199 , \8423 );
and \U$17530 ( \18200 , \18198 , \18199 );
not \U$17531 ( \18201 , RIaaa4808_448);
nor \U$17532 ( \18202 , \18201 , \17508 );
nor \U$17533 ( \18203 , \18200 , \18202 );
not \U$17534 ( \18204 , \18059 );
not \U$17535 ( \18205 , \13760 );
and \U$17536 ( \18206 , \18204 , \18205 );
nor \U$17537 ( \18207 , \17475 , \8405 );
nor \U$17538 ( \18208 , \18206 , \18207 );
nand \U$17539 ( \18209 , \11953 , RIaaa4970_451);
nand \U$17540 ( \18210 , \18203 , \18208 , \18209 );
not \U$17541 ( \18211 , \17518 );
not \U$17542 ( \18212 , RIaaa44c0_441);
not \U$17543 ( \18213 , \18212 );
and \U$17544 ( \18214 , \18211 , \18213 );
and \U$17545 ( \18215 , \12221 , RIaaa4790_447);
nor \U$17546 ( \18216 , \18214 , \18215 );
not \U$17547 ( \18217 , RIaaa4628_444);
not \U$17548 ( \18218 , \11948 );
nor \U$17549 ( \18219 , \18217 , \18218 );
nor \U$17550 ( \18220 , \12196 , \3138 );
nor \U$17551 ( \18221 , \18219 , \18220 );
nand \U$17552 ( \18222 , \18216 , \18221 );
nor \U$17553 ( \18223 , \18210 , \18222 );
and \U$17554 ( \18224 , \12209 , RIaaa43d0_439);
not \U$17555 ( \18225 , RIaaa46a0_445);
nor \U$17556 ( \18226 , \18225 , \17690 );
nor \U$17557 ( \18227 , \18224 , \18226 );
and \U$17558 ( \18228 , \12233 , RIaaa4448_440);
and \U$17559 ( \18229 , \17493 , RIaaa4358_438);
and \U$17560 ( \18230 , \17487 , RIaaa42e0_437);
nor \U$17561 ( \18231 , \18228 , \18229 , \18230 );
nand \U$17562 ( \18232 , \18227 , \18231 );
nand \U$17563 ( \18233 , \12231 , RIaaa4880_449);
nand \U$17564 ( \18234 , \17684 , RIaaa4718_446);
nand \U$17565 ( \18235 , \18233 , \18234 , \13755 );
nor \U$17566 ( \18236 , \18232 , \18235 );
nand \U$17567 ( \18237 , \18223 , \18236 );
not \U$17568 ( \18238 , \18237 );
or \U$17569 ( \18239 , \18197 , \18238 );
not \U$17570 ( \18240 , \18192 );
nand \U$17571 ( \18241 , \18240 , \18194 );
not \U$17572 ( \18242 , \18241 );
not \U$17573 ( \18243 , \18238 );
not \U$17574 ( \18244 , \18243 );
nand \U$17575 ( \18245 , \18242 , \18244 );
not \U$17576 ( \18246 , \12214 );
not \U$17577 ( \18247 , \8215 );
and \U$17578 ( \18248 , \18246 , \18247 );
and \U$17579 ( \18249 , \17686 , RIaaa3980_417);
nor \U$17580 ( \18250 , \18248 , \18249 );
not \U$17581 ( \18251 , \17499 );
not \U$17582 ( \18252 , RIaaa37a0_413);
not \U$17583 ( \18253 , \18252 );
and \U$17584 ( \18254 , \18251 , \18253 );
not \U$17585 ( \18255 , RIaaa36b0_411);
nor \U$17586 ( \18256 , \18255 , \18008 );
nor \U$17587 ( \18257 , \18254 , \18256 );
nand \U$17588 ( \18258 , \18250 , \18257 );
not \U$17589 ( \18259 , \12106 );
not \U$17590 ( \18260 , RIaaa33e0_405);
not \U$17591 ( \18261 , \18260 );
and \U$17592 ( \18262 , \18259 , \18261 );
and \U$17593 ( \18263 , \11969 , RIaaa3458_406);
nor \U$17594 ( \18264 , \18262 , \18263 );
not \U$17595 ( \18265 , \12206 );
not \U$17596 ( \18266 , RIaaa3908_416);
not \U$17597 ( \18267 , \18266 );
and \U$17598 ( \18268 , \18265 , \18267 );
and \U$17599 ( \18269 , \17775 , RIaaa3890_415);
nor \U$17600 ( \18270 , \18268 , \18269 );
nand \U$17601 ( \18271 , \18264 , \18270 );
nor \U$17602 ( \18272 , \18258 , \18271 );
not \U$17603 ( \18273 , \17518 );
and \U$17604 ( \18274 , \18273 , RIaaa32f0_403);
not \U$17605 ( \18275 , RIaaa3818_414);
nor \U$17606 ( \18276 , \18275 , \18218 );
nor \U$17607 ( \18277 , \18274 , \18276 );
not \U$17608 ( \18278 , \18059 );
not \U$17609 ( \18279 , \8199 );
and \U$17610 ( \18280 , \18278 , \18279 );
and \U$17611 ( \18281 , \12209 , RIaaa3278_402);
nor \U$17612 ( \18282 , \18280 , \18281 );
nand \U$17613 ( \18283 , \18277 , \18282 );
and \U$17614 ( \18284 , \12233 , RIaaa3368_404);
and \U$17615 ( \18285 , RIaaa35c0_409, \17493 );
and \U$17616 ( \18286 , \17487 , RIaaa3548_408);
nor \U$17617 ( \18287 , \18284 , \18285 , \18286 );
nand \U$17618 ( \18288 , \11985 , RIaaa3728_412);
nand \U$17619 ( \18289 , \18287 , \18288 , \13667 );
nor \U$17620 ( \18290 , \18283 , \18289 );
nand \U$17621 ( \18291 , \18272 , \18290 );
not \U$17622 ( \18292 , \18291 );
not \U$17623 ( \18293 , \18191 );
nand \U$17624 ( \18294 , \18293 , \18194 );
not \U$17625 ( \18295 , \18294 );
and \U$17626 ( \18296 , \18292 , \18295 );
not \U$17627 ( \18297 , \18292 );
not \U$17628 ( \18298 , \18193 );
nor \U$17629 ( \18299 , \18298 , \18191 );
buf \U$17630 ( \18300 , \18299 );
and \U$17631 ( \18301 , \18297 , \18300 );
nor \U$17632 ( \18302 , \18296 , \18301 );
nand \U$17633 ( \18303 , \18239 , \18245 , \18302 );
nor \U$17634 ( \18304 , \18171 , \18303 );
not \U$17635 ( \18305 , \18304 );
nand \U$17636 ( \18306 , \18303 , \18171 );
nand \U$17637 ( \18307 , \18305 , \18306 );
not \U$17638 ( \18308 , \18307 );
or \U$17639 ( \18309 , \17940 , \18308 );
or \U$17640 ( \18310 , \18307 , \17939 );
nand \U$17641 ( \18311 , \18309 , \18310 );
and \U$17642 ( \18312 , \17684 , RIaaa68d8_518);
and \U$17643 ( \18313 , \17775 , RIaaa67e8_516);
nor \U$17644 ( \18314 , \18312 , \18313 );
and \U$17645 ( \18315 , \17686 , RIaaa6950_519);
and \U$17646 ( \18316 , \17861 , RIaaa64a0_509);
nor \U$17647 ( \18317 , \18315 , \18316 );
nand \U$17648 ( \18318 , \18314 , \18317 );
not \U$17649 ( \18319 , \18318 );
and \U$17650 ( \18320 , RIaaa6590_511, \12227 );
and \U$17651 ( \18321 , \12057 , RIaaa6248_504);
nor \U$17652 ( \18322 , \18218 , \8522 );
nor \U$17653 ( \18323 , \18320 , \18321 , \18322 );
and \U$17654 ( \18324 , \12215 , RIaaa66f8_514);
and \U$17655 ( \18325 , \11985 , RIaaa6680_513);
nor \U$17656 ( \18326 , \18324 , \18325 );
nand \U$17657 ( \18327 , \12209 , RIaaa63b0_507);
not \U$17658 ( \18328 , \12196 );
nand \U$17659 ( \18329 , \18328 , RIaaa6518_510);
nand \U$17660 ( \18330 , \12233 , RIaaa6428_508);
and \U$17661 ( \18331 , \17493 , RIaaa6338_506);
and \U$17662 ( \18332 , \17487 , RIaaa62c0_505);
nor \U$17663 ( \18333 , \18331 , \18332 );
nand \U$17664 ( \18334 , \18327 , \18329 , \18330 , \18333 );
nand \U$17665 ( \18335 , \12231 , RIaaa6608_512);
nand \U$17666 ( \18336 , \11953 , RIaaa6770_515);
nand \U$17667 ( \18337 , \18335 , \18336 , \14036 );
nor \U$17668 ( \18338 , \18334 , \18337 );
nand \U$17669 ( \18339 , \18319 , \18323 , \18326 , \18338 );
buf \U$17670 ( \18340 , \18339 );
and \U$17671 ( \18341 , \18340 , \18196 );
not \U$17672 ( \18342 , \18340 );
and \U$17673 ( \18343 , \18342 , \18242 );
nor \U$17674 ( \18344 , \18341 , \18343 );
and \U$17675 ( \18345 , \18243 , \18299 );
not \U$17676 ( \18346 , \18243 );
and \U$17677 ( \18347 , \18346 , \18295 );
nor \U$17678 ( \18348 , \18345 , \18347 );
nand \U$17679 ( \18349 , \18344 , \18348 );
not \U$17680 ( \18350 , \18349 );
not \U$17681 ( \18351 , \18291 );
not \U$17682 ( \18352 , \18123 );
or \U$17683 ( \18353 , \18351 , \18352 );
not \U$17684 ( \18354 , \18127 );
not \U$17685 ( \18355 , \18291 );
and \U$17686 ( \18356 , \18354 , \18355 );
or \U$17687 ( \18357 , \18084 , \18161 );
not \U$17688 ( \18358 , \18083 );
nor \U$17689 ( \18359 , \18164 , \18121 );
nand \U$17690 ( \18360 , \18358 , \18359 );
nand \U$17691 ( \18361 , \18357 , \18360 );
nor \U$17692 ( \18362 , \18356 , \18361 );
nand \U$17693 ( \18363 , \18353 , \18362 );
not \U$17694 ( \18364 , \18363 );
buf \U$17695 ( \18365 , \18042 );
and \U$17696 ( \18366 , \17982 , \17988 );
and \U$17697 ( \18367 , \18365 , \18366 );
not \U$17698 ( \18368 , \17993 );
not \U$17699 ( \18369 , \18159 );
not \U$17700 ( \18370 , \18369 );
or \U$17701 ( \18371 , \18368 , \18370 );
not \U$17702 ( \18372 , \18042 );
or \U$17703 ( \18373 , \17981 , \17989 );
not \U$17704 ( \18374 , \18373 );
nand \U$17705 ( \18375 , \18372 , \18374 );
nand \U$17706 ( \18376 , \18371 , \18375 );
nor \U$17707 ( \18377 , \18367 , \18376 );
not \U$17708 ( \18378 , \18377 );
and \U$17709 ( \18379 , \18364 , \18378 );
and \U$17710 ( \18380 , \18363 , \18377 );
nor \U$17711 ( \18381 , \18379 , \18380 );
not \U$17712 ( \18382 , \18381 );
and \U$17713 ( \18383 , \18350 , \18382 );
and \U$17714 ( \18384 , \18349 , \18381 );
nor \U$17715 ( \18385 , \18383 , \18384 );
and \U$17716 ( \18386 , \17684 , RIaaa86d8_582);
and \U$17717 ( \18387 , \17775 , RIaaa8660_581);
nor \U$17718 ( \18388 , \18386 , \18387 );
and \U$17719 ( \18389 , \17686 , RIaaa8750_583);
and \U$17720 ( \18390 , \12215 , RIaaa88b8_586);
nor \U$17721 ( \18391 , \18389 , \18390 );
and \U$17722 ( \18392 , \11953 , RIaaa8930_587);
and \U$17723 ( \18393 , \12231 , RIaaa8840_585);
nor \U$17724 ( \18394 , \18392 , \18393 );
not \U$17725 ( \18395 , \17475 );
not \U$17726 ( \18396 , RIaaa84f8_578);
not \U$17727 ( \18397 , \18396 );
and \U$17728 ( \18398 , \18395 , \18397 );
and \U$17729 ( \18399 , \17501 , RIaaa8570_579);
nor \U$17730 ( \18400 , \18398 , \18399 );
and \U$17731 ( \18401 , \18388 , \18391 , \18394 , \18400 );
and \U$17732 ( \18402 , \17853 , RIaaa8228_572);
and \U$17733 ( \18403 , \17493 , RIaaa8318_574);
and \U$17734 ( \18404 , \17487 , RIaaa82a0_573);
nor \U$17735 ( \18405 , \18402 , \18403 , \18404 );
nand \U$17736 ( \18406 , \11985 , RIaaa87c8_584);
and \U$17737 ( \18407 , \18405 , \18406 , \15339 );
and \U$17738 ( \18408 , \17506 , RIaaa85e8_580);
and \U$17739 ( \18409 , \17861 , RIaaa8408_576);
nor \U$17740 ( \18410 , \18408 , \18409 );
and \U$17741 ( \18411 , \12209 , RIaaa8390_575);
and \U$17742 ( \18412 , \12233 , RIaaa8480_577);
nor \U$17743 ( \18413 , \18411 , \18412 );
nand \U$17744 ( \18414 , \18401 , \18407 , \18410 , \18413 );
buf \U$17745 ( \18415 , \18414 );
not \U$17746 ( \18416 , \18415 );
not \U$17747 ( \18417 , \18416 );
nor \U$17748 ( \18418 , \17738 , \17742 );
not \U$17749 ( \18419 , \18418 );
or \U$17750 ( \18420 , \18417 , \18419 );
and \U$17751 ( \18421 , \12221 , RIaaa7760_549);
and \U$17752 ( \18422 , \12231 , RIaaa7850_551);
nor \U$17753 ( \18423 , \18421 , \18422 );
and \U$17754 ( \18424 , \11953 , RIaaa7940_553);
and \U$17755 ( \18425 , \12215 , RIaaa78c8_552);
nor \U$17756 ( \18426 , \18424 , \18425 );
nand \U$17757 ( \18427 , \18423 , \18426 );
and \U$17758 ( \18428 , \11966 , RIaaa76e8_548);
and \U$17759 ( \18429 , \11951 , RIaaa7670_547);
nor \U$17760 ( \18430 , \18428 , \18429 );
not \U$17761 ( \18431 , \17475 );
not \U$17762 ( \18432 , \4566 );
and \U$17763 ( \18433 , \18431 , \18432 );
and \U$17764 ( \18434 , \11969 , RIaaa7580_545);
nor \U$17765 ( \18435 , \18433 , \18434 );
nand \U$17766 ( \18436 , \18430 , \18435 );
nor \U$17767 ( \18437 , \18427 , \18436 );
and \U$17768 ( \18438 , \17506 , RIaaa75f8_546);
and \U$17769 ( \18439 , \17919 , RIaaa7490_543);
nor \U$17770 ( \18440 , \18438 , \18439 );
and \U$17771 ( \18441 , \12209 , RIaaa73a0_541);
and \U$17772 ( \18442 , \12233 , RIaaa7418_542);
nor \U$17773 ( \18443 , \18441 , \18442 );
nand \U$17774 ( \18444 , \18440 , \18443 );
and \U$17775 ( \18445 , \17853 , RIaaa7238_538);
and \U$17776 ( \18446 , \17493 , RIaaa7328_540);
and \U$17777 ( \18447 , \17487 , RIaaa72b0_539);
nor \U$17778 ( \18448 , \18446 , \18447 );
not \U$17779 ( \18449 , \18448 );
nor \U$17780 ( \18450 , \18445 , \18449 );
nand \U$17781 ( \18451 , \11985 , RIaaa77d8_550);
nand \U$17782 ( \18452 , \18450 , \18451 , \15242 );
nor \U$17783 ( \18453 , \18444 , \18452 );
nand \U$17784 ( \18454 , \18437 , \18453 );
buf \U$17785 ( \18455 , \18454 );
not \U$17786 ( \18456 , \17740 );
nand \U$17787 ( \18457 , \17633 , \18456 );
not \U$17788 ( \18458 , \18457 );
and \U$17789 ( \18459 , \18455 , \18458 );
not \U$17790 ( \18460 , \18455 );
buf \U$17791 ( \18461 , \17890 );
and \U$17792 ( \18462 , \18460 , \18461 );
nor \U$17793 ( \18463 , \18459 , \18462 );
nand \U$17794 ( \18464 , \18420 , \18463 );
not \U$17795 ( \18465 , \17842 );
not \U$17796 ( \18466 , \18465 );
nor \U$17797 ( \18467 , \18466 , \18416 );
nor \U$17798 ( \18468 , \18464 , \18467 );
xor \U$17799 ( \18469 , \18385 , \18468 );
not \U$17800 ( \18470 , \17518 );
not \U$17801 ( \18471 , \4153 );
and \U$17802 ( \18472 , \18470 , \18471 );
and \U$17803 ( \18473 , \12215 , RIaaa5ca8_492);
nor \U$17804 ( \18474 , \18472 , \18473 );
and \U$17805 ( \18475 , \12227 , RIaaa6068_500);
and \U$17806 ( \18476 , \12057 , RIaaa5e10_495);
nor \U$17807 ( \18477 , \18475 , \18476 );
nand \U$17808 ( \18478 , \11985 , RIaaa60e0_501);
nand \U$17809 ( \18479 , \18474 , \18477 , \18478 );
and \U$17810 ( \18480 , \12221 , RIaaa5f78_498);
and \U$17811 ( \18481 , \11953 , RIaaa5d20_493);
nor \U$17812 ( \18482 , \18480 , \18481 );
not \U$17813 ( \18483 , \18218 );
not \U$17814 ( \18484 , \4144 );
and \U$17815 ( \18485 , \18483 , \18484 );
nor \U$17816 ( \18486 , \12206 , \4179 );
nor \U$17817 ( \18487 , \18485 , \18486 );
nand \U$17818 ( \18488 , \18482 , \18487 );
nor \U$17819 ( \18489 , \18479 , \18488 );
and \U$17820 ( \18490 , \11969 , RIaaa5ac8_488);
and \U$17821 ( \18491 , \17775 , RIaaa5a50_487);
nor \U$17822 ( \18492 , \18490 , \18491 );
and \U$17823 ( \18493 , \12209 , RIaaa5bb8_490);
and \U$17824 ( \18494 , \12231 , RIaaa6158_502);
nor \U$17825 ( \18495 , \18493 , \18494 );
and \U$17826 ( \18496 , \12233 , RIaaa5c30_491);
and \U$17827 ( \18497 , \17493 , RIaaa5f00_497);
and \U$17828 ( \18498 , \17487 , RIaaa5e88_496);
nor \U$17829 ( \18499 , \18496 , \18497 , \18498 );
and \U$17830 ( \18500 , \18492 , \18495 , \18499 , \14762 );
nand \U$17831 ( \18501 , \18489 , \18500 );
buf \U$17832 ( \18502 , \18501 );
not \U$17833 ( \18503 , \18502 );
not \U$17834 ( \18504 , \17548 );
not \U$17835 ( \18505 , \17550 );
not \U$17836 ( \18506 , \18178 );
or \U$17837 ( \18507 , \18505 , \18506 );
nand \U$17838 ( \18508 , \18507 , \17577 );
not \U$17839 ( \18509 , \18508 );
or \U$17840 ( \18510 , \18504 , \18509 );
nand \U$17841 ( \18511 , \18510 , \17581 );
not \U$17842 ( \18512 , \17585 );
nand \U$17843 ( \18513 , \18512 , \17545 );
and \U$17844 ( \18514 , \18511 , \18513 );
not \U$17845 ( \18515 , \18511 );
not \U$17846 ( \18516 , \18513 );
and \U$17847 ( \18517 , \18515 , \18516 );
nor \U$17848 ( \18518 , \18514 , \18517 );
not \U$17849 ( \18519 , \18518 );
not \U$17850 ( \18520 , \18519 );
not \U$17851 ( \18521 , \17545 );
not \U$17852 ( \18522 , \18511 );
or \U$17853 ( \18523 , \18521 , \18522 );
nand \U$17854 ( \18524 , \18523 , \18512 );
nand \U$17855 ( \18525 , \17546 , \17589 );
not \U$17856 ( \18526 , \18525 );
and \U$17857 ( \18527 , \18524 , \18526 );
not \U$17858 ( \18528 , \18524 );
and \U$17859 ( \18529 , \18528 , \18525 );
nor \U$17860 ( \18530 , \18527 , \18529 );
not \U$17861 ( \18531 , \18530 );
not \U$17862 ( \18532 , \18531 );
or \U$17863 ( \18533 , \18520 , \18532 );
nand \U$17864 ( \18534 , \18530 , \18518 );
nand \U$17865 ( \18535 , \18533 , \18534 );
buf \U$17866 ( \18536 , \17730 );
nand \U$17867 ( \18537 , \18535 , \18536 );
not \U$17868 ( \18538 , \18537 );
not \U$17869 ( \18539 , \18538 );
or \U$17870 ( \18540 , \18503 , \18539 );
and \U$17871 ( \18541 , \11953 , RIaaa6f68_532);
and \U$17872 ( \18542 , \11978 , RIaaa6e00_529);
nor \U$17873 ( \18543 , \18541 , \18542 );
and \U$17874 ( \18544 , \12221 , RIaaa6d10_527);
and \U$17875 ( \18545 , \12215 , RIaaa6ef0_531);
nor \U$17876 ( \18546 , \18544 , \18545 );
nand \U$17877 ( \18547 , \18543 , \18546 );
not \U$17878 ( \18548 , \12206 );
not \U$17879 ( \18549 , \4324 );
and \U$17880 ( \18550 , \18548 , \18549 );
and \U$17881 ( \18551 , \17775 , RIaaa6ab8_522);
nor \U$17882 ( \18552 , \18550 , \18551 );
not \U$17883 ( \18553 , \12106 );
not \U$17884 ( \18554 , RIaaa6e78_530);
not \U$17885 ( \18555 , \18554 );
and \U$17886 ( \18556 , \18553 , \18555 );
and \U$17887 ( \18557 , \17501 , RIaaa6a40_521);
nor \U$17888 ( \18558 , \18556 , \18557 );
nand \U$17889 ( \18559 , \18552 , \18558 );
nor \U$17890 ( \18560 , \18547 , \18559 );
not \U$17891 ( \18561 , \12210 );
not \U$17892 ( \18562 , \4337 );
and \U$17893 ( \18563 , \18561 , \18562 );
and \U$17894 ( \18564 , \17506 , RIaaa6b30_523);
nor \U$17895 ( \18565 , \18563 , \18564 );
and \U$17896 ( \18566 , \12057 , RIaaa6fe0_533);
and \U$17897 ( \18567 , \17919 , RIaaa69c8_520);
nor \U$17898 ( \18568 , \18566 , \18567 );
nand \U$17899 ( \18569 , \18565 , \18568 );
and \U$17900 ( \18570 , \12233 , RIaaa6ba8_524);
not \U$17901 ( \18571 , RIaaa7058_534);
not \U$17902 ( \18572 , \17487 );
or \U$17903 ( \18573 , \18571 , \18572 );
or \U$17904 ( \18574 , \17494 , \4334 );
nand \U$17905 ( \18575 , \18573 , \18574 );
nor \U$17906 ( \18576 , \18570 , \18575 );
nand \U$17907 ( \18577 , \11985 , RIaaa6d88_528);
nand \U$17908 ( \18578 , \18576 , \18577 , \15010 );
nor \U$17909 ( \18579 , \18569 , \18578 );
nand \U$17910 ( \18580 , \18560 , \18579 );
buf \U$17911 ( \18581 , \18580 );
nand \U$17912 ( \18582 , \18530 , \18519 , \18536 );
not \U$17913 ( \18583 , \18582 );
and \U$17914 ( \18584 , \18581 , \18583 );
not \U$17915 ( \18585 , \18581 );
not \U$17916 ( \18586 , \18530 );
not \U$17917 ( \18587 , \18519 );
not \U$17918 ( \18588 , \18536 );
nand \U$17919 ( \18589 , \18586 , \18587 , \18588 );
not \U$17920 ( \18590 , \18589 );
and \U$17921 ( \18591 , \18585 , \18590 );
nor \U$17922 ( \18592 , \18584 , \18591 );
nand \U$17923 ( \18593 , \18540 , \18592 );
nand \U$17924 ( \18594 , \18535 , \18588 );
nor \U$17925 ( \18595 , \18594 , \18502 );
nor \U$17926 ( \18596 , \18593 , \18595 );
and \U$17927 ( \18597 , \18469 , \18596 );
and \U$17928 ( \18598 , \18385 , \18468 );
or \U$17929 ( \18599 , \18597 , \18598 );
xor \U$17930 ( \18600 , \18311 , \18599 );
not \U$17931 ( \18601 , \18381 );
not \U$17932 ( \18602 , \18601 );
not \U$17933 ( \18603 , \18349 );
or \U$17934 ( \18604 , \18602 , \18603 );
not \U$17935 ( \18605 , \18377 );
nand \U$17936 ( \18606 , \18605 , \18363 );
nand \U$17937 ( \18607 , \18604 , \18606 );
not \U$17938 ( \18608 , \18455 );
not \U$17939 ( \18609 , \18465 );
or \U$17940 ( \18610 , \18608 , \18609 );
not \U$17941 ( \18611 , \18455 );
and \U$17942 ( \18612 , \17848 , \18611 );
not \U$17943 ( \18613 , \18458 );
and \U$17944 ( \18614 , \18581 , \18613 );
not \U$17945 ( \18615 , \18581 );
and \U$17946 ( \18616 , \18615 , \17891 );
nor \U$17947 ( \18617 , \18614 , \18616 );
nor \U$17948 ( \18618 , \18612 , \18617 );
nand \U$17949 ( \18619 , \18610 , \18618 );
xor \U$17950 ( \18620 , \18607 , \18619 );
not \U$17951 ( \18621 , \18508 );
nand \U$17952 ( \18622 , \17548 , \17581 );
not \U$17953 ( \18623 , \18622 );
and \U$17954 ( \18624 , \18621 , \18623 );
and \U$17955 ( \18625 , \18508 , \18622 );
nor \U$17956 ( \18626 , \18624 , \18625 );
not \U$17957 ( \18627 , \18626 );
not \U$17958 ( \18628 , \18627 );
not \U$17959 ( \18629 , \18519 );
or \U$17960 ( \18630 , \18628 , \18629 );
and \U$17961 ( \18631 , \18518 , \18626 );
not \U$17962 ( \18632 , \18184 );
not \U$17963 ( \18633 , \18626 );
or \U$17964 ( \18634 , \18632 , \18633 );
or \U$17965 ( \18635 , \18626 , \18194 );
nand \U$17966 ( \18636 , \18634 , \18635 );
nor \U$17967 ( \18637 , \18631 , \18636 );
nand \U$17968 ( \18638 , \18630 , \18637 );
buf \U$17969 ( \18639 , \18519 );
nor \U$17970 ( \18640 , \18638 , \18639 );
buf \U$17971 ( \18641 , \18640 );
not \U$17972 ( \18642 , \17508 );
not \U$17973 ( \18643 , \8925 );
and \U$17974 ( \18644 , \18642 , \18643 );
and \U$17975 ( \18645 , \11948 , RIaaa5618_478);
nor \U$17976 ( \18646 , \18644 , \18645 );
and \U$17977 ( \18647 , \11969 , RIaaa5438_474);
and \U$17978 ( \18648 , \12057 , RIaaa54b0_475);
nor \U$17979 ( \18649 , \18647 , \18648 );
nand \U$17980 ( \18650 , \12215 , RIaaa57f8_482);
nand \U$17981 ( \18651 , \18646 , \18649 , \18650 );
not \U$17982 ( \18652 , \18008 );
not \U$17983 ( \18653 , \14437 );
and \U$17984 ( \18654 , \18652 , \18653 );
nor \U$17985 ( \18655 , \12220 , \8943 );
nor \U$17986 ( \18656 , \18654 , \18655 );
not \U$17987 ( \18657 , \12206 );
not \U$17988 ( \18658 , \8937 );
and \U$17989 ( \18659 , \18657 , \18658 );
and \U$17990 ( \18660 , \17919 , RIaaa52d0_471);
nor \U$17991 ( \18661 , \18659 , \18660 );
nand \U$17992 ( \18662 , \18656 , \18661 );
nor \U$17993 ( \18663 , \18651 , \18662 );
and \U$17994 ( \18664 , \11978 , RIaaa5780_481);
and \U$17995 ( \18665 , \11951 , RIaaa5690_479);
not \U$17996 ( \18666 , \14447 );
nor \U$17997 ( \18667 , \18664 , \18665 , \18666 );
and \U$17998 ( \18668 , \12209 , RIaaa5258_470);
and \U$17999 ( \18669 , \12227 , RIaaa53c0_473);
nor \U$18000 ( \18670 , \18668 , \18669 );
and \U$18001 ( \18671 , \12233 , RIaaa5348_472);
and \U$18002 ( \18672 , \17493 , RIaaa5528_476);
and \U$18003 ( \18673 , \17487 , RIaaa55a0_477);
nor \U$18004 ( \18674 , \18671 , \18672 , \18673 );
nand \U$18005 ( \18675 , \18663 , \18667 , \18670 , \18674 );
not \U$18006 ( \18676 , \18675 );
not \U$18007 ( \18677 , \18676 );
not \U$18008 ( \18678 , \18677 );
buf \U$18009 ( \18679 , \18678 );
not \U$18010 ( \18680 , \18679 );
and \U$18011 ( \18681 , \18641 , \18680 );
buf \U$18012 ( \18682 , \18519 );
buf \U$18013 ( \18683 , \18636 );
nand \U$18014 ( \18684 , \18682 , \18683 );
buf \U$18015 ( \18685 , \18684 );
buf \U$18016 ( \18686 , \18340 );
or \U$18017 ( \18687 , \18685 , \18686 );
not \U$18018 ( \18688 , \18519 );
nand \U$18019 ( \18689 , \18688 , \18683 );
not \U$18020 ( \18690 , \18689 );
nand \U$18021 ( \18691 , \18690 , \18686 );
nand \U$18022 ( \18692 , \18687 , \18691 );
nor \U$18023 ( \18693 , \18681 , \18692 );
nor \U$18024 ( \18694 , \18638 , \18587 );
buf \U$18025 ( \18695 , \18694 );
nand \U$18026 ( \18696 , \18695 , \18679 );
nand \U$18027 ( \18697 , \18693 , \18696 );
xnor \U$18028 ( \18698 , \18620 , \18697 );
xor \U$18029 ( \18699 , \18600 , \18698 );
not \U$18030 ( \18700 , \18699 );
and \U$18031 ( \18701 , \18415 , \17643 );
not \U$18032 ( \18702 , \18415 );
and \U$18033 ( \18703 , \18702 , \17642 );
nor \U$18034 ( \18704 , \18701 , \18703 );
not \U$18035 ( \18705 , \18704 );
not \U$18036 ( \18706 , \17653 );
not \U$18037 ( \18707 , \18706 );
and \U$18038 ( \18708 , \18705 , \18707 );
not \U$18039 ( \18709 , \17806 );
not \U$18040 ( \18710 , \17936 );
not \U$18041 ( \18711 , \17642 );
or \U$18042 ( \18712 , \18710 , \18711 );
buf \U$18043 ( \18713 , \17935 );
not \U$18044 ( \18714 , \18713 );
or \U$18045 ( \18715 , \17642 , \18714 );
nand \U$18046 ( \18716 , \18712 , \18715 );
and \U$18047 ( \18717 , \18709 , \18716 );
nor \U$18048 ( \18718 , \18708 , \18717 );
or \U$18049 ( \18719 , \17475 , \8793 );
or \U$18050 ( \18720 , \17852 , \8768 );
nand \U$18051 ( \18721 , \18719 , \18720 );
not \U$18052 ( \18722 , RIaaa50f0_467);
nor \U$18053 ( \18723 , \18722 , \17508 );
nor \U$18054 ( \18724 , \18721 , \18723 );
not \U$18055 ( \18725 , \12220 );
not \U$18056 ( \18726 , RIaaa4cb8_458);
not \U$18057 ( \18727 , \18726 );
and \U$18058 ( \18728 , \18725 , \18727 );
and \U$18059 ( \18729 , \17861 , RIaaa4f88_464);
nor \U$18060 ( \18730 , \18728 , \18729 );
and \U$18061 ( \18731 , \17501 , RIaaa4f10_463);
and \U$18062 ( \18732 , \11982 , RIaaa49e8_452);
nor \U$18063 ( \18733 , \18731 , \18732 );
and \U$18064 ( \18734 , \11953 , RIaaa4a60_453);
and \U$18065 ( \18735 , \17506 , RIaaa4e98_462);
nor \U$18066 ( \18736 , \18734 , \18735 );
nand \U$18067 ( \18737 , \18724 , \18730 , \18733 , \18736 );
not \U$18068 ( \18738 , \17690 );
not \U$18069 ( \18739 , \8771 );
and \U$18070 ( \18740 , \18738 , \18739 );
and \U$18071 ( \18741 , \17870 , RIaaa4d30_459);
nor \U$18072 ( \18742 , \18740 , \18741 );
not \U$18073 ( \18743 , \17499 );
not \U$18074 ( \18744 , RIaaa5168_468);
not \U$18075 ( \18745 , \18744 );
and \U$18076 ( \18746 , \18743 , \18745 );
and \U$18077 ( \18747 , \12209 , RIaaa5000_465);
nor \U$18078 ( \18748 , \18746 , \18747 );
and \U$18079 ( \18749 , \12233 , RIaaa5078_466);
and \U$18080 ( \18750 , \17493 , RIaaa4c40_457);
and \U$18081 ( \18751 , \17487 , RIaaa4bc8_456);
nor \U$18082 ( \18752 , \18749 , \18750 , \18751 );
nand \U$18083 ( \18753 , \18742 , \18748 , \18752 , \14493 );
or \U$18084 ( \18754 , \18737 , \18753 );
buf \U$18085 ( \18755 , \18754 );
not \U$18086 ( \18756 , \18755 );
not \U$18087 ( \18757 , \18538 );
not \U$18088 ( \18758 , \18757 );
not \U$18089 ( \18759 , \18758 );
or \U$18090 ( \18760 , \18756 , \18759 );
not \U$18091 ( \18761 , \18502 );
and \U$18092 ( \18762 , \18590 , \18761 );
not \U$18093 ( \18763 , \18583 );
nor \U$18094 ( \18764 , \18763 , \18761 );
nor \U$18095 ( \18765 , \18762 , \18764 );
nand \U$18096 ( \18766 , \18760 , \18765 );
buf \U$18097 ( \18767 , \18594 );
nor \U$18098 ( \18768 , \18767 , \18755 );
nor \U$18099 ( \18769 , \18766 , \18768 );
xor \U$18100 ( \18770 , \18718 , \18769 );
not \U$18101 ( \18771 , \17717 );
nand \U$18102 ( \18772 , \18771 , \18536 );
and \U$18103 ( \18773 , \18772 , \18713 );
nor \U$18104 ( \18774 , \18771 , \18536 );
nor \U$18105 ( \18775 , \18773 , \18774 );
nand \U$18106 ( \18776 , \17634 , \18775 );
not \U$18107 ( \18777 , \18369 );
and \U$18108 ( \18778 , \18777 , \18366 );
or \U$18109 ( \18779 , \18085 , \17992 );
or \U$18110 ( \18780 , \18777 , \18373 );
nand \U$18111 ( \18781 , \18779 , \18780 );
nor \U$18112 ( \18782 , \18778 , \18781 );
nor \U$18113 ( \18783 , \18776 , \18782 );
not \U$18114 ( \18784 , \18783 );
not \U$18115 ( \18785 , \18784 );
nand \U$18116 ( \18786 , \17652 , \18713 );
not \U$18117 ( \18787 , \18786 );
or \U$18118 ( \18788 , \18785 , \18787 );
not \U$18119 ( \18789 , \18783 );
not \U$18120 ( \18790 , \18786 );
or \U$18121 ( \18791 , \18789 , \18790 );
or \U$18122 ( \18792 , \18786 , \18783 );
nand \U$18123 ( \18793 , \18791 , \18792 );
not \U$18124 ( \18794 , \18683 );
not \U$18125 ( \18795 , \18794 );
not \U$18126 ( \18796 , \18755 );
and \U$18127 ( \18797 , \18639 , \18796 );
not \U$18128 ( \18798 , \18639 );
and \U$18129 ( \18799 , \18798 , \18755 );
nor \U$18130 ( \18800 , \18797 , \18799 );
not \U$18131 ( \18801 , \18800 );
or \U$18132 ( \18802 , \18795 , \18801 );
not \U$18133 ( \18803 , \18680 );
not \U$18134 ( \18804 , \18639 );
or \U$18135 ( \18805 , \18803 , \18804 );
not \U$18136 ( \18806 , \18639 );
and \U$18137 ( \18807 , \18806 , \18679 );
nor \U$18138 ( \18808 , \18807 , \18794 );
nand \U$18139 ( \18809 , \18805 , \18808 );
buf \U$18140 ( \18810 , \18638 );
nand \U$18141 ( \18811 , \18809 , \18810 );
nand \U$18142 ( \18812 , \18802 , \18811 );
nand \U$18143 ( \18813 , \18793 , \18812 );
nand \U$18144 ( \18814 , \18788 , \18813 );
xor \U$18145 ( \18815 , \18770 , \18814 );
not \U$18146 ( \18816 , \18815 );
and \U$18147 ( \18817 , \18123 , \18243 );
or \U$18148 ( \18818 , \18161 , \18292 );
or \U$18149 ( \18819 , \18127 , \18243 );
not \U$18150 ( \18820 , \18292 );
or \U$18151 ( \18821 , \18166 , \18820 );
nand \U$18152 ( \18822 , \18818 , \18819 , \18821 );
nor \U$18153 ( \18823 , \18817 , \18822 );
not \U$18154 ( \18824 , \18242 );
not \U$18155 ( \18825 , \18824 );
and \U$18156 ( \18826 , \18825 , \18679 );
not \U$18157 ( \18827 , \18677 );
not \U$18158 ( \18828 , \18196 );
or \U$18159 ( \18829 , \18827 , \18828 );
and \U$18160 ( \18830 , \18686 , \18300 );
not \U$18161 ( \18831 , \18686 );
not \U$18162 ( \18832 , \18294 );
and \U$18163 ( \18833 , \18831 , \18832 );
nor \U$18164 ( \18834 , \18830 , \18833 );
nand \U$18165 ( \18835 , \18829 , \18834 );
nor \U$18166 ( \18836 , \18826 , \18835 );
xor \U$18167 ( \18837 , \18823 , \18836 );
not \U$18168 ( \18838 , \18782 );
not \U$18169 ( \18839 , \18776 );
or \U$18170 ( \18840 , \18838 , \18839 );
nand \U$18171 ( \18841 , \18840 , \18784 );
and \U$18172 ( \18842 , \18837 , \18841 );
and \U$18173 ( \18843 , \18823 , \18836 );
or \U$18174 ( \18844 , \18842 , \18843 );
not \U$18175 ( \18845 , \18366 );
not \U$18176 ( \18846 , \18085 );
or \U$18177 ( \18847 , \18845 , \18846 );
and \U$18178 ( \18848 , \18292 , \17993 );
and \U$18179 ( \18849 , \18358 , \18374 );
nor \U$18180 ( \18850 , \18848 , \18849 );
nand \U$18181 ( \18851 , \18847 , \18850 );
not \U$18182 ( \18852 , \18340 );
not \U$18183 ( \18853 , \18123 );
or \U$18184 ( \18854 , \18852 , \18853 );
not \U$18185 ( \18855 , \18340 );
and \U$18186 ( \18856 , \18855 , \18128 );
and \U$18187 ( \18857 , \18237 , \18161 );
not \U$18188 ( \18858 , \18237 );
and \U$18189 ( \18859 , \18858 , \18166 );
nor \U$18190 ( \18860 , \18857 , \18859 );
nor \U$18191 ( \18861 , \18856 , \18860 );
nand \U$18192 ( \18862 , \18854 , \18861 );
xor \U$18193 ( \18863 , \18851 , \18862 );
nor \U$18194 ( \18864 , \17740 , \17936 );
and \U$18195 ( \18865 , \18863 , \18864 );
and \U$18196 ( \18866 , \18851 , \18862 );
nor \U$18197 ( \18867 , \18865 , \18866 );
nor \U$18198 ( \18868 , \18638 , \18587 );
and \U$18199 ( \18869 , \18868 , \18761 );
not \U$18200 ( \18870 , \18502 );
nor \U$18201 ( \18871 , \18638 , \18639 );
not \U$18202 ( \18872 , \18871 );
or \U$18203 ( \18873 , \18870 , \18872 );
and \U$18204 ( \18874 , \18682 , \18683 );
and \U$18205 ( \18875 , \18796 , \18874 );
not \U$18206 ( \18876 , \18796 );
not \U$18207 ( \18877 , \18689 );
and \U$18208 ( \18878 , \18876 , \18877 );
nor \U$18209 ( \18879 , \18875 , \18878 );
nand \U$18210 ( \18880 , \18873 , \18879 );
nor \U$18211 ( \18881 , \18869 , \18880 );
xor \U$18212 ( \18882 , \18867 , \18881 );
not \U$18213 ( \18883 , \18714 );
not \U$18214 ( \18884 , \17848 );
or \U$18215 ( \18885 , \18883 , \18884 );
not \U$18216 ( \18886 , \18414 );
not \U$18217 ( \18887 , \18886 );
not \U$18218 ( \18888 , \18613 );
and \U$18219 ( \18889 , \18887 , \18888 );
not \U$18220 ( \18890 , \18887 );
and \U$18221 ( \18891 , \18890 , \18461 );
nor \U$18222 ( \18892 , \18889 , \18891 );
nand \U$18223 ( \18893 , \18885 , \18892 );
nor \U$18224 ( \18894 , \18466 , \18714 );
nor \U$18225 ( \18895 , \18893 , \18894 );
and \U$18226 ( \18896 , \18882 , \18895 );
and \U$18227 ( \18897 , \18867 , \18881 );
or \U$18228 ( \18898 , \18896 , \18897 );
xor \U$18229 ( \18899 , \18844 , \18898 );
not \U$18230 ( \18900 , \18812 );
not \U$18231 ( \18901 , \18793 );
not \U$18232 ( \18902 , \18901 );
or \U$18233 ( \18903 , \18900 , \18902 );
or \U$18234 ( \18904 , \18901 , \18812 );
nand \U$18235 ( \18905 , \18903 , \18904 );
and \U$18236 ( \18906 , \18899 , \18905 );
and \U$18237 ( \18907 , \18844 , \18898 );
nor \U$18238 ( \18908 , \18906 , \18907 );
not \U$18239 ( \18909 , \18908 );
or \U$18240 ( \18910 , \18816 , \18909 );
or \U$18241 ( \18911 , \18908 , \18815 );
nand \U$18242 ( \18912 , \18910 , \18911 );
not \U$18243 ( \18913 , \18912 );
not \U$18244 ( \18914 , \18913 );
or \U$18245 ( \18915 , \18700 , \18914 );
not \U$18246 ( \18916 , \18699 );
nand \U$18247 ( \18917 , \18916 , \18912 );
nand \U$18248 ( \18918 , \18915 , \18917 );
xor \U$18249 ( \18919 , \18385 , \18468 );
xor \U$18250 ( \18920 , \18919 , \18596 );
xor \U$18251 ( \18921 , \18823 , \18836 );
xor \U$18252 ( \18922 , \18921 , \18841 );
not \U$18253 ( \18923 , \18581 );
not \U$18254 ( \18924 , \18758 );
or \U$18255 ( \18925 , \18923 , \18924 );
buf \U$18256 ( \18926 , \18582 );
not \U$18257 ( \18927 , \18926 );
and \U$18258 ( \18928 , \18455 , \18927 );
not \U$18259 ( \18929 , \18455 );
not \U$18260 ( \18930 , \18590 );
not \U$18261 ( \18931 , \18930 );
and \U$18262 ( \18932 , \18929 , \18931 );
nor \U$18263 ( \18933 , \18928 , \18932 );
nand \U$18264 ( \18934 , \18925 , \18933 );
nor \U$18265 ( \18935 , \18767 , \18581 );
nor \U$18266 ( \18936 , \18934 , \18935 );
xor \U$18267 ( \18937 , \18922 , \18936 );
not \U$18268 ( \18938 , \18755 );
not \U$18269 ( \18939 , \18196 );
or \U$18270 ( \18940 , \18938 , \18939 );
and \U$18271 ( \18941 , \18678 , \18832 );
not \U$18272 ( \18942 , \18678 );
and \U$18273 ( \18943 , \18942 , \18300 );
nor \U$18274 ( \18944 , \18941 , \18943 );
nand \U$18275 ( \18945 , \18940 , \18944 );
and \U$18276 ( \18946 , \18825 , \18796 );
nor \U$18277 ( \18947 , \18945 , \18946 );
not \U$18278 ( \18948 , \18947 );
not \U$18279 ( \18949 , \17993 );
not \U$18280 ( \18950 , \18238 );
or \U$18281 ( \18951 , \18949 , \18950 );
and \U$18282 ( \18952 , \18292 , \18374 );
and \U$18283 ( \18953 , \18291 , \18366 );
nor \U$18284 ( \18954 , \18952 , \18953 );
nand \U$18285 ( \18955 , \18951 , \18954 );
not \U$18286 ( \18956 , \18677 );
not \U$18287 ( \18957 , \18123 );
or \U$18288 ( \18958 , \18956 , \18957 );
and \U$18289 ( \18959 , \18128 , \18676 );
and \U$18290 ( \18960 , \18339 , \18161 );
not \U$18291 ( \18961 , \18339 );
and \U$18292 ( \18962 , \18961 , \18166 );
nor \U$18293 ( \18963 , \18960 , \18962 );
nor \U$18294 ( \18964 , \18959 , \18963 );
nand \U$18295 ( \18965 , \18958 , \18964 );
and \U$18296 ( \18966 , \18955 , \18965 );
not \U$18297 ( \18967 , \18966 );
not \U$18298 ( \18968 , \18967 );
and \U$18299 ( \18969 , \18948 , \18968 );
not \U$18300 ( \18970 , \18581 );
not \U$18301 ( \18971 , \18970 );
not \U$18302 ( \18972 , \18695 );
or \U$18303 ( \18973 , \18971 , \18972 );
and \U$18304 ( \18974 , \18641 , \18581 );
or \U$18305 ( \18975 , \18685 , \18502 );
buf \U$18306 ( \18976 , \18690 );
nand \U$18307 ( \18977 , \18976 , \18502 );
nand \U$18308 ( \18978 , \18975 , \18977 );
nor \U$18309 ( \18979 , \18974 , \18978 );
nand \U$18310 ( \18980 , \18973 , \18979 );
and \U$18311 ( \18981 , \18947 , \18966 );
not \U$18312 ( \18982 , \18947 );
and \U$18313 ( \18983 , \18982 , \18967 );
nor \U$18314 ( \18984 , \18981 , \18983 );
not \U$18315 ( \18985 , \18984 );
and \U$18316 ( \18986 , \18980 , \18985 );
nor \U$18317 ( \18987 , \18969 , \18986 );
and \U$18318 ( \18988 , \18937 , \18987 );
and \U$18319 ( \18989 , \18922 , \18936 );
or \U$18320 ( \18990 , \18988 , \18989 );
xor \U$18321 ( \18991 , \18920 , \18990 );
xor \U$18322 ( \18992 , \18899 , \18905 );
and \U$18323 ( \18993 , \18991 , \18992 );
and \U$18324 ( \18994 , \18920 , \18990 );
or \U$18325 ( \18995 , \18993 , \18994 );
nand \U$18326 ( \18996 , \18918 , \18995 );
xor \U$18327 ( \18997 , \18920 , \18990 );
xor \U$18328 ( \18998 , \18997 , \18992 );
xor \U$18329 ( \18999 , \18867 , \18881 );
xor \U$18330 ( \19000 , \18999 , \18895 );
xnor \U$18331 ( \19001 , \18863 , \18864 );
not \U$18332 ( \19002 , \19001 );
not \U$18333 ( \19003 , \19002 );
not \U$18334 ( \19004 , \18611 );
and \U$18335 ( \19005 , \18535 , \18588 );
not \U$18336 ( \19006 , \19005 );
or \U$18337 ( \19007 , \19004 , \19006 );
buf \U$18338 ( \19008 , \18538 );
and \U$18339 ( \19009 , \18455 , \19008 );
not \U$18340 ( \19010 , \18886 );
not \U$18341 ( \19011 , \18590 );
or \U$18342 ( \19012 , \19010 , \19011 );
not \U$18343 ( \19013 , \18416 );
nand \U$18344 ( \19014 , \18583 , \19013 );
nand \U$18345 ( \19015 , \19012 , \19014 );
nor \U$18346 ( \19016 , \19009 , \19015 );
nand \U$18347 ( \19017 , \19007 , \19016 );
xor \U$18348 ( \19018 , \18955 , \18965 );
not \U$18349 ( \19019 , \18502 );
not \U$18350 ( \19020 , \19019 );
not \U$18351 ( \19021 , \18825 );
or \U$18352 ( \19022 , \19020 , \19021 );
and \U$18353 ( \19023 , \18196 , \18502 );
not \U$18354 ( \19024 , \18300 );
and \U$18355 ( \19025 , \18755 , \19024 );
not \U$18356 ( \19026 , \18755 );
not \U$18357 ( \19027 , \18832 );
and \U$18358 ( \19028 , \19026 , \19027 );
nor \U$18359 ( \19029 , \19025 , \19028 );
nor \U$18360 ( \19030 , \19023 , \19029 );
nand \U$18361 ( \19031 , \19022 , \19030 );
xor \U$18362 ( \19032 , \19018 , \19031 );
not \U$18363 ( \19033 , \18586 );
not \U$18364 ( \19034 , \19033 );
nand \U$18365 ( \19035 , \19034 , \18587 );
not \U$18366 ( \19036 , \17936 );
and \U$18367 ( \19037 , \19035 , \19036 );
not \U$18368 ( \19038 , \19033 );
not \U$18369 ( \19039 , \18587 );
not \U$18370 ( \19040 , \19039 );
or \U$18371 ( \19041 , \19038 , \19040 );
nand \U$18372 ( \19042 , \19041 , \18588 );
nor \U$18373 ( \19043 , \19037 , \19042 );
and \U$18374 ( \19044 , \19032 , \19043 );
and \U$18375 ( \19045 , \19018 , \19031 );
nor \U$18376 ( \19046 , \19044 , \19045 );
and \U$18377 ( \19047 , \19017 , \19046 );
not \U$18378 ( \19048 , \19017 );
not \U$18379 ( \19049 , \19046 );
and \U$18380 ( \19050 , \19048 , \19049 );
or \U$18381 ( \19051 , \19047 , \19050 );
not \U$18382 ( \19052 , \19051 );
or \U$18383 ( \19053 , \19003 , \19052 );
nand \U$18384 ( \19054 , \19017 , \19049 );
nand \U$18385 ( \19055 , \19053 , \19054 );
not \U$18386 ( \19056 , \19055 );
xor \U$18387 ( \19057 , \19000 , \19056 );
xor \U$18388 ( \19058 , \18922 , \18936 );
xor \U$18389 ( \19059 , \19058 , \18987 );
and \U$18390 ( \19060 , \19057 , \19059 );
and \U$18391 ( \19061 , \19000 , \19056 );
or \U$18392 ( \19062 , \19060 , \19061 );
nor \U$18393 ( \19063 , \18998 , \19062 );
nand \U$18394 ( \19064 , \18996 , \19063 );
not \U$18395 ( \19065 , \19064 );
nor \U$18396 ( \19066 , \18918 , \18995 );
not \U$18397 ( \19067 , \17747 );
not \U$18398 ( \19068 , \18714 );
and \U$18399 ( \19069 , \19067 , \19068 );
and \U$18400 ( \19070 , \18641 , \18686 );
not \U$18401 ( \19071 , \18877 );
or \U$18402 ( \19072 , \19071 , \18244 );
not \U$18403 ( \19073 , \18244 );
or \U$18404 ( \19074 , \18685 , \19073 );
nand \U$18405 ( \19075 , \19072 , \19074 );
nor \U$18406 ( \19076 , \19070 , \19075 );
not \U$18407 ( \19077 , \18686 );
nand \U$18408 ( \19078 , \18695 , \19077 );
nand \U$18409 ( \19079 , \19076 , \19078 );
not \U$18410 ( \19080 , \19079 );
and \U$18411 ( \19081 , \18050 , \18170 );
and \U$18412 ( \19082 , \19080 , \19081 );
nor \U$18413 ( \19083 , \19069 , \19082 );
not \U$18414 ( \19084 , \19081 );
nand \U$18415 ( \19085 , \19084 , \19079 );
nand \U$18416 ( \19086 , \19083 , \19085 );
not \U$18417 ( \19087 , \18123 );
not \U$18418 ( \19088 , \18777 );
or \U$18419 ( \19089 , \19087 , \19088 );
not \U$18420 ( \19090 , \18127 );
and \U$18421 ( \19091 , \19090 , \18369 );
and \U$18422 ( \19092 , \18042 , \18160 );
not \U$18423 ( \19093 , \18042 );
and \U$18424 ( \19094 , \19093 , \18359 );
or \U$18425 ( \19095 , \19092 , \19094 );
nor \U$18426 ( \19096 , \19091 , \19095 );
nand \U$18427 ( \19097 , \19089 , \19096 );
not \U$18428 ( \19098 , \19097 );
not \U$18429 ( \19099 , \18001 );
not \U$18430 ( \19100 , \13105 );
and \U$18431 ( \19101 , \19099 , \19100 );
and \U$18432 ( \19102 , \17501 , RIaaa1dd8_358);
nor \U$18433 ( \19103 , \19101 , \19102 );
not \U$18434 ( \19104 , \12214 );
not \U$18435 ( \19105 , \7197 );
and \U$18436 ( \19106 , \19104 , \19105 );
and \U$18437 ( \19107 , \11953 , RIaaa2198_366);
nor \U$18438 ( \19108 , \19106 , \19107 );
nand \U$18439 ( \19109 , \19103 , \19108 );
not \U$18440 ( \19110 , \12220 );
not \U$18441 ( \19111 , \13102 );
and \U$18442 ( \19112 , \19110 , \19111 );
and \U$18443 ( \19113 , \12209 , RIaaa1bf8_354);
nor \U$18444 ( \19114 , \19112 , \19113 );
and \U$18445 ( \19115 , \17474 , RIaaa1d60_357);
and \U$18446 ( \19116 , \12057 , RIaaa1a90_351);
nor \U$18447 ( \19117 , \19115 , \19116 );
nand \U$18448 ( \19118 , \19114 , \19117 );
nor \U$18449 ( \19119 , \19109 , \19118 );
not \U$18450 ( \19120 , RIaaa2030_363);
not \U$18451 ( \19121 , \11985 );
or \U$18452 ( \19122 , \19120 , \19121 );
and \U$18453 ( \19123 , \12233 , RIaaa1c70_355);
and \U$18454 ( \19124 , \17493 , RIaaa1b80_353);
and \U$18455 ( \19125 , \17487 , RIaaa1b08_352);
nor \U$18456 ( \19126 , \19123 , \19124 , \19125 );
nand \U$18457 ( \19127 , \19122 , \19126 );
not \U$18458 ( \19128 , RIaaa1e50_359);
not \U$18459 ( \19129 , \11948 );
or \U$18460 ( \19130 , \19128 , \19129 );
nand \U$18461 ( \19131 , \17919 , RIaaa1ce8_356);
nand \U$18462 ( \19132 , \19130 , \19131 );
nor \U$18463 ( \19133 , \19127 , \19132 );
nand \U$18464 ( \19134 , \11966 , RIaaa1f40_361);
nand \U$18465 ( \19135 , \11951 , RIaaa1ec8_360);
and \U$18466 ( \19136 , \19134 , \19135 , \13096 );
nand \U$18467 ( \19137 , \19119 , \19133 , \19136 );
not \U$18468 ( \19138 , \19137 );
nand \U$18469 ( \19139 , \19138 , \18374 );
nand \U$18470 ( \19140 , \19137 , \18366 );
not \U$18471 ( \19141 , \17970 );
nand \U$18472 ( \19142 , \19141 , \17993 );
and \U$18473 ( \19143 , \19139 , \19140 , \19142 );
not \U$18474 ( \19144 , \19143 );
and \U$18475 ( \19145 , \19098 , \19144 );
and \U$18476 ( \19146 , \19097 , \19143 );
nor \U$18477 ( \19147 , \19145 , \19146 );
not \U$18478 ( \19148 , \19147 );
not \U$18479 ( \19149 , \18820 );
not \U$18480 ( \19150 , \18195 );
or \U$18481 ( \19151 , \19149 , \19150 );
buf \U$18482 ( \19152 , \18358 );
and \U$18483 ( \19153 , \19152 , \18295 );
not \U$18484 ( \19154 , \19152 );
and \U$18485 ( \19155 , \19154 , \18299 );
nor \U$18486 ( \19156 , \19153 , \19155 );
nand \U$18487 ( \19157 , \19151 , \19156 );
not \U$18488 ( \19158 , \19157 );
nand \U$18489 ( \19159 , \18242 , \18292 );
nand \U$18490 ( \19160 , \19158 , \19159 );
not \U$18491 ( \19161 , \19160 );
and \U$18492 ( \19162 , \19148 , \19161 );
and \U$18493 ( \19163 , \19160 , \19147 );
nor \U$18494 ( \19164 , \19162 , \19163 );
not \U$18495 ( \19165 , \19164 );
not \U$18496 ( \19166 , \18581 );
not \U$18497 ( \19167 , \18465 );
or \U$18498 ( \19168 , \19166 , \19167 );
not \U$18499 ( \19169 , \18581 );
and \U$18500 ( \19170 , \18418 , \19169 );
or \U$18501 ( \19171 , \17891 , \18502 );
nand \U$18502 ( \19172 , \18458 , \18502 );
nand \U$18503 ( \19173 , \19171 , \19172 );
nor \U$18504 ( \19174 , \19170 , \19173 );
nand \U$18505 ( \19175 , \19168 , \19174 );
not \U$18506 ( \19176 , \19175 );
or \U$18507 ( \19177 , \19165 , \19176 );
or \U$18508 ( \19178 , \19175 , \19164 );
nand \U$18509 ( \19179 , \19177 , \19178 );
not \U$18510 ( \19180 , \19179 );
not \U$18511 ( \19181 , \18680 );
not \U$18512 ( \19182 , \18538 );
or \U$18513 ( \19183 , \19181 , \19182 );
and \U$18514 ( \19184 , \18755 , \18583 );
not \U$18515 ( \19185 , \18755 );
buf \U$18516 ( \19186 , \18589 );
not \U$18517 ( \19187 , \19186 );
and \U$18518 ( \19188 , \19185 , \19187 );
nor \U$18519 ( \19189 , \19184 , \19188 );
nand \U$18520 ( \19190 , \19183 , \19189 );
nor \U$18521 ( \19191 , \18594 , \18680 );
nor \U$18522 ( \19192 , \19190 , \19191 );
not \U$18523 ( \19193 , \19192 );
or \U$18524 ( \19194 , \19180 , \19193 );
or \U$18525 ( \19195 , \19192 , \19179 );
nand \U$18526 ( \19196 , \19194 , \19195 );
xor \U$18527 ( \19197 , \19086 , \19196 );
not \U$18528 ( \19198 , \18607 );
not \U$18529 ( \19199 , \18697 );
or \U$18530 ( \19200 , \19198 , \19199 );
or \U$18531 ( \19201 , \18697 , \18607 );
nand \U$18532 ( \19202 , \19201 , \18619 );
nand \U$18533 ( \19203 , \19200 , \19202 );
or \U$18534 ( \19204 , \17939 , \18304 );
nand \U$18535 ( \19205 , \19204 , \18306 );
not \U$18536 ( \19206 , \19205 );
not \U$18537 ( \19207 , \18611 );
not \U$18538 ( \19208 , \17642 );
or \U$18539 ( \19209 , \19207 , \19208 );
or \U$18540 ( \19210 , \17642 , \18611 );
nand \U$18541 ( \19211 , \19209 , \19210 );
not \U$18542 ( \19212 , \19211 );
not \U$18543 ( \19213 , \17653 );
or \U$18544 ( \19214 , \19212 , \19213 );
not \U$18545 ( \19215 , \18704 );
nand \U$18546 ( \19216 , \19215 , \17641 );
nand \U$18547 ( \19217 , \19214 , \19216 );
not \U$18548 ( \19218 , \19217 );
not \U$18549 ( \19219 , \19218 );
or \U$18550 ( \19220 , \19206 , \19219 );
not \U$18551 ( \19221 , \19205 );
nand \U$18552 ( \19222 , \19221 , \19217 );
nand \U$18553 ( \19223 , \19220 , \19222 );
and \U$18554 ( \19224 , \19203 , \19223 );
not \U$18555 ( \19225 , \19203 );
not \U$18556 ( \19226 , \19223 );
and \U$18557 ( \19227 , \19225 , \19226 );
nor \U$18558 ( \19228 , \19224 , \19227 );
xnor \U$18559 ( \19229 , \19197 , \19228 );
not \U$18560 ( \19230 , \19229 );
xor \U$18561 ( \19231 , \18718 , \18769 );
and \U$18562 ( \19232 , \19231 , \18814 );
and \U$18563 ( \19233 , \18718 , \18769 );
or \U$18564 ( \19234 , \19232 , \19233 );
not \U$18565 ( \19235 , \19234 );
and \U$18566 ( \19236 , \18600 , \18698 );
and \U$18567 ( \19237 , \18311 , \18599 );
nor \U$18568 ( \19238 , \19236 , \19237 );
nor \U$18569 ( \19239 , \19235 , \19238 );
not \U$18570 ( \19240 , \19239 );
not \U$18571 ( \19241 , \19234 );
nand \U$18572 ( \19242 , \19241 , \19238 );
nand \U$18573 ( \19243 , \19240 , \19242 );
not \U$18574 ( \19244 , \19243 );
or \U$18575 ( \19245 , \19230 , \19244 );
or \U$18576 ( \19246 , \19243 , \19229 );
nand \U$18577 ( \19247 , \19245 , \19246 );
not \U$18578 ( \19248 , \18699 );
not \U$18579 ( \19249 , \18912 );
or \U$18580 ( \19250 , \19248 , \19249 );
not \U$18581 ( \19251 , \18908 );
nand \U$18582 ( \19252 , \19251 , \18815 );
nand \U$18583 ( \19253 , \19250 , \19252 );
nor \U$18584 ( \19254 , \19247 , \19253 );
nor \U$18585 ( \19255 , \19066 , \19254 );
not \U$18586 ( \19256 , \19197 );
not \U$18587 ( \19257 , \19228 );
or \U$18588 ( \19258 , \19256 , \19257 );
nand \U$18589 ( \19259 , \19196 , \19086 );
nand \U$18590 ( \19260 , \19258 , \19259 );
not \U$18591 ( \19261 , \19152 );
and \U$18592 ( \19262 , \18196 , \19261 );
or \U$18593 ( \19263 , \18777 , \19027 );
nand \U$18594 ( \19264 , \18300 , \18777 );
nand \U$18595 ( \19265 , \19263 , \19264 );
nor \U$18596 ( \19266 , \19262 , \19265 );
nand \U$18597 ( \19267 , \18825 , \19152 );
nand \U$18598 ( \19268 , \19266 , \19267 );
not \U$18599 ( \19269 , \19268 );
not \U$18600 ( \19270 , \18365 );
not \U$18601 ( \19271 , \18123 );
or \U$18602 ( \19272 , \19270 , \19271 );
not \U$18603 ( \19273 , \18365 );
and \U$18604 ( \19274 , \18128 , \19273 );
or \U$18605 ( \19275 , \18161 , \19141 );
nand \U$18606 ( \19276 , \18359 , \19141 );
nand \U$18607 ( \19277 , \19275 , \19276 );
nor \U$18608 ( \19278 , \19274 , \19277 );
nand \U$18609 ( \19279 , \19272 , \19278 );
not \U$18610 ( \19280 , \19279 );
and \U$18611 ( \19281 , \19138 , \17993 );
and \U$18612 ( \19282 , \17684 , RIaaa0de8_324);
and \U$18613 ( \19283 , \12231 , RIaaa0d70_323);
nor \U$18614 ( \19284 , \19282 , \19283 );
not \U$18615 ( \19285 , \12214 );
not \U$18616 ( \19286 , \1946 );
and \U$18617 ( \19287 , \19285 , \19286 );
and \U$18618 ( \19288 , \17686 , RIaaa0e60_325);
nor \U$18619 ( \19289 , \19287 , \19288 );
not \U$18620 ( \19290 , \17690 );
not \U$18621 ( \19291 , \13181 );
and \U$18622 ( \19292 , \19290 , \19291 );
and \U$18623 ( \19293 , \11969 , RIaaa0aa0_317);
nor \U$18624 ( \19294 , \19292 , \19293 );
nand \U$18625 ( \19295 , \19284 , \19289 , \19294 , \13220 );
not \U$18626 ( \19296 , RIaaa0c08_320);
or \U$18627 ( \19297 , \17669 , \19296 );
and \U$18628 ( \19298 , \17493 , RIaaa1040_329);
and \U$18629 ( \19299 , \17487 , RIaaa0fc8_328);
nor \U$18630 ( \19300 , \19298 , \19299 );
nand \U$18631 ( \19301 , \19297 , \19300 );
not \U$18632 ( \19302 , RIaaa0cf8_322);
nor \U$18633 ( \19303 , \19302 , \17508 );
nor \U$18634 ( \19304 , \19301 , \19303 );
not \U$18635 ( \19305 , \12210 );
not \U$18636 ( \19306 , RIaaa0c80_321);
not \U$18637 ( \19307 , \19306 );
and \U$18638 ( \19308 , \19305 , \19307 );
and \U$18639 ( \19309 , \11953 , RIaaa10b8_330);
nor \U$18640 ( \19310 , \19308 , \19309 );
and \U$18641 ( \19311 , \11948 , RIaaa0b18_318);
and \U$18642 ( \19312 , \17861 , RIaaa0a28_316);
nor \U$18643 ( \19313 , \19311 , \19312 );
and \U$18644 ( \19314 , \17474 , RIaaa0ed8_326);
and \U$18645 ( \19315 , \12057 , RIaaa0f50_327);
nor \U$18646 ( \19316 , \19314 , \19315 );
nand \U$18647 ( \19317 , \19304 , \19310 , \19313 , \19316 );
nor \U$18648 ( \19318 , \19295 , \19317 );
and \U$18649 ( \19319 , \19318 , \18374 );
nor \U$18650 ( \19320 , \19281 , \19319 );
not \U$18651 ( \19321 , \19318 );
nand \U$18652 ( \19322 , \19321 , \18366 );
and \U$18653 ( \19323 , \19320 , \19322 );
not \U$18654 ( \19324 , \19323 );
and \U$18655 ( \19325 , \19280 , \19324 );
and \U$18656 ( \19326 , \19279 , \19323 );
nor \U$18657 ( \19327 , \19325 , \19326 );
not \U$18658 ( \19328 , \19327 );
and \U$18659 ( \19329 , \19269 , \19328 );
and \U$18660 ( \19330 , \19268 , \19327 );
nor \U$18661 ( \19331 , \19329 , \19330 );
and \U$18662 ( \19332 , \19079 , \19081 );
xor \U$18663 ( \19333 , \19331 , \19332 );
not \U$18664 ( \19334 , \18502 );
not \U$18665 ( \19335 , \17844 );
or \U$18666 ( \19336 , \19334 , \19335 );
and \U$18667 ( \19337 , \17848 , \18761 );
and \U$18668 ( \19338 , \18755 , \18613 );
not \U$18669 ( \19339 , \18755 );
and \U$18670 ( \19340 , \19339 , \17891 );
nor \U$18671 ( \19341 , \19338 , \19340 );
nor \U$18672 ( \19342 , \19337 , \19341 );
nand \U$18673 ( \19343 , \19336 , \19342 );
not \U$18674 ( \19344 , \19343 );
not \U$18675 ( \19345 , \19344 );
not \U$18676 ( \19346 , \19147 );
not \U$18677 ( \19347 , \19346 );
not \U$18678 ( \19348 , \19160 );
or \U$18679 ( \19349 , \19347 , \19348 );
not \U$18680 ( \19350 , \19143 );
nand \U$18681 ( \19351 , \19350 , \19097 );
nand \U$18682 ( \19352 , \19349 , \19351 );
not \U$18683 ( \19353 , \19352 );
not \U$18684 ( \19354 , \19353 );
and \U$18685 ( \19355 , \19073 , \18871 );
and \U$18686 ( \19356 , \18292 , \18684 );
not \U$18687 ( \19357 , \18292 );
and \U$18688 ( \19358 , \19357 , \18689 );
nor \U$18689 ( \19359 , \19356 , \19358 );
nor \U$18690 ( \19360 , \19355 , \19359 );
nand \U$18691 ( \19361 , \18868 , \18244 );
nand \U$18692 ( \19362 , \19360 , \19361 );
not \U$18693 ( \19363 , \19362 );
or \U$18694 ( \19364 , \19354 , \19363 );
nand \U$18695 ( \19365 , \19352 , \19361 , \19360 );
nand \U$18696 ( \19366 , \19364 , \19365 );
buf \U$18697 ( \19367 , \19366 );
not \U$18698 ( \19368 , \19367 );
or \U$18699 ( \19369 , \19345 , \19368 );
or \U$18700 ( \19370 , \19367 , \19344 );
nand \U$18701 ( \19371 , \19369 , \19370 );
xnor \U$18702 ( \19372 , \19333 , \19371 );
xor \U$18703 ( \19373 , \19260 , \19372 );
not \U$18704 ( \19374 , \19192 );
not \U$18705 ( \19375 , \19374 );
not \U$18706 ( \19376 , \19179 );
or \U$18707 ( \19377 , \19375 , \19376 );
not \U$18708 ( \19378 , \19164 );
nand \U$18709 ( \19379 , \19378 , \19175 );
nand \U$18710 ( \19380 , \19377 , \19379 );
and \U$18711 ( \19381 , \18680 , \18927 );
not \U$18712 ( \19382 , \18680 );
and \U$18713 ( \19383 , \19382 , \18590 );
nor \U$18714 ( \19384 , \19381 , \19383 );
buf \U$18715 ( \19385 , \18535 );
or \U$18716 ( \19386 , \19077 , \18588 );
not \U$18717 ( \19387 , \18588 );
or \U$18718 ( \19388 , \18686 , \19387 );
nand \U$18719 ( \19389 , \19386 , \19388 );
and \U$18720 ( \19390 , \19385 , \19389 );
and \U$18721 ( \19391 , \17746 , \19013 );
nor \U$18722 ( \19392 , \19390 , \19391 );
nand \U$18723 ( \19393 , \19384 , \19392 );
not \U$18724 ( \19394 , \19393 );
or \U$18725 ( \19395 , \18970 , \17655 );
not \U$18726 ( \19396 , \18581 );
nand \U$18727 ( \19397 , \19396 , \17705 );
nand \U$18728 ( \19398 , \19395 , \19397 );
not \U$18729 ( \19399 , \19211 );
nor \U$18730 ( \19400 , \19399 , \17807 );
nor \U$18731 ( \19401 , \19398 , \19400 );
not \U$18732 ( \19402 , \19401 );
or \U$18733 ( \19403 , \19394 , \19402 );
or \U$18734 ( \19404 , \19401 , \19393 );
nand \U$18735 ( \19405 , \19403 , \19404 );
xor \U$18736 ( \19406 , \19380 , \19405 );
not \U$18737 ( \19407 , \19223 );
not \U$18738 ( \19408 , \19203 );
or \U$18739 ( \19409 , \19407 , \19408 );
nand \U$18740 ( \19410 , \19217 , \19205 );
nand \U$18741 ( \19411 , \19409 , \19410 );
xor \U$18742 ( \19412 , \19406 , \19411 );
xor \U$18743 ( \19413 , \19373 , \19412 );
or \U$18744 ( \19414 , \19229 , \19239 );
nand \U$18745 ( \19415 , \19414 , \19242 );
nand \U$18746 ( \19416 , \19413 , \19415 );
nand \U$18747 ( \19417 , \19255 , \19416 );
nor \U$18748 ( \19418 , \19065 , \19417 );
not \U$18749 ( \19419 , \19418 );
not \U$18750 ( \19420 , \18695 );
not \U$18751 ( \19421 , \19420 );
not \U$18752 ( \19422 , \19013 );
and \U$18753 ( \19423 , \19421 , \19422 );
not \U$18754 ( \19424 , \18887 );
not \U$18755 ( \19425 , \18641 );
or \U$18756 ( \19426 , \19424 , \19425 );
and \U$18757 ( \19427 , \18611 , \18874 );
not \U$18758 ( \19428 , \18611 );
and \U$18759 ( \19429 , \19428 , \18877 );
nor \U$18760 ( \19430 , \19427 , \19429 );
nand \U$18761 ( \19431 , \19426 , \19430 );
nor \U$18762 ( \19432 , \19423 , \19431 );
not \U$18763 ( \19433 , \18122 );
not \U$18764 ( \19434 , \19019 );
and \U$18765 ( \19435 , \19433 , \19434 );
or \U$18766 ( \19436 , \18127 , \18502 );
and \U$18767 ( \19437 , \18754 , \18160 );
not \U$18768 ( \19438 , \18754 );
and \U$18769 ( \19439 , \19438 , \18359 );
nor \U$18770 ( \19440 , \19437 , \19439 );
nand \U$18771 ( \19441 , \19436 , \19440 );
nor \U$18772 ( \19442 , \19435 , \19441 );
not \U$18773 ( \19443 , \19442 );
nand \U$18774 ( \19444 , \18193 , \17936 );
and \U$18775 ( \19445 , \19444 , \18627 );
and \U$18776 ( \19446 , \18713 , \18194 );
nor \U$18777 ( \19447 , \19445 , \19446 );
and \U$18778 ( \19448 , \18639 , \19447 );
nand \U$18779 ( \19449 , \19443 , \19448 );
nand \U$18780 ( \19450 , \19385 , \18713 );
and \U$18781 ( \19451 , \19449 , \19450 );
or \U$18782 ( \19452 , \19432 , \19451 );
or \U$18783 ( \19453 , \19449 , \19450 );
nand \U$18784 ( \19454 , \19452 , \19453 );
not \U$18785 ( \19455 , \19454 );
xnor \U$18786 ( \19456 , \19043 , \19032 );
not \U$18787 ( \19457 , \19456 );
and \U$18788 ( \19458 , \19455 , \19457 );
and \U$18789 ( \19459 , \19454 , \19456 );
nor \U$18790 ( \19460 , \19458 , \19459 );
not \U$18791 ( \19461 , \19460 );
not \U$18792 ( \19462 , \19461 );
and \U$18793 ( \19463 , \18243 , \18366 );
and \U$18794 ( \19464 , \18855 , \17993 );
and \U$18795 ( \19465 , \18238 , \18374 );
nor \U$18796 ( \19466 , \19463 , \19464 , \19465 );
not \U$18797 ( \19467 , \18121 );
and \U$18798 ( \19468 , \18755 , \19467 );
not \U$18799 ( \19469 , \18755 );
and \U$18800 ( \19470 , \19469 , \18121 );
nor \U$18801 ( \19471 , \19468 , \19470 );
and \U$18802 ( \19472 , \19471 , \18119 );
nor \U$18803 ( \19473 , \19472 , \18165 );
and \U$18804 ( \19474 , \18678 , \18121 );
and \U$18805 ( \19475 , \18677 , \19467 );
nor \U$18806 ( \19476 , \19474 , \19475 );
nor \U$18807 ( \19477 , \19476 , \18119 );
or \U$18808 ( \19478 , \19473 , \19477 );
xor \U$18809 ( \19479 , \19466 , \19478 );
not \U$18810 ( \19480 , \18824 );
not \U$18811 ( \19481 , \18581 );
and \U$18812 ( \19482 , \19480 , \19481 );
not \U$18813 ( \19483 , \18581 );
not \U$18814 ( \19484 , \18196 );
or \U$18815 ( \19485 , \19483 , \19484 );
and \U$18816 ( \19486 , \18502 , \18300 );
not \U$18817 ( \19487 , \18502 );
and \U$18818 ( \19488 , \19487 , \18295 );
nor \U$18819 ( \19489 , \19486 , \19488 );
nand \U$18820 ( \19490 , \19485 , \19489 );
nor \U$18821 ( \19491 , \19482 , \19490 );
and \U$18822 ( \19492 , \19479 , \19491 );
and \U$18823 ( \19493 , \19466 , \19478 );
or \U$18824 ( \19494 , \19492 , \19493 );
not \U$18825 ( \19495 , \19494 );
and \U$18826 ( \19496 , \18641 , \18455 );
not \U$18827 ( \19497 , \18690 );
or \U$18828 ( \19498 , \19497 , \19169 );
nand \U$18829 ( \19499 , \18874 , \19169 );
nand \U$18830 ( \19500 , \19498 , \19499 );
nor \U$18831 ( \19501 , \19496 , \19500 );
nand \U$18832 ( \19502 , \18695 , \18611 );
nand \U$18833 ( \19503 , \19501 , \19502 );
not \U$18834 ( \19504 , \18887 );
not \U$18835 ( \19505 , \18538 );
or \U$18836 ( \19506 , \19504 , \19505 );
and \U$18837 ( \19507 , \18713 , \18583 );
not \U$18838 ( \19508 , \18713 );
and \U$18839 ( \19509 , \19508 , \18590 );
nor \U$18840 ( \19510 , \19507 , \19509 );
nand \U$18841 ( \19511 , \19506 , \19510 );
nor \U$18842 ( \19512 , \18594 , \18415 );
nor \U$18843 ( \19513 , \19511 , \19512 );
xnor \U$18844 ( \19514 , \19503 , \19513 );
not \U$18845 ( \19515 , \19514 );
or \U$18846 ( \19516 , \19495 , \19515 );
or \U$18847 ( \19517 , \19514 , \19494 );
nand \U$18848 ( \19518 , \19516 , \19517 );
not \U$18849 ( \19519 , \19518 );
or \U$18850 ( \19520 , \19462 , \19519 );
not \U$18851 ( \19521 , \19456 );
nand \U$18852 ( \19522 , \19521 , \19454 );
nand \U$18853 ( \19523 , \19520 , \19522 );
xor \U$18854 ( \19524 , \19051 , \19001 );
not \U$18855 ( \19525 , \18984 );
not \U$18856 ( \19526 , \18980 );
or \U$18857 ( \19527 , \19525 , \19526 );
or \U$18858 ( \19528 , \18980 , \18984 );
nand \U$18859 ( \19529 , \19527 , \19528 );
not \U$18860 ( \19530 , \19494 );
not \U$18861 ( \19531 , \19530 );
not \U$18862 ( \19532 , \19514 );
or \U$18863 ( \19533 , \19531 , \19532 );
not \U$18864 ( \19534 , \19513 );
nand \U$18865 ( \19535 , \19534 , \19503 );
nand \U$18866 ( \19536 , \19533 , \19535 );
xor \U$18867 ( \19537 , \19529 , \19536 );
xnor \U$18868 ( \19538 , \19524 , \19537 );
xor \U$18869 ( \19539 , \19523 , \19538 );
not \U$18870 ( \19540 , \19460 );
not \U$18871 ( \19541 , \19518 );
or \U$18872 ( \19542 , \19540 , \19541 );
or \U$18873 ( \19543 , \19518 , \19460 );
nand \U$18874 ( \19544 , \19542 , \19543 );
not \U$18875 ( \19545 , \19544 );
xor \U$18876 ( \19546 , \19466 , \19478 );
xor \U$18877 ( \19547 , \19546 , \19491 );
not \U$18878 ( \19548 , \19442 );
not \U$18879 ( \19549 , \19448 );
or \U$18880 ( \19550 , \19548 , \19549 );
or \U$18881 ( \19551 , \19448 , \19442 );
nand \U$18882 ( \19552 , \19550 , \19551 );
not \U$18883 ( \19553 , \18241 );
not \U$18884 ( \19554 , \18455 );
and \U$18885 ( \19555 , \19553 , \19554 );
not \U$18886 ( \19556 , \18196 );
not \U$18887 ( \19557 , \18455 );
or \U$18888 ( \19558 , \19556 , \19557 );
and \U$18889 ( \19559 , \19169 , \18295 );
not \U$18890 ( \19560 , \19169 );
and \U$18891 ( \19561 , \19560 , \18300 );
nor \U$18892 ( \19562 , \19559 , \19561 );
nand \U$18893 ( \19563 , \19558 , \19562 );
nor \U$18894 ( \19564 , \19555 , \19563 );
and \U$18895 ( \19565 , \18340 , \18366 );
not \U$18896 ( \19566 , \18340 );
and \U$18897 ( \19567 , \19566 , \18374 );
nor \U$18898 ( \19568 , \19565 , \19567 );
nand \U$18899 ( \19569 , \18678 , \17993 );
and \U$18900 ( \19570 , \19568 , \19569 );
nor \U$18901 ( \19571 , \19564 , \19570 );
or \U$18902 ( \19572 , \19552 , \19571 );
nand \U$18903 ( \19573 , \19564 , \19570 );
nand \U$18904 ( \19574 , \19572 , \19573 );
xor \U$18905 ( \19575 , \19547 , \19574 );
xor \U$18906 ( \19576 , \19450 , \19449 );
xor \U$18907 ( \19577 , \19432 , \19576 );
and \U$18908 ( \19578 , \19575 , \19577 );
and \U$18909 ( \19579 , \19547 , \19574 );
or \U$18910 ( \19580 , \19578 , \19579 );
not \U$18911 ( \19581 , \19580 );
and \U$18912 ( \19582 , \19545 , \19581 );
and \U$18913 ( \19583 , \19580 , \19544 );
nor \U$18914 ( \19584 , \19582 , \19583 );
not \U$18915 ( \19585 , \19571 );
nand \U$18916 ( \19586 , \19585 , \19573 );
not \U$18917 ( \19587 , \19586 );
not \U$18918 ( \19588 , \19552 );
or \U$18919 ( \19589 , \19587 , \19588 );
or \U$18920 ( \19590 , \19552 , \19586 );
nand \U$18921 ( \19591 , \19589 , \19590 );
not \U$18922 ( \19592 , \18416 );
not \U$18923 ( \19593 , \18242 );
or \U$18924 ( \19594 , \19592 , \19593 );
and \U$18925 ( \19595 , \18196 , \18887 );
and \U$18926 ( \19596 , \18455 , \19024 );
not \U$18927 ( \19597 , \18455 );
and \U$18928 ( \19598 , \19597 , \19027 );
nor \U$18929 ( \19599 , \19596 , \19598 );
nor \U$18930 ( \19600 , \19595 , \19599 );
nand \U$18931 ( \19601 , \19594 , \19600 );
not \U$18932 ( \19602 , \19601 );
not \U$18933 ( \19603 , \18581 );
not \U$18934 ( \19604 , \18123 );
or \U$18935 ( \19605 , \19603 , \19604 );
not \U$18936 ( \19606 , \18127 );
and \U$18937 ( \19607 , \19606 , \19169 );
not \U$18938 ( \19608 , \18501 );
or \U$18939 ( \19609 , \19608 , \18161 );
or \U$18940 ( \19610 , \18501 , \18166 );
nand \U$18941 ( \19611 , \19609 , \19610 );
nor \U$18942 ( \19612 , \19607 , \19611 );
nand \U$18943 ( \19613 , \19605 , \19612 );
not \U$18944 ( \19614 , \19613 );
nand \U$18945 ( \19615 , \18683 , \18713 );
not \U$18946 ( \19616 , \19615 );
or \U$18947 ( \19617 , \19614 , \19616 );
or \U$18948 ( \19618 , \19615 , \19613 );
nand \U$18949 ( \19619 , \19617 , \19618 );
not \U$18950 ( \19620 , \19619 );
or \U$18951 ( \19621 , \19602 , \19620 );
not \U$18952 ( \19622 , \19615 );
nand \U$18953 ( \19623 , \19622 , \19613 );
nand \U$18954 ( \19624 , \19621 , \19623 );
not \U$18955 ( \19625 , \19624 );
and \U$18956 ( \19626 , \18415 , \18976 );
not \U$18957 ( \19627 , \18415 );
and \U$18958 ( \19628 , \19627 , \18874 );
nor \U$18959 ( \19629 , \19626 , \19628 );
and \U$18960 ( \19630 , \17936 , \18639 );
not \U$18961 ( \19631 , \17936 );
and \U$18962 ( \19632 , \19631 , \18806 );
nor \U$18963 ( \19633 , \19630 , \19632 );
or \U$18964 ( \19634 , \19633 , \18810 );
and \U$18965 ( \19635 , \19629 , \19634 );
not \U$18966 ( \19636 , \19635 );
or \U$18967 ( \19637 , \19625 , \19636 );
or \U$18968 ( \19638 , \19635 , \19624 );
nand \U$18969 ( \19639 , \19637 , \19638 );
xor \U$18970 ( \19640 , \19591 , \19639 );
and \U$18971 ( \19641 , \18678 , \18374 );
and \U$18972 ( \19642 , \18677 , \18366 );
nor \U$18973 ( \19643 , \19641 , \19642 );
nand \U$18974 ( \19644 , \18796 , \17993 );
and \U$18975 ( \19645 , \19643 , \19644 );
not \U$18976 ( \19646 , \18123 );
not \U$18977 ( \19647 , \18454 );
or \U$18978 ( \19648 , \19646 , \19647 );
not \U$18979 ( \19649 , \18127 );
not \U$18980 ( \19650 , \18454 );
and \U$18981 ( \19651 , \19649 , \19650 );
and \U$18982 ( \19652 , \18580 , \18161 );
not \U$18983 ( \19653 , \18580 );
and \U$18984 ( \19654 , \19653 , \18166 );
nor \U$18985 ( \19655 , \19652 , \19654 );
nor \U$18986 ( \19656 , \19651 , \19655 );
nand \U$18987 ( \19657 , \19648 , \19656 );
and \U$18988 ( \19658 , \18190 , \17935 );
not \U$18989 ( \19659 , \18189 );
nor \U$18990 ( \19660 , \19658 , \19659 );
and \U$18991 ( \19661 , \19660 , \18194 );
nand \U$18992 ( \19662 , \19657 , \19661 );
xor \U$18993 ( \19663 , \19645 , \19662 );
not \U$18994 ( \19664 , \19663 );
xor \U$18995 ( \19665 , \19619 , \19601 );
not \U$18996 ( \19666 , \19665 );
or \U$18997 ( \19667 , \19664 , \19666 );
or \U$18998 ( \19668 , \19662 , \19645 );
nand \U$18999 ( \19669 , \19667 , \19668 );
nor \U$19000 ( \19670 , \19640 , \19669 );
or \U$19001 ( \19671 , \18197 , \18714 );
nand \U$19002 ( \19672 , \18242 , \18714 );
and \U$19003 ( \19673 , \18886 , \18832 );
not \U$19004 ( \19674 , \18886 );
and \U$19005 ( \19675 , \19674 , \18300 );
nor \U$19006 ( \19676 , \19673 , \19675 );
nand \U$19007 ( \19677 , \19671 , \19672 , \19676 );
or \U$19008 ( \19678 , \18796 , \17982 );
nand \U$19009 ( \19679 , \19678 , \17988 );
and \U$19010 ( \19680 , \19679 , \17992 );
or \U$19011 ( \19681 , \19019 , \17992 );
or \U$19012 ( \19682 , \18755 , \17983 );
nand \U$19013 ( \19683 , \19681 , \19682 );
nor \U$19014 ( \19684 , \19680 , \19683 );
nand \U$19015 ( \19685 , \19677 , \19684 );
or \U$19016 ( \19686 , \19677 , \19684 );
nand \U$19017 ( \19687 , \19685 , \19686 );
not \U$19018 ( \19688 , \19661 );
not \U$19019 ( \19689 , \19657 );
not \U$19020 ( \19690 , \19689 );
or \U$19021 ( \19691 , \19688 , \19690 );
or \U$19022 ( \19692 , \19689 , \19661 );
nand \U$19023 ( \19693 , \19691 , \19692 );
not \U$19024 ( \19694 , \19693 );
and \U$19025 ( \19695 , \19687 , \19694 );
not \U$19026 ( \19696 , \19687 );
and \U$19027 ( \19697 , \19696 , \19693 );
nor \U$19028 ( \19698 , \19695 , \19697 );
not \U$19029 ( \19699 , \19698 );
nor \U$19030 ( \19700 , \18191 , \17936 );
not \U$19031 ( \19701 , \17993 );
not \U$19032 ( \19702 , \19169 );
or \U$19033 ( \19703 , \19701 , \19702 );
and \U$19034 ( \19704 , \19608 , \18374 );
and \U$19035 ( \19705 , \18501 , \18366 );
nor \U$19036 ( \19706 , \19704 , \19705 );
nand \U$19037 ( \19707 , \19703 , \19706 );
xor \U$19038 ( \19708 , \19700 , \19707 );
not \U$19039 ( \19709 , \18415 );
not \U$19040 ( \19710 , \18123 );
or \U$19041 ( \19711 , \19709 , \19710 );
and \U$19042 ( \19712 , \19606 , \18886 );
not \U$19043 ( \19713 , \18359 );
not \U$19044 ( \19714 , \18454 );
not \U$19045 ( \19715 , \19714 );
or \U$19046 ( \19716 , \19713 , \19715 );
or \U$19047 ( \19717 , \19714 , \18161 );
nand \U$19048 ( \19718 , \19716 , \19717 );
nor \U$19049 ( \19719 , \19712 , \19718 );
nand \U$19050 ( \19720 , \19711 , \19719 );
and \U$19051 ( \19721 , \19708 , \19720 );
and \U$19052 ( \19722 , \19700 , \19707 );
or \U$19053 ( \19723 , \19721 , \19722 );
not \U$19054 ( \19724 , \19723 );
and \U$19055 ( \19725 , \19699 , \19724 );
and \U$19056 ( \19726 , \19665 , \19663 );
not \U$19057 ( \19727 , \19665 );
not \U$19058 ( \19728 , \19663 );
and \U$19059 ( \19729 , \19727 , \19728 );
or \U$19060 ( \19730 , \19726 , \19729 );
and \U$19061 ( \19731 , \19686 , \19693 );
not \U$19062 ( \19732 , \19685 );
nor \U$19063 ( \19733 , \19731 , \19732 );
and \U$19064 ( \19734 , \19730 , \19733 );
nor \U$19065 ( \19735 , \19725 , \19734 );
nand \U$19066 ( \19736 , \19698 , \19723 );
xor \U$19067 ( \19737 , \19700 , \19707 );
xor \U$19068 ( \19738 , \19737 , \19720 );
nand \U$19069 ( \19739 , \18098 , \17982 );
and \U$19070 ( \19740 , \17935 , \19739 );
not \U$19071 ( \19741 , \18098 );
nand \U$19072 ( \19742 , \19741 , \17983 );
nand \U$19073 ( \19743 , \19467 , \19742 );
nor \U$19074 ( \19744 , \19740 , \19743 );
not \U$19075 ( \19745 , \19744 );
and \U$19076 ( \19746 , \18581 , \18366 );
or \U$19077 ( \19747 , \18454 , \17992 );
or \U$19078 ( \19748 , \18580 , \18373 );
nand \U$19079 ( \19749 , \19747 , \19748 );
nor \U$19080 ( \19750 , \19746 , \19749 );
nor \U$19081 ( \19751 , \19745 , \19750 );
and \U$19082 ( \19752 , \19738 , \19751 );
not \U$19083 ( \19753 , \19750 );
not \U$19084 ( \19754 , \19744 );
and \U$19085 ( \19755 , \19753 , \19754 );
and \U$19086 ( \19756 , \19750 , \19744 );
nor \U$19087 ( \19757 , \19755 , \19756 );
nor \U$19088 ( \19758 , \19714 , \18366 );
not \U$19089 ( \19759 , \19758 );
nand \U$19090 ( \19760 , \19714 , \18373 );
nand \U$19091 ( \19761 , \19759 , \19760 , \18713 );
nand \U$19092 ( \19762 , \19761 , \18415 );
not \U$19093 ( \19763 , \19760 );
or \U$19094 ( \19764 , \19763 , \19758 );
nand \U$19095 ( \19765 , \19764 , \17992 );
and \U$19096 ( \19766 , \19036 , \18164 );
and \U$19097 ( \19767 , \18714 , \17982 );
nor \U$19098 ( \19768 , \19766 , \19767 );
nand \U$19099 ( \19769 , \19762 , \19765 , \19768 );
and \U$19100 ( \19770 , \19757 , \19769 );
nor \U$19101 ( \19771 , \19738 , \19751 );
and \U$19102 ( \19772 , \18123 , \18713 );
nor \U$19103 ( \19773 , \19757 , \19769 );
or \U$19104 ( \19774 , \18161 , \18886 );
not \U$19105 ( \19775 , \19606 );
or \U$19106 ( \19776 , \19775 , \18713 );
or \U$19107 ( \19777 , \18166 , \18887 );
nand \U$19108 ( \19778 , \19774 , \19776 , \19777 );
nor \U$19109 ( \19779 , \19772 , \19773 , \19778 );
nor \U$19110 ( \19780 , \19770 , \19771 , \19779 );
nor \U$19111 ( \19781 , \19752 , \19780 );
nand \U$19112 ( \19782 , \19736 , \19781 );
and \U$19113 ( \19783 , \19735 , \19782 );
nor \U$19114 ( \19784 , \19730 , \19733 );
nor \U$19115 ( \19785 , \19783 , \19784 );
or \U$19116 ( \19786 , \19670 , \19785 );
nand \U$19117 ( \19787 , \19640 , \19669 );
nand \U$19118 ( \19788 , \19786 , \19787 );
xor \U$19119 ( \19789 , \19547 , \19574 );
xor \U$19120 ( \19790 , \19789 , \19577 );
nand \U$19121 ( \19791 , \19639 , \19591 );
not \U$19122 ( \19792 , \19635 );
nand \U$19123 ( \19793 , \19792 , \19624 );
and \U$19124 ( \19794 , \19791 , \19793 );
nand \U$19125 ( \19795 , \19790 , \19794 );
and \U$19126 ( \19796 , \19788 , \19795 );
nor \U$19127 ( \19797 , \19790 , \19794 );
nor \U$19128 ( \19798 , \19796 , \19797 );
or \U$19129 ( \19799 , \19584 , \19798 );
not \U$19130 ( \19800 , \19580 );
nand \U$19131 ( \19801 , \19800 , \19544 );
nand \U$19132 ( \19802 , \19799 , \19801 );
and \U$19133 ( \19803 , \19539 , \19802 );
and \U$19134 ( \19804 , \19523 , \19538 );
nor \U$19135 ( \19805 , \19803 , \19804 );
not \U$19136 ( \19806 , \19524 );
and \U$19137 ( \19807 , \19537 , \19806 );
and \U$19138 ( \19808 , \19529 , \19536 );
nor \U$19139 ( \19809 , \19807 , \19808 );
xor \U$19140 ( \19810 , \19000 , \19056 );
xor \U$19141 ( \19811 , \19810 , \19059 );
not \U$19142 ( \19812 , \19811 );
and \U$19143 ( \19813 , \19809 , \19812 );
not \U$19144 ( \19814 , \19809 );
and \U$19145 ( \19815 , \19814 , \19811 );
nor \U$19146 ( \19816 , \19813 , \19815 );
or \U$19147 ( \19817 , \19805 , \19816 );
not \U$19148 ( \19818 , \19809 );
nand \U$19149 ( \19819 , \19818 , \19812 );
nand \U$19150 ( \19820 , \19817 , \19819 );
and \U$19151 ( \19821 , \18918 , \18995 );
and \U$19152 ( \19822 , \18998 , \19062 );
nor \U$19153 ( \19823 , \19821 , \19822 );
nand \U$19154 ( \19824 , \19820 , \19823 );
not \U$19155 ( \19825 , \19824 );
or \U$19156 ( \19826 , \19419 , \19825 );
not \U$19157 ( \19827 , \19415 );
not \U$19158 ( \19828 , \19827 );
not \U$19159 ( \19829 , \19413 );
not \U$19160 ( \19830 , \19829 );
or \U$19161 ( \19831 , \19828 , \19830 );
nand \U$19162 ( \19832 , \19247 , \19253 );
nand \U$19163 ( \19833 , \19831 , \19832 );
buf \U$19164 ( \19834 , \19416 );
and \U$19165 ( \19835 , \19833 , \19834 );
xor \U$19166 ( \19836 , \19380 , \19405 );
and \U$19167 ( \19837 , \19836 , \19411 );
and \U$19168 ( \19838 , \19380 , \19405 );
or \U$19169 ( \19839 , \19837 , \19838 );
not \U$19170 ( \19840 , \19323 );
and \U$19171 ( \19841 , \19279 , \19840 );
not \U$19172 ( \19842 , \18366 );
not \U$19173 ( \19843 , \17886 );
or \U$19174 ( \19844 , \19842 , \19843 );
and \U$19175 ( \19845 , \19318 , \17993 );
not \U$19176 ( \19846 , \17886 );
and \U$19177 ( \19847 , \19846 , \18374 );
nor \U$19178 ( \19848 , \19845 , \19847 );
nand \U$19179 ( \19849 , \19844 , \19848 );
buf \U$19180 ( \19850 , \17970 );
not \U$19181 ( \19851 , \19850 );
not \U$19182 ( \19852 , \18123 );
or \U$19183 ( \19853 , \19851 , \19852 );
not \U$19184 ( \19854 , \19850 );
and \U$19185 ( \19855 , \19606 , \19854 );
and \U$19186 ( \19856 , \19137 , \18161 );
not \U$19187 ( \19857 , \19137 );
and \U$19188 ( \19858 , \19857 , \18166 );
nor \U$19189 ( \19859 , \19856 , \19858 );
nor \U$19190 ( \19860 , \19855 , \19859 );
nand \U$19191 ( \19861 , \19853 , \19860 );
xor \U$19192 ( \19862 , \19849 , \19861 );
xor \U$19193 ( \19863 , \19841 , \19862 );
not \U$19194 ( \19864 , \18777 );
not \U$19195 ( \19865 , \19864 );
not \U$19196 ( \19866 , \18825 );
or \U$19197 ( \19867 , \19865 , \19866 );
and \U$19198 ( \19868 , \18196 , \18777 );
and \U$19199 ( \19869 , \19273 , \19027 );
not \U$19200 ( \19870 , \19273 );
and \U$19201 ( \19871 , \19870 , \19024 );
nor \U$19202 ( \19872 , \19869 , \19871 );
nor \U$19203 ( \19873 , \19868 , \19872 );
nand \U$19204 ( \19874 , \19867 , \19873 );
not \U$19205 ( \19875 , \19874 );
xor \U$19206 ( \19876 , \19863 , \19875 );
not \U$19207 ( \19877 , \18244 );
not \U$19208 ( \19878 , \19005 );
or \U$19209 ( \19879 , \19877 , \19878 );
not \U$19210 ( \19880 , \18757 );
not \U$19211 ( \19881 , \18244 );
and \U$19212 ( \19882 , \19880 , \19881 );
nand \U$19213 ( \19883 , \19186 , \18926 );
and \U$19214 ( \19884 , \19883 , \19389 );
nor \U$19215 ( \19885 , \19882 , \19884 );
nand \U$19216 ( \19886 , \19879 , \19885 );
not \U$19217 ( \19887 , \18796 );
not \U$19218 ( \19888 , \18418 );
or \U$19219 ( \19889 , \19887 , \19888 );
and \U$19220 ( \19890 , \18677 , \18458 );
not \U$19221 ( \19891 , \18677 );
and \U$19222 ( \19892 , \19891 , \17892 );
nor \U$19223 ( \19893 , \19890 , \19892 );
nand \U$19224 ( \19894 , \19889 , \19893 );
and \U$19225 ( \19895 , \18465 , \18755 );
nor \U$19226 ( \19896 , \19894 , \19895 );
not \U$19227 ( \19897 , \19896 );
buf \U$19228 ( \19898 , \18820 );
not \U$19229 ( \19899 , \19898 );
not \U$19230 ( \19900 , \19899 );
not \U$19231 ( \19901 , \18868 );
or \U$19232 ( \19902 , \19900 , \19901 );
and \U$19233 ( \19903 , \18871 , \18820 );
and \U$19234 ( \19904 , \19261 , \18689 );
not \U$19235 ( \19905 , \19261 );
and \U$19236 ( \19906 , \19905 , \18684 );
nor \U$19237 ( \19907 , \19904 , \19906 );
nor \U$19238 ( \19908 , \19903 , \19907 );
nand \U$19239 ( \19909 , \19902 , \19908 );
not \U$19240 ( \19910 , \19909 );
or \U$19241 ( \19911 , \19897 , \19910 );
or \U$19242 ( \19912 , \19909 , \19896 );
nand \U$19243 ( \19913 , \19911 , \19912 );
xor \U$19244 ( \19914 , \19886 , \19913 );
xor \U$19245 ( \19915 , \19876 , \19914 );
not \U$19246 ( \19916 , \19343 );
not \U$19247 ( \19917 , \19366 );
or \U$19248 ( \19918 , \19916 , \19917 );
nand \U$19249 ( \19919 , \19362 , \19352 );
nand \U$19250 ( \19920 , \19918 , \19919 );
not \U$19251 ( \19921 , \19920 );
xnor \U$19252 ( \19922 , \19915 , \19921 );
xnor \U$19253 ( \19923 , \19839 , \19922 );
not \U$19254 ( \19924 , \19332 );
xor \U$19255 ( \19925 , \19331 , \19343 );
xnor \U$19256 ( \19926 , \19925 , \19366 );
not \U$19257 ( \19927 , \19926 );
or \U$19258 ( \19928 , \19924 , \19927 );
not \U$19259 ( \19929 , \19331 );
nand \U$19260 ( \19930 , \19929 , \19371 );
nand \U$19261 ( \19931 , \19928 , \19930 );
not \U$19262 ( \19932 , \18581 );
not \U$19263 ( \19933 , \17645 );
or \U$19264 ( \19934 , \19932 , \19933 );
and \U$19265 ( \19935 , \17650 , \18970 );
or \U$19266 ( \19936 , \17655 , \18761 );
nand \U$19267 ( \19937 , \17705 , \18761 );
nand \U$19268 ( \19938 , \19936 , \19937 );
nor \U$19269 ( \19939 , \19935 , \19938 );
nand \U$19270 ( \19940 , \19934 , \19939 );
not \U$19271 ( \19941 , \19940 );
not \U$19272 ( \19942 , \17747 );
not \U$19273 ( \19943 , \18611 );
and \U$19274 ( \19944 , \19942 , \19943 );
not \U$19275 ( \19945 , \19327 );
and \U$19276 ( \19946 , \19268 , \19945 );
nor \U$19277 ( \19947 , \19944 , \19946 );
not \U$19278 ( \19948 , \19947 );
and \U$19279 ( \19949 , \19941 , \19948 );
and \U$19280 ( \19950 , \19940 , \19947 );
nor \U$19281 ( \19951 , \19949 , \19950 );
not \U$19282 ( \19952 , \19951 );
not \U$19283 ( \19953 , \19952 );
not \U$19284 ( \19954 , \19401 );
nand \U$19285 ( \19955 , \19954 , \19393 );
not \U$19286 ( \19956 , \19955 );
and \U$19287 ( \19957 , \19953 , \19956 );
and \U$19288 ( \19958 , \19952 , \19955 );
nor \U$19289 ( \19959 , \19957 , \19958 );
and \U$19290 ( \19960 , \19931 , \19959 );
not \U$19291 ( \19961 , \19931 );
not \U$19292 ( \19962 , \19959 );
and \U$19293 ( \19963 , \19961 , \19962 );
nor \U$19294 ( \19964 , \19960 , \19963 );
and \U$19295 ( \19965 , \19923 , \19964 );
not \U$19296 ( \19966 , \19923 );
not \U$19297 ( \19967 , \19964 );
and \U$19298 ( \19968 , \19966 , \19967 );
or \U$19299 ( \19969 , \19965 , \19968 );
xor \U$19300 ( \19970 , \19260 , \19372 );
and \U$19301 ( \19971 , \19970 , \19412 );
and \U$19302 ( \19972 , \19260 , \19372 );
or \U$19303 ( \19973 , \19971 , \19972 );
nor \U$19304 ( \19974 , \19969 , \19973 );
nor \U$19305 ( \19975 , \19835 , \19974 );
nand \U$19306 ( \19976 , \19826 , \19975 );
not \U$19307 ( \19977 , \19947 );
nand \U$19308 ( \19978 , \19977 , \19940 );
not \U$19309 ( \19979 , \18502 );
not \U$19310 ( \19980 , \17645 );
or \U$19311 ( \19981 , \19979 , \19980 );
and \U$19312 ( \19982 , \17650 , \18761 );
or \U$19313 ( \19983 , \18796 , \17655 );
nand \U$19314 ( \19984 , \17705 , \18796 );
nand \U$19315 ( \19985 , \19983 , \19984 );
nor \U$19316 ( \19986 , \19982 , \19985 );
nand \U$19317 ( \19987 , \19981 , \19986 );
not \U$19318 ( \19988 , \19862 );
xor \U$19319 ( \19989 , \19841 , \19874 );
not \U$19320 ( \19990 , \19989 );
or \U$19321 ( \19991 , \19988 , \19990 );
and \U$19322 ( \19992 , \19874 , \19841 );
and \U$19323 ( \19993 , \17746 , \18581 );
nor \U$19324 ( \19994 , \19992 , \19993 );
nand \U$19325 ( \19995 , \19991 , \19994 );
nor \U$19326 ( \19996 , \19987 , \19995 );
not \U$19327 ( \19997 , \19996 );
nand \U$19328 ( \19998 , \19987 , \19995 );
nand \U$19329 ( \19999 , \19997 , \19998 );
xor \U$19330 ( \20000 , \19978 , \19999 );
not \U$19331 ( \20001 , \19921 );
not \U$19332 ( \20002 , \19876 );
and \U$19333 ( \20003 , \20001 , \20002 );
not \U$19334 ( \20004 , \19876 );
not \U$19335 ( \20005 , \19920 );
or \U$19336 ( \20006 , \20004 , \20005 );
or \U$19337 ( \20007 , \19920 , \19876 );
nand \U$19338 ( \20008 , \20006 , \20007 );
and \U$19339 ( \20009 , \20008 , \19914 );
nor \U$19340 ( \20010 , \20003 , \20009 );
xor \U$19341 ( \20011 , \20000 , \20010 );
not \U$19342 ( \20012 , \20011 );
and \U$19343 ( \20013 , \19849 , \19861 );
and \U$19344 ( \20014 , \19846 , \17993 );
and \U$19345 ( \20015 , \17789 , \18374 );
nor \U$19346 ( \20016 , \20014 , \20015 );
not \U$19347 ( \20017 , \17789 );
nand \U$19348 ( \20018 , \20017 , \18366 );
and \U$19349 ( \20019 , \20016 , \20018 );
not \U$19350 ( \20020 , \20019 );
not \U$19351 ( \20021 , \19138 );
not \U$19352 ( \20022 , \20021 );
not \U$19353 ( \20023 , \18123 );
or \U$19354 ( \20024 , \20022 , \20023 );
and \U$19355 ( \20025 , \19321 , \18160 );
not \U$19356 ( \20026 , \19321 );
buf \U$19357 ( \20027 , \18359 );
and \U$19358 ( \20028 , \20026 , \20027 );
nor \U$19359 ( \20029 , \20025 , \20028 );
nand \U$19360 ( \20030 , \18128 , \19138 );
and \U$19361 ( \20031 , \20029 , \20030 );
nand \U$19362 ( \20032 , \20024 , \20031 );
not \U$19363 ( \20033 , \20032 );
or \U$19364 ( \20034 , \20020 , \20033 );
or \U$19365 ( \20035 , \20032 , \20019 );
nand \U$19366 ( \20036 , \20034 , \20035 );
xor \U$19367 ( \20037 , \20013 , \20036 );
not \U$19368 ( \20038 , \19273 );
not \U$19369 ( \20039 , \18825 );
or \U$19370 ( \20040 , \20038 , \20039 );
not \U$19371 ( \20041 , \19273 );
and \U$19372 ( \20042 , \18196 , \20041 );
buf \U$19373 ( \20043 , \19850 );
and \U$19374 ( \20044 , \20043 , \19024 );
not \U$19375 ( \20045 , \20043 );
and \U$19376 ( \20046 , \20045 , \19027 );
nor \U$19377 ( \20047 , \20044 , \20046 );
nor \U$19378 ( \20048 , \20042 , \20047 );
nand \U$19379 ( \20049 , \20040 , \20048 );
xor \U$19380 ( \20050 , \20037 , \20049 );
not \U$19381 ( \20051 , \20050 );
not \U$19382 ( \20052 , \19886 );
not \U$19383 ( \20053 , \19913 );
or \U$19384 ( \20054 , \20052 , \20053 );
not \U$19385 ( \20055 , \19896 );
nand \U$19386 ( \20056 , \20055 , \19909 );
nand \U$19387 ( \20057 , \20054 , \20056 );
not \U$19388 ( \20058 , \20057 );
not \U$19389 ( \20059 , \20058 );
or \U$19390 ( \20060 , \20051 , \20059 );
not \U$19391 ( \20061 , \20050 );
nand \U$19392 ( \20062 , \20061 , \20057 );
nand \U$19393 ( \20063 , \20060 , \20062 );
not \U$19394 ( \20064 , \18680 );
not \U$19395 ( \20065 , \17844 );
or \U$19396 ( \20066 , \20064 , \20065 );
and \U$19397 ( \20067 , \18679 , \17848 );
and \U$19398 ( \20068 , \18686 , \18613 );
not \U$19399 ( \20069 , \18686 );
not \U$19400 ( \20070 , \18461 );
and \U$19401 ( \20071 , \20069 , \20070 );
nor \U$19402 ( \20072 , \20068 , \20071 );
nor \U$19403 ( \20073 , \20067 , \20072 );
nand \U$19404 ( \20074 , \20066 , \20073 );
not \U$19405 ( \20075 , \19899 );
not \U$19406 ( \20076 , \19005 );
or \U$19407 ( \20077 , \20075 , \20076 );
and \U$19408 ( \20078 , \18538 , \19898 );
and \U$19409 ( \20079 , \18243 , \18583 );
not \U$19410 ( \20080 , \18243 );
and \U$19411 ( \20081 , \20080 , \18590 );
or \U$19412 ( \20082 , \20079 , \20081 );
nor \U$19413 ( \20083 , \20078 , \20082 );
nand \U$19414 ( \20084 , \20077 , \20083 );
xor \U$19415 ( \20085 , \20074 , \20084 );
not \U$19416 ( \20086 , \19261 );
not \U$19417 ( \20087 , \20086 );
not \U$19418 ( \20088 , \18695 );
or \U$19419 ( \20089 , \20087 , \20088 );
and \U$19420 ( \20090 , \18641 , \19261 );
not \U$19421 ( \20091 , \18976 );
or \U$19422 ( \20092 , \20091 , \19864 );
or \U$19423 ( \20093 , \18685 , \18777 );
nand \U$19424 ( \20094 , \20092 , \20093 );
nor \U$19425 ( \20095 , \20090 , \20094 );
nand \U$19426 ( \20096 , \20089 , \20095 );
xor \U$19427 ( \20097 , \20085 , \20096 );
not \U$19428 ( \20098 , \20097 );
and \U$19429 ( \20099 , \20063 , \20098 );
not \U$19430 ( \20100 , \20063 );
and \U$19431 ( \20101 , \20100 , \20097 );
nor \U$19432 ( \20102 , \20099 , \20101 );
not \U$19433 ( \20103 , \20102 );
nand \U$19434 ( \20104 , \19951 , \19955 );
not \U$19435 ( \20105 , \20104 );
not \U$19436 ( \20106 , \19931 );
or \U$19437 ( \20107 , \20105 , \20106 );
not \U$19438 ( \20108 , \19955 );
nand \U$19439 ( \20109 , \20108 , \19952 );
nand \U$19440 ( \20110 , \20107 , \20109 );
not \U$19441 ( \20111 , \20110 );
or \U$19442 ( \20112 , \20103 , \20111 );
or \U$19443 ( \20113 , \20110 , \20102 );
nand \U$19444 ( \20114 , \20112 , \20113 );
not \U$19445 ( \20115 , \20114 );
or \U$19446 ( \20116 , \20012 , \20115 );
or \U$19447 ( \20117 , \20114 , \20011 );
nand \U$19448 ( \20118 , \20116 , \20117 );
not \U$19449 ( \20119 , \20118 );
not \U$19450 ( \20120 , \19967 );
not \U$19451 ( \20121 , \19923 );
or \U$19452 ( \20122 , \20120 , \20121 );
not \U$19453 ( \20123 , \19922 );
nand \U$19454 ( \20124 , \20123 , \19839 );
nand \U$19455 ( \20125 , \20122 , \20124 );
not \U$19456 ( \20126 , \20125 );
nand \U$19457 ( \20127 , \20119 , \20126 );
not \U$19458 ( \20128 , \20127 );
nor \U$19459 ( \20129 , \19976 , \20128 );
or \U$19460 ( \20130 , \18594 , \20043 );
nand \U$19461 ( \20131 , \18538 , \20043 );
buf \U$19462 ( \20132 , \18365 );
and \U$19463 ( \20133 , \20132 , \18927 );
not \U$19464 ( \20134 , \20132 );
and \U$19465 ( \20135 , \20134 , \19187 );
nor \U$19466 ( \20136 , \20133 , \20135 );
nand \U$19467 ( \20137 , \20130 , \20131 , \20136 );
not \U$19468 ( \20138 , \20137 );
not \U$19469 ( \20139 , \17887 );
not \U$19470 ( \20140 , \18196 );
or \U$19471 ( \20141 , \20139 , \20140 );
and \U$19472 ( \20142 , \17790 , \18832 );
not \U$19473 ( \20143 , \17790 );
and \U$19474 ( \20144 , \20143 , \18300 );
nor \U$19475 ( \20145 , \20142 , \20144 );
nand \U$19476 ( \20146 , \20141 , \20145 );
nor \U$19477 ( \20147 , \18824 , \17887 );
nor \U$19478 ( \20148 , \20146 , \20147 );
nor \U$19479 ( \20149 , \20148 , \17983 );
not \U$19480 ( \20150 , \20149 );
nand \U$19481 ( \20151 , \20148 , \17983 );
nand \U$19482 ( \20152 , \20150 , \20151 );
not \U$19483 ( \20153 , \20152 );
not \U$19484 ( \20154 , \20153 );
not \U$19485 ( \20155 , \17843 );
not \U$19486 ( \20156 , \20086 );
and \U$19487 ( \20157 , \20155 , \20156 );
not \U$19488 ( \20158 , \20086 );
not \U$19489 ( \20159 , \17848 );
or \U$19490 ( \20160 , \20158 , \20159 );
and \U$19491 ( \20161 , \18777 , \18458 );
not \U$19492 ( \20162 , \18777 );
and \U$19493 ( \20163 , \20162 , \18461 );
nor \U$19494 ( \20164 , \20161 , \20163 );
nand \U$19495 ( \20165 , \20160 , \20164 );
nor \U$19496 ( \20166 , \20157 , \20165 );
not \U$19497 ( \20167 , \20166 );
not \U$19498 ( \20168 , \20167 );
or \U$19499 ( \20169 , \20154 , \20168 );
nand \U$19500 ( \20170 , \20166 , \20152 );
nand \U$19501 ( \20171 , \20169 , \20170 );
not \U$19502 ( \20172 , \20171 );
or \U$19503 ( \20173 , \20138 , \20172 );
nand \U$19504 ( \20174 , \20167 , \20152 );
nand \U$19505 ( \20175 , \20173 , \20174 );
not \U$19506 ( \20176 , \17791 );
not \U$19507 ( \20177 , \20176 );
not \U$19508 ( \20178 , \20177 );
not \U$19509 ( \20179 , \18242 );
or \U$19510 ( \20180 , \20178 , \20179 );
and \U$19511 ( \20181 , \18196 , \20176 );
not \U$19512 ( \20182 , \18295 );
and \U$19513 ( \20183 , \17533 , \20182 );
not \U$19514 ( \20184 , \17533 );
and \U$19515 ( \20185 , \20184 , \19024 );
nor \U$19516 ( \20186 , \20183 , \20185 );
nor \U$19517 ( \20187 , \20181 , \20186 );
nand \U$19518 ( \20188 , \20180 , \20187 );
not \U$19519 ( \20189 , \20151 );
xor \U$19520 ( \20190 , \20188 , \20189 );
not \U$19521 ( \20191 , \17702 );
not \U$19522 ( \20192 , \18123 );
or \U$19523 ( \20193 , \20191 , \20192 );
and \U$19524 ( \20194 , \19606 , \17706 );
nor \U$19525 ( \20195 , \20194 , \20027 );
nand \U$19526 ( \20196 , \20193 , \20195 );
not \U$19527 ( \20197 , \20196 );
xor \U$19528 ( \20198 , \20190 , \20197 );
and \U$19529 ( \20199 , \20175 , \20198 );
not \U$19530 ( \20200 , \20175 );
not \U$19531 ( \20201 , \20198 );
and \U$19532 ( \20202 , \20200 , \20201 );
or \U$19533 ( \20203 , \20199 , \20202 );
not \U$19534 ( \20204 , \20021 );
not \U$19535 ( \20205 , \20204 );
or \U$19536 ( \20206 , \18767 , \20205 );
nand \U$19537 ( \20207 , \18758 , \20205 );
not \U$19538 ( \20208 , \18763 );
not \U$19539 ( \20209 , \20043 );
not \U$19540 ( \20210 , \20209 );
and \U$19541 ( \20211 , \20208 , \20210 );
and \U$19542 ( \20212 , \18931 , \20209 );
nor \U$19543 ( \20213 , \20211 , \20212 );
nand \U$19544 ( \20214 , \20206 , \20207 , \20213 );
and \U$19545 ( \20215 , \17849 , \19864 );
not \U$19546 ( \20216 , \18888 );
not \U$19547 ( \20217 , \20041 );
or \U$19548 ( \20218 , \20216 , \20217 );
or \U$19549 ( \20219 , \20070 , \20041 );
nand \U$19550 ( \20220 , \20218 , \20219 );
nor \U$19551 ( \20221 , \20215 , \20220 );
not \U$19552 ( \20222 , \18466 );
nand \U$19553 ( \20223 , \20222 , \18777 );
nand \U$19554 ( \20224 , \20221 , \20223 );
buf \U$19555 ( \20225 , \19318 );
not \U$19556 ( \20226 , \20225 );
and \U$19557 ( \20227 , \18641 , \20226 );
or \U$19558 ( \20228 , \18685 , \17887 );
nand \U$19559 ( \20229 , \18690 , \17887 );
nand \U$19560 ( \20230 , \20228 , \20229 );
nor \U$19561 ( \20231 , \20227 , \20230 );
not \U$19562 ( \20232 , \20226 );
nand \U$19563 ( \20233 , \18695 , \20232 );
nand \U$19564 ( \20234 , \20231 , \20233 );
xor \U$19565 ( \20235 , \20224 , \20234 );
xor \U$19566 ( \20236 , \20214 , \20235 );
not \U$19567 ( \20237 , \20236 );
and \U$19568 ( \20238 , \20203 , \20237 );
not \U$19569 ( \20239 , \20203 );
and \U$19570 ( \20240 , \20239 , \20236 );
nor \U$19571 ( \20241 , \20238 , \20240 );
not \U$19572 ( \20242 , \20241 );
not \U$19573 ( \20243 , \17993 );
not \U$19574 ( \20244 , \17532 );
or \U$19575 ( \20245 , \20243 , \20244 );
and \U$19576 ( \20246 , \17700 , \18374 );
not \U$19577 ( \20247 , \17700 );
and \U$19578 ( \20248 , \20247 , \18366 );
nor \U$19579 ( \20249 , \20246 , \20248 );
nand \U$19580 ( \20250 , \20245 , \20249 );
not \U$19581 ( \20251 , \17887 );
not \U$19582 ( \20252 , \18123 );
or \U$19583 ( \20253 , \20251 , \20252 );
and \U$19584 ( \20254 , \19606 , \19846 );
and \U$19585 ( \20255 , \17789 , \18166 );
not \U$19586 ( \20256 , \17789 );
and \U$19587 ( \20257 , \20256 , \18161 );
nor \U$19588 ( \20258 , \20255 , \20257 );
nor \U$19589 ( \20259 , \20254 , \20258 );
nand \U$19590 ( \20260 , \20253 , \20259 );
xor \U$19591 ( \20261 , \20250 , \20260 );
not \U$19592 ( \20262 , \20261 );
not \U$19593 ( \20263 , \20225 );
not \U$19594 ( \20264 , \18128 );
or \U$19595 ( \20265 , \20263 , \20264 );
and \U$19596 ( \20266 , \17886 , \18160 );
not \U$19597 ( \20267 , \17886 );
and \U$19598 ( \20268 , \20267 , \20027 );
nor \U$19599 ( \20269 , \20266 , \20268 );
nand \U$19600 ( \20270 , \20265 , \20269 );
and \U$19601 ( \20271 , \18123 , \19321 );
nor \U$19602 ( \20272 , \20270 , \20271 );
not \U$19603 ( \20273 , \17532 );
nand \U$19604 ( \20274 , \20273 , \18366 );
nand \U$19605 ( \20275 , \17532 , \18374 );
nand \U$19606 ( \20276 , \17789 , \17993 );
and \U$19607 ( \20277 , \20274 , \20275 , \20276 );
nor \U$19608 ( \20278 , \20272 , \20277 );
not \U$19609 ( \20279 , \20278 );
not \U$19610 ( \20280 , \20021 );
not \U$19611 ( \20281 , \18196 );
or \U$19612 ( \20282 , \20280 , \20281 );
and \U$19613 ( \20283 , \20226 , \18300 );
not \U$19614 ( \20284 , \20226 );
and \U$19615 ( \20285 , \20284 , \18832 );
nor \U$19616 ( \20286 , \20283 , \20285 );
nand \U$19617 ( \20287 , \20282 , \20286 );
nor \U$19618 ( \20288 , \18824 , \20021 );
nor \U$19619 ( \20289 , \20287 , \20288 );
not \U$19620 ( \20290 , \20289 );
or \U$19621 ( \20291 , \20279 , \20290 );
or \U$19622 ( \20292 , \20289 , \20278 );
nand \U$19623 ( \20293 , \20291 , \20292 );
not \U$19624 ( \20294 , \20293 );
or \U$19625 ( \20295 , \20262 , \20294 );
not \U$19626 ( \20296 , \20289 );
and \U$19627 ( \20297 , \20296 , \20278 );
and \U$19628 ( \20298 , \17746 , \18680 );
nor \U$19629 ( \20299 , \20297 , \20298 );
nand \U$19630 ( \20300 , \20295 , \20299 );
and \U$19631 ( \20301 , \17650 , \19077 );
nand \U$19632 ( \20302 , \17653 , \17654 );
or \U$19633 ( \20303 , \20302 , \18244 );
nand \U$19634 ( \20304 , \17705 , \18244 );
nand \U$19635 ( \20305 , \20303 , \20304 );
nor \U$19636 ( \20306 , \20301 , \20305 );
not \U$19637 ( \20307 , \19077 );
nand \U$19638 ( \20308 , \20307 , \17645 );
nand \U$19639 ( \20309 , \20306 , \20308 );
and \U$19640 ( \20310 , \20300 , \20309 );
and \U$19641 ( \20311 , \17701 , \17993 );
nor \U$19642 ( \20312 , \20311 , \17982 );
not \U$19643 ( \20313 , \17790 );
not \U$19644 ( \20314 , \20313 );
not \U$19645 ( \20315 , \18123 );
or \U$19646 ( \20316 , \20314 , \20315 );
not \U$19647 ( \20317 , \20017 );
and \U$19648 ( \20318 , \19606 , \20317 );
and \U$19649 ( \20319 , \17532 , \18166 );
not \U$19650 ( \20320 , \17532 );
and \U$19651 ( \20321 , \20320 , \18161 );
nor \U$19652 ( \20322 , \20319 , \20321 );
nor \U$19653 ( \20323 , \20318 , \20322 );
nand \U$19654 ( \20324 , \20316 , \20323 );
xor \U$19655 ( \20325 , \20312 , \20324 );
not \U$19656 ( \20326 , \20325 );
and \U$19657 ( \20327 , \20250 , \20260 );
not \U$19658 ( \20328 , \20226 );
not \U$19659 ( \20329 , \18196 );
or \U$19660 ( \20330 , \20328 , \20329 );
not \U$19661 ( \20331 , \17887 );
and \U$19662 ( \20332 , \20331 , \18832 );
not \U$19663 ( \20333 , \20331 );
and \U$19664 ( \20334 , \20333 , \18300 );
nor \U$19665 ( \20335 , \20332 , \20334 );
nand \U$19666 ( \20336 , \20330 , \20335 );
nor \U$19667 ( \20337 , \20226 , \18824 );
nor \U$19668 ( \20338 , \20336 , \20337 );
xnor \U$19669 ( \20339 , \20327 , \20338 );
not \U$19670 ( \20340 , \20339 );
or \U$19671 ( \20341 , \20326 , \20340 );
not \U$19672 ( \20342 , \17747 );
not \U$19673 ( \20343 , \19077 );
and \U$19674 ( \20344 , \20342 , \20343 );
not \U$19675 ( \20345 , \20338 );
and \U$19676 ( \20346 , \20345 , \20327 );
nor \U$19677 ( \20347 , \20344 , \20346 );
nand \U$19678 ( \20348 , \20341 , \20347 );
not \U$19679 ( \20349 , \19073 );
not \U$19680 ( \20350 , \17645 );
or \U$19681 ( \20351 , \20349 , \20350 );
and \U$19682 ( \20352 , \17650 , \18244 );
not \U$19683 ( \20353 , \18820 );
or \U$19684 ( \20354 , \20302 , \20353 );
not \U$19685 ( \20355 , \17704 );
nand \U$19686 ( \20356 , \20355 , \20353 );
nand \U$19687 ( \20357 , \20354 , \20356 );
nor \U$19688 ( \20358 , \20352 , \20357 );
nand \U$19689 ( \20359 , \20351 , \20358 );
xor \U$19690 ( \20360 , \20348 , \20359 );
xor \U$19691 ( \20361 , \20310 , \20360 );
not \U$19692 ( \20362 , \20361 );
not \U$19693 ( \20363 , \18583 );
not \U$19694 ( \20364 , \19261 );
or \U$19695 ( \20365 , \20363 , \20364 );
or \U$19696 ( \20366 , \18930 , \19261 );
nand \U$19697 ( \20367 , \20365 , \20366 );
not \U$19698 ( \20368 , \20367 );
not \U$19699 ( \20369 , \19864 );
nand \U$19700 ( \20370 , \20369 , \19008 );
nand \U$19701 ( \20371 , \19005 , \19864 );
nand \U$19702 ( \20372 , \20368 , \20370 , \20371 );
not \U$19703 ( \20373 , \20372 );
not \U$19704 ( \20374 , \19073 );
not \U$19705 ( \20375 , \20222 );
or \U$19706 ( \20376 , \20374 , \20375 );
and \U$19707 ( \20377 , \17849 , \18244 );
not \U$19708 ( \20378 , \18888 );
not \U$19709 ( \20379 , \19898 );
or \U$19710 ( \20380 , \20378 , \20379 );
or \U$19711 ( \20381 , \20070 , \18820 );
nand \U$19712 ( \20382 , \20380 , \20381 );
nor \U$19713 ( \20383 , \20377 , \20382 );
nand \U$19714 ( \20384 , \20376 , \20383 );
not \U$19715 ( \20385 , \19273 );
not \U$19716 ( \20386 , \18695 );
or \U$19717 ( \20387 , \20385 , \20386 );
and \U$19718 ( \20388 , \18641 , \20132 );
and \U$19719 ( \20389 , \20043 , \19497 );
not \U$19720 ( \20390 , \20043 );
and \U$19721 ( \20391 , \20390 , \18685 );
nor \U$19722 ( \20392 , \20389 , \20391 );
nor \U$19723 ( \20393 , \20388 , \20392 );
nand \U$19724 ( \20394 , \20387 , \20393 );
xor \U$19725 ( \20395 , \20384 , \20394 );
not \U$19726 ( \20396 , \20395 );
or \U$19727 ( \20397 , \20373 , \20396 );
nand \U$19728 ( \20398 , \20394 , \20384 );
nand \U$19729 ( \20399 , \20397 , \20398 );
not \U$19730 ( \20400 , \20399 );
xor \U$19731 ( \20401 , \20327 , \20325 );
xnor \U$19732 ( \20402 , \20401 , \20345 );
not \U$19733 ( \20403 , \17842 );
not \U$19734 ( \20404 , \20353 );
and \U$19735 ( \20405 , \20403 , \20404 );
not \U$19736 ( \20406 , \20353 );
not \U$19737 ( \20407 , \18418 );
or \U$19738 ( \20408 , \20406 , \20407 );
and \U$19739 ( \20409 , \19261 , \18458 );
not \U$19740 ( \20410 , \19261 );
and \U$19741 ( \20411 , \20410 , \17890 );
nor \U$19742 ( \20412 , \20409 , \20411 );
nand \U$19743 ( \20413 , \20408 , \20412 );
nor \U$19744 ( \20414 , \20405 , \20413 );
not \U$19745 ( \20415 , \20132 );
not \U$19746 ( \20416 , \20415 );
not \U$19747 ( \20417 , \19005 );
or \U$19748 ( \20418 , \20416 , \20417 );
not \U$19749 ( \20419 , \18537 );
not \U$19750 ( \20420 , \19273 );
and \U$19751 ( \20421 , \20419 , \20420 );
and \U$19752 ( \20422 , \18777 , \18582 );
not \U$19753 ( \20423 , \18777 );
and \U$19754 ( \20424 , \20423 , \18589 );
nor \U$19755 ( \20425 , \20422 , \20424 );
nor \U$19756 ( \20426 , \20421 , \20425 );
nand \U$19757 ( \20427 , \20418 , \20426 );
xor \U$19758 ( \20428 , \20414 , \20427 );
and \U$19759 ( \20429 , \18641 , \20043 );
not \U$19760 ( \20430 , \18690 );
not \U$19761 ( \20431 , \20205 );
or \U$19762 ( \20432 , \20430 , \20431 );
or \U$19763 ( \20433 , \18685 , \20021 );
nand \U$19764 ( \20434 , \20432 , \20433 );
nor \U$19765 ( \20435 , \20429 , \20434 );
nand \U$19766 ( \20436 , \18695 , \20209 );
nand \U$19767 ( \20437 , \20435 , \20436 );
xnor \U$19768 ( \20438 , \20428 , \20437 );
xnor \U$19769 ( \20439 , \20402 , \20438 );
not \U$19770 ( \20440 , \20439 );
or \U$19771 ( \20441 , \20400 , \20440 );
not \U$19772 ( \20442 , \20402 );
nand \U$19773 ( \20443 , \20442 , \20438 );
nand \U$19774 ( \20444 , \20441 , \20443 );
not \U$19775 ( \20445 , \20444 );
or \U$19776 ( \20446 , \20362 , \20445 );
nand \U$19777 ( \20447 , \20310 , \20360 );
nand \U$19778 ( \20448 , \20446 , \20447 );
not \U$19779 ( \20449 , \20448 );
or \U$19780 ( \20450 , \20242 , \20449 );
or \U$19781 ( \20451 , \20448 , \20241 );
nand \U$19782 ( \20452 , \20450 , \20451 );
nand \U$19783 ( \20453 , \20359 , \20348 );
and \U$19784 ( \20454 , \17650 , \20353 );
not \U$19785 ( \20455 , \20086 );
not \U$19786 ( \20456 , \17812 );
or \U$19787 ( \20457 , \20455 , \20456 );
or \U$19788 ( \20458 , \17812 , \20086 );
nand \U$19789 ( \20459 , \20457 , \20458 );
not \U$19790 ( \20460 , \20459 );
nor \U$19791 ( \20461 , \20460 , \17809 );
nor \U$19792 ( \20462 , \20454 , \20461 );
nand \U$19793 ( \20463 , \17645 , \18820 );
nand \U$19794 ( \20464 , \20462 , \20463 );
nand \U$19795 ( \20465 , \20324 , \20312 );
and \U$19796 ( \20466 , \18123 , \17534 );
or \U$19797 ( \20467 , \19775 , \20273 );
and \U$19798 ( \20468 , \17700 , \20027 );
not \U$19799 ( \20469 , \17700 );
and \U$19800 ( \20470 , \20469 , \18160 );
nor \U$19801 ( \20471 , \20468 , \20470 );
nand \U$19802 ( \20472 , \20467 , \20471 );
nor \U$19803 ( \20473 , \20466 , \20472 );
nand \U$19804 ( \20474 , \20465 , \20473 );
not \U$19805 ( \20475 , \20474 );
not \U$19806 ( \20476 , \20204 );
not \U$19807 ( \20477 , \18695 );
or \U$19808 ( \20478 , \20476 , \20477 );
and \U$19809 ( \20479 , \18641 , \20205 );
or \U$19810 ( \20480 , \18685 , \20226 );
nand \U$19811 ( \20481 , \18690 , \20226 );
nand \U$19812 ( \20482 , \20480 , \20481 );
nor \U$19813 ( \20483 , \20479 , \20482 );
nand \U$19814 ( \20484 , \20478 , \20483 );
not \U$19815 ( \20485 , \20484 );
or \U$19816 ( \20486 , \20475 , \20485 );
and \U$19817 ( \20487 , \17746 , \19073 );
nor \U$19818 ( \20488 , \20465 , \20473 );
nor \U$19819 ( \20489 , \20487 , \20488 );
nand \U$19820 ( \20490 , \20486 , \20489 );
xor \U$19821 ( \20491 , \20464 , \20490 );
xor \U$19822 ( \20492 , \20453 , \20491 );
not \U$19823 ( \20493 , \20474 );
nor \U$19824 ( \20494 , \20493 , \20488 );
xnor \U$19825 ( \20495 , \20494 , \20484 );
not \U$19826 ( \20496 , \20495 );
not \U$19827 ( \20497 , \20427 );
not \U$19828 ( \20498 , \20437 );
or \U$19829 ( \20499 , \20497 , \20498 );
nand \U$19830 ( \20500 , \20499 , \20414 );
or \U$19831 ( \20501 , \20437 , \20427 );
nand \U$19832 ( \20502 , \20500 , \20501 );
not \U$19833 ( \20503 , \20502 );
or \U$19834 ( \20504 , \20496 , \20503 );
xor \U$19835 ( \20505 , \20137 , \20171 );
nand \U$19836 ( \20506 , \20504 , \20505 );
not \U$19837 ( \20507 , \20502 );
not \U$19838 ( \20508 , \20495 );
nand \U$19839 ( \20509 , \20507 , \20508 );
nand \U$19840 ( \20510 , \20506 , \20509 );
xnor \U$19841 ( \20511 , \20492 , \20510 );
nand \U$19842 ( \20512 , \20452 , \20511 );
not \U$19843 ( \20513 , \20452 );
not \U$19844 ( \20514 , \20511 );
nand \U$19845 ( \20515 , \20513 , \20514 );
nand \U$19846 ( \20516 , \20512 , \20515 );
xor \U$19847 ( \20517 , \20502 , \20508 );
xor \U$19848 ( \20518 , \20517 , \20505 );
xor \U$19849 ( \20519 , \20278 , \20261 );
xnor \U$19850 ( \20520 , \20519 , \20289 );
not \U$19851 ( \20521 , \18465 );
not \U$19852 ( \20522 , \18686 );
or \U$19853 ( \20523 , \20521 , \20522 );
and \U$19854 ( \20524 , \17848 , \19077 );
and \U$19855 ( \20525 , \18243 , \18613 );
not \U$19856 ( \20526 , \18243 );
and \U$19857 ( \20527 , \20526 , \17891 );
nor \U$19858 ( \20528 , \20525 , \20527 );
nor \U$19859 ( \20529 , \20524 , \20528 );
nand \U$19860 ( \20530 , \20523 , \20529 );
not \U$19861 ( \20531 , \19883 );
and \U$19862 ( \20532 , \19261 , \18588 );
not \U$19863 ( \20533 , \19261 );
and \U$19864 ( \20534 , \20533 , \18536 );
nor \U$19865 ( \20535 , \20532 , \20534 );
nand \U$19866 ( \20536 , \19385 , \20535 );
and \U$19867 ( \20537 , \20531 , \20536 );
and \U$19868 ( \20538 , \20353 , \19387 );
and \U$19869 ( \20539 , \18820 , \18588 );
nor \U$19870 ( \20540 , \20538 , \20539 );
nor \U$19871 ( \20541 , \19385 , \20540 );
nor \U$19872 ( \20542 , \20537 , \20541 );
xor \U$19873 ( \20543 , \20530 , \20542 );
not \U$19874 ( \20544 , \19864 );
not \U$19875 ( \20545 , \18695 );
or \U$19876 ( \20546 , \20544 , \20545 );
and \U$19877 ( \20547 , \18641 , \18777 );
or \U$19878 ( \20548 , \20091 , \20415 );
or \U$19879 ( \20549 , \18685 , \20132 );
nand \U$19880 ( \20550 , \20548 , \20549 );
nor \U$19881 ( \20551 , \20547 , \20550 );
nand \U$19882 ( \20552 , \20546 , \20551 );
and \U$19883 ( \20553 , \20543 , \20552 );
and \U$19884 ( \20554 , \20530 , \20542 );
or \U$19885 ( \20555 , \20553 , \20554 );
xor \U$19886 ( \20556 , \20520 , \20555 );
and \U$19887 ( \20557 , \20395 , \20372 );
not \U$19888 ( \20558 , \20395 );
not \U$19889 ( \20559 , \20372 );
and \U$19890 ( \20560 , \20558 , \20559 );
nor \U$19891 ( \20561 , \20557 , \20560 );
and \U$19892 ( \20562 , \20556 , \20561 );
and \U$19893 ( \20563 , \20520 , \20555 );
nor \U$19894 ( \20564 , \20562 , \20563 );
not \U$19895 ( \20565 , \20564 );
not \U$19896 ( \20566 , \20019 );
nand \U$19897 ( \20567 , \20566 , \20032 );
not \U$19898 ( \20568 , \20209 );
not \U$19899 ( \20569 , \18825 );
or \U$19900 ( \20570 , \20568 , \20569 );
and \U$19901 ( \20571 , \18196 , \20043 );
or \U$19902 ( \20572 , \19024 , \20204 );
or \U$19903 ( \20573 , \19027 , \20021 );
nand \U$19904 ( \20574 , \20572 , \20573 );
nor \U$19905 ( \20575 , \20571 , \20574 );
nand \U$19906 ( \20576 , \20570 , \20575 );
not \U$19907 ( \20577 , \20576 );
xor \U$19908 ( \20578 , \20567 , \20577 );
xor \U$19909 ( \20579 , \20277 , \20272 );
and \U$19910 ( \20580 , \20578 , \20579 );
not \U$19911 ( \20581 , \20567 );
not \U$19912 ( \20582 , \20581 );
not \U$19913 ( \20583 , \20576 );
or \U$19914 ( \20584 , \20582 , \20583 );
nand \U$19915 ( \20585 , \17746 , \18755 );
nand \U$19916 ( \20586 , \20584 , \20585 );
nor \U$19917 ( \20587 , \20580 , \20586 );
not \U$19918 ( \20588 , \20587 );
not \U$19919 ( \20589 , \18680 );
not \U$19920 ( \20590 , \17645 );
or \U$19921 ( \20591 , \20589 , \20590 );
and \U$19922 ( \20592 , \17650 , \18679 );
or \U$19923 ( \20593 , \20302 , \19077 );
nand \U$19924 ( \20594 , \20355 , \19077 );
nand \U$19925 ( \20595 , \20593 , \20594 );
nor \U$19926 ( \20596 , \20592 , \20595 );
nand \U$19927 ( \20597 , \20591 , \20596 );
nand \U$19928 ( \20598 , \20588 , \20597 );
not \U$19929 ( \20599 , \20598 );
xor \U$19930 ( \20600 , \20300 , \20309 );
not \U$19931 ( \20601 , \20600 );
or \U$19932 ( \20602 , \20599 , \20601 );
or \U$19933 ( \20603 , \20598 , \20600 );
nand \U$19934 ( \20604 , \20602 , \20603 );
nand \U$19935 ( \20605 , \20565 , \20604 );
not \U$19936 ( \20606 , \20598 );
nand \U$19937 ( \20607 , \20606 , \20600 );
and \U$19938 ( \20608 , \20605 , \20607 );
xor \U$19939 ( \20609 , \20518 , \20608 );
xnor \U$19940 ( \20610 , \20444 , \20361 );
and \U$19941 ( \20611 , \20609 , \20610 );
and \U$19942 ( \20612 , \20518 , \20608 );
or \U$19943 ( \20613 , \20611 , \20612 );
and \U$19944 ( \20614 , \20516 , \20613 );
xor \U$19945 ( \20615 , \20518 , \20608 );
xor \U$19946 ( \20616 , \20615 , \20610 );
buf \U$19947 ( \20617 , \20439 );
not \U$19948 ( \20618 , \20399 );
and \U$19949 ( \20619 , \20617 , \20618 );
not \U$19950 ( \20620 , \20617 );
and \U$19951 ( \20621 , \20620 , \20399 );
nor \U$19952 ( \20622 , \20619 , \20621 );
xor \U$19953 ( \20623 , \20567 , \20579 );
xnor \U$19954 ( \20624 , \20623 , \20576 );
xor \U$19955 ( \20625 , \20074 , \20084 );
and \U$19956 ( \20626 , \20625 , \20096 );
and \U$19957 ( \20627 , \20074 , \20084 );
or \U$19958 ( \20628 , \20626 , \20627 );
xor \U$19959 ( \20629 , \20624 , \20628 );
xor \U$19960 ( \20630 , \20530 , \20542 );
xor \U$19961 ( \20631 , \20630 , \20552 );
and \U$19962 ( \20632 , \20629 , \20631 );
and \U$19963 ( \20633 , \20624 , \20628 );
or \U$19964 ( \20634 , \20632 , \20633 );
xnor \U$19965 ( \20635 , \20597 , \20587 );
not \U$19966 ( \20636 , \20635 );
not \U$19967 ( \20637 , \17747 );
not \U$19968 ( \20638 , \18761 );
and \U$19969 ( \20639 , \20637 , \20638 );
xor \U$19970 ( \20640 , \20013 , \20036 );
and \U$19971 ( \20641 , \20640 , \20049 );
and \U$19972 ( \20642 , \20013 , \20036 );
or \U$19973 ( \20643 , \20641 , \20642 );
nor \U$19974 ( \20644 , \20639 , \20643 );
not \U$19975 ( \20645 , \20644 );
or \U$19976 ( \20646 , \17655 , \18679 );
nand \U$19977 ( \20647 , \17705 , \18679 );
nand \U$19978 ( \20648 , \20646 , \20647 );
not \U$19979 ( \20649 , \20648 );
and \U$19980 ( \20650 , \18796 , \17650 );
not \U$19981 ( \20651 , \18796 );
and \U$19982 ( \20652 , \20651 , \17645 );
nor \U$19983 ( \20653 , \20650 , \20652 );
nand \U$19984 ( \20654 , \20649 , \20653 );
nand \U$19985 ( \20655 , \20645 , \20654 );
nand \U$19986 ( \20656 , \20636 , \20655 );
nand \U$19987 ( \20657 , \20634 , \20656 );
not \U$19988 ( \20658 , \20655 );
nand \U$19989 ( \20659 , \20658 , \20635 );
and \U$19990 ( \20660 , \20657 , \20659 );
xor \U$19991 ( \20661 , \20622 , \20660 );
not \U$19992 ( \20662 , \20564 );
not \U$19993 ( \20663 , \20604 );
and \U$19994 ( \20664 , \20662 , \20663 );
and \U$19995 ( \20665 , \20564 , \20604 );
nor \U$19996 ( \20666 , \20664 , \20665 );
and \U$19997 ( \20667 , \20661 , \20666 );
and \U$19998 ( \20668 , \20622 , \20660 );
or \U$19999 ( \20669 , \20667 , \20668 );
nand \U$20000 ( \20670 , \20616 , \20669 );
not \U$20001 ( \20671 , \20644 );
nor \U$20002 ( \20672 , \20671 , \20654 );
not \U$20003 ( \20673 , \20672 );
nand \U$20004 ( \20674 , \20673 , \20655 );
not \U$20005 ( \20675 , \20674 );
not \U$20006 ( \20676 , \20675 );
not \U$20007 ( \20677 , \19998 );
not \U$20008 ( \20678 , \20677 );
or \U$20009 ( \20679 , \20676 , \20678 );
not \U$20010 ( \20680 , \20674 );
not \U$20011 ( \20681 , \19998 );
or \U$20012 ( \20682 , \20680 , \20681 );
not \U$20013 ( \20683 , \20097 );
not \U$20014 ( \20684 , \20063 );
or \U$20015 ( \20685 , \20683 , \20684 );
nand \U$20016 ( \20686 , \20057 , \20050 );
nand \U$20017 ( \20687 , \20685 , \20686 );
nand \U$20018 ( \20688 , \20682 , \20687 );
nand \U$20019 ( \20689 , \20679 , \20688 );
xor \U$20020 ( \20690 , \20556 , \20561 );
nor \U$20021 ( \20691 , \20689 , \20690 );
nand \U$20022 ( \20692 , \20656 , \20659 );
and \U$20023 ( \20693 , \20692 , \20634 );
not \U$20024 ( \20694 , \20692 );
not \U$20025 ( \20695 , \20634 );
and \U$20026 ( \20696 , \20694 , \20695 );
nor \U$20027 ( \20697 , \20693 , \20696 );
or \U$20028 ( \20698 , \20691 , \20697 );
nand \U$20029 ( \20699 , \20689 , \20690 );
nand \U$20030 ( \20700 , \20698 , \20699 );
not \U$20031 ( \20701 , \20700 );
xor \U$20032 ( \20702 , \20622 , \20660 );
xor \U$20033 ( \20703 , \20702 , \20666 );
nand \U$20034 ( \20704 , \20701 , \20703 );
nand \U$20035 ( \20705 , \20670 , \20704 );
nor \U$20036 ( \20706 , \20614 , \20705 );
xor \U$20037 ( \20707 , \20677 , \20675 );
xnor \U$20038 ( \20708 , \20707 , \20687 );
xor \U$20039 ( \20709 , \20624 , \20628 );
xor \U$20040 ( \20710 , \20709 , \20631 );
not \U$20041 ( \20711 , \20710 );
xor \U$20042 ( \20712 , \19978 , \19999 );
and \U$20043 ( \20713 , \20712 , \20010 );
and \U$20044 ( \20714 , \19978 , \19999 );
or \U$20045 ( \20715 , \20713 , \20714 );
not \U$20046 ( \20716 , \20715 );
or \U$20047 ( \20717 , \20711 , \20716 );
or \U$20048 ( \20718 , \20715 , \20710 );
nand \U$20049 ( \20719 , \20717 , \20718 );
xor \U$20050 ( \20720 , \20708 , \20719 );
not \U$20051 ( \20721 , \20102 );
not \U$20052 ( \20722 , \20110 );
not \U$20053 ( \20723 , \20722 );
or \U$20054 ( \20724 , \20721 , \20723 );
not \U$20055 ( \20725 , \20102 );
not \U$20056 ( \20726 , \20725 );
not \U$20057 ( \20727 , \20110 );
or \U$20058 ( \20728 , \20726 , \20727 );
nand \U$20059 ( \20729 , \20728 , \20011 );
nand \U$20060 ( \20730 , \20724 , \20729 );
nand \U$20061 ( \20731 , \20720 , \20730 );
not \U$20062 ( \20732 , \20708 );
not \U$20063 ( \20733 , \20719 );
or \U$20064 ( \20734 , \20732 , \20733 );
not \U$20065 ( \20735 , \20710 );
nand \U$20066 ( \20736 , \20735 , \20715 );
nand \U$20067 ( \20737 , \20734 , \20736 );
xor \U$20068 ( \20738 , \20690 , \20689 );
xor \U$20069 ( \20739 , \20738 , \20697 );
nand \U$20070 ( \20740 , \20737 , \20739 );
nand \U$20071 ( \20741 , \20731 , \20740 );
not \U$20072 ( \20742 , \20741 );
nand \U$20073 ( \20743 , \20129 , \20706 , \20742 );
nand \U$20074 ( \20744 , \20118 , \20125 );
not \U$20075 ( \20745 , \20744 );
nand \U$20076 ( \20746 , \19969 , \19973 );
not \U$20077 ( \20747 , \20746 );
or \U$20078 ( \20748 , \20745 , \20747 );
nand \U$20079 ( \20749 , \20748 , \20127 );
or \U$20080 ( \20750 , \20749 , \20741 );
nor \U$20081 ( \20751 , \20720 , \20730 );
and \U$20082 ( \20752 , \20751 , \20740 );
nor \U$20083 ( \20753 , \20737 , \20739 );
nor \U$20084 ( \20754 , \20752 , \20753 );
nand \U$20085 ( \20755 , \20750 , \20754 );
not \U$20086 ( \20756 , \20241 );
not \U$20087 ( \20757 , \20756 );
not \U$20088 ( \20758 , \20448 );
or \U$20089 ( \20759 , \20757 , \20758 );
nand \U$20090 ( \20760 , \20759 , \20512 );
not \U$20091 ( \20761 , \20760 );
not \U$20092 ( \20762 , \20236 );
not \U$20093 ( \20763 , \20203 );
or \U$20094 ( \20764 , \20762 , \20763 );
nand \U$20095 ( \20765 , \20175 , \20201 );
nand \U$20096 ( \20766 , \20764 , \20765 );
and \U$20097 ( \20767 , \20464 , \20490 );
and \U$20098 ( \20768 , \17746 , \19898 );
not \U$20099 ( \20769 , \17641 );
not \U$20100 ( \20770 , \20459 );
or \U$20101 ( \20771 , \20769 , \20770 );
and \U$20102 ( \20772 , \19864 , \17813 );
not \U$20103 ( \20773 , \19864 );
and \U$20104 ( \20774 , \20773 , \17642 );
nor \U$20105 ( \20775 , \20772 , \20774 );
nand \U$20106 ( \20776 , \20775 , \17808 );
nand \U$20107 ( \20777 , \20771 , \20776 );
xor \U$20108 ( \20778 , \20768 , \20777 );
xor \U$20109 ( \20779 , \19743 , \20188 );
not \U$20110 ( \20780 , \20779 );
and \U$20111 ( \20781 , \18196 , \17534 );
or \U$20112 ( \20782 , \19027 , \17702 );
nand \U$20113 ( \20783 , \18300 , \17702 );
nand \U$20114 ( \20784 , \20782 , \20783 );
nor \U$20115 ( \20785 , \20781 , \20784 );
nand \U$20116 ( \20786 , \18825 , \17533 );
and \U$20117 ( \20787 , \20785 , \20786 );
not \U$20118 ( \20788 , \20787 );
and \U$20119 ( \20789 , \20780 , \20788 );
and \U$20120 ( \20790 , \20779 , \20787 );
nor \U$20121 ( \20791 , \20789 , \20790 );
xnor \U$20122 ( \20792 , \20778 , \20791 );
xor \U$20123 ( \20793 , \20767 , \20792 );
xnor \U$20124 ( \20794 , \20766 , \20793 );
not \U$20125 ( \20795 , \20794 );
xor \U$20126 ( \20796 , \20188 , \20189 );
not \U$20127 ( \20797 , \20196 );
and \U$20128 ( \20798 , \20796 , \20797 );
and \U$20129 ( \20799 , \20188 , \20189 );
or \U$20130 ( \20800 , \20798 , \20799 );
not \U$20131 ( \20801 , \20800 );
not \U$20132 ( \20802 , \20801 );
not \U$20133 ( \20803 , \20214 );
not \U$20134 ( \20804 , \20235 );
or \U$20135 ( \20805 , \20803 , \20804 );
nand \U$20136 ( \20806 , \20234 , \20224 );
nand \U$20137 ( \20807 , \20805 , \20806 );
not \U$20138 ( \20808 , \20807 );
not \U$20139 ( \20809 , \20808 );
or \U$20140 ( \20810 , \20802 , \20809 );
nand \U$20141 ( \20811 , \20807 , \20800 );
nand \U$20142 ( \20812 , \20810 , \20811 );
not \U$20143 ( \20813 , \20812 );
not \U$20144 ( \20814 , \20331 );
not \U$20145 ( \20815 , \18695 );
or \U$20146 ( \20816 , \20814 , \20815 );
and \U$20147 ( \20817 , \18641 , \17887 );
or \U$20148 ( \20818 , \20091 , \17792 );
not \U$20149 ( \20819 , \20177 );
or \U$20150 ( \20820 , \18685 , \20819 );
nand \U$20151 ( \20821 , \20818 , \20820 );
nor \U$20152 ( \20822 , \20817 , \20821 );
nand \U$20153 ( \20823 , \20816 , \20822 );
not \U$20154 ( \20824 , \20041 );
not \U$20155 ( \20825 , \17844 );
or \U$20156 ( \20826 , \20824 , \20825 );
and \U$20157 ( \20827 , \17849 , \19273 );
or \U$20158 ( \20828 , \20070 , \20043 );
nand \U$20159 ( \20829 , \18888 , \20043 );
nand \U$20160 ( \20830 , \20828 , \20829 );
nor \U$20161 ( \20831 , \20827 , \20830 );
nand \U$20162 ( \20832 , \20826 , \20831 );
not \U$20163 ( \20833 , \20832 );
and \U$20164 ( \20834 , \20823 , \20833 );
not \U$20165 ( \20835 , \20823 );
and \U$20166 ( \20836 , \20835 , \20832 );
or \U$20167 ( \20837 , \20834 , \20836 );
nor \U$20168 ( \20838 , \18767 , \20226 );
not \U$20169 ( \20839 , \20838 );
not \U$20170 ( \20840 , \18763 );
not \U$20171 ( \20841 , \20204 );
and \U$20172 ( \20842 , \20840 , \20841 );
and \U$20173 ( \20843 , \18931 , \20204 );
nor \U$20174 ( \20844 , \20842 , \20843 );
nand \U$20175 ( \20845 , \19008 , \20226 );
nand \U$20176 ( \20846 , \20839 , \20844 , \20845 );
xor \U$20177 ( \20847 , \20837 , \20846 );
not \U$20178 ( \20848 , \20847 );
not \U$20179 ( \20849 , \20848 );
and \U$20180 ( \20850 , \20813 , \20849 );
and \U$20181 ( \20851 , \20812 , \20848 );
nor \U$20182 ( \20852 , \20850 , \20851 );
not \U$20183 ( \20853 , \20852 );
not \U$20184 ( \20854 , \20853 );
not \U$20185 ( \20855 , \20491 );
not \U$20186 ( \20856 , \20453 );
not \U$20187 ( \20857 , \20510 );
or \U$20188 ( \20858 , \20856 , \20857 );
or \U$20189 ( \20859 , \20510 , \20453 );
nand \U$20190 ( \20860 , \20858 , \20859 );
not \U$20191 ( \20861 , \20860 );
or \U$20192 ( \20862 , \20855 , \20861 );
not \U$20193 ( \20863 , \20453 );
nand \U$20194 ( \20864 , \20863 , \20510 );
nand \U$20195 ( \20865 , \20862 , \20864 );
not \U$20196 ( \20866 , \20865 );
not \U$20197 ( \20867 , \20866 );
or \U$20198 ( \20868 , \20854 , \20867 );
nand \U$20199 ( \20869 , \20865 , \20852 );
nand \U$20200 ( \20870 , \20868 , \20869 );
not \U$20201 ( \20871 , \20870 );
or \U$20202 ( \20872 , \20795 , \20871 );
or \U$20203 ( \20873 , \20870 , \20794 );
nand \U$20204 ( \20874 , \20872 , \20873 );
not \U$20205 ( \20875 , \20874 );
or \U$20206 ( \20876 , \20761 , \20875 );
nand \U$20207 ( \20877 , \20876 , \20614 );
not \U$20208 ( \20878 , \20705 );
nand \U$20209 ( \20879 , \20755 , \20877 , \20878 );
not \U$20210 ( \20880 , \20760 );
not \U$20211 ( \20881 , \20874 );
or \U$20212 ( \20882 , \20880 , \20881 );
not \U$20213 ( \20883 , \20613 );
nand \U$20214 ( \20884 , \20883 , \20512 , \20515 );
nand \U$20215 ( \20885 , \20882 , \20884 );
not \U$20216 ( \20886 , \20670 );
not \U$20217 ( \20887 , \20703 );
nand \U$20218 ( \20888 , \20700 , \20887 );
or \U$20219 ( \20889 , \20886 , \20888 );
or \U$20220 ( \20890 , \20616 , \20669 );
nand \U$20221 ( \20891 , \20889 , \20890 );
or \U$20222 ( \20892 , \20885 , \20891 );
nand \U$20223 ( \20893 , \20892 , \20877 );
nand \U$20224 ( \20894 , \20743 , \20879 , \20893 );
or \U$20225 ( \20895 , \20874 , \20760 );
nand \U$20226 ( \20896 , \20894 , \20895 );
not \U$20227 ( \20897 , \20896 );
not \U$20228 ( \20898 , \20226 );
not \U$20229 ( \20899 , \17743 );
or \U$20230 ( \20900 , \20898 , \20899 );
or \U$20231 ( \20901 , \17634 , \20226 );
nand \U$20232 ( \20902 , \20900 , \20901 );
nand \U$20233 ( \20903 , \20902 , \17739 );
not \U$20234 ( \20904 , \20204 );
not \U$20235 ( \20905 , \17634 );
not \U$20236 ( \20906 , \20905 );
or \U$20237 ( \20907 , \20904 , \20906 );
or \U$20238 ( \20908 , \17742 , \19138 );
nand \U$20239 ( \20909 , \20907 , \20908 );
nand \U$20240 ( \20910 , \20909 , \17740 );
nand \U$20241 ( \20911 , \20903 , \17741 , \20910 );
not \U$20242 ( \20912 , \20911 );
nand \U$20243 ( \20913 , \18241 , \20182 );
not \U$20244 ( \20914 , \20913 );
not \U$20245 ( \20915 , \18192 );
nor \U$20246 ( \20916 , \20915 , \18832 );
or \U$20247 ( \20917 , \17701 , \18194 );
nand \U$20248 ( \20918 , \18194 , \18191 , \17701 );
nand \U$20249 ( \20919 , \20917 , \20918 );
nor \U$20250 ( \20920 , \20916 , \20919 );
not \U$20251 ( \20921 , \20920 );
and \U$20252 ( \20922 , \20914 , \20921 );
and \U$20253 ( \20923 , \20913 , \20920 );
nor \U$20254 ( \20924 , \20922 , \20923 );
not \U$20255 ( \20925 , \20924 );
not \U$20256 ( \20926 , \20925 );
or \U$20257 ( \20927 , \20912 , \20926 );
buf \U$20258 ( \20928 , \20920 );
not \U$20259 ( \20929 , \20928 );
nand \U$20260 ( \20930 , \20913 , \20929 );
nand \U$20261 ( \20931 , \20927 , \20930 );
not \U$20262 ( \20932 , \20232 );
not \U$20263 ( \20933 , \17849 );
or \U$20264 ( \20934 , \20932 , \20933 );
and \U$20265 ( \20935 , \17887 , \18888 );
not \U$20266 ( \20936 , \17887 );
and \U$20267 ( \20937 , \20936 , \17892 );
nor \U$20268 ( \20938 , \20935 , \20937 );
nand \U$20269 ( \20939 , \20934 , \20938 );
and \U$20270 ( \20940 , \20222 , \20226 );
nor \U$20271 ( \20941 , \20939 , \20940 );
xor \U$20272 ( \20942 , \20931 , \20941 );
and \U$20273 ( \20943 , \20204 , \17812 );
not \U$20274 ( \20944 , \20204 );
and \U$20275 ( \20945 , \20944 , \17813 );
nor \U$20276 ( \20946 , \20943 , \20945 );
and \U$20277 ( \20947 , \17807 , \20946 );
not \U$20278 ( \20948 , \20209 );
not \U$20279 ( \20949 , \17643 );
or \U$20280 ( \20950 , \20948 , \20949 );
or \U$20281 ( \20951 , \17813 , \20209 );
nand \U$20282 ( \20952 , \20950 , \20951 );
and \U$20283 ( \20953 , \20952 , \17809 );
nor \U$20284 ( \20954 , \20947 , \20953 );
nand \U$20285 ( \20955 , \20954 , \17810 );
xor \U$20286 ( \20956 , \20942 , \20955 );
not \U$20287 ( \20957 , \20956 );
nand \U$20288 ( \20958 , \17746 , \19261 );
not \U$20289 ( \20959 , \20958 );
and \U$20290 ( \20960 , \18931 , \20232 );
and \U$20291 ( \20961 , \18536 , \20331 );
and \U$20292 ( \20962 , \17887 , \18588 );
nor \U$20293 ( \20963 , \20961 , \20962 );
not \U$20294 ( \20964 , \20963 );
not \U$20295 ( \20965 , \19385 );
or \U$20296 ( \20966 , \20964 , \20965 );
or \U$20297 ( \20967 , \18763 , \20232 );
nand \U$20298 ( \20968 , \20966 , \20967 );
nor \U$20299 ( \20969 , \20960 , \20968 );
not \U$20300 ( \20970 , \20969 );
or \U$20301 ( \20971 , \20959 , \20970 );
not \U$20302 ( \20972 , \20787 );
and \U$20303 ( \20973 , \20779 , \20972 );
and \U$20304 ( \20974 , \19743 , \20188 );
nor \U$20305 ( \20975 , \20973 , \20974 );
not \U$20306 ( \20976 , \20975 );
nand \U$20307 ( \20977 , \20971 , \20976 );
not \U$20308 ( \20978 , \20977 );
and \U$20309 ( \20979 , \18641 , \17534 );
and \U$20310 ( \20980 , \17702 , \20091 );
not \U$20311 ( \20981 , \17702 );
and \U$20312 ( \20982 , \20981 , \18685 );
nor \U$20313 ( \20983 , \20980 , \20982 );
nor \U$20314 ( \20984 , \20979 , \20983 );
nand \U$20315 ( \20985 , \18695 , \17533 );
nand \U$20316 ( \20986 , \20984 , \20985 );
not \U$20317 ( \20987 , \18767 );
not \U$20318 ( \20988 , \17829 );
and \U$20319 ( \20989 , \20987 , \20988 );
and \U$20320 ( \20990 , \19008 , \20819 );
nor \U$20321 ( \20991 , \20989 , \20990 );
and \U$20322 ( \20992 , \19883 , \20963 );
and \U$20323 ( \20993 , \17746 , \18777 );
nor \U$20324 ( \20994 , \20992 , \20993 );
nand \U$20325 ( \20995 , \20991 , \20994 );
xor \U$20326 ( \20996 , \20986 , \20995 );
nand \U$20327 ( \20997 , \20978 , \20996 );
not \U$20328 ( \20998 , \20997 );
and \U$20329 ( \20999 , \20911 , \20924 );
not \U$20330 ( \21000 , \20911 );
and \U$20331 ( \21001 , \21000 , \20925 );
or \U$20332 ( \21002 , \20999 , \21001 );
nand \U$20333 ( \21003 , \17807 , \20952 );
not \U$20334 ( \21004 , \20041 );
not \U$20335 ( \21005 , \17812 );
or \U$20336 ( \21006 , \21004 , \21005 );
or \U$20337 ( \21007 , \17812 , \20132 );
nand \U$20338 ( \21008 , \21006 , \21007 );
and \U$20339 ( \21009 , \21008 , \17809 );
nor \U$20340 ( \21010 , \20043 , \20132 );
not \U$20341 ( \21011 , \21010 );
not \U$20342 ( \21012 , \17643 );
or \U$20343 ( \21013 , \21011 , \21012 );
nand \U$20344 ( \21014 , \20043 , \20041 );
or \U$20345 ( \21015 , \17813 , \21014 );
nand \U$20346 ( \21016 , \21013 , \21015 );
nor \U$20347 ( \21017 , \21009 , \21016 );
and \U$20348 ( \21018 , \17810 , \21003 , \21017 );
xor \U$20349 ( \21019 , \21002 , \21018 );
not \U$20350 ( \21020 , \20929 );
and \U$20351 ( \21021 , \18641 , \20819 );
or \U$20352 ( \21022 , \18685 , \17534 );
nand \U$20353 ( \21023 , \18877 , \17534 );
nand \U$20354 ( \21024 , \21022 , \21023 );
nor \U$20355 ( \21025 , \21021 , \21024 );
nand \U$20356 ( \21026 , \18695 , \20177 );
nand \U$20357 ( \21027 , \21025 , \21026 );
not \U$20358 ( \21028 , \21027 );
or \U$20359 ( \21029 , \21020 , \21028 );
not \U$20360 ( \21030 , \20209 );
not \U$20361 ( \21031 , \17848 );
or \U$20362 ( \21032 , \21030 , \21031 );
and \U$20363 ( \21033 , \20204 , \17892 );
not \U$20364 ( \21034 , \20204 );
and \U$20365 ( \21035 , \21034 , \18888 );
nor \U$20366 ( \21036 , \21033 , \21035 );
nand \U$20367 ( \21037 , \21032 , \21036 );
nor \U$20368 ( \21038 , \17845 , \20209 );
nor \U$20369 ( \21039 , \21037 , \21038 );
nand \U$20370 ( \21040 , \21029 , \21039 );
not \U$20371 ( \21041 , \21027 );
nand \U$20372 ( \21042 , \21041 , \20928 );
nand \U$20373 ( \21043 , \21040 , \21042 );
xor \U$20374 ( \21044 , \21019 , \21043 );
not \U$20375 ( \21045 , \21044 );
not \U$20376 ( \21046 , \21045 );
or \U$20377 ( \21047 , \20998 , \21046 );
not \U$20378 ( \21048 , \20996 );
nand \U$20379 ( \21049 , \21048 , \20977 );
nand \U$20380 ( \21050 , \21047 , \21049 );
xor \U$20381 ( \21051 , \20957 , \21050 );
not \U$20382 ( \21052 , \21018 );
not \U$20383 ( \21053 , \21052 );
or \U$20384 ( \21054 , \21043 , \21002 );
not \U$20385 ( \21055 , \21054 );
or \U$20386 ( \21056 , \21053 , \21055 );
nand \U$20387 ( \21057 , \21043 , \21002 );
nand \U$20388 ( \21058 , \21056 , \21057 );
and \U$20389 ( \21059 , \19387 , \17533 );
and \U$20390 ( \21060 , \17534 , \18588 );
nor \U$20391 ( \21061 , \21059 , \21060 );
and \U$20392 ( \21062 , \19385 , \21061 );
or \U$20393 ( \21063 , \19883 , \21062 );
and \U$20394 ( \21064 , \19387 , \17791 );
and \U$20395 ( \21065 , \20176 , \18588 );
nor \U$20396 ( \21066 , \21064 , \21065 );
or \U$20397 ( \21067 , \19385 , \21066 );
nand \U$20398 ( \21068 , \21063 , \21067 );
not \U$20399 ( \21069 , \21068 );
and \U$20400 ( \21070 , \18685 , \18810 );
or \U$20401 ( \21071 , \18639 , \17702 );
nand \U$20402 ( \21072 , \18639 , \18794 , \17702 );
nand \U$20403 ( \21073 , \21071 , \21072 );
nor \U$20404 ( \21074 , \21070 , \21073 );
not \U$20405 ( \21075 , \21074 );
and \U$20406 ( \21076 , \21069 , \21075 );
and \U$20407 ( \21077 , \21068 , \21074 );
nor \U$20408 ( \21078 , \21076 , \21077 );
nand \U$20409 ( \21079 , \17746 , \20041 );
and \U$20410 ( \21080 , \21078 , \21079 );
and \U$20411 ( \21081 , \20986 , \20995 );
and \U$20412 ( \21082 , \21080 , \21081 );
not \U$20413 ( \21083 , \21080 );
not \U$20414 ( \21084 , \21081 );
and \U$20415 ( \21085 , \21083 , \21084 );
nor \U$20416 ( \21086 , \21082 , \21085 );
not \U$20417 ( \21087 , \21086 );
and \U$20418 ( \21088 , \21058 , \21087 );
not \U$20419 ( \21089 , \21058 );
and \U$20420 ( \21090 , \21089 , \21086 );
nor \U$20421 ( \21091 , \21088 , \21090 );
and \U$20422 ( \21092 , \21051 , \21091 );
and \U$20423 ( \21093 , \20957 , \21050 );
nor \U$20424 ( \21094 , \21092 , \21093 );
not \U$20425 ( \21095 , \21094 );
not \U$20426 ( \21096 , \20955 );
not \U$20427 ( \21097 , \20942 );
not \U$20428 ( \21098 , \21097 );
or \U$20429 ( \21099 , \21096 , \21098 );
not \U$20430 ( \21100 , \20941 );
nand \U$20431 ( \21101 , \21100 , \20931 );
nand \U$20432 ( \21102 , \21099 , \21101 );
not \U$20433 ( \21103 , \21078 );
nor \U$20434 ( \21104 , \21103 , \21068 );
nand \U$20435 ( \21105 , \19420 , \18685 );
not \U$20436 ( \21106 , \21105 );
not \U$20437 ( \21107 , \20331 );
not \U$20438 ( \21108 , \17849 );
or \U$20439 ( \21109 , \21107 , \21108 );
and \U$20440 ( \21110 , \20819 , \18888 );
not \U$20441 ( \21111 , \20819 );
and \U$20442 ( \21112 , \21111 , \18461 );
nor \U$20443 ( \21113 , \21110 , \21112 );
nand \U$20444 ( \21114 , \21109 , \21113 );
and \U$20445 ( \21115 , \20222 , \17887 );
nor \U$20446 ( \21116 , \21114 , \21115 );
not \U$20447 ( \21117 , \21116 );
not \U$20448 ( \21118 , \21117 );
or \U$20449 ( \21119 , \21106 , \21118 );
not \U$20450 ( \21120 , \21105 );
nand \U$20451 ( \21121 , \21120 , \21116 );
nand \U$20452 ( \21122 , \21119 , \21121 );
not \U$20453 ( \21123 , \17702 );
not \U$20454 ( \21124 , \18758 );
or \U$20455 ( \21125 , \21123 , \21124 );
not \U$20456 ( \21126 , \18926 );
not \U$20457 ( \21127 , \17533 );
and \U$20458 ( \21128 , \21126 , \21127 );
and \U$20459 ( \21129 , \17533 , \18931 );
nor \U$20460 ( \21130 , \21128 , \21129 );
nand \U$20461 ( \21131 , \21125 , \21130 );
nor \U$20462 ( \21132 , \18767 , \17702 );
nor \U$20463 ( \21133 , \21131 , \21132 );
buf \U$20464 ( \21134 , \21133 );
xor \U$20465 ( \21135 , \21122 , \21134 );
xnor \U$20466 ( \21136 , \21104 , \21135 );
xor \U$20467 ( \21137 , \21102 , \21136 );
not \U$20468 ( \21138 , \21087 );
not \U$20469 ( \21139 , \21058 );
or \U$20470 ( \21140 , \21138 , \21139 );
nand \U$20471 ( \21141 , \21080 , \21084 );
nand \U$20472 ( \21142 , \21140 , \21141 );
not \U$20473 ( \21143 , \20226 );
not \U$20474 ( \21144 , \17812 );
or \U$20475 ( \21145 , \21143 , \21144 );
or \U$20476 ( \21146 , \17812 , \20226 );
nand \U$20477 ( \21147 , \21145 , \21146 );
nand \U$20478 ( \21148 , \17807 , \21147 );
nand \U$20479 ( \21149 , \20946 , \17809 );
nand \U$20480 ( \21150 , \17810 , \21148 , \21149 );
nand \U$20481 ( \21151 , \17746 , \20043 );
and \U$20482 ( \21152 , \20941 , \21151 );
and \U$20483 ( \21153 , \21150 , \21152 );
nor \U$20484 ( \21154 , \21150 , \21152 );
nor \U$20485 ( \21155 , \21153 , \21154 );
and \U$20486 ( \21156 , \21142 , \21155 );
not \U$20487 ( \21157 , \21142 );
not \U$20488 ( \21158 , \21155 );
and \U$20489 ( \21159 , \21157 , \21158 );
or \U$20490 ( \21160 , \21156 , \21159 );
xor \U$20491 ( \21161 , \21137 , \21160 );
nand \U$20492 ( \21162 , \21095 , \21161 );
xor \U$20493 ( \21163 , \20956 , \21091 );
xor \U$20494 ( \21164 , \21163 , \21050 );
not \U$20495 ( \21165 , \21164 );
and \U$20496 ( \21166 , \17657 , \20041 );
and \U$20497 ( \21167 , \17705 , \19273 );
nor \U$20498 ( \21168 , \21166 , \21167 );
not \U$20499 ( \21169 , \17807 );
nand \U$20500 ( \21170 , \21169 , \20775 );
nand \U$20501 ( \21171 , \21168 , \21170 );
xor \U$20502 ( \21172 , \20929 , \21039 );
xnor \U$20503 ( \21173 , \21172 , \21027 );
xor \U$20504 ( \21174 , \21171 , \21173 );
not \U$20505 ( \21175 , \20846 );
not \U$20506 ( \21176 , \20837 );
or \U$20507 ( \21177 , \21175 , \21176 );
not \U$20508 ( \21178 , \20833 );
nand \U$20509 ( \21179 , \21178 , \20823 );
nand \U$20510 ( \21180 , \21177 , \21179 );
and \U$20511 ( \21181 , \21174 , \21180 );
and \U$20512 ( \21182 , \21171 , \21173 );
nor \U$20513 ( \21183 , \21181 , \21182 );
not \U$20514 ( \21184 , \21183 );
not \U$20515 ( \21185 , \20977 );
not \U$20516 ( \21186 , \20996 );
or \U$20517 ( \21187 , \21185 , \21186 );
or \U$20518 ( \21188 , \20996 , \20977 );
nand \U$20519 ( \21189 , \21187 , \21188 );
not \U$20520 ( \21190 , \21189 );
not \U$20521 ( \21191 , \21045 );
or \U$20522 ( \21192 , \21190 , \21191 );
not \U$20523 ( \21193 , \21189 );
nand \U$20524 ( \21194 , \21193 , \21044 );
nand \U$20525 ( \21195 , \21192 , \21194 );
not \U$20526 ( \21196 , \21195 );
or \U$20527 ( \21197 , \21184 , \21196 );
or \U$20528 ( \21198 , \21195 , \21183 );
nand \U$20529 ( \21199 , \21197 , \21198 );
not \U$20530 ( \21200 , \20847 );
not \U$20531 ( \21201 , \20812 );
or \U$20532 ( \21202 , \21200 , \21201 );
nand \U$20533 ( \21203 , \20807 , \20801 );
nand \U$20534 ( \21204 , \21202 , \21203 );
not \U$20535 ( \21205 , \21204 );
not \U$20536 ( \21206 , \21205 );
not \U$20537 ( \21207 , \20768 );
not \U$20538 ( \21208 , \20777 );
nand \U$20539 ( \21209 , \21208 , \20791 );
not \U$20540 ( \21210 , \21209 );
or \U$20541 ( \21211 , \21207 , \21210 );
not \U$20542 ( \21212 , \20791 );
nand \U$20543 ( \21213 , \21212 , \20777 );
nand \U$20544 ( \21214 , \21211 , \21213 );
nand \U$20545 ( \21215 , \20975 , \20958 );
and \U$20546 ( \21216 , \21215 , \20969 );
not \U$20547 ( \21217 , \21215 );
not \U$20548 ( \21218 , \20969 );
and \U$20549 ( \21219 , \21217 , \21218 );
nor \U$20550 ( \21220 , \21216 , \21219 );
xor \U$20551 ( \21221 , \21214 , \21220 );
not \U$20552 ( \21222 , \21221 );
and \U$20553 ( \21223 , \21206 , \21222 );
not \U$20554 ( \21224 , \21214 );
nor \U$20555 ( \21225 , \21224 , \21220 );
nor \U$20556 ( \21226 , \21223 , \21225 );
not \U$20557 ( \21227 , \21226 );
nand \U$20558 ( \21228 , \21199 , \21227 );
not \U$20559 ( \21229 , \21183 );
nand \U$20560 ( \21230 , \21229 , \21195 );
nand \U$20561 ( \21231 , \21165 , \21228 , \21230 );
and \U$20562 ( \21232 , \21162 , \21231 );
not \U$20563 ( \21233 , \21227 );
not \U$20564 ( \21234 , \21199 );
not \U$20565 ( \21235 , \21234 );
or \U$20566 ( \21236 , \21233 , \21235 );
nand \U$20567 ( \21237 , \21199 , \21226 );
nand \U$20568 ( \21238 , \21236 , \21237 );
and \U$20569 ( \21239 , \20766 , \20793 );
and \U$20570 ( \21240 , \20767 , \20792 );
nor \U$20571 ( \21241 , \21239 , \21240 );
not \U$20572 ( \21242 , \21241 );
xor \U$20573 ( \21243 , \21180 , \21174 );
not \U$20574 ( \21244 , \21243 );
or \U$20575 ( \21245 , \21242 , \21244 );
or \U$20576 ( \21246 , \21241 , \21243 );
nand \U$20577 ( \21247 , \21245 , \21246 );
not \U$20578 ( \21248 , \21247 );
not \U$20579 ( \21249 , \21204 );
not \U$20580 ( \21250 , \21221 );
and \U$20581 ( \21251 , \21249 , \21250 );
and \U$20582 ( \21252 , \21204 , \21221 );
nor \U$20583 ( \21253 , \21251 , \21252 );
not \U$20584 ( \21254 , \21253 );
not \U$20585 ( \21255 , \21254 );
or \U$20586 ( \21256 , \21248 , \21255 );
not \U$20587 ( \21257 , \21241 );
nand \U$20588 ( \21258 , \21257 , \21243 );
nand \U$20589 ( \21259 , \21256 , \21258 );
nor \U$20590 ( \21260 , \21238 , \21259 );
not \U$20591 ( \21261 , \21247 );
not \U$20592 ( \21262 , \21261 );
not \U$20593 ( \21263 , \21254 );
or \U$20594 ( \21264 , \21262 , \21263 );
nand \U$20595 ( \21265 , \21247 , \21253 );
nand \U$20596 ( \21266 , \21264 , \21265 );
not \U$20597 ( \21267 , \20794 );
not \U$20598 ( \21268 , \21267 );
not \U$20599 ( \21269 , \20870 );
or \U$20600 ( \21270 , \21268 , \21269 );
nand \U$20601 ( \21271 , \20865 , \20853 );
nand \U$20602 ( \21272 , \21270 , \21271 );
nor \U$20603 ( \21273 , \21266 , \21272 );
nor \U$20604 ( \21274 , \21260 , \21273 );
nand \U$20605 ( \21275 , \21232 , \21274 );
not \U$20606 ( \21276 , \17894 );
not \U$20607 ( \21277 , \17840 );
or \U$20608 ( \21278 , \21276 , \21277 );
nand \U$20609 ( \21279 , \21278 , \17895 );
not \U$20610 ( \21280 , \21279 );
not \U$20611 ( \21281 , \17534 );
not \U$20612 ( \21282 , \17844 );
or \U$20613 ( \21283 , \21281 , \21282 );
and \U$20614 ( \21284 , \17849 , \17533 );
and \U$20615 ( \21285 , \17706 , \18461 );
and \U$20616 ( \21286 , \18888 , \17702 );
nor \U$20617 ( \21287 , \21284 , \21285 , \21286 );
nand \U$20618 ( \21288 , \21283 , \21287 );
not \U$20619 ( \21289 , \17829 );
not \U$20620 ( \21290 , \17844 );
or \U$20621 ( \21291 , \21289 , \21290 );
and \U$20622 ( \21292 , \17849 , \20177 );
and \U$20623 ( \21293 , \17533 , \18461 );
and \U$20624 ( \21294 , \18888 , \17534 );
nor \U$20625 ( \21295 , \21292 , \21293 , \21294 );
nand \U$20626 ( \21296 , \21291 , \21295 );
not \U$20627 ( \21297 , \21296 );
and \U$20628 ( \21298 , \21288 , \21297 );
not \U$20629 ( \21299 , \21288 );
and \U$20630 ( \21300 , \21299 , \21296 );
or \U$20631 ( \21301 , \21298 , \21300 );
and \U$20632 ( \21302 , \21301 , \19042 );
and \U$20633 ( \21303 , \21288 , \21296 );
nor \U$20634 ( \21304 , \21302 , \21303 );
or \U$20635 ( \21305 , \21280 , \21304 );
and \U$20636 ( \21306 , \21304 , \21279 );
not \U$20637 ( \21307 , \21304 );
and \U$20638 ( \21308 , \21307 , \21280 );
or \U$20639 ( \21309 , \21306 , \21308 );
not \U$20640 ( \21310 , \21309 );
and \U$20641 ( \21311 , \18931 , \17706 );
or \U$20642 ( \21312 , \18763 , \17706 );
or \U$20643 ( \21313 , \17747 , \20204 );
nand \U$20644 ( \21314 , \21312 , \21313 );
nor \U$20645 ( \21315 , \21311 , \21314 );
nand \U$20646 ( \21316 , \21315 , \18767 );
nand \U$20647 ( \21317 , \21297 , \21316 );
not \U$20648 ( \21318 , \21317 );
not \U$20649 ( \21319 , \17887 );
not \U$20650 ( \21320 , \17645 );
or \U$20651 ( \21321 , \21319 , \21320 );
and \U$20652 ( \21322 , \17650 , \20331 );
not \U$20653 ( \21323 , \17705 );
not \U$20654 ( \21324 , \17792 );
or \U$20655 ( \21325 , \21323 , \21324 );
or \U$20656 ( \21326 , \17656 , \17792 );
nand \U$20657 ( \21327 , \21325 , \21326 );
nor \U$20658 ( \21328 , \21322 , \21327 );
nand \U$20659 ( \21329 , \21321 , \21328 );
not \U$20660 ( \21330 , \21329 );
nand \U$20661 ( \21331 , \17746 , \20226 );
not \U$20662 ( \21332 , \21331 );
and \U$20663 ( \21333 , \21330 , \21332 );
and \U$20664 ( \21334 , \21329 , \21331 );
nor \U$20665 ( \21335 , \21333 , \21334 );
not \U$20666 ( \21336 , \21335 );
nand \U$20667 ( \21337 , \21318 , \21336 );
not \U$20668 ( \21338 , \21331 );
nand \U$20669 ( \21339 , \21338 , \21329 );
and \U$20670 ( \21340 , \21337 , \21339 );
or \U$20671 ( \21341 , \21310 , \21340 );
nand \U$20672 ( \21342 , \21305 , \21341 );
not \U$20673 ( \21343 , \17895 );
not \U$20674 ( \21344 , \17827 );
or \U$20675 ( \21345 , \21343 , \21344 );
or \U$20676 ( \21346 , \17827 , \17895 );
nand \U$20677 ( \21347 , \21345 , \21346 );
nor \U$20678 ( \21348 , \21342 , \21347 );
not \U$20679 ( \21349 , \21348 );
not \U$20680 ( \21350 , \21309 );
not \U$20681 ( \21351 , \21340 );
and \U$20682 ( \21352 , \21350 , \21351 );
and \U$20683 ( \21353 , \21340 , \21309 );
nor \U$20684 ( \21354 , \21352 , \21353 );
and \U$20685 ( \21355 , \21301 , \19042 );
not \U$20686 ( \21356 , \21301 );
not \U$20687 ( \21357 , \19042 );
and \U$20688 ( \21358 , \21356 , \21357 );
nor \U$20689 ( \21359 , \21355 , \21358 );
not \U$20690 ( \21360 , \21359 );
and \U$20691 ( \21361 , \21147 , \17809 );
or \U$20692 ( \21362 , \17812 , \20226 , \17887 );
nand \U$20693 ( \21363 , \17812 , \20226 , \17887 );
nand \U$20694 ( \21364 , \21362 , \21363 );
nor \U$20695 ( \21365 , \21361 , \21364 );
not \U$20696 ( \21366 , \17887 );
not \U$20697 ( \21367 , \17812 );
or \U$20698 ( \21368 , \21366 , \21367 );
or \U$20699 ( \21369 , \17812 , \17887 );
nand \U$20700 ( \21370 , \21368 , \21369 );
nand \U$20701 ( \21371 , \17807 , \21370 );
and \U$20702 ( \21372 , \21365 , \17810 , \21371 );
not \U$20703 ( \21373 , \21105 );
not \U$20704 ( \21374 , \21133 );
or \U$20705 ( \21375 , \21373 , \21374 );
nand \U$20706 ( \21376 , \21375 , \21117 );
or \U$20707 ( \21377 , \21105 , \21133 );
nand \U$20708 ( \21378 , \21376 , \21377 );
xor \U$20709 ( \21379 , \21372 , \21378 );
and \U$20710 ( \21380 , \21379 , \21154 );
and \U$20711 ( \21381 , \21372 , \21378 );
or \U$20712 ( \21382 , \21380 , \21381 );
not \U$20713 ( \21383 , \21382 );
or \U$20714 ( \21384 , \21360 , \21383 );
or \U$20715 ( \21385 , \21382 , \21359 );
and \U$20716 ( \21386 , \21317 , \21336 );
not \U$20717 ( \21387 , \21317 );
and \U$20718 ( \21388 , \21387 , \21335 );
or \U$20719 ( \21389 , \21386 , \21388 );
nand \U$20720 ( \21390 , \21385 , \21389 );
nand \U$20721 ( \21391 , \21384 , \21390 );
not \U$20722 ( \21392 , \21391 );
nand \U$20723 ( \21393 , \21354 , \21392 );
not \U$20724 ( \21394 , \21393 );
not \U$20725 ( \21395 , \21137 );
not \U$20726 ( \21396 , \21160 );
or \U$20727 ( \21397 , \21395 , \21396 );
nand \U$20728 ( \21398 , \21142 , \21158 );
nand \U$20729 ( \21399 , \21397 , \21398 );
not \U$20730 ( \21400 , \21102 );
not \U$20731 ( \21401 , \21136 );
or \U$20732 ( \21402 , \21400 , \21401 );
not \U$20733 ( \21403 , \21104 );
nand \U$20734 ( \21404 , \21403 , \21135 );
nand \U$20735 ( \21405 , \21402 , \21404 );
not \U$20736 ( \21406 , \21296 );
not \U$20737 ( \21407 , \21316 );
and \U$20738 ( \21408 , \21406 , \21407 );
and \U$20739 ( \21409 , \21296 , \21316 );
nor \U$20740 ( \21410 , \21408 , \21409 );
not \U$20741 ( \21411 , \21410 );
xor \U$20742 ( \21412 , \21372 , \21378 );
xor \U$20743 ( \21413 , \21412 , \21154 );
not \U$20744 ( \21414 , \21413 );
or \U$20745 ( \21415 , \21411 , \21414 );
or \U$20746 ( \21416 , \21413 , \21410 );
nand \U$20747 ( \21417 , \21415 , \21416 );
xor \U$20748 ( \21418 , \21405 , \21417 );
nand \U$20749 ( \21419 , \21399 , \21418 );
not \U$20750 ( \21420 , \21405 );
not \U$20751 ( \21421 , \21417 );
or \U$20752 ( \21422 , \21420 , \21421 );
not \U$20753 ( \21423 , \21413 );
nand \U$20754 ( \21424 , \21423 , \21410 );
nand \U$20755 ( \21425 , \21422 , \21424 );
xor \U$20756 ( \21426 , \21359 , \21382 );
xnor \U$20757 ( \21427 , \21426 , \21389 );
nand \U$20758 ( \21428 , \21425 , \21427 );
nand \U$20759 ( \21429 , \21419 , \21428 );
nor \U$20760 ( \21430 , \21394 , \21429 );
nand \U$20761 ( \21431 , \21349 , \21430 );
nor \U$20762 ( \21432 , \21275 , \21431 );
and \U$20763 ( \21433 , \20897 , \21432 );
not \U$20764 ( \21434 , \21231 );
nand \U$20765 ( \21435 , \21266 , \21272 );
or \U$20766 ( \21436 , \21260 , \21435 );
nand \U$20767 ( \21437 , \21238 , \21259 );
nand \U$20768 ( \21438 , \21436 , \21437 );
not \U$20769 ( \21439 , \21438 );
or \U$20770 ( \21440 , \21434 , \21439 );
not \U$20771 ( \21441 , \21230 );
not \U$20772 ( \21442 , \21228 );
or \U$20773 ( \21443 , \21441 , \21442 );
nand \U$20774 ( \21444 , \21443 , \21164 );
not \U$20775 ( \21445 , \21161 );
nand \U$20776 ( \21446 , \21445 , \21094 );
and \U$20777 ( \21447 , \21444 , \21446 );
nand \U$20778 ( \21448 , \21440 , \21447 );
buf \U$20779 ( \21449 , \21162 );
nand \U$20780 ( \21450 , \21448 , \21430 , \21449 );
not \U$20781 ( \21451 , \21428 );
nor \U$20782 ( \21452 , \21399 , \21418 );
not \U$20783 ( \21453 , \21452 );
or \U$20784 ( \21454 , \21451 , \21453 );
or \U$20785 ( \21455 , \21425 , \21427 );
nand \U$20786 ( \21456 , \21454 , \21455 );
nor \U$20787 ( \21457 , \21354 , \21392 );
or \U$20788 ( \21458 , \21456 , \21457 );
nand \U$20789 ( \21459 , \21458 , \21393 );
nand \U$20790 ( \21460 , \21342 , \21347 );
and \U$20791 ( \21461 , \21459 , \21460 );
and \U$20792 ( \21462 , \21450 , \21461 );
nor \U$20793 ( \21463 , \21462 , \21348 );
nor \U$20794 ( \21464 , \21433 , \21463 );
not \U$20795 ( \21465 , \21464 );
not \U$20796 ( \21466 , \21465 );
or \U$20797 ( \21467 , \17903 , \21466 );
not \U$20798 ( \21468 , \17896 );
nand \U$20799 ( \21469 , \21468 , \17898 );
nand \U$20800 ( \21470 , \21467 , \21469 );
not \U$20801 ( \21471 , \21470 );
or \U$20802 ( \21472 , \17826 , \21471 );
or \U$20803 ( \21473 , \21470 , \17825 );
nand \U$20804 ( \21474 , \21472 , \21473 );
not \U$20805 ( \21475 , \17471 );
nand \U$20806 ( \21476 , \21474 , \21475 );
nand \U$20807 ( \21477 , \17473 , \21476 );
buf \U$20808 ( \21478 , \21477 );
not \U$20809 ( \21479 , \16763 );
not \U$20810 ( \21480 , \21479 );
nand \U$20811 ( \21481 , \16784 , \12715 );
not \U$20812 ( \21482 , \21481 );
nand \U$20813 ( \21483 , \21482 , \17471 );
nor \U$20814 ( \21484 , \16779 , \21483 );
nand \U$20815 ( \21485 , \21480 , \21484 , \14371 );
and \U$20816 ( \21486 , \21481 , \17471 );
and \U$20817 ( \21487 , \21479 , \21486 );
not \U$20818 ( \21488 , \21486 );
not \U$20819 ( \21489 , \16779 );
or \U$20820 ( \21490 , \21488 , \21489 );
not \U$20821 ( \21491 , \17902 );
not \U$20822 ( \21492 , \21464 );
or \U$20823 ( \21493 , \21491 , \21492 );
or \U$20824 ( \21494 , \21464 , \17902 );
nand \U$20825 ( \21495 , \21493 , \21494 );
nand \U$20826 ( \21496 , \21495 , \17470 );
nand \U$20827 ( \21497 , \21490 , \21496 );
nor \U$20828 ( \21498 , \21487 , \21497 );
not \U$20829 ( \21499 , \14371 );
nand \U$20830 ( \21500 , \21499 , \21486 );
nand \U$20831 ( \21501 , \21485 , \21498 , \21500 );
buf \U$20832 ( \21502 , \21501 );
not \U$20833 ( \21503 , \16761 );
not \U$20834 ( \21504 , \16366 );
and \U$20835 ( \21505 , \16735 , \16173 , \16281 );
not \U$20836 ( \21506 , \21505 );
or \U$20837 ( \21507 , \21504 , \21506 );
not \U$20838 ( \21508 , \16276 );
nand \U$20839 ( \21509 , \21507 , \21508 );
nor \U$20840 ( \21510 , \15953 , \16738 );
and \U$20841 ( \21511 , \21510 , \15670 );
and \U$20842 ( \21512 , \21509 , \21511 );
not \U$20843 ( \21513 , \15824 );
nor \U$20844 ( \21514 , \21512 , \21513 );
not \U$20845 ( \21515 , \15875 );
or \U$20846 ( \21516 , \21514 , \21515 );
nand \U$20847 ( \21517 , \21516 , \15885 );
not \U$20848 ( \21518 , \15187 );
nand \U$20849 ( \21519 , \21518 , \14197 );
not \U$20850 ( \21520 , \15147 );
nand \U$20851 ( \21521 , \21520 , \16758 );
nor \U$20852 ( \21522 , \21519 , \21521 , \16757 );
and \U$20853 ( \21523 , \21517 , \21522 );
not \U$20854 ( \21524 , \16754 );
not \U$20855 ( \21525 , \16760 );
or \U$20856 ( \21526 , \21524 , \21525 );
nand \U$20857 ( \21527 , \21526 , \13467 );
nor \U$20858 ( \21528 , \21523 , \21527 );
nand \U$20859 ( \21529 , \21528 , \14225 );
not \U$20860 ( \21530 , \21529 );
or \U$20861 ( \21531 , \21503 , \21530 );
not \U$20862 ( \21532 , \16775 );
nand \U$20863 ( \21533 , \21531 , \21532 );
and \U$20864 ( \21534 , \16778 , \14369 );
nand \U$20865 ( \21535 , \21534 , \17471 );
or \U$20866 ( \21536 , \21533 , \21535 );
not \U$20867 ( \21537 , \21430 );
not \U$20868 ( \21538 , \20706 );
not \U$20869 ( \21539 , \20742 );
not \U$20870 ( \21540 , \20129 );
or \U$20871 ( \21541 , \21539 , \21540 );
not \U$20872 ( \21542 , \20755 );
nand \U$20873 ( \21543 , \21541 , \21542 );
not \U$20874 ( \21544 , \21543 );
or \U$20875 ( \21545 , \21538 , \21544 );
nand \U$20876 ( \21546 , \21545 , \20893 );
not \U$20877 ( \21547 , \21546 );
not \U$20878 ( \21548 , \20895 );
nor \U$20879 ( \21549 , \21548 , \21275 );
not \U$20880 ( \21550 , \21549 );
or \U$20881 ( \21551 , \21547 , \21550 );
nand \U$20882 ( \21552 , \21448 , \21449 );
nand \U$20883 ( \21553 , \21551 , \21552 );
not \U$20884 ( \21554 , \21553 );
or \U$20885 ( \21555 , \21537 , \21554 );
nand \U$20886 ( \21556 , \21555 , \21459 );
not \U$20887 ( \21557 , \21556 );
not \U$20888 ( \21558 , \21460 );
nor \U$20889 ( \21559 , \21558 , \21348 );
not \U$20890 ( \21560 , \17471 );
nand \U$20891 ( \21561 , \21559 , \21560 );
not \U$20892 ( \21562 , \21561 );
and \U$20893 ( \21563 , \21557 , \21562 );
nor \U$20894 ( \21564 , \21559 , \17471 );
and \U$20895 ( \21565 , \21556 , \21564 );
nor \U$20896 ( \21566 , \21563 , \21565 );
nor \U$20897 ( \21567 , \21534 , \17470 );
nand \U$20898 ( \21568 , \21533 , \21567 );
nand \U$20899 ( \21569 , \21536 , \21566 , \21568 );
buf \U$20900 ( \21570 , \21569 );
and \U$20901 ( \21571 , \14285 , \14355 );
not \U$20902 ( \21572 , \21571 );
not \U$20903 ( \21573 , \21529 );
or \U$20904 ( \21574 , \21572 , \21573 );
not \U$20905 ( \21575 , \16771 );
nand \U$20906 ( \21576 , \21574 , \21575 );
and \U$20907 ( \21577 , \14348 , \16774 );
buf \U$20908 ( \21578 , \17471 );
nand \U$20909 ( \21579 , \21577 , \21578 );
or \U$20910 ( \21580 , \21576 , \21579 );
not \U$20911 ( \21581 , \21429 );
not \U$20912 ( \21582 , \21581 );
not \U$20913 ( \21583 , \21553 );
or \U$20914 ( \21584 , \21582 , \21583 );
not \U$20915 ( \21585 , \21456 );
nand \U$20916 ( \21586 , \21584 , \21585 );
not \U$20917 ( \21587 , \21586 );
not \U$20918 ( \21588 , \21391 );
not \U$20919 ( \21589 , \21354 );
or \U$20920 ( \21590 , \21588 , \21589 );
or \U$20921 ( \21591 , \21354 , \21391 );
nand \U$20922 ( \21592 , \21590 , \21591 );
nand \U$20923 ( \21593 , \21592 , \21560 );
not \U$20924 ( \21594 , \21593 );
and \U$20925 ( \21595 , \21587 , \21594 );
nor \U$20926 ( \21596 , \21592 , \17471 );
and \U$20927 ( \21597 , \21586 , \21596 );
nor \U$20928 ( \21598 , \21595 , \21597 );
nor \U$20929 ( \21599 , \21577 , \17470 );
nand \U$20930 ( \21600 , \21576 , \21599 );
nand \U$20931 ( \21601 , \21580 , \21598 , \21600 );
buf \U$20932 ( \21602 , \21601 );
not \U$20933 ( \21603 , \14285 );
not \U$20934 ( \21604 , \21529 );
or \U$20935 ( \21605 , \21603 , \21604 );
buf \U$20936 ( \21606 , \16767 );
not \U$20937 ( \21607 , \21606 );
nand \U$20938 ( \21608 , \21605 , \21607 );
nand \U$20939 ( \21609 , \16770 , \14355 );
not \U$20940 ( \21610 , \21609 );
nand \U$20941 ( \21611 , \21610 , \17471 );
or \U$20942 ( \21612 , \21608 , \21611 );
not \U$20943 ( \21613 , \21419 );
not \U$20944 ( \21614 , \21553 );
or \U$20945 ( \21615 , \21613 , \21614 );
not \U$20946 ( \21616 , \21452 );
nand \U$20947 ( \21617 , \21615 , \21616 );
not \U$20948 ( \21618 , \21617 );
and \U$20949 ( \21619 , \21455 , \21428 );
nand \U$20950 ( \21620 , \21619 , \17470 );
not \U$20951 ( \21621 , \21620 );
and \U$20952 ( \21622 , \21618 , \21621 );
nor \U$20953 ( \21623 , \21619 , \21578 );
and \U$20954 ( \21624 , \21617 , \21623 );
nor \U$20955 ( \21625 , \21622 , \21624 );
and \U$20956 ( \21626 , \21609 , \17471 );
nand \U$20957 ( \21627 , \21608 , \21626 );
nand \U$20958 ( \21628 , \21612 , \21625 , \21627 );
buf \U$20959 ( \21629 , \21628 );
not \U$20960 ( \21630 , \21606 );
nand \U$20961 ( \21631 , \21630 , \14285 );
and \U$20962 ( \21632 , \21529 , \21631 );
not \U$20963 ( \21633 , \21529 );
not \U$20964 ( \21634 , \21631 );
and \U$20965 ( \21635 , \21633 , \21634 );
nor \U$20966 ( \21636 , \21632 , \21635 );
or \U$20967 ( \21637 , \21636 , \21475 );
not \U$20968 ( \21638 , \21553 );
nand \U$20969 ( \21639 , \21616 , \21419 );
not \U$20970 ( \21640 , \21639 );
and \U$20971 ( \21641 , \21638 , \21640 );
and \U$20972 ( \21642 , \21553 , \21639 );
nor \U$20973 ( \21643 , \21641 , \21642 );
or \U$20974 ( \21644 , \21643 , \17471 );
nand \U$20975 ( \21645 , \21637 , \21644 );
buf \U$20976 ( \21646 , \21645 );
not \U$20977 ( \21647 , \14218 );
not \U$20978 ( \21648 , \16759 );
not \U$20979 ( \21649 , \21648 );
not \U$20980 ( \21650 , \16756 );
or \U$20981 ( \21651 , \21649 , \21650 );
buf \U$20982 ( \21652 , \14198 );
nand \U$20983 ( \21653 , \21651 , \21652 );
not \U$20984 ( \21654 , \21653 );
or \U$20985 ( \21655 , \21647 , \21654 );
and \U$20986 ( \21656 , \14224 , \13467 );
and \U$20987 ( \21657 , \21656 , \14221 , \17471 );
nand \U$20988 ( \21658 , \21655 , \21657 );
nor \U$20989 ( \21659 , \21656 , \21560 );
nand \U$20990 ( \21660 , \21653 , \21659 , \14218 );
not \U$20991 ( \21661 , \21444 );
not \U$20992 ( \21662 , \20897 );
not \U$20993 ( \21663 , \21662 );
buf \U$20994 ( \21664 , \21274 );
and \U$20995 ( \21665 , \21663 , \21664 );
buf \U$20996 ( \21666 , \21438 );
nor \U$20997 ( \21667 , \21665 , \21666 );
not \U$20998 ( \21668 , \21667 );
buf \U$20999 ( \21669 , \21231 );
nand \U$21000 ( \21670 , \21668 , \21669 );
not \U$21001 ( \21671 , \21670 );
or \U$21002 ( \21672 , \21661 , \21671 );
nand \U$21003 ( \21673 , \21449 , \21446 );
and \U$21004 ( \21674 , \21673 , \21560 );
nand \U$21005 ( \21675 , \21672 , \21674 );
nor \U$21006 ( \21676 , \21673 , \17471 );
and \U$21007 ( \21677 , \21670 , \21676 , \21444 );
not \U$21008 ( \21678 , \14221 );
nand \U$21009 ( \21679 , \21678 , \17471 );
nor \U$21010 ( \21680 , \21656 , \21679 );
nor \U$21011 ( \21681 , \21677 , \21680 );
nand \U$21012 ( \21682 , \21658 , \21660 , \21675 , \21681 );
buf \U$21013 ( \21683 , \21682 );
not \U$21014 ( \21684 , \21653 );
not \U$21015 ( \21685 , \21678 );
nand \U$21016 ( \21686 , \21685 , \14218 );
not \U$21017 ( \21687 , \21686 );
and \U$21018 ( \21688 , \21684 , \21687 );
and \U$21019 ( \21689 , \21653 , \21686 );
nor \U$21020 ( \21690 , \21688 , \21689 );
and \U$21021 ( \21691 , \17471 , \21690 );
not \U$21022 ( \21692 , \17471 );
nand \U$21023 ( \21693 , \21669 , \21444 );
xnor \U$21024 ( \21694 , \21667 , \21693 );
and \U$21025 ( \21695 , \21692 , \21694 );
nor \U$21026 ( \21696 , \21691 , \21695 );
buf \U$21027 ( \21697 , \21696 );
buf \U$21028 ( \21698 , \21273 );
not \U$21029 ( \21699 , \21698 );
and \U$21030 ( \21700 , \21663 , \21699 );
not \U$21031 ( \21701 , \21435 );
nor \U$21032 ( \21702 , \21700 , \21701 );
not \U$21033 ( \21703 , \21260 );
nand \U$21034 ( \21704 , \21703 , \21437 );
xnor \U$21035 ( \21705 , \21702 , \21704 );
and \U$21036 ( \21706 , \17470 , \21705 );
not \U$21037 ( \21707 , \17470 );
not \U$21038 ( \21708 , \16758 );
not \U$21039 ( \21709 , \16756 );
or \U$21040 ( \21710 , \21708 , \21709 );
nand \U$21041 ( \21711 , \21710 , \14193 );
nand \U$21042 ( \21712 , \14197 , \13976 );
and \U$21043 ( \21713 , \21711 , \21712 );
not \U$21044 ( \21714 , \21711 );
not \U$21045 ( \21715 , \21712 );
and \U$21046 ( \21716 , \21714 , \21715 );
nor \U$21047 ( \21717 , \21713 , \21716 );
and \U$21048 ( \21718 , \21707 , \21717 );
nor \U$21049 ( \21719 , \21706 , \21718 );
buf \U$21050 ( \21720 , \21719 );
and \U$21051 ( \21721 , \16758 , \14193 );
xnor \U$21052 ( \21722 , \21721 , \16756 );
not \U$21053 ( \21723 , \21578 );
or \U$21054 ( \21724 , \21722 , \21723 );
not \U$21055 ( \21725 , \21698 );
nand \U$21056 ( \21726 , \21725 , \21435 );
xnor \U$21057 ( \21727 , \21662 , \21726 );
or \U$21058 ( \21728 , \21727 , \21578 );
nand \U$21059 ( \21729 , \21724 , \21728 );
buf \U$21060 ( \21730 , \21729 );
not \U$21061 ( \21731 , \21520 );
not \U$21062 ( \21732 , \16366 );
not \U$21063 ( \21733 , \21505 );
or \U$21064 ( \21734 , \21732 , \21733 );
nand \U$21065 ( \21735 , \21734 , \21508 );
nand \U$21066 ( \21736 , \21735 , \15875 , \21511 );
nand \U$21067 ( \21737 , \21736 , \15876 , \15885 );
not \U$21068 ( \21738 , \21737 );
or \U$21069 ( \21739 , \21731 , \21738 );
buf \U$21070 ( \21740 , \14919 );
and \U$21071 ( \21741 , \21740 , \16749 );
not \U$21072 ( \21742 , \16744 );
nor \U$21073 ( \21743 , \21741 , \21742 );
nand \U$21074 ( \21744 , \21739 , \21743 );
buf \U$21075 ( \21745 , \15177 );
and \U$21076 ( \21746 , \21744 , \21745 );
buf \U$21077 ( \21747 , \16743 );
not \U$21078 ( \21748 , \21747 );
nor \U$21079 ( \21749 , \21746 , \21748 );
not \U$21080 ( \21750 , \21749 );
and \U$21081 ( \21751 , \16752 , \15186 );
not \U$21082 ( \21752 , \21751 );
and \U$21083 ( \21753 , \21750 , \21752 );
and \U$21084 ( \21754 , \21749 , \21751 );
nor \U$21085 ( \21755 , \21753 , \21754 );
and \U$21086 ( \21756 , \17471 , \21755 );
not \U$21087 ( \21757 , \17471 );
and \U$21088 ( \21758 , \21543 , \20878 );
nor \U$21089 ( \21759 , \21758 , \20891 );
or \U$21090 ( \21760 , \21759 , \20614 );
buf \U$21091 ( \21761 , \20884 );
nand \U$21092 ( \21762 , \21760 , \21761 );
not \U$21093 ( \21763 , \21762 );
not \U$21094 ( \21764 , \20760 );
not \U$21095 ( \21765 , \20874 );
or \U$21096 ( \21766 , \21764 , \21765 );
nand \U$21097 ( \21767 , \21766 , \20895 );
not \U$21098 ( \21768 , \21767 );
and \U$21099 ( \21769 , \21763 , \21768 );
and \U$21100 ( \21770 , \21762 , \21767 );
nor \U$21101 ( \21771 , \21769 , \21770 );
and \U$21102 ( \21772 , \21757 , \21771 );
nor \U$21103 ( \21773 , \21756 , \21772 );
buf \U$21104 ( \21774 , \21773 );
nand \U$21105 ( \21775 , \21747 , \21745 );
and \U$21106 ( \21776 , \21744 , \21775 );
not \U$21107 ( \21777 , \21744 );
not \U$21108 ( \21778 , \21775 );
and \U$21109 ( \21779 , \21777 , \21778 );
nor \U$21110 ( \21780 , \21776 , \21779 );
and \U$21111 ( \21781 , \17471 , \21780 );
not \U$21112 ( \21782 , \17471 );
not \U$21113 ( \21783 , \20614 );
nand \U$21114 ( \21784 , \21783 , \21761 );
xnor \U$21115 ( \21785 , \21759 , \21784 );
and \U$21116 ( \21786 , \21782 , \21785 );
nor \U$21117 ( \21787 , \21781 , \21786 );
buf \U$21118 ( \21788 , \21787 );
buf \U$21119 ( \21789 , \15146 );
not \U$21120 ( \21790 , \21789 );
not \U$21121 ( \21791 , \21737 );
or \U$21122 ( \21792 , \21790 , \21791 );
not \U$21123 ( \21793 , \16749 );
nand \U$21124 ( \21794 , \21792 , \21793 );
nand \U$21125 ( \21795 , \21740 , \16744 );
and \U$21126 ( \21796 , \21794 , \21795 );
not \U$21127 ( \21797 , \21794 );
not \U$21128 ( \21798 , \21795 );
and \U$21129 ( \21799 , \21797 , \21798 );
nor \U$21130 ( \21800 , \21796 , \21799 );
or \U$21131 ( \21801 , \21800 , \21723 );
not \U$21132 ( \21802 , \20704 );
not \U$21133 ( \21803 , \21543 );
or \U$21134 ( \21804 , \21802 , \21803 );
nand \U$21135 ( \21805 , \21804 , \20888 );
not \U$21136 ( \21806 , \21805 );
not \U$21137 ( \21807 , \20886 );
nand \U$21138 ( \21808 , \21807 , \20890 );
not \U$21139 ( \21809 , \21808 );
and \U$21140 ( \21810 , \21806 , \21809 );
and \U$21141 ( \21811 , \21805 , \21808 );
nor \U$21142 ( \21812 , \21810 , \21811 );
or \U$21143 ( \21813 , \21812 , \17471 );
nand \U$21144 ( \21814 , \21801 , \21813 );
buf \U$21145 ( \21815 , \21814 );
nand \U$21146 ( \21816 , \21789 , \21793 );
and \U$21147 ( \21817 , \21737 , \21816 );
not \U$21148 ( \21818 , \21737 );
not \U$21149 ( \21819 , \21816 );
and \U$21150 ( \21820 , \21818 , \21819 );
nor \U$21151 ( \21821 , \21817 , \21820 );
or \U$21152 ( \21822 , \21821 , \17470 );
not \U$21153 ( \21823 , \21543 );
nand \U$21154 ( \21824 , \20704 , \20888 );
not \U$21155 ( \21825 , \21824 );
and \U$21156 ( \21826 , \21823 , \21825 );
and \U$21157 ( \21827 , \21543 , \21824 );
nor \U$21158 ( \21828 , \21826 , \21827 );
or \U$21159 ( \21829 , \21828 , \21578 );
nand \U$21160 ( \21830 , \21822 , \21829 );
buf \U$21161 ( \21831 , \21830 );
not \U$21162 ( \21832 , \15857 );
not \U$21163 ( \21833 , \16740 );
not \U$21164 ( \21834 , \21833 );
not \U$21165 ( \21835 , \16737 );
or \U$21166 ( \21836 , \21834 , \21835 );
not \U$21167 ( \21837 , \21513 );
nand \U$21168 ( \21838 , \21836 , \21837 );
not \U$21169 ( \21839 , \21838 );
or \U$21170 ( \21840 , \21832 , \21839 );
buf \U$21171 ( \21841 , \15880 );
nand \U$21172 ( \21842 , \21840 , \21841 );
not \U$21173 ( \21843 , \21842 );
not \U$21174 ( \21844 , \15877 );
nand \U$21175 ( \21845 , \21844 , \15883 );
not \U$21176 ( \21846 , \21845 );
and \U$21177 ( \21847 , \21843 , \21846 );
and \U$21178 ( \21848 , \21842 , \21845 );
nor \U$21179 ( \21849 , \21847 , \21848 );
and \U$21180 ( \21850 , \21578 , \21849 );
not \U$21181 ( \21851 , \21578 );
buf \U$21182 ( \21852 , \20129 );
not \U$21183 ( \21853 , \20749 );
nor \U$21184 ( \21854 , \21852 , \21853 );
not \U$21185 ( \21855 , \21854 );
and \U$21186 ( \21856 , \21855 , \20731 );
nor \U$21187 ( \21857 , \21856 , \20751 );
not \U$21188 ( \21858 , \21857 );
not \U$21189 ( \21859 , \20740 );
nor \U$21190 ( \21860 , \21859 , \20753 );
not \U$21191 ( \21861 , \21860 );
and \U$21192 ( \21862 , \21858 , \21861 );
and \U$21193 ( \21863 , \21857 , \21860 );
nor \U$21194 ( \21864 , \21862 , \21863 );
and \U$21195 ( \21865 , \21851 , \21864 );
nor \U$21196 ( \21866 , \21850 , \21865 );
buf \U$21197 ( \21867 , \21866 );
nand \U$21198 ( \21868 , \15857 , \21841 );
xor \U$21199 ( \21869 , \21838 , \21868 );
and \U$21200 ( \21870 , \21578 , \21869 );
not \U$21201 ( \21871 , \21578 );
xnor \U$21202 ( \21872 , \20720 , \20730 );
xnor \U$21203 ( \21873 , \21854 , \21872 );
and \U$21204 ( \21874 , \21871 , \21873 );
nor \U$21205 ( \21875 , \21870 , \21874 );
buf \U$21206 ( \21876 , \21875 );
not \U$21207 ( \21877 , \16739 );
not \U$21208 ( \21878 , \16737 );
or \U$21209 ( \21879 , \21877 , \21878 );
nand \U$21210 ( \21880 , \21879 , \15822 );
not \U$21211 ( \21881 , \21880 );
nor \U$21212 ( \21882 , \15423 , \15669 );
not \U$21213 ( \21883 , \21882 );
nand \U$21214 ( \21884 , \21883 , \15670 );
not \U$21215 ( \21885 , \21884 );
and \U$21216 ( \21886 , \21881 , \21885 );
and \U$21217 ( \21887 , \21880 , \21884 );
nor \U$21218 ( \21888 , \21886 , \21887 );
and \U$21219 ( \21889 , \21578 , \21888 );
not \U$21220 ( \21890 , \21578 );
nand \U$21221 ( \21891 , \19976 , \20746 );
nand \U$21222 ( \21892 , \20744 , \20127 );
xor \U$21223 ( \21893 , \21891 , \21892 );
and \U$21224 ( \21894 , \21890 , \21893 );
nor \U$21225 ( \21895 , \21889 , \21894 );
buf \U$21226 ( \21896 , \21895 );
nand \U$21227 ( \21897 , \16739 , \15822 );
xor \U$21228 ( \21898 , \16737 , \21897 );
or \U$21229 ( \21899 , \21898 , \17470 );
not \U$21230 ( \21900 , \19066 );
and \U$21231 ( \21901 , \21900 , \19064 );
nand \U$21232 ( \21902 , \19824 , \21901 );
buf \U$21233 ( \21903 , \19254 );
nor \U$21234 ( \21904 , \21902 , \21903 );
or \U$21235 ( \21905 , \21904 , \19833 );
nand \U$21236 ( \21906 , \21905 , \19834 );
not \U$21237 ( \21907 , \19974 );
nand \U$21238 ( \21908 , \21907 , \20746 );
xor \U$21239 ( \21909 , \21906 , \21908 );
or \U$21240 ( \21910 , \21909 , \17471 );
nand \U$21241 ( \21911 , \21899 , \21910 );
buf \U$21242 ( \21912 , \21911 );
buf \U$21243 ( \21913 , \16270 );
not \U$21244 ( \21914 , \21913 );
not \U$21245 ( \21915 , \16365 );
not \U$21246 ( \21916 , \16425 );
not \U$21247 ( \21917 , \16731 );
or \U$21248 ( \21918 , \21916 , \21917 );
nand \U$21249 ( \21919 , \21918 , \16734 );
not \U$21250 ( \21920 , \21919 );
or \U$21251 ( \21921 , \21915 , \21920 );
nand \U$21252 ( \21922 , \21921 , \16733 );
not \U$21253 ( \21923 , \21922 );
not \U$21254 ( \21924 , \16282 );
or \U$21255 ( \21925 , \21923 , \21924 );
nand \U$21256 ( \21926 , \21925 , \16256 );
not \U$21257 ( \21927 , \21926 );
or \U$21258 ( \21928 , \21914 , \21927 );
not \U$21259 ( \21929 , \16274 );
nand \U$21260 ( \21930 , \21928 , \21929 );
not \U$21261 ( \21931 , \15952 );
not \U$21262 ( \21932 , \15893 );
or \U$21263 ( \21933 , \21931 , \21932 );
nand \U$21264 ( \21934 , \21933 , \15954 );
and \U$21265 ( \21935 , \21930 , \21934 );
not \U$21266 ( \21936 , \21930 );
not \U$21267 ( \21937 , \21934 );
and \U$21268 ( \21938 , \21936 , \21937 );
nor \U$21269 ( \21939 , \21935 , \21938 );
and \U$21270 ( \21940 , \17471 , \21939 );
not \U$21271 ( \21941 , \17471 );
not \U$21272 ( \21942 , \19832 );
not \U$21273 ( \21943 , \21902 );
or \U$21274 ( \21944 , \21942 , \21943 );
not \U$21275 ( \21945 , \21903 );
nand \U$21276 ( \21946 , \21944 , \21945 );
not \U$21277 ( \21947 , \21946 );
not \U$21278 ( \21948 , \19829 );
nor \U$21279 ( \21949 , \21948 , \19415 );
not \U$21280 ( \21950 , \21949 );
nand \U$21281 ( \21951 , \21950 , \19834 );
not \U$21282 ( \21952 , \21951 );
and \U$21283 ( \21953 , \21947 , \21952 );
and \U$21284 ( \21954 , \21946 , \21951 );
nor \U$21285 ( \21955 , \21953 , \21954 );
and \U$21286 ( \21956 , \21941 , \21955 );
nor \U$21287 ( \21957 , \21940 , \21956 );
buf \U$21288 ( \21958 , \21957 );
not \U$21289 ( \21959 , \21902 );
not \U$21290 ( \21960 , \21959 );
not \U$21291 ( \21961 , \19832 );
nor \U$21292 ( \21962 , \21961 , \21903 );
not \U$21293 ( \21963 , \21962 );
and \U$21294 ( \21964 , \21960 , \21963 );
and \U$21295 ( \21965 , \21904 , \19832 );
nor \U$21296 ( \21966 , \21964 , \21965 );
and \U$21297 ( \21967 , \17470 , \21966 );
not \U$21298 ( \21968 , \17470 );
not \U$21299 ( \21969 , \16274 );
nand \U$21300 ( \21970 , \21969 , \21913 );
and \U$21301 ( \21971 , \21926 , \21970 );
not \U$21302 ( \21972 , \21926 );
not \U$21303 ( \21973 , \21970 );
and \U$21304 ( \21974 , \21972 , \21973 );
nor \U$21305 ( \21975 , \21971 , \21974 );
and \U$21306 ( \21976 , \21968 , \21975 );
nor \U$21307 ( \21977 , \21967 , \21976 );
buf \U$21308 ( \21978 , \21977 );
not \U$21309 ( \21979 , \21922 );
not \U$21310 ( \21980 , \16281 );
or \U$21311 ( \21981 , \21979 , \21980 );
buf \U$21312 ( \21982 , \16254 );
nand \U$21313 ( \21983 , \21981 , \21982 );
not \U$21314 ( \21984 , \21983 );
nor \U$21315 ( \21985 , \16070 , \16172 );
not \U$21316 ( \21986 , \21985 );
nand \U$21317 ( \21987 , \21986 , \16173 );
not \U$21318 ( \21988 , \21987 );
and \U$21319 ( \21989 , \21984 , \21988 );
and \U$21320 ( \21990 , \21983 , \21987 );
nor \U$21321 ( \21991 , \21989 , \21990 );
or \U$21322 ( \21992 , \21991 , \17470 );
buf \U$21323 ( \21993 , \19820 );
or \U$21324 ( \21994 , \21993 , \19063 );
nand \U$21325 ( \21995 , \18998 , \19062 );
nand \U$21326 ( \21996 , \21994 , \21995 );
and \U$21327 ( \21997 , \21900 , \18996 );
xor \U$21328 ( \21998 , \21996 , \21997 );
or \U$21329 ( \21999 , \21998 , \17471 );
nand \U$21330 ( \22000 , \21992 , \21999 );
buf \U$21331 ( \22001 , \22000 );
nand \U$21332 ( \22002 , \16281 , \16254 );
xnor \U$21333 ( \22003 , \21979 , \22002 );
and \U$21334 ( \22004 , \17471 , \22003 );
not \U$21335 ( \22005 , \17471 );
not \U$21336 ( \22006 , \21993 );
not \U$21337 ( \22007 , \19063 );
nand \U$21338 ( \22008 , \22007 , \21995 );
not \U$21339 ( \22009 , \22008 );
and \U$21340 ( \22010 , \22006 , \22009 );
and \U$21341 ( \22011 , \21993 , \22008 );
nor \U$21342 ( \22012 , \22010 , \22011 );
and \U$21343 ( \22013 , \22005 , \22012 );
nor \U$21344 ( \22014 , \22004 , \22013 );
buf \U$21345 ( \22015 , \22014 );
buf \U$21346 ( \22016 , \19805 );
not \U$21347 ( \22017 , \22016 );
not \U$21348 ( \22018 , \19816 );
not \U$21349 ( \22019 , \22018 );
and \U$21350 ( \22020 , \22017 , \22019 );
and \U$21351 ( \22021 , \22016 , \22018 );
nor \U$21352 ( \22022 , \22020 , \22021 );
and \U$21353 ( \22023 , \17470 , \22022 );
not \U$21354 ( \22024 , \17470 );
nand \U$21355 ( \22025 , \16365 , \16733 );
xor \U$21356 ( \22026 , \21919 , \22025 );
and \U$21357 ( \22027 , \22024 , \22026 );
nor \U$21358 ( \22028 , \22023 , \22027 );
buf \U$21359 ( \22029 , \22028 );
nand \U$21360 ( \22030 , \16734 , \16425 );
xor \U$21361 ( \22031 , \22030 , \16731 );
or \U$21362 ( \22032 , \22031 , \17470 );
xnor \U$21363 ( \22033 , \19802 , \19539 );
or \U$21364 ( \22034 , \22033 , \17469 );
nand \U$21365 ( \22035 , \22032 , \22034 );
buf \U$21366 ( \22036 , \22035 );
xnor \U$21367 ( \22037 , \16726 , \16706 );
and \U$21368 ( \22038 , \17469 , \22037 );
not \U$21369 ( \22039 , \17469 );
xnor \U$21370 ( \22040 , \19798 , \19584 );
and \U$21371 ( \22041 , \22039 , \22040 );
nor \U$21372 ( \22042 , \22038 , \22041 );
buf \U$21373 ( \22043 , \22042 );
not \U$21374 ( \22044 , \19797 );
nand \U$21375 ( \22045 , \22044 , \19795 );
xor \U$21376 ( \22046 , \22045 , \19788 );
and \U$21377 ( \22047 , \17468 , \22046 );
not \U$21378 ( \22048 , \17468 );
nand \U$21379 ( \22049 , \16519 , \16705 );
xor \U$21380 ( \22050 , \22049 , \16700 );
and \U$21381 ( \22051 , \22048 , \22050 );
nor \U$21382 ( \22052 , \22047 , \22051 );
buf \U$21383 ( \22053 , \22052 );
and \U$21384 ( \22054 , \16528 , \16565 );
not \U$21385 ( \22055 , \16528 );
and \U$21386 ( \22056 , \22055 , \16564 );
nor \U$21387 ( \22057 , \22054 , \22056 );
xnor \U$21388 ( \22058 , \16698 , \22057 );
or \U$21389 ( \22059 , \22058 , \17468 );
not \U$21390 ( \22060 , \19670 );
nand \U$21391 ( \22061 , \22060 , \19787 );
xnor \U$21392 ( \22062 , \22061 , \19785 );
or \U$21393 ( \22063 , \22062 , \17467 );
nand \U$21394 ( \22064 , \22059 , \22063 );
buf \U$21395 ( \22065 , \22064 );
endmodule

