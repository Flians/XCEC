//
// Conformal-LEC Version 20.10-d214 (03-Sep-2020)
//
module top(RIaa97c98_14,RIaa9e7f0_243,RIaa9e868_244,RIaa9e778_242,RIaa9e9d0_247,RIaa97d88_16,RIaa97d10_15,RIaa97e00_17,RIaa97c20_13,
        RIaa9e688_240,RIaa9e700_241,RIaa9e8e0_245,RIaa9e958_246,RIaa9cf90_191,RIaa9d170_195,RIaa9cea0_189,RIaa9d1e8_196,RIaa9d080_193,RIaa9d0f8_194,
        RIaa9d5a8_204,RIaa9d620_205,RIaa9d2d8_198,RIaa9d008_192,RIaa9d3c8_200,RIaa9d4b8_202,RIaa9d260_197,RIaa9d350_199,RIaa9cf18_190,RIaa9d530_203,
        RIaa9d440_201,RIaa97860_5,RIaa976f8_2,RIaa97770_3,RIaa977e8_4,RIaa9ba00_145,RIaa9b640_137,RIaa9b910_143,RIaa9bd48_152,RIaa9ba78_146,
        RIaa9bb68_148,RIaa9b7a8_140,RIaa9bdc0_153,RIaa9baf0_147,RIaa9b730_139,RIaa9bc58_150,RIaa9b6b8_138,RIaa9b898_142,RIaa9bcd0_151,RIaa9b988_144,
        RIaa9b820_141,RIaa9bbe0_149,RIaa9b370_131,RIaa9b0a0_125,RIaa9b5c8_136,RIaa9b3e8_132,RIaa9ae48_120,RIaa9b460_133,RIaa9b190_127,RIaa9b118_126,
        RIaa9b4d8_134,RIaa9b280_129,RIaa9b028_124,RIaa9af38_122,RIaa9b2f8_130,RIaa9aec0_121,RIaa9b550_135,RIaa9afb0_123,RIaa9b208_128,RIaa9c2e8_164,
        RIaa9c4c8_168,RIaa9c018_158,RIaa9c3d8_166,RIaa9c450_167,RIaa9be38_154,RIaa9bfa0_157,RIaa9beb0_155,RIaa9c270_163,RIaa9c090_159,RIaa9c108_160,
        RIaa9c180_161,RIaa9bf28_156,RIaa9c5b8_170,RIaa9c1f8_162,RIaa9c360_165,RIaa9c540_169,RIaa9ce28_188,RIaa9c978_178,RIaa9c9f0_179,RIaa9c900_177,
        RIaa9cdb0_187,RIaa9c810_175,RIaa9c720_173,RIaa9cb58_182,RIaa9cae0_181,RIaa9c630_171,RIaa9ca68_180,RIaa9cc48_184,RIaa9ccc0_185,RIaa9c888_176,
        RIaa9c6a8_172,RIaa9c798_174,RIaa9cbd0_183,RIaa9cd38_186,RIaa9ab78_114,RIaa9aa10_111,RIaa9ac68_116,RIaa9a7b8_106,RIaa9a6c8_104,RIaa9add0_119,
        RIaa9abf0_115,RIaa9a8a8_108,RIaa9a998_110,RIaa9a920_109,RIaa9a830_107,RIaa9ad58_118,RIaa9a740_105,RIaa9ab00_113,RIaa9aa88_112,RIaa9a650_103,
        RIaa9ace0_117,RIaa978d8_6,RIaa9a308_96,RIaa9a218_94,RIaa9a380_97,RIaa9a038_90,RIaa99ed0_87,RIaa9a290_95,RIaa9a0b0_91,RIaa99fc0_89,
        RIaa9a470_99,RIaa99f48_88,RIaa9a4e8_100,RIaa9a1a0_93,RIaa9a3f8_98,RIaa99e58_86,RIaa9a560_101,RIaa9a128_92,RIaa9a5d8_102,RIaa97950_7,
        RIaa99b10_79,RIaa999a8_76,RIaa99a20_77,RIaa996d8_70,RIaa99930_75,RIaa99d68_84,RIaa99b88_80,RIaa99660_69,RIaa99cf0_83,RIaa99c00_81,
        RIaa998b8_74,RIaa99de0_85,RIaa99a98_78,RIaa99c78_82,RIaa997c8_72,RIaa99840_73,RIaa99750_71,RIaa979c8_8,RIaa9f6f0_275,RIaa9f768_276,
        RIaa9f3a8_268,RIaa9f600_273,RIaa9f2b8_266,RIaa9f330_267,RIaa9f420_269,RIaa9f9c0_281,RIaa9f948_280,RIaa9f678_274,RIaa9f8d0_279,RIaa9f588_272,
        RIaa9f240_265,RIaa9f510_271,RIaa9f7e0_277,RIaa9f858_278,RIaa9f498_270,RIaa9eca0_253,RIaa9ee08_256,RIaa9eef8_258,RIaa9ed90_255,RIaa9f1c8_264,
        RIaa9efe8_260,RIaa9ef70_259,RIaa9ed18_254,RIaa9eb38_250,RIaa9ebb0_251,RIaa9ea48_248,RIaa9f0d8_262,RIaa9ee80_257,RIaa9eac0_249,RIaa9f150_263,
        RIaa9f060_261,RIaa9ec28_252,RIaa97b30_11,RIaa97ba8_12,RIaa9de18_222,RIaa9db48_216,RIaa9d968_212,RIaa9dbc0_217,RIaa9dda0_221,RIaa9dd28_220,
        RIaa9dad0_215,RIaa9d800_209,RIaa9dc38_218,RIaa9d710_207,RIaa9dcb0_219,RIaa9d788_208,RIaa9d698_206,RIaa9da58_214,RIaa9d9e0_213,RIaa9d878_210,
        RIaa9d8f0_211,RIaa994f8_66,RIaa99048_56,RIaa98f58_54,RIaa99570_67,RIaa990c0_57,RIaa99138_58,RIaa99390_63,RIaa98ee0_53,RIaa99480_65,
        RIaa98fd0_55,RIaa995e8_68,RIaa99318_62,RIaa991b0_59,RIaa99408_64,RIaa992a0_61,RIaa98e68_52,RIaa99228_60,RIaa9e160_229,RIaa9df80_225,
        RIaa9e3b8_234,RIaa9de90_223,RIaa9e610_239,RIaa9e2c8_232,RIaa9e598_238,RIaa9e1d8_230,RIaa9df08_224,RIaa9e520_237,RIaa9e340_233,RIaa9e250_231,
        RIaa9e430_235,RIaa9e0e8_228,RIaa9dff8_226,RIaa9e4a8_236,RIaa9e070_227,RIaa97ab8_10,RIaa97a40_9,RIaa98b20_45,RIaa989b8_42,RIaa98c88_48,
        RIaa98a30_43,RIaa98aa8_44,RIaa98df0_51,RIaa98940_41,RIaa98c10_47,RIaa98670_35,RIaa98850_39,RIaa98760_37,RIaa986e8_36,RIaa98d00_49,
        RIaa98b98_46,RIaa987d8_38,RIaa988c8_40,RIaa98d78_50,RIaaa1ce8_356,RIaaa1e50_359,RIaaa2030_363,RIaaa1fb8_362,RIaaa1f40_361,RIaaa1c70_355,
        RIaaa1d60_357,RIaaa1ec8_360,RIaaa1b80_353,RIaaa1bf8_354,RIaaa20a8_364,RIaaa1a90_351,RIaaa2120_365,RIaaa1dd8_358,RIaaa2198_366,RIaaa1b08_352,
        RIaaa1a18_350,RIaaa1130_331,RIaaa0f50_327,RIaaa0a28_316,RIaaa0b90_319,RIaaa0b18_318,RIaaa1040_329,RIaaa0c80_321,RIaaa0cf8_322,RIaaa0c08_320,
        RIaaa0ed8_326,RIaaa0d70_323,RIaaa0aa0_317,RIaaa0fc8_328,RIaaa11a8_332,RIaaa10b8_330,RIaaa0e60_325,RIaaa0de8_324,RIaa97680_1,RIaa98508_32,
        RIaa98328_28,RIaa98238_26,RIaa98418_30,RIaa97e78_18,RIaa981c0_25,RIaa985f8_34,RIaa982b0_27,RIaa98580_33,RIaa97ef0_19,RIaa98058_22,
        RIaa98148_24,RIaa97f68_20,RIaa97fe0_21,RIaa983a0_29,RIaa980d0_23,RIaa98490_31,RIaaa2cd8_390,RIaaa2af8_386,RIaaa3110_399,RIaaa3188_400,
        RIaaa2f30_395,RIaaa2c60_389,RIaaa2eb8_394,RIaaa2dc8_392,RIaaa2e40_393,RIaaa2fa8_396,RIaaa3020_397,RIaaa2a08_384,RIaaa3098_398,RIaaa2be8_388,
        RIaaa2b70_387,RIaaa2a80_385,RIaaa2d50_391,RIaaa1298_334,RIaaa16d0_343,RIaaa1928_348,RIaaa1658_342,RIaaa1838_346,RIaaa14f0_339,RIaaa1388_336,
        RIaaa1400_337,RIaaa19a0_349,RIaaa1748_344,RIaaa15e0_341,RIaaa1310_335,RIaaa1220_333,RIaaa1478_338,RIaaa1568_340,RIaaa17c0_345,RIaaa18b0_347,
        RIaa9ff60_293,RIaa9fba0_285,RIaa9fa38_282,RIaaa0050_295,RIaa9ffd8_294,RIaa9fe70_291,RIaa9fc90_287,RIaaa01b8_298,RIaaa0140_297,RIaa9fdf8_290,
        RIaa9fab0_283,RIaa9fc18_286,RIaa9fb28_284,RIaa9fd08_288,RIaaa00c8_296,RIaa9fee8_292,RIaa9fd80_289,RIaaa05f0_307,RIaaa0938_314,RIaaa0758_310,
        RIaaa0488_304,RIaaa0578_306,RIaaa0230_299,RIaaa06e0_309,RIaaa0848_312,RIaaa0398_302,RIaaa0320_301,RIaaa0668_308,RIaaa0410_303,RIaaa02a8_300,
        RIaaa08c0_313,RIaaa0500_305,RIaaa07d0_311,RIaaa09b0_315,RIaaa24e0_373,RIaaa2558_374,RIaaa2738_378,RIaaa2828_380,RIaaa2300_369,RIaaa26c0_377,
        RIaaa2918_382,RIaaa2468_372,RIaaa2378_370,RIaaa2288_368,RIaaa2648_376,RIaaa23f0_371,RIaaa2210_367,RIaaa25d0_375,RIaaa27b0_379,RIaaa28a0_381,
        RIaaa2990_383,RIaaa3f20_429,RIaaa3f98_430,RIaaa3cc8_424,RIaaa3c50_423,RIaaa4010_431,RIaaa4100_433,RIaaa3db8_426,RIaaa3b60_421,RIaaa3d40_425,
        RIaaa3ae8_420,RIaaa3a70_419,RIaaa39f8_418,RIaaa4178_434,RIaaa3e30_427,RIaaa3bd8_422,RIaaa4088_432,RIaaa3ea8_428,RIaaa32f0_403,RIaaa3890_415,
        RIaaa34d0_407,RIaaa3638_410,RIaaa3728_412,RIaaa35c0_409,RIaaa3278_402,RIaaa3818_414,RIaaa33e0_405,RIaaa3368_404,RIaaa37a0_413,RIaaa3980_417,
        RIaaa3908_416,RIaaa36b0_411,RIaaa3458_406,RIaaa3548_408,RIaaa3200_401,RIaaa4448_440,RIaaa4538_442,RIaaa4268_436,RIaaa43d0_439,RIaaa42e0_437,
        RIaaa41f0_435,RIaaa4628_444,RIaaa4808_448,RIaaa45b0_443,RIaaa4718_446,RIaaa44c0_441,RIaaa48f8_450,RIaaa4358_438,RIaaa4970_451,RIaaa4880_449,
        RIaaa4790_447,RIaaa46a0_445,RIaaa6248_504,RIaaa66f8_514,RIaaa6860_517,RIaaa67e8_516,RIaaa6680_513,RIaaa64a0_509,RIaaa6338_506,RIaaa63b0_507,
        RIaaa6950_519,RIaaa6608_512,RIaaa6590_511,RIaaa6428_508,RIaaa6770_515,RIaaa68d8_518,RIaaa6518_510,RIaaa62c0_505,RIaaa61d0_503,RIaaa57f8_482,
        RIaaa54b0_475,RIaaa5618_478,RIaaa52d0_471,RIaaa5528_476,RIaaa5258_470,RIaaa5708_480,RIaaa5690_479,RIaaa5348_472,RIaaa53c0_473,RIaaa58e8_484,
        RIaaa5960_485,RIaaa5780_481,RIaaa5438_474,RIaaa5870_483,RIaaa55a0_477,RIaaa51e0_469,RIaaa4e98_462,RIaaa49e8_452,RIaaa4b50_455,RIaaa4e20_461,
        RIaaa50f0_467,RIaaa4f88_464,RIaaa5000_465,RIaaa4c40_457,RIaaa4cb8_458,RIaaa4a60_453,RIaaa4f10_463,RIaaa4bc8_456,RIaaa4ad8_454,RIaaa5168_468,
        RIaaa4d30_459,RIaaa4da8_460,RIaaa5078_466,RIaaa5e10_495,RIaaa5ca8_492,RIaaa59d8_486,RIaaa60e0_501,RIaaa5b40_489,RIaaa5a50_487,RIaaa5f00_497,
        RIaaa5bb8_490,RIaaa6158_502,RIaaa5f78_498,RIaaa5ac8_488,RIaaa5e88_496,RIaaa5d98_494,RIaaa5ff0_499,RIaaa5d20_493,RIaaa6068_500,RIaaa5c30_491,
        RIaaa6d10_527,RIaaa6a40_521,RIaaa7058_534,RIaaa7148_536,RIaaa6e00_529,RIaaa6ba8_524,RIaaa6e78_530,RIaaa6c98_526,RIaaa6f68_532,RIaaa6ab8_522,
        RIaaa70d0_535,RIaaa6c20_525,RIaaa69c8_520,RIaaa6d88_528,RIaaa6fe0_533,RIaaa6ef0_531,RIaaa6b30_523,RIaaa8408_576,RIaaa87c8_584,RIaaa84f8_578,
        RIaaa8390_575,RIaaa8318_574,RIaaa8660_581,RIaaa8228_572,RIaaa88b8_586,RIaaa8930_587,RIaaa8750_583,RIaaa8480_577,RIaaa8840_585,RIaaa86d8_582,
        RIaaa85e8_580,RIaaa8570_579,RIaaa82a0_573,RIaaa81b0_571,RIaaa7670_547,RIaaa7238_538,RIaaa7490_543,RIaaa75f8_546,RIaaa78c8_552,RIaaa7328_540,
        RIaaa73a0_541,RIaaa77d8_550,RIaaa7850_551,RIaaa76e8_548,RIaaa7580_545,RIaaa72b0_539,RIaaa71c0_537,RIaaa7508_544,RIaaa7418_542,RIaaa7940_553,
        RIaaa7760_549,RIaaa7d00_561,RIaaa7f58_566,RIaaa7fd0_567,RIaaa7b98_558,RIaaa7b20_557,RIaaa7df0_563,RIaaa7c88_560,RIaaa7e68_564,RIaaa7ee0_565,
        RIaaa7d78_562,RIaaa8048_568,RIaaa7c10_559,RIaaa8138_570,RIaaa80c0_569,RIaaa7aa8_556,RIaaa7a30_555,RIaaa79b8_554,RIaaa89a8_588,RIaaa95d8_614,
        RIaaa9218_606,RIaaa90b0_603,RIaaa9128_604,RIaaa91a0_605,RIaaa9380_609,RIaaa9308_608,RIaaa9290_607,RIaaa9038_602,RIaaa93f8_610,RIaaa9470_611,
        RIaaa94e8_612,RIaaa8c78_594,RIaaa8cf0_595,RIaaa8a98_590,RIaaa8b10_591,RIaaa8a20_589,RIaaa8b88_592,RIaaa8c00_593,RIaaa8d68_596,RIaaa8de0_597,
        RIaaa8e58_598,RIaaa8ed0_599,RIaaa8f48_600,RIaaa8fc0_601,RIaaa9560_613,R_267_b0ecd58,R_268_b0ece00,R_269_b0ecea8,R_26a_b0ecf50,R_26b_b0ecff8,
        R_26c_b0ed0a0,R_26d_b0ed148,R_26e_b0ed1f0,R_26f_b0ed298,R_270_b0ed340,R_271_b0ed3e8,R_272_b0ed490,R_273_b0ed538,R_274_b0ed5e0,R_275_b0ed688,
        R_276_b0ed730,R_277_b0ed7d8,R_278_b0ed880,R_279_b0ed928,R_27a_b0ed9d0,R_27b_b0eda78,R_27c_b0edb20,R_27d_b0edbc8,R_27e_b0edc70,R_27f_b0edd18,
        R_280_b0eddc0,R_281_b0ede68,R_282_b0edf10,R_283_b0edfb8,R_284_b0ee060,R_285_b0ee108,R_286_b0ee1b0,R_287_b0ee258,R_288_b0ee300,R_289_b0ee3a8,
        R_28a_b0ee450,R_28b_b0ee4f8,R_28c_b0ee5a0,R_28d_b0ee648,R_28e_b0ee6f0,R_28f_b0ee798,R_290_b0ee840,R_291_b0ee8e8,R_292_b0ee990,R_293_b0eea38,
        R_294_b0eeae0,R_295_b0eeb88,R_296_b0eec30,R_297_b0eecd8,R_298_b0eed80,R_299_b0eee28,R_29a_b0eeed0,R_29b_b0eef78,R_29c_b0ef020);
input RIaa97c98_14,RIaa9e7f0_243,RIaa9e868_244,RIaa9e778_242,RIaa9e9d0_247,RIaa97d88_16,RIaa97d10_15,RIaa97e00_17,RIaa97c20_13,
        RIaa9e688_240,RIaa9e700_241,RIaa9e8e0_245,RIaa9e958_246,RIaa9cf90_191,RIaa9d170_195,RIaa9cea0_189,RIaa9d1e8_196,RIaa9d080_193,RIaa9d0f8_194,
        RIaa9d5a8_204,RIaa9d620_205,RIaa9d2d8_198,RIaa9d008_192,RIaa9d3c8_200,RIaa9d4b8_202,RIaa9d260_197,RIaa9d350_199,RIaa9cf18_190,RIaa9d530_203,
        RIaa9d440_201,RIaa97860_5,RIaa976f8_2,RIaa97770_3,RIaa977e8_4,RIaa9ba00_145,RIaa9b640_137,RIaa9b910_143,RIaa9bd48_152,RIaa9ba78_146,
        RIaa9bb68_148,RIaa9b7a8_140,RIaa9bdc0_153,RIaa9baf0_147,RIaa9b730_139,RIaa9bc58_150,RIaa9b6b8_138,RIaa9b898_142,RIaa9bcd0_151,RIaa9b988_144,
        RIaa9b820_141,RIaa9bbe0_149,RIaa9b370_131,RIaa9b0a0_125,RIaa9b5c8_136,RIaa9b3e8_132,RIaa9ae48_120,RIaa9b460_133,RIaa9b190_127,RIaa9b118_126,
        RIaa9b4d8_134,RIaa9b280_129,RIaa9b028_124,RIaa9af38_122,RIaa9b2f8_130,RIaa9aec0_121,RIaa9b550_135,RIaa9afb0_123,RIaa9b208_128,RIaa9c2e8_164,
        RIaa9c4c8_168,RIaa9c018_158,RIaa9c3d8_166,RIaa9c450_167,RIaa9be38_154,RIaa9bfa0_157,RIaa9beb0_155,RIaa9c270_163,RIaa9c090_159,RIaa9c108_160,
        RIaa9c180_161,RIaa9bf28_156,RIaa9c5b8_170,RIaa9c1f8_162,RIaa9c360_165,RIaa9c540_169,RIaa9ce28_188,RIaa9c978_178,RIaa9c9f0_179,RIaa9c900_177,
        RIaa9cdb0_187,RIaa9c810_175,RIaa9c720_173,RIaa9cb58_182,RIaa9cae0_181,RIaa9c630_171,RIaa9ca68_180,RIaa9cc48_184,RIaa9ccc0_185,RIaa9c888_176,
        RIaa9c6a8_172,RIaa9c798_174,RIaa9cbd0_183,RIaa9cd38_186,RIaa9ab78_114,RIaa9aa10_111,RIaa9ac68_116,RIaa9a7b8_106,RIaa9a6c8_104,RIaa9add0_119,
        RIaa9abf0_115,RIaa9a8a8_108,RIaa9a998_110,RIaa9a920_109,RIaa9a830_107,RIaa9ad58_118,RIaa9a740_105,RIaa9ab00_113,RIaa9aa88_112,RIaa9a650_103,
        RIaa9ace0_117,RIaa978d8_6,RIaa9a308_96,RIaa9a218_94,RIaa9a380_97,RIaa9a038_90,RIaa99ed0_87,RIaa9a290_95,RIaa9a0b0_91,RIaa99fc0_89,
        RIaa9a470_99,RIaa99f48_88,RIaa9a4e8_100,RIaa9a1a0_93,RIaa9a3f8_98,RIaa99e58_86,RIaa9a560_101,RIaa9a128_92,RIaa9a5d8_102,RIaa97950_7,
        RIaa99b10_79,RIaa999a8_76,RIaa99a20_77,RIaa996d8_70,RIaa99930_75,RIaa99d68_84,RIaa99b88_80,RIaa99660_69,RIaa99cf0_83,RIaa99c00_81,
        RIaa998b8_74,RIaa99de0_85,RIaa99a98_78,RIaa99c78_82,RIaa997c8_72,RIaa99840_73,RIaa99750_71,RIaa979c8_8,RIaa9f6f0_275,RIaa9f768_276,
        RIaa9f3a8_268,RIaa9f600_273,RIaa9f2b8_266,RIaa9f330_267,RIaa9f420_269,RIaa9f9c0_281,RIaa9f948_280,RIaa9f678_274,RIaa9f8d0_279,RIaa9f588_272,
        RIaa9f240_265,RIaa9f510_271,RIaa9f7e0_277,RIaa9f858_278,RIaa9f498_270,RIaa9eca0_253,RIaa9ee08_256,RIaa9eef8_258,RIaa9ed90_255,RIaa9f1c8_264,
        RIaa9efe8_260,RIaa9ef70_259,RIaa9ed18_254,RIaa9eb38_250,RIaa9ebb0_251,RIaa9ea48_248,RIaa9f0d8_262,RIaa9ee80_257,RIaa9eac0_249,RIaa9f150_263,
        RIaa9f060_261,RIaa9ec28_252,RIaa97b30_11,RIaa97ba8_12,RIaa9de18_222,RIaa9db48_216,RIaa9d968_212,RIaa9dbc0_217,RIaa9dda0_221,RIaa9dd28_220,
        RIaa9dad0_215,RIaa9d800_209,RIaa9dc38_218,RIaa9d710_207,RIaa9dcb0_219,RIaa9d788_208,RIaa9d698_206,RIaa9da58_214,RIaa9d9e0_213,RIaa9d878_210,
        RIaa9d8f0_211,RIaa994f8_66,RIaa99048_56,RIaa98f58_54,RIaa99570_67,RIaa990c0_57,RIaa99138_58,RIaa99390_63,RIaa98ee0_53,RIaa99480_65,
        RIaa98fd0_55,RIaa995e8_68,RIaa99318_62,RIaa991b0_59,RIaa99408_64,RIaa992a0_61,RIaa98e68_52,RIaa99228_60,RIaa9e160_229,RIaa9df80_225,
        RIaa9e3b8_234,RIaa9de90_223,RIaa9e610_239,RIaa9e2c8_232,RIaa9e598_238,RIaa9e1d8_230,RIaa9df08_224,RIaa9e520_237,RIaa9e340_233,RIaa9e250_231,
        RIaa9e430_235,RIaa9e0e8_228,RIaa9dff8_226,RIaa9e4a8_236,RIaa9e070_227,RIaa97ab8_10,RIaa97a40_9,RIaa98b20_45,RIaa989b8_42,RIaa98c88_48,
        RIaa98a30_43,RIaa98aa8_44,RIaa98df0_51,RIaa98940_41,RIaa98c10_47,RIaa98670_35,RIaa98850_39,RIaa98760_37,RIaa986e8_36,RIaa98d00_49,
        RIaa98b98_46,RIaa987d8_38,RIaa988c8_40,RIaa98d78_50,RIaaa1ce8_356,RIaaa1e50_359,RIaaa2030_363,RIaaa1fb8_362,RIaaa1f40_361,RIaaa1c70_355,
        RIaaa1d60_357,RIaaa1ec8_360,RIaaa1b80_353,RIaaa1bf8_354,RIaaa20a8_364,RIaaa1a90_351,RIaaa2120_365,RIaaa1dd8_358,RIaaa2198_366,RIaaa1b08_352,
        RIaaa1a18_350,RIaaa1130_331,RIaaa0f50_327,RIaaa0a28_316,RIaaa0b90_319,RIaaa0b18_318,RIaaa1040_329,RIaaa0c80_321,RIaaa0cf8_322,RIaaa0c08_320,
        RIaaa0ed8_326,RIaaa0d70_323,RIaaa0aa0_317,RIaaa0fc8_328,RIaaa11a8_332,RIaaa10b8_330,RIaaa0e60_325,RIaaa0de8_324,RIaa97680_1,RIaa98508_32,
        RIaa98328_28,RIaa98238_26,RIaa98418_30,RIaa97e78_18,RIaa981c0_25,RIaa985f8_34,RIaa982b0_27,RIaa98580_33,RIaa97ef0_19,RIaa98058_22,
        RIaa98148_24,RIaa97f68_20,RIaa97fe0_21,RIaa983a0_29,RIaa980d0_23,RIaa98490_31,RIaaa2cd8_390,RIaaa2af8_386,RIaaa3110_399,RIaaa3188_400,
        RIaaa2f30_395,RIaaa2c60_389,RIaaa2eb8_394,RIaaa2dc8_392,RIaaa2e40_393,RIaaa2fa8_396,RIaaa3020_397,RIaaa2a08_384,RIaaa3098_398,RIaaa2be8_388,
        RIaaa2b70_387,RIaaa2a80_385,RIaaa2d50_391,RIaaa1298_334,RIaaa16d0_343,RIaaa1928_348,RIaaa1658_342,RIaaa1838_346,RIaaa14f0_339,RIaaa1388_336,
        RIaaa1400_337,RIaaa19a0_349,RIaaa1748_344,RIaaa15e0_341,RIaaa1310_335,RIaaa1220_333,RIaaa1478_338,RIaaa1568_340,RIaaa17c0_345,RIaaa18b0_347,
        RIaa9ff60_293,RIaa9fba0_285,RIaa9fa38_282,RIaaa0050_295,RIaa9ffd8_294,RIaa9fe70_291,RIaa9fc90_287,RIaaa01b8_298,RIaaa0140_297,RIaa9fdf8_290,
        RIaa9fab0_283,RIaa9fc18_286,RIaa9fb28_284,RIaa9fd08_288,RIaaa00c8_296,RIaa9fee8_292,RIaa9fd80_289,RIaaa05f0_307,RIaaa0938_314,RIaaa0758_310,
        RIaaa0488_304,RIaaa0578_306,RIaaa0230_299,RIaaa06e0_309,RIaaa0848_312,RIaaa0398_302,RIaaa0320_301,RIaaa0668_308,RIaaa0410_303,RIaaa02a8_300,
        RIaaa08c0_313,RIaaa0500_305,RIaaa07d0_311,RIaaa09b0_315,RIaaa24e0_373,RIaaa2558_374,RIaaa2738_378,RIaaa2828_380,RIaaa2300_369,RIaaa26c0_377,
        RIaaa2918_382,RIaaa2468_372,RIaaa2378_370,RIaaa2288_368,RIaaa2648_376,RIaaa23f0_371,RIaaa2210_367,RIaaa25d0_375,RIaaa27b0_379,RIaaa28a0_381,
        RIaaa2990_383,RIaaa3f20_429,RIaaa3f98_430,RIaaa3cc8_424,RIaaa3c50_423,RIaaa4010_431,RIaaa4100_433,RIaaa3db8_426,RIaaa3b60_421,RIaaa3d40_425,
        RIaaa3ae8_420,RIaaa3a70_419,RIaaa39f8_418,RIaaa4178_434,RIaaa3e30_427,RIaaa3bd8_422,RIaaa4088_432,RIaaa3ea8_428,RIaaa32f0_403,RIaaa3890_415,
        RIaaa34d0_407,RIaaa3638_410,RIaaa3728_412,RIaaa35c0_409,RIaaa3278_402,RIaaa3818_414,RIaaa33e0_405,RIaaa3368_404,RIaaa37a0_413,RIaaa3980_417,
        RIaaa3908_416,RIaaa36b0_411,RIaaa3458_406,RIaaa3548_408,RIaaa3200_401,RIaaa4448_440,RIaaa4538_442,RIaaa4268_436,RIaaa43d0_439,RIaaa42e0_437,
        RIaaa41f0_435,RIaaa4628_444,RIaaa4808_448,RIaaa45b0_443,RIaaa4718_446,RIaaa44c0_441,RIaaa48f8_450,RIaaa4358_438,RIaaa4970_451,RIaaa4880_449,
        RIaaa4790_447,RIaaa46a0_445,RIaaa6248_504,RIaaa66f8_514,RIaaa6860_517,RIaaa67e8_516,RIaaa6680_513,RIaaa64a0_509,RIaaa6338_506,RIaaa63b0_507,
        RIaaa6950_519,RIaaa6608_512,RIaaa6590_511,RIaaa6428_508,RIaaa6770_515,RIaaa68d8_518,RIaaa6518_510,RIaaa62c0_505,RIaaa61d0_503,RIaaa57f8_482,
        RIaaa54b0_475,RIaaa5618_478,RIaaa52d0_471,RIaaa5528_476,RIaaa5258_470,RIaaa5708_480,RIaaa5690_479,RIaaa5348_472,RIaaa53c0_473,RIaaa58e8_484,
        RIaaa5960_485,RIaaa5780_481,RIaaa5438_474,RIaaa5870_483,RIaaa55a0_477,RIaaa51e0_469,RIaaa4e98_462,RIaaa49e8_452,RIaaa4b50_455,RIaaa4e20_461,
        RIaaa50f0_467,RIaaa4f88_464,RIaaa5000_465,RIaaa4c40_457,RIaaa4cb8_458,RIaaa4a60_453,RIaaa4f10_463,RIaaa4bc8_456,RIaaa4ad8_454,RIaaa5168_468,
        RIaaa4d30_459,RIaaa4da8_460,RIaaa5078_466,RIaaa5e10_495,RIaaa5ca8_492,RIaaa59d8_486,RIaaa60e0_501,RIaaa5b40_489,RIaaa5a50_487,RIaaa5f00_497,
        RIaaa5bb8_490,RIaaa6158_502,RIaaa5f78_498,RIaaa5ac8_488,RIaaa5e88_496,RIaaa5d98_494,RIaaa5ff0_499,RIaaa5d20_493,RIaaa6068_500,RIaaa5c30_491,
        RIaaa6d10_527,RIaaa6a40_521,RIaaa7058_534,RIaaa7148_536,RIaaa6e00_529,RIaaa6ba8_524,RIaaa6e78_530,RIaaa6c98_526,RIaaa6f68_532,RIaaa6ab8_522,
        RIaaa70d0_535,RIaaa6c20_525,RIaaa69c8_520,RIaaa6d88_528,RIaaa6fe0_533,RIaaa6ef0_531,RIaaa6b30_523,RIaaa8408_576,RIaaa87c8_584,RIaaa84f8_578,
        RIaaa8390_575,RIaaa8318_574,RIaaa8660_581,RIaaa8228_572,RIaaa88b8_586,RIaaa8930_587,RIaaa8750_583,RIaaa8480_577,RIaaa8840_585,RIaaa86d8_582,
        RIaaa85e8_580,RIaaa8570_579,RIaaa82a0_573,RIaaa81b0_571,RIaaa7670_547,RIaaa7238_538,RIaaa7490_543,RIaaa75f8_546,RIaaa78c8_552,RIaaa7328_540,
        RIaaa73a0_541,RIaaa77d8_550,RIaaa7850_551,RIaaa76e8_548,RIaaa7580_545,RIaaa72b0_539,RIaaa71c0_537,RIaaa7508_544,RIaaa7418_542,RIaaa7940_553,
        RIaaa7760_549,RIaaa7d00_561,RIaaa7f58_566,RIaaa7fd0_567,RIaaa7b98_558,RIaaa7b20_557,RIaaa7df0_563,RIaaa7c88_560,RIaaa7e68_564,RIaaa7ee0_565,
        RIaaa7d78_562,RIaaa8048_568,RIaaa7c10_559,RIaaa8138_570,RIaaa80c0_569,RIaaa7aa8_556,RIaaa7a30_555,RIaaa79b8_554,RIaaa89a8_588,RIaaa95d8_614,
        RIaaa9218_606,RIaaa90b0_603,RIaaa9128_604,RIaaa91a0_605,RIaaa9380_609,RIaaa9308_608,RIaaa9290_607,RIaaa9038_602,RIaaa93f8_610,RIaaa9470_611,
        RIaaa94e8_612,RIaaa8c78_594,RIaaa8cf0_595,RIaaa8a98_590,RIaaa8b10_591,RIaaa8a20_589,RIaaa8b88_592,RIaaa8c00_593,RIaaa8d68_596,RIaaa8de0_597,
        RIaaa8e58_598,RIaaa8ed0_599,RIaaa8f48_600,RIaaa8fc0_601,RIaaa9560_613;
output R_267_b0ecd58,R_268_b0ece00,R_269_b0ecea8,R_26a_b0ecf50,R_26b_b0ecff8,R_26c_b0ed0a0,R_26d_b0ed148,R_26e_b0ed1f0,R_26f_b0ed298,
        R_270_b0ed340,R_271_b0ed3e8,R_272_b0ed490,R_273_b0ed538,R_274_b0ed5e0,R_275_b0ed688,R_276_b0ed730,R_277_b0ed7d8,R_278_b0ed880,R_279_b0ed928,
        R_27a_b0ed9d0,R_27b_b0eda78,R_27c_b0edb20,R_27d_b0edbc8,R_27e_b0edc70,R_27f_b0edd18,R_280_b0eddc0,R_281_b0ede68,R_282_b0edf10,R_283_b0edfb8,
        R_284_b0ee060,R_285_b0ee108,R_286_b0ee1b0,R_287_b0ee258,R_288_b0ee300,R_289_b0ee3a8,R_28a_b0ee450,R_28b_b0ee4f8,R_28c_b0ee5a0,R_28d_b0ee648,
        R_28e_b0ee6f0,R_28f_b0ee798,R_290_b0ee840,R_291_b0ee8e8,R_292_b0ee990,R_293_b0eea38,R_294_b0eeae0,R_295_b0eeb88,R_296_b0eec30,R_297_b0eecd8,
        R_298_b0eed80,R_299_b0eee28,R_29a_b0eeed0,R_29b_b0eef78,R_29c_b0ef020;

wire \649_ZERO , \650_ONE , \651 , \652 , \653 , \654 , \655 , \656 , \657 ,
         \658 , \659 , \660 , \661 , \662 , \663 , \664 , \665 , \666 , \667 ,
         \668 , \669 , \670 , \671 , \672 , \673 , \674 , \675 , \676 , \677 ,
         \678 , \679 , \680 , \681 , \682 , \683 , \684 , \685 , \686 , \687 ,
         \688 , \689 , \690 , \691 , \692 , \693 , \694 , \695 , \696 , \697 ,
         \698 , \699 , \700 , \701 , \702 , \703 , \704 , \705 , \706 , \707 ,
         \708 , \709 , \710 , \711 , \712 , \713 , \714 , \715 , \716 , \717 ,
         \718 , \719 , \720 , \721 , \722 , \723 , \724 , \725 , \726 , \727 ,
         \728 , \729 , \730 , \731 , \732 , \733 , \734 , \735 , \736 , \737 ,
         \738 , \739 , \740 , \741 , \742 , \743 , \744 , \745 , \746 , \747 ,
         \748 , \749 , \750 , \751_nG11a6 , \752 , \753 , \754 , \755 , \756 , \757 ,
         \758 , \759 , \760 , \761 , \762 , \763 , \764 , \765 , \766 , \767 ,
         \768 , \769 , \770 , \771 , \772 , \773 , \774 , \775 , \776 , \777 ,
         \778 , \779 , \780 , \781 , \782 , \783 , \784 , \785 , \786 , \787_nGfc6 ,
         \788 , \789 , \790 , \791 , \792 , \793 , \794 , \795 , \796 , \797 ,
         \798 , \799 , \800 , \801 , \802 , \803 , \804 , \805 , \806 , \807 ,
         \808 , \809 , \810 , \811 , \812 , \813 , \814 , \815 , \816 , \817 ,
         \818 , \819 , \820 , \821 , \822 , \823_nGfc4 , \824 , \825 , \826 , \827 ,
         \828 , \829 , \830 , \831 , \832 , \833 , \834 , \835 , \836 , \837 ,
         \838 , \839 , \840 , \841 , \842 , \843 , \844 , \845 , \846 , \847 ,
         \848 , \849 , \850 , \851 , \852 , \853 , \854 , \855 , \856 , \857 ,
         \858 , \859 , \860 , \861_nGe1a , \862 , \863 , \864 , \865 , \866 , \867 ,
         \868 , \869 , \870 , \871 , \872 , \873 , \874 , \875 , \876 , \877 ,
         \878 , \879 , \880 , \881 , \882 , \883 , \884 , \885 , \886 , \887 ,
         \888 , \889 , \890 , \891 , \892 , \893 , \894 , \895 , \896 , \897 ,
         \898 , \899_nGe18 , \900 , \901 , \902 , \903 , \904 , \905 , \906 , \907 ,
         \908 , \909 , \910 , \911 , \912 , \913 , \914 , \915 , \916 , \917 ,
         \918 , \919 , \920 , \921 , \922 , \923 , \924 , \925 , \926 , \927 ,
         \928 , \929 , \930 , \931 , \932 , \933 , \934 , \935 , \936 , \937_nGa83 ,
         \938 , \939 , \940 , \941 , \942 , \943 , \944 , \945 , \946 , \947 ,
         \948 , \949 , \950 , \951 , \952 , \953 , \954 , \955 , \956 , \957 ,
         \958 , \959 , \960 , \961 , \962 , \963 , \964 , \965 , \966 , \967 ,
         \968 , \969 , \970 , \971 , \972 , \973 , \974 , \975_nGa81 , \976 , \977 ,
         \978 , \979 , \980 , \981 , \982 , \983 , \984 , \985 , \986 , \987 ,
         \988 , \989 , \990 , \991 , \992 , \993 , \994 , \995 , \996 , \997 ,
         \998 , \999 , \1000 , \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 ,
         \1008 , \1009 , \1010 , \1011_nGa12 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 ,
         \1018 , \1019 , \1020 , \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 ,
         \1028 , \1029 , \1030 , \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 ,
         \1038 , \1039 , \1040 , \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 ,
         \1048 , \1049_nGa10 , \1050 , \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 ,
         \1058 , \1059 , \1060 , \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 ,
         \1068 , \1069 , \1070 , \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 ,
         \1078 , \1079 , \1080 , \1081_nG9bb , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 ,
         \1088 , \1089 , \1090 , \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 ,
         \1098 , \1099 , \1100 , \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 ,
         \1108 , \1109 , \1110 , \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117_nG9bd ,
         \1118 , \1119 , \1120 , \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 ,
         \1128 , \1129 , \1130 , \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 ,
         \1138 , \1139 , \1140 , \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 ,
         \1148_nG949 , \1149 , \1150 , \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 ,
         \1158 , \1159 , \1160 , \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 ,
         \1168 , \1169 , \1170 , \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 ,
         \1178 , \1179 , \1180 , \1181_nG947 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 ,
         \1188 , \1189 , \1190 , \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 ,
         \1198 , \1199 , \1200 , \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 ,
         \1208 , \1209 , \1210 , \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 ,
         \1218 , \1219 , \1220 , \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 ,
         \1228 , \1229 , \1230 , \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 ,
         \1238 , \1239 , \1240 , \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 ,
         \1248 , \1249 , \1250 , \1251 , \1252 , \1253_nG17dd , \1254 , \1255 , \1256 , \1257 ,
         \1258 , \1259 , \1260 , \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 ,
         \1268 , \1269 , \1270 , \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 ,
         \1278 , \1279 , \1280 , \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 ,
         \1288 , \1289 , \1290 , \1291 , \1292 , \1293_nG18eb , \1294 , \1295 , \1296 , \1297 ,
         \1298 , \1299 , \1300 , \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 ,
         \1308 , \1309 , \1310 , \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 ,
         \1318 , \1319 , \1320 , \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 ,
         \1328 , \1329 , \1330 , \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 ,
         \1338 , \1339 , \1340 , \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 ,
         \1348_nG16d6 , \1349 , \1350 , \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 ,
         \1358 , \1359 , \1360 , \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 ,
         \1368 , \1369 , \1370 , \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 ,
         \1378 , \1379 , \1380 , \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 ,
         \1388 , \1389 , \1390 , \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 ,
         \1398 , \1399 , \1400 , \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 ,
         \1408 , \1409 , \1410 , \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 ,
         \1418 , \1419 , \1420 , \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 ,
         \1428 , \1429 , \1430 , \1431 , \1432 , \1433 , \1434 , \1435_nG15b1 , \1436 , \1437 ,
         \1438 , \1439 , \1440 , \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 ,
         \1448 , \1449 , \1450 , \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 ,
         \1458 , \1459 , \1460 , \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 ,
         \1468 , \1469 , \1470 , \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 ,
         \1478 , \1479 , \1480 , \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 ,
         \1488 , \1489 , \1490 , \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 ,
         \1498 , \1499 , \1500 , \1501 , \1502_nG14c8 , \1503 , \1504 , \1505 , \1506 , \1507 ,
         \1508 , \1509 , \1510 , \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 ,
         \1518 , \1519 , \1520 , \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 ,
         \1528 , \1529 , \1530 , \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 ,
         \1538 , \1539 , \1540 , \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 ,
         \1548 , \1549 , \1550 , \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 ,
         \1558 , \1559_nG13c8 , \1560 , \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 ,
         \1568 , \1569 , \1570 , \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 ,
         \1578 , \1579 , \1580 , \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 ,
         \1588 , \1589 , \1590 , \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 ,
         \1598 , \1599 , \1600 , \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 ,
         \1608 , \1609 , \1610 , \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 ,
         \1618 , \1619 , \1620 , \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 ,
         \1628 , \1629 , \1630 , \1631_nG12c9 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 ,
         \1638 , \1639 , \1640 , \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 ,
         \1648 , \1649 , \1650 , \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 ,
         \1658 , \1659 , \1660 , \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 ,
         \1668 , \1669 , \1670 , \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 ,
         \1678 , \1679 , \1680 , \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 ,
         \1688 , \1689 , \1690 , \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 ,
         \1698 , \1699 , \1700 , \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 ,
         \1708 , \1709 , \1710_nG11c1 , \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 ,
         \1718 , \1719 , \1720 , \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 ,
         \1728 , \1729 , \1730 , \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 ,
         \1738 , \1739 , \1740 , \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 ,
         \1748 , \1749 , \1750 , \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 ,
         \1758 , \1759 , \1760 , \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 ,
         \1768 , \1769 , \1770 , \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 ,
         \1778 , \1779 , \1780 , \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787_nG10e2 ,
         \1788 , \1789 , \1790 , \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 ,
         \1798 , \1799 , \1800 , \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 ,
         \1808 , \1809 , \1810 , \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 ,
         \1818 , \1819 , \1820 , \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 ,
         \1828 , \1829 , \1830 , \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 ,
         \1838 , \1839 , \1840 , \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 ,
         \1848 , \1849 , \1850 , \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 ,
         \1858 , \1859 , \1860 , \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 ,
         \1868 , \1869 , \1870 , \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 ,
         \1878 , \1879 , \1880 , \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 ,
         \1888 , \1889 , \1890 , \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 ,
         \1898 , \1899 , \1900 , \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 ,
         \1908 , \1909 , \1910 , \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 ,
         \1918 , \1919 , \1920 , \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 ,
         \1928 , \1929 , \1930 , \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 ,
         \1938 , \1939 , \1940 , \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 ,
         \1948 , \1949 , \1950 , \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 ,
         \1958 , \1959 , \1960 , \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 ,
         \1968 , \1969 , \1970 , \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 ,
         \1978 , \1979 , \1980 , \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 ,
         \1988 , \1989 , \1990 , \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 ,
         \1998 , \1999 , \2000 , \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 ,
         \2008 , \2009 , \2010 , \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 ,
         \2018 , \2019 , \2020 , \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 ,
         \2028 , \2029 , \2030 , \2031 , \2032 , \2033 , \2034_nGfe1 , \2035 , \2036 , \2037 ,
         \2038 , \2039 , \2040 , \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 ,
         \2048 , \2049 , \2050 , \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 ,
         \2058 , \2059 , \2060 , \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 ,
         \2068 , \2069 , \2070 , \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 ,
         \2078 , \2079 , \2080 , \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 ,
         \2088 , \2089 , \2090 , \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 ,
         \2098 , \2099 , \2100 , \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 ,
         \2108 , \2109 , \2110 , \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 ,
         \2118 , \2119 , \2120 , \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 ,
         \2128 , \2129 , \2130 , \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 ,
         \2138 , \2139 , \2140 , \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 ,
         \2148 , \2149 , \2150 , \2151 , \2152 , \2153 , \2154 , \2155 , \2156_nGf08 , \2157 ,
         \2158 , \2159 , \2160 , \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 ,
         \2168 , \2169 , \2170 , \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 ,
         \2178 , \2179 , \2180 , \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 ,
         \2188 , \2189 , \2190 , \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 ,
         \2198 , \2199 , \2200 , \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 ,
         \2208 , \2209 , \2210 , \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 ,
         \2218 , \2219 , \2220 , \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 ,
         \2228 , \2229_nGe35 , \2230 , \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 ,
         \2238 , \2239 , \2240 , \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 ,
         \2248 , \2249 , \2250 , \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 ,
         \2258 , \2259 , \2260 , \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 ,
         \2268 , \2269 , \2270 , \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 ,
         \2278 , \2279 , \2280 , \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 ,
         \2288 , \2289 , \2290 , \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 ,
         \2298 , \2299 , \2300 , \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 ,
         \2308 , \2309 , \2310 , \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 ,
         \2318 , \2319 , \2320 , \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 ,
         \2328 , \2329 , \2330 , \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 ,
         \2338 , \2339 , \2340 , \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 ,
         \2348 , \2349 , \2350 , \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 ,
         \2358 , \2359 , \2360 , \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 ,
         \2368 , \2369 , \2370 , \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 ,
         \2378 , \2379 , \2380 , \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 ,
         \2388 , \2389 , \2390 , \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 ,
         \2398 , \2399 , \2400 , \2401 , \2402 , \2403 , \2404_nGad6 , \2405 , \2406 , \2407 ,
         \2408 , \2409 , \2410 , \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 ,
         \2418 , \2419 , \2420 , \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 ,
         \2428 , \2429 , \2430 , \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 ,
         \2438 , \2439 , \2440 , \2441 , \2442 , \2443 , \2444 , \2445 , \2446_nGa9e , \2447 ,
         \2448 , \2449 , \2450 , \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 ,
         \2458 , \2459 , \2460 , \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 ,
         \2468 , \2469 , \2470 , \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 ,
         \2478 , \2479 , \2480 , \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 ,
         \2488 , \2489 , \2490 , \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 ,
         \2498 , \2499 , \2500 , \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 ,
         \2508 , \2509 , \2510 , \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 ,
         \2518 , \2519 , \2520 , \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 ,
         \2528 , \2529 , \2530 , \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 ,
         \2538 , \2539 , \2540 , \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 ,
         \2548 , \2549 , \2550 , \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 ,
         \2558 , \2559 , \2560 , \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 ,
         \2568 , \2569 , \2570 , \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 ,
         \2578 , \2579 , \2580 , \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 ,
         \2588 , \2589 , \2590 , \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 ,
         \2598 , \2599 , \2600 , \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 ,
         \2608 , \2609 , \2610 , \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 ,
         \2618 , \2619 , \2620 , \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 ,
         \2628 , \2629 , \2630 , \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 ,
         \2638 , \2639 , \2640 , \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 ,
         \2648 , \2649 , \2650 , \2651 , \2652 , \2653_nGa66 , \2654 , \2655 , \2656 , \2657 ,
         \2658 , \2659 , \2660 , \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 ,
         \2668 , \2669 , \2670 , \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 ,
         \2678 , \2679 , \2680 , \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 ,
         \2688 , \2689 , \2690 , \2691 , \2692 , \2693 , \2694 , \2695_nGa2d , \2696 , \2697 ,
         \2698 , \2699 , \2700 , \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 ,
         \2708 , \2709 , \2710 , \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 ,
         \2718 , \2719 , \2720 , \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 ,
         \2728 , \2729 , \2730 , \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 ,
         \2738 , \2739 , \2740 , \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 ,
         \2748 , \2749 , \2750 , \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 ,
         \2758 , \2759 , \2760 , \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 ,
         \2768 , \2769 , \2770 , \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 ,
         \2778 , \2779 , \2780 , \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 ,
         \2788 , \2789 , \2790 , \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 ,
         \2798 , \2799 , \2800 , \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 ,
         \2808 , \2809 , \2810 , \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 ,
         \2818 , \2819 , \2820 , \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 ,
         \2828 , \2829 , \2830 , \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 ,
         \2838 , \2839 , \2840 , \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 ,
         \2848 , \2849 , \2850 , \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 ,
         \2858 , \2859 , \2860 , \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 ,
         \2868 , \2869 , \2870 , \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 ,
         \2878 , \2879 , \2880 , \2881 , \2882 , \2883 , \2884 , \2885 , \2886_nG9f5 , \2887 ,
         \2888 , \2889 , \2890 , \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 ,
         \2898 , \2899 , \2900 , \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 ,
         \2908 , \2909 , \2910 , \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 ,
         \2918 , \2919 , \2920 , \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 ,
         \2928 , \2929 , \2930 , \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 ,
         \2938 , \2939 , \2940 , \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 ,
         \2948 , \2949 , \2950 , \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 ,
         \2958 , \2959 , \2960 , \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 ,
         \2968 , \2969 , \2970 , \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 ,
         \2978 , \2979 , \2980 , \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 ,
         \2988 , \2989 , \2990 , \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 ,
         \2998 , \2999 , \3000 , \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 ,
         \3008_nG9b9 , \3009 , \3010 , \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 ,
         \3018 , \3019 , \3020 , \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 ,
         \3028 , \3029 , \3030 , \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 ,
         \3038 , \3039 , \3040 , \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 ,
         \3048 , \3049 , \3050 , \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 ,
         \3058 , \3059 , \3060 , \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 ,
         \3068 , \3069 , \3070 , \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 ,
         \3078 , \3079 , \3080 , \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 ,
         \3088 , \3089 , \3090 , \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 ,
         \3098 , \3099 , \3100 , \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 ,
         \3108 , \3109 , \3110 , \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 ,
         \3118 , \3119 , \3120 , \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 ,
         \3128 , \3129 , \3130 , \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 ,
         \3138 , \3139 , \3140 , \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 ,
         \3148 , \3149 , \3150 , \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 ,
         \3158 , \3159 , \3160 , \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 ,
         \3168 , \3169 , \3170 , \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 ,
         \3178 , \3179 , \3180 , \3181 , \3182_nG984 , \3183 , \3184 , \3185 , \3186 , \3187 ,
         \3188 , \3189 , \3190 , \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 ,
         \3198 , \3199 , \3200 , \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 ,
         \3208 , \3209 , \3210 , \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 ,
         \3218 , \3219 , \3220 , \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 ,
         \3228 , \3229 , \3230 , \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 ,
         \3238 , \3239 , \3240 , \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 ,
         \3248 , \3249 , \3250 , \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 ,
         \3258 , \3259 , \3260 , \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 ,
         \3268 , \3269 , \3270 , \3271 , \3272 , \3273_nG944 , \3274 , \3275 , \3276 , \3277 ,
         \3278 , \3279 , \3280 , \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 ,
         \3288 , \3289 , \3290 , \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 ,
         \3298 , \3299 , \3300 , \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 ,
         \3308 , \3309 , \3310 , \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 ,
         \3318 , \3319 , \3320 , \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 ,
         \3328 , \3329 , \3330 , \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 ,
         \3338 , \3339 , \3340 , \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 ,
         \3348 , \3349 , \3350 , \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 ,
         \3358 , \3359 , \3360 , \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 ,
         \3368 , \3369 , \3370 , \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 ,
         \3378 , \3379 , \3380 , \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 ,
         \3388 , \3389 , \3390 , \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 ,
         \3398 , \3399 , \3400 , \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 ,
         \3408 , \3409 , \3410 , \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 ,
         \3418 , \3419 , \3420 , \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 ,
         \3428 , \3429 , \3430 , \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 ,
         \3438 , \3439 , \3440 , \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 ,
         \3448 , \3449 , \3450 , \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 ,
         \3458 , \3459 , \3460 , \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 ,
         \3468 , \3469 , \3470 , \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 ,
         \3478 , \3479 , \3480 , \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 ,
         \3488 , \3489 , \3490 , \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 ,
         \3498 , \3499 , \3500 , \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 ,
         \3508 , \3509 , \3510 , \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 ,
         \3518 , \3519 , \3520 , \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 ,
         \3528 , \3529 , \3530 , \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 ,
         \3538 , \3539 , \3540 , \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 ,
         \3548 , \3549 , \3550 , \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 ,
         \3558 , \3559 , \3560 , \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 ,
         \3568 , \3569 , \3570 , \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 ,
         \3578 , \3579 , \3580 , \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 ,
         \3588 , \3589 , \3590 , \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 ,
         \3598 , \3599 , \3600 , \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 ,
         \3608 , \3609 , \3610 , \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 ,
         \3618 , \3619 , \3620 , \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 ,
         \3628 , \3629 , \3630 , \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 ,
         \3638 , \3639 , \3640 , \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 ,
         \3648 , \3649 , \3650 , \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 ,
         \3658 , \3659 , \3660 , \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 ,
         \3668 , \3669 , \3670 , \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 ,
         \3678 , \3679 , \3680 , \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 ,
         \3688 , \3689 , \3690 , \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 ,
         \3698 , \3699 , \3700 , \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 ,
         \3708 , \3709 , \3710 , \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 ,
         \3718 , \3719 , \3720 , \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 ,
         \3728 , \3729 , \3730 , \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 ,
         \3738 , \3739 , \3740 , \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 ,
         \3748 , \3749 , \3750 , \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 ,
         \3758 , \3759 , \3760 , \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 ,
         \3768 , \3769 , \3770 , \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 ,
         \3778 , \3779 , \3780 , \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 ,
         \3788 , \3789 , \3790 , \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 ,
         \3798 , \3799 , \3800 , \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 ,
         \3808 , \3809 , \3810 , \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 ,
         \3818 , \3819 , \3820 , \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 ,
         \3828 , \3829 , \3830 , \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 ,
         \3838 , \3839 , \3840 , \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 ,
         \3848 , \3849 , \3850 , \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 ,
         \3858 , \3859 , \3860 , \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 ,
         \3868 , \3869 , \3870 , \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 ,
         \3878 , \3879 , \3880 , \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 ,
         \3888 , \3889 , \3890 , \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 ,
         \3898 , \3899 , \3900 , \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 ,
         \3908 , \3909 , \3910 , \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 ,
         \3918 , \3919 , \3920 , \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 ,
         \3928 , \3929 , \3930 , \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 ,
         \3938 , \3939 , \3940 , \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 ,
         \3948 , \3949 , \3950 , \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 ,
         \3958 , \3959 , \3960 , \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 ,
         \3968 , \3969 , \3970 , \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 ,
         \3978 , \3979 , \3980 , \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 ,
         \3988 , \3989 , \3990 , \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 ,
         \3998 , \3999 , \4000 , \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 ,
         \4008 , \4009 , \4010 , \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 ,
         \4018 , \4019 , \4020 , \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 ,
         \4028 , \4029 , \4030 , \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 ,
         \4038 , \4039 , \4040 , \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 ,
         \4048 , \4049 , \4050 , \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 ,
         \4058 , \4059 , \4060 , \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 ,
         \4068 , \4069 , \4070 , \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 ,
         \4078 , \4079 , \4080 , \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 ,
         \4088 , \4089 , \4090 , \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 ,
         \4098 , \4099 , \4100 , \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 ,
         \4108 , \4109 , \4110 , \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 ,
         \4118 , \4119 , \4120 , \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 ,
         \4128 , \4129 , \4130 , \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 ,
         \4138 , \4139 , \4140 , \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 ,
         \4148 , \4149 , \4150 , \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 ,
         \4158 , \4159 , \4160 , \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 ,
         \4168 , \4169 , \4170 , \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 ,
         \4178 , \4179 , \4180_nG11c3 , \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 ,
         \4188 , \4189 , \4190 , \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 ,
         \4198 , \4199 , \4200 , \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 ,
         \4208 , \4209_nGfe5 , \4210 , \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 ,
         \4218 , \4219 , \4220 , \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 ,
         \4228 , \4229 , \4230 , \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 ,
         \4238_nGfe3 , \4239 , \4240 , \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 ,
         \4248 , \4249 , \4250 , \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 ,
         \4258 , \4259 , \4260 , \4261 , \4262 , \4263 , \4264 , \4265 , \4266_nGe39 , \4267 ,
         \4268 , \4269 , \4270 , \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 ,
         \4278 , \4279 , \4280 , \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 ,
         \4288 , \4289 , \4290 , \4291 , \4292 , \4293 , \4294 , \4295_nGe37 , \4296 , \4297 ,
         \4298 , \4299 , \4300 , \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 ,
         \4308 , \4309 , \4310 , \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 ,
         \4318 , \4319 , \4320 , \4321 , \4322 , \4323 , \4324_nGaa2 , \4325 , \4326 , \4327 ,
         \4328 , \4329 , \4330 , \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 ,
         \4338 , \4339 , \4340 , \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 ,
         \4348 , \4349 , \4350 , \4351 , \4352 , \4353_nGaa0 , \4354 , \4355 , \4356 , \4357 ,
         \4358 , \4359 , \4360 , \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 ,
         \4368 , \4369 , \4370 , \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 ,
         \4378 , \4379 , \4380 , \4381 , \4382_nGa31 , \4383 , \4384 , \4385 , \4386 , \4387 ,
         \4388 , \4389 , \4390 , \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 ,
         \4398 , \4399 , \4400 , \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 ,
         \4408 , \4409 , \4410 , \4411_nGa2f , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 ,
         \4418 , \4419 , \4420 , \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 ,
         \4428 , \4429 , \4430 , \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 ,
         \4438 , \4439 , \4440_nG9d8 , \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 ,
         \4448 , \4449 , \4450 , \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 ,
         \4458 , \4459 , \4460 , \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 ,
         \4468 , \4469_nG9da , \4470 , \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 ,
         \4478 , \4479 , \4480 , \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 ,
         \4488 , \4489 , \4490 , \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 ,
         \4498_nG969 , \4499 , \4500 , \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 ,
         \4508 , \4509 , \4510 , \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 ,
         \4518 , \4519 , \4520 , \4521 , \4522 , \4523 , \4524 , \4525 , \4526_nG967 , \4527 ,
         \4528 , \4529 , \4530 , \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 ,
         \4538 , \4539 , \4540 , \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 ,
         \4548 , \4549 , \4550 , \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 ,
         \4558 , \4559 , \4560 , \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 ,
         \4568 , \4569 , \4570 , \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 ,
         \4578 , \4579 , \4580 , \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 ,
         \4588 , \4589 , \4590 , \4591 , \4592 , \4593_nG17f6 , \4594 , \4595 , \4596 , \4597 ,
         \4598 , \4599 , \4600 , \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 ,
         \4608 , \4609 , \4610 , \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 ,
         \4618 , \4619 , \4620 , \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 ,
         \4628 , \4629 , \4630 , \4631 , \4632_nG1905 , \4633 , \4634 , \4635 , \4636 , \4637 ,
         \4638 , \4639 , \4640 , \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 ,
         \4648 , \4649 , \4650 , \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 ,
         \4658 , \4659 , \4660 , \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 ,
         \4668 , \4669 , \4670 , \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 ,
         \4678 , \4679 , \4680 , \4681 , \4682 , \4683 , \4684 , \4685 , \4686_nG16f0 , \4687 ,
         \4688 , \4689 , \4690 , \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 ,
         \4698 , \4699 , \4700 , \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 ,
         \4708 , \4709 , \4710 , \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 ,
         \4718 , \4719 , \4720 , \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 ,
         \4728 , \4729 , \4730 , \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 ,
         \4738 , \4739 , \4740 , \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 ,
         \4748 , \4749 , \4750 , \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757_nG15ca ,
         \4758 , \4759 , \4760 , \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 ,
         \4768 , \4769 , \4770 , \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 ,
         \4778 , \4779 , \4780 , \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 ,
         \4788 , \4789 , \4790 , \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 ,
         \4798 , \4799 , \4800 , \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 ,
         \4808 , \4809 , \4810 , \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 ,
         \4818 , \4819 , \4820 , \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 ,
         \4828 , \4829 , \4830 , \4831 , \4832 , \4833 , \4834 , \4835 , \4836_nG14e1 , \4837 ,
         \4838 , \4839 , \4840 , \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 ,
         \4848 , \4849 , \4850 , \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 ,
         \4858 , \4859 , \4860 , \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 ,
         \4868 , \4869 , \4870 , \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 ,
         \4878 , \4879 , \4880 , \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 ,
         \4888 , \4889 , \4890 , \4891_nG13e1 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 ,
         \4898 , \4899 , \4900 , \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 ,
         \4908 , \4909 , \4910 , \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 ,
         \4918 , \4919 , \4920 , \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 ,
         \4928 , \4929 , \4930 , \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 ,
         \4938 , \4939 , \4940 , \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 ,
         \4948 , \4949 , \4950 , \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 ,
         \4958 , \4959 , \4960_nG12e2 , \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 ,
         \4968 , \4969 , \4970 , \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 ,
         \4978 , \4979 , \4980 , \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 ,
         \4988 , \4989 , \4990 , \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 ,
         \4998 , \4999 , \5000 , \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 ,
         \5008 , \5009 , \5010 , \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 ,
         \5018 , \5019 , \5020 , \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 ,
         \5028 , \5029 , \5030 , \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 ,
         \5038 , \5039 , \5040 , \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 ,
         \5048 , \5049 , \5050 , \5051 , \5052 , \5053 , \5054 , \5055_nG11dc , \5056 , \5057 ,
         \5058 , \5059 , \5060 , \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 ,
         \5068 , \5069 , \5070 , \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 ,
         \5078 , \5079 , \5080 , \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 ,
         \5088 , \5089 , \5090 , \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 ,
         \5098 , \5099 , \5100 , \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 ,
         \5108 , \5109 , \5110 , \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 ,
         \5118 , \5119_nG10fb , \5120 , \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 ,
         \5128 , \5129 , \5130 , \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 ,
         \5138 , \5139 , \5140 , \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 ,
         \5148 , \5149 , \5150 , \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 ,
         \5158 , \5159 , \5160 , \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 ,
         \5168 , \5169 , \5170 , \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 ,
         \5178 , \5179 , \5180 , \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 ,
         \5188 , \5189 , \5190 , \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 ,
         \5198 , \5199 , \5200 , \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 ,
         \5208 , \5209 , \5210 , \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 ,
         \5218 , \5219 , \5220 , \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 ,
         \5228 , \5229 , \5230 , \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 ,
         \5238 , \5239 , \5240 , \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 ,
         \5248 , \5249 , \5250 , \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 ,
         \5258 , \5259 , \5260 , \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 ,
         \5268 , \5269 , \5270 , \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 ,
         \5278 , \5279 , \5280 , \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 ,
         \5288 , \5289 , \5290 , \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 ,
         \5298 , \5299 , \5300 , \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 ,
         \5308 , \5309 , \5310 , \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 ,
         \5318 , \5319 , \5320 , \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 ,
         \5328 , \5329 , \5330 , \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 ,
         \5338 , \5339 , \5340 , \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 ,
         \5348 , \5349 , \5350 , \5351_nGffe , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 ,
         \5358 , \5359 , \5360 , \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 ,
         \5368 , \5369 , \5370 , \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 ,
         \5378 , \5379 , \5380 , \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 ,
         \5388 , \5389 , \5390 , \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 ,
         \5398 , \5399 , \5400 , \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 ,
         \5408 , \5409 , \5410 , \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 ,
         \5418 , \5419 , \5420 , \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 ,
         \5428 , \5429 , \5430 , \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 ,
         \5438 , \5439 , \5440 , \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 ,
         \5448 , \5449 , \5450 , \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 ,
         \5458 , \5459 , \5460 , \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 ,
         \5468 , \5469 , \5470 , \5471_nGf21 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 ,
         \5478 , \5479 , \5480 , \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 ,
         \5488 , \5489 , \5490 , \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 ,
         \5498 , \5499 , \5500 , \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 ,
         \5508 , \5509 , \5510 , \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 ,
         \5518 , \5519 , \5520 , \5521 , \5522 , \5523 , \5524 , \5525 , \5526_nGe53 , \5527 ,
         \5528 , \5529 , \5530 , \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 ,
         \5538 , \5539 , \5540 , \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 ,
         \5548 , \5549 , \5550 , \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 ,
         \5558 , \5559 , \5560 , \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 ,
         \5568 , \5569 , \5570 , \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 ,
         \5578 , \5579 , \5580 , \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 ,
         \5588 , \5589 , \5590 , \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 ,
         \5598 , \5599 , \5600 , \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 ,
         \5608 , \5609 , \5610 , \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 ,
         \5618 , \5619 , \5620 , \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 ,
         \5628 , \5629 , \5630 , \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 ,
         \5638 , \5639 , \5640 , \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 ,
         \5648 , \5649 , \5650 , \5651 , \5652 , \5653 , \5654 , \5655 , \5656_nGaf0 , \5657 ,
         \5658 , \5659 , \5660 , \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 ,
         \5668 , \5669 , \5670 , \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 ,
         \5678 , \5679 , \5680 , \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 ,
         \5688 , \5689 , \5690 , \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 ,
         \5698 , \5699 , \5700 , \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 ,
         \5708 , \5709 , \5710 , \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 ,
         \5718 , \5719 , \5720 , \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 ,
         \5728 , \5729 , \5730 , \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 ,
         \5738 , \5739 , \5740 , \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 ,
         \5748 , \5749 , \5750 , \5751_nGabb , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 ,
         \5758 , \5759 , \5760 , \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 ,
         \5768 , \5769 , \5770 , \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 ,
         \5778 , \5779 , \5780 , \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 ,
         \5788 , \5789 , \5790 , \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 ,
         \5798 , \5799 , \5800 , \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 ,
         \5808 , \5809 , \5810 , \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 ,
         \5818 , \5819 , \5820 , \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 ,
         \5828 , \5829 , \5830 , \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 ,
         \5838 , \5839 , \5840 , \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 ,
         \5848 , \5849 , \5850 , \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 ,
         \5858 , \5859 , \5860 , \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 ,
         \5868 , \5869 , \5870 , \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 ,
         \5878 , \5879 , \5880 , \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 ,
         \5888 , \5889 , \5890 , \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 ,
         \5898 , \5899 , \5900 , \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 ,
         \5908 , \5909 , \5910 , \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 ,
         \5918 , \5919 , \5920 , \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 ,
         \5928 , \5929 , \5930 , \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 ,
         \5938 , \5939 , \5940 , \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 ,
         \5948 , \5949 , \5950_nGa4b , \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 ,
         \5958 , \5959 , \5960 , \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 ,
         \5968 , \5969 , \5970 , \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 ,
         \5978_nGa7f , \5979 , \5980 , \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 ,
         \5988 , \5989 , \5990 , \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 ,
         \5998 , \5999 , \6000 , \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 ,
         \6008 , \6009 , \6010 , \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 ,
         \6018 , \6019 , \6020 , \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 ,
         \6028 , \6029 , \6030 , \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 ,
         \6038 , \6039 , \6040 , \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 ,
         \6048 , \6049 , \6050 , \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 ,
         \6058 , \6059 , \6060 , \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 ,
         \6068 , \6069 , \6070 , \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 ,
         \6078 , \6079 , \6080 , \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 ,
         \6088 , \6089 , \6090 , \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 ,
         \6098 , \6099 , \6100 , \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 ,
         \6108 , \6109 , \6110 , \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 ,
         \6118 , \6119 , \6120 , \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 ,
         \6128 , \6129 , \6130 , \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 ,
         \6138 , \6139 , \6140 , \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 ,
         \6148 , \6149 , \6150 , \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 ,
         \6158 , \6159 , \6160 , \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 ,
         \6168 , \6169 , \6170 , \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 ,
         \6178 , \6179 , \6180 , \6181_nGa0e , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 ,
         \6188 , \6189 , \6190 , \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 ,
         \6198 , \6199 , \6200 , \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 ,
         \6208 , \6209 , \6210 , \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 ,
         \6218 , \6219 , \6220 , \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 ,
         \6228 , \6229 , \6230 , \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 ,
         \6238 , \6239 , \6240 , \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 ,
         \6248 , \6249 , \6250 , \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 ,
         \6258 , \6259 , \6260 , \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 ,
         \6268 , \6269 , \6270 , \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 ,
         \6278 , \6279 , \6280 , \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 ,
         \6288 , \6289 , \6290 , \6291 , \6292 , \6293 , \6294 , \6295_nG9d6 , \6296 , \6297 ,
         \6298 , \6299 , \6300 , \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 ,
         \6308 , \6309 , \6310 , \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 ,
         \6318 , \6319 , \6320 , \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 ,
         \6328 , \6329 , \6330 , \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 ,
         \6338 , \6339 , \6340 , \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 ,
         \6348 , \6349 , \6350 , \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 ,
         \6358 , \6359 , \6360 , \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 ,
         \6368 , \6369 , \6370 , \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 ,
         \6378 , \6379 , \6380 , \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 ,
         \6388 , \6389 , \6390 , \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 ,
         \6398 , \6399 , \6400 , \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 ,
         \6408 , \6409 , \6410 , \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 ,
         \6418 , \6419 , \6420 , \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 ,
         \6428 , \6429 , \6430 , \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 ,
         \6438 , \6439 , \6440 , \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 ,
         \6448 , \6449 , \6450 , \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 ,
         \6458 , \6459 , \6460 , \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467_nG99e ,
         \6468 , \6469 , \6470 , \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 ,
         \6478 , \6479 , \6480 , \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 ,
         \6488 , \6489 , \6490 , \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 ,
         \6498 , \6499 , \6500 , \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 ,
         \6508 , \6509 , \6510 , \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 ,
         \6518 , \6519 , \6520 , \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 ,
         \6528 , \6529 , \6530 , \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 ,
         \6538 , \6539 , \6540 , \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 ,
         \6548 , \6549 , \6550 , \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 ,
         \6558 , \6559 , \6560 , \6561 , \6562_nG964 , \6563 , \6564 , \6565 , \6566 , \6567 ,
         \6568 , \6569 , \6570 , \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 ,
         \6578 , \6579 , \6580 , \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 ,
         \6588 , \6589 , \6590 , \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 ,
         \6598 , \6599 , \6600 , \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 ,
         \6608 , \6609 , \6610 , \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 ,
         \6618 , \6619 , \6620 , \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 ,
         \6628 , \6629 , \6630 , \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 ,
         \6638 , \6639 , \6640 , \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 ,
         \6648 , \6649 , \6650 , \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 ,
         \6658 , \6659 , \6660 , \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 ,
         \6668 , \6669 , \6670 , \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 ,
         \6678 , \6679 , \6680 , \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 ,
         \6688 , \6689 , \6690 , \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 ,
         \6698 , \6699 , \6700 , \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 ,
         \6708 , \6709 , \6710 , \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 ,
         \6718 , \6719 , \6720 , \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 ,
         \6728 , \6729 , \6730 , \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 ,
         \6738 , \6739 , \6740 , \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 ,
         \6748 , \6749 , \6750 , \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 ,
         \6758 , \6759 , \6760 , \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 ,
         \6768 , \6769 , \6770 , \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 ,
         \6778 , \6779 , \6780 , \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 ,
         \6788 , \6789 , \6790 , \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 ,
         \6798 , \6799 , \6800 , \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 ,
         \6808 , \6809 , \6810 , \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 ,
         \6818 , \6819 , \6820 , \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 ,
         \6828 , \6829 , \6830 , \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 ,
         \6838 , \6839 , \6840 , \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 ,
         \6848 , \6849 , \6850 , \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 ,
         \6858 , \6859 , \6860 , \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 ,
         \6868 , \6869 , \6870 , \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 ,
         \6878 , \6879 , \6880 , \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 ,
         \6888 , \6889 , \6890 , \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 ,
         \6898 , \6899 , \6900 , \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 ,
         \6908 , \6909 , \6910 , \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 ,
         \6918 , \6919 , \6920 , \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 ,
         \6928 , \6929 , \6930 , \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 ,
         \6938 , \6939 , \6940 , \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 ,
         \6948 , \6949 , \6950 , \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 ,
         \6958 , \6959 , \6960 , \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 ,
         \6968 , \6969 , \6970 , \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 ,
         \6978 , \6979 , \6980 , \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 ,
         \6988 , \6989 , \6990 , \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 ,
         \6998 , \6999 , \7000 , \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 ,
         \7008 , \7009 , \7010 , \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 ,
         \7018 , \7019 , \7020 , \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 ,
         \7028 , \7029 , \7030 , \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 ,
         \7038 , \7039 , \7040 , \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 ,
         \7048 , \7049 , \7050 , \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 ,
         \7058 , \7059 , \7060 , \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 ,
         \7068 , \7069 , \7070 , \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 ,
         \7078 , \7079 , \7080 , \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 ,
         \7088 , \7089 , \7090 , \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 ,
         \7098 , \7099 , \7100 , \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 ,
         \7108 , \7109 , \7110 , \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 ,
         \7118 , \7119 , \7120 , \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 ,
         \7128 , \7129 , \7130 , \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 ,
         \7138 , \7139 , \7140 , \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 ,
         \7148 , \7149 , \7150 , \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 ,
         \7158 , \7159 , \7160 , \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 ,
         \7168 , \7169 , \7170 , \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 ,
         \7178 , \7179 , \7180 , \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 ,
         \7188 , \7189 , \7190 , \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 ,
         \7198 , \7199 , \7200 , \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 ,
         \7208 , \7209 , \7210 , \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 ,
         \7218 , \7219 , \7220 , \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 ,
         \7228 , \7229 , \7230 , \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 ,
         \7238 , \7239 , \7240 , \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 ,
         \7248 , \7249 , \7250 , \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 ,
         \7258 , \7259 , \7260 , \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 ,
         \7268 , \7269 , \7270 , \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 ,
         \7278 , \7279 , \7280 , \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 ,
         \7288 , \7289 , \7290 , \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 ,
         \7298 , \7299 , \7300 , \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 ,
         \7308 , \7309 , \7310 , \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 ,
         \7318 , \7319 , \7320 , \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 ,
         \7328 , \7329 , \7330 , \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 ,
         \7338 , \7339 , \7340 , \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 ,
         \7348 , \7349 , \7350 , \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 ,
         \7358 , \7359 , \7360 , \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 ,
         \7368 , \7369 , \7370 , \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 ,
         \7378 , \7379 , \7380 , \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 ,
         \7388 , \7389 , \7390 , \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 ,
         \7398 , \7399 , \7400 , \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407_nG4e5 ,
         \7408 , \7409 , \7410_nG506 , \7411 , \7412 , \7413 , \7414_nG5c2 , \7415 , \7416 , \7417 ,
         \7418_nG5c4 , \7419 , \7420 , \7421 , \7422_nG5e3 , \7423 , \7424 , \7425_nG5e5 , \7426 , \7427 ,
         \7428 , \7429 , \7430_nG5a5 , \7431 , \7432 , \7433 , \7434_nG5a3 , \7435 , \7436 , \7437 ,
         \7438 , \7439_nG586 , \7440 , \7441 , \7442 , \7443 , \7444 , \7445_nG584 , \7446 , \7447 ,
         \7448 , \7449_nG567 , \7450 , \7451 , \7452_nG565 , \7453 , \7454 , \7455 , \7456 , \7457 ,
         \7458_nG546 , \7459 , \7460 , \7461 , \7462 , \7463 , \7464_nG544 , \7465 , \7466 , \7467 ,
         \7468_nG527 , \7469 , \7470 , \7471_nG525 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 ,
         \7478 , \7479 , \7480_nG504 , \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487_nG4e3 ,
         \7488 , \7489 , \7490 , \7491_nG4c4 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497_nG4c2 ,
         \7498 , \7499 , \7500 , \7501_nG4a3 , \7502 , \7503 , \7504_nG4a1 , \7505 , \7506 , \7507 ,
         \7508 , \7509 , \7510_nG484 , \7511 , \7512 , \7513 , \7514 , \7515 , \7516_nG482 , \7517 ,
         \7518 , \7519 , \7520_nG465 , \7521 , \7522 , \7523_nG462 , \7524 , \7525 , \7526 , \7527 ,
         \7528 , \7529 , \7530 , \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 ,
         \7538 , \7539 , \7540 , \7541 , \7542 , \7543 , \7544 , \7545 , \7546_nG301 , \7547 ,
         \7548 , \7549 , \7550 , \7551_nG33a , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 ,
         \7558 , \7559 , \7560 , \7561 , \7562_nG357 , \7563 , \7564 , \7565 , \7566 , \7567 ,
         \7568 , \7569 , \7570_nG391 , \7571 , \7572 , \7573_nG3ae , \7574 , \7575 , \7576 , \7577_nG3cb ,
         \7578 , \7579 , \7580 , \7581 , \7582 , \7583 , \7584_nG3e8 , \7585 , \7586 , \7587_nG405 ,
         \7588 , \7589 , \7590 , \7591 , \7592 , \7593 , \7594_nG422 , \7595 , \7596_nG43e , \7597 ,
         \7598 , \7599 , \7600 , \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 ,
         \7608 , \7609 , \7610 , \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 ,
         \7618 , \7619 , \7620 , \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 ,
         \7628 , \7629 , \7630 , \7631 , \7632_nG374 , \7633 , \7634 , \7635 , \7636 , \7637 ,
         \7638 , \7639 , \7640 , \7641 , \7642 , \7643 , \7644 , \7645 , \7646_nG31e , \7647 ,
         \7648 , \7649 , \7650 , \7651 , \7652_nG2e4 , \7653 , \7654 , \7655 , \7656 , \7657 ,
         \7658 , \7659 , \7660 , \7661 , \7662 , \7663 , \7664 , \7665_nG21fd , \7666 , \7667 ,
         \7668 , \7669 , \7670_nG21c3 , \7671 , \7672 , \7673 , \7674 , \7675 , \7676_nG2194 , \7677 ,
         \7678 , \7679 , \7680 , \7681 , \7682_nG215b , \7683 , \7684 , \7685 , \7686 , \7687 ,
         \7688_nG20f7 , \7689 , \7690 , \7691 , \7692 , \7693 , \7694_nG208a , \7695 , \7696 , \7697 ,
         \7698 , \7699 , \7700_nG2017 , \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707_nG1f99 ,
         \7708 , \7709 , \7710 , \7711 , \7712 , \7713 , \7714 , \7715 , \7716_nG1eee , \7717 ,
         \7718 , \7719 , \7720 , \7721 , \7722 , \7723 , \7724 , \7725 , \7726_nG1e36 , \7727 ,
         \7728 , \7729 , \7730 , \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 ,
         \7738 , \7739 , \7740 , \7741 , \7742_nG1d83 , \7743 , \7744 , \7745 , \7746 , \7747 ,
         \7748_nG1ca7 , \7749 , \7750 , \7751 , \7752 , \7753 , \7754 , \7755 , \7756_nG1bcd , \7757 ,
         \7758 , \7759 , \7760 , \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 ,
         \7768 , \7769 , \7770 , \7771 , \7772_nG1af9 , \7773 , \7774 , \7775 , \7776 , \7777 ,
         \7778_nG19e9 , \7779 , \7780 , \7781 , \7782 , \7783 , \7784_nG18d0 , \7785 , \7786 , \7787 ,
         \7788 , \7789 , \7790 , \7791_nG17c2 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 ,
         \7798 , \7799 , \7800 , \7801 , \7802 , \7803_nG16bb , \7804 , \7805 , \7806 , \7807 ,
         \7808 , \7809 , \7810 , \7811 , \7812 , \7813 , \7814 , \7815_nG1596 , \7816 , \7817 ,
         \7818 , \7819 , \7820 , \7821 , \7822 , \7823 , \7824 , \7825 , \7826 , \7827 ,
         \7828 , \7829 , \7830 , \7831_nG14ad , \7832 , \7833 , \7834 , \7835 , \7836 , \7837_nG13ad ,
         \7838 , \7839 , \7840 , \7841 , \7842 , \7843_nG12ae , \7844 , \7845 , \7846 , \7847 ,
         \7848 , \7849_nG11a4 , \7850 , \7851 , \7852 , \7853 , \7854 , \7855_nG10c7 , \7856 , \7857 ,
         \7858 , \7859 , \7860 , \7861_nGfc2 , \7862 , \7863 , \7864 , \7865 , \7866 , \7867_nGeed ,
         \7868 , \7869 , \7870 , \7871 , \7872 , \7873_nGe16 , \7874 , \7875 , \7876 , \7877 ,
         \7878 , \7879 , \7880 , \7881 , \7882 , \7883 , \7884 , \7885 , \7886 , \7887 ,
         \7888 , \7889 , \7890 , \7891 , \7892 , \7893 , \7894 , \7895 , \7896 , \7897 ,
         \7898 , \7899 , \7900 , \7901 , \7902 , \7903 , \7904 , \7905 , \7906 , \7907 ,
         \7908 , \7909 , \7910 , \7911 , \7912 , \7913 , \7914 , \7915 , \7916 , \7917 ,
         \7918 , \7919 , \7920 , \7921 , \7922 , \7923 , \7924 , \7925 , \7926 , \7927 ,
         \7928 , \7929 , \7930 , \7931 , \7932 , \7933 , \7934 , \7935 , \7936 , \7937 ,
         \7938 , \7939 , \7940 , \7941 , \7942 , \7943 , \7944 , \7945 , \7946 , \7947 ,
         \7948 , \7949 , \7950 , \7951 , \7952 , \7953 , \7954 , \7955 , \7956 , \7957 ,
         \7958 , \7959 , \7960 , \7961 , \7962 , \7963 , \7964 , \7965 , \7966 , \7967 ,
         \7968 , \7969 , \7970 , \7971 , \7972 , \7973 , \7974_nG2a78 , \7975 , \7976 , \7977 ,
         \7978 , \7979 , \7980 , \7981 , \7982 , \7983 , \7984 , \7985 , \7986 , \7987 ,
         \7988 , \7989 , \7990 , \7991 , \7992 , \7993 , \7994 , \7995 , \7996 , \7997 ,
         \7998 , \7999 , \8000 , \8001 , \8002 , \8003 , \8004 , \8005 , \8006 , \8007 ,
         \8008 , \8009 , \8010 , \8011 , \8012_nG2898 , \8013 , \8014 , \8015 , \8016 , \8017 ,
         \8018 , \8019 , \8020 , \8021 , \8022 , \8023 , \8024 , \8025 , \8026 , \8027 ,
         \8028 , \8029 , \8030 , \8031 , \8032 , \8033 , \8034 , \8035 , \8036 , \8037 ,
         \8038 , \8039 , \8040 , \8041 , \8042 , \8043 , \8044 , \8045 , \8046 , \8047 ,
         \8048 , \8049 , \8050_nG2896 , \8051 , \8052 , \8053 , \8054 , \8055 , \8056 , \8057 ,
         \8058 , \8059 , \8060 , \8061 , \8062 , \8063 , \8064 , \8065 , \8066 , \8067 ,
         \8068 , \8069 , \8070 , \8071 , \8072 , \8073 , \8074 , \8075 , \8076 , \8077 ,
         \8078 , \8079 , \8080 , \8081 , \8082 , \8083 , \8084 , \8085 , \8086 , \8087 ,
         \8088_nG26eb , \8089 , \8090 , \8091 , \8092 , \8093 , \8094 , \8095 , \8096 , \8097 ,
         \8098 , \8099 , \8100 , \8101 , \8102 , \8103 , \8104 , \8105 , \8106 , \8107 ,
         \8108 , \8109 , \8110 , \8111 , \8112 , \8113 , \8114 , \8115 , \8116 , \8117 ,
         \8118 , \8119 , \8120 , \8121 , \8122 , \8123 , \8124_nG26e9 , \8125 , \8126 , \8127 ,
         \8128 , \8129 , \8130 , \8131 , \8132 , \8133 , \8134 , \8135 , \8136 , \8137 ,
         \8138 , \8139 , \8140 , \8141 , \8142 , \8143 , \8144 , \8145 , \8146 , \8147 ,
         \8148 , \8149 , \8150 , \8151 , \8152 , \8153 , \8154 , \8155 , \8156 , \8157 ,
         \8158 , \8159 , \8160 , \8161 , \8162_nG2358 , \8163 , \8164 , \8165 , \8166 , \8167 ,
         \8168 , \8169 , \8170 , \8171 , \8172 , \8173 , \8174 , \8175 , \8176 , \8177 ,
         \8178 , \8179 , \8180 , \8181 , \8182 , \8183 , \8184 , \8185 , \8186 , \8187 ,
         \8188 , \8189 , \8190 , \8191 , \8192 , \8193 , \8194 , \8195 , \8196 , \8197 ,
         \8198_nG2356 , \8199 , \8200 , \8201 , \8202 , \8203 , \8204 , \8205 , \8206 , \8207 ,
         \8208 , \8209 , \8210 , \8211 , \8212 , \8213 , \8214 , \8215 , \8216 , \8217 ,
         \8218 , \8219 , \8220 , \8221 , \8222 , \8223 , \8224 , \8225 , \8226 , \8227 ,
         \8228 , \8229 , \8230 , \8231 , \8232 , \8233 , \8234_nG22e8 , \8235 , \8236 , \8237 ,
         \8238 , \8239 , \8240 , \8241 , \8242 , \8243 , \8244 , \8245 , \8246 , \8247 ,
         \8248 , \8249 , \8250 , \8251 , \8252 , \8253 , \8254 , \8255 , \8256 , \8257 ,
         \8258 , \8259 , \8260 , \8261 , \8262 , \8263 , \8264 , \8265 , \8266 , \8267 ,
         \8268 , \8269 , \8270_nG22e6 , \8271 , \8272 , \8273 , \8274 , \8275 , \8276 , \8277 ,
         \8278 , \8279 , \8280 , \8281 , \8282 , \8283 , \8284 , \8285 , \8286 , \8287 ,
         \8288 , \8289 , \8290 , \8291 , \8292 , \8293 , \8294 , \8295 , \8296 , \8297 ,
         \8298 , \8299 , \8300 , \8301 , \8302_nG2290 , \8303 , \8304 , \8305 , \8306 , \8307 ,
         \8308 , \8309 , \8310 , \8311 , \8312 , \8313 , \8314 , \8315 , \8316 , \8317 ,
         \8318 , \8319 , \8320 , \8321 , \8322 , \8323 , \8324 , \8325 , \8326 , \8327 ,
         \8328 , \8329 , \8330 , \8331 , \8332 , \8333 , \8334 , \8335 , \8336 , \8337 ,
         \8338_nG2292 , \8339 , \8340 , \8341 , \8342 , \8343 , \8344 , \8345 , \8346 , \8347 ,
         \8348 , \8349 , \8350 , \8351 , \8352 , \8353 , \8354 , \8355 , \8356 , \8357 ,
         \8358 , \8359 , \8360 , \8361 , \8362 , \8363 , \8364 , \8365 , \8366 , \8367 ,
         \8368 , \8369 , \8370 , \8371_nG221f , \8372 , \8373 , \8374 , \8375 , \8376 , \8377 ,
         \8378 , \8379 , \8380 , \8381 , \8382 , \8383 , \8384 , \8385 , \8386 , \8387 ,
         \8388 , \8389 , \8390 , \8391 , \8392 , \8393 , \8394 , \8395 , \8396 , \8397 ,
         \8398 , \8399 , \8400 , \8401 , \8402_nG221d , \8403 , \8404 , \8405 , \8406 , \8407 ,
         \8408 , \8409 , \8410 , \8411 , \8412 , \8413 , \8414 , \8415 , \8416 , \8417 ,
         \8418 , \8419 , \8420 , \8421 , \8422 , \8423 , \8424 , \8425 , \8426 , \8427 ,
         \8428 , \8429 , \8430 , \8431 , \8432 , \8433 , \8434 , \8435 , \8436 , \8437 ,
         \8438 , \8439 , \8440 , \8441 , \8442 , \8443 , \8444 , \8445 , \8446 , \8447 ,
         \8448 , \8449 , \8450 , \8451 , \8452 , \8453 , \8454 , \8455 , \8456 , \8457 ,
         \8458 , \8459 , \8460 , \8461 , \8462 , \8463 , \8464 , \8465 , \8466 , \8467 ,
         \8468 , \8469 , \8470 , \8471 , \8472 , \8473 , \8474_nG30a2 , \8475 , \8476 , \8477 ,
         \8478 , \8479 , \8480 , \8481 , \8482 , \8483 , \8484 , \8485 , \8486 , \8487 ,
         \8488 , \8489 , \8490 , \8491 , \8492 , \8493 , \8494 , \8495 , \8496 , \8497 ,
         \8498 , \8499 , \8500 , \8501 , \8502 , \8503 , \8504 , \8505 , \8506 , \8507 ,
         \8508 , \8509 , \8510 , \8511 , \8512 , \8513 , \8514_nG31b0 , \8515 , \8516 , \8517 ,
         \8518 , \8519 , \8520 , \8521 , \8522 , \8523 , \8524 , \8525 , \8526 , \8527 ,
         \8528 , \8529 , \8530 , \8531 , \8532 , \8533 , \8534 , \8535 , \8536 , \8537 ,
         \8538 , \8539 , \8540 , \8541 , \8542 , \8543 , \8544 , \8545 , \8546 , \8547 ,
         \8548 , \8549 , \8550 , \8551 , \8552 , \8553 , \8554 , \8555 , \8556 , \8557 ,
         \8558 , \8559 , \8560 , \8561 , \8562 , \8563 , \8564 , \8565 , \8566 , \8567 ,
         \8568_nG2f9c , \8569 , \8570 , \8571 , \8572 , \8573 , \8574 , \8575 , \8576 , \8577 ,
         \8578 , \8579 , \8580 , \8581 , \8582 , \8583 , \8584 , \8585 , \8586 , \8587 ,
         \8588 , \8589 , \8590 , \8591 , \8592 , \8593 , \8594 , \8595 , \8596 , \8597 ,
         \8598 , \8599 , \8600 , \8601 , \8602 , \8603 , \8604 , \8605 , \8606 , \8607 ,
         \8608 , \8609 , \8610 , \8611 , \8612 , \8613 , \8614 , \8615 , \8616 , \8617 ,
         \8618 , \8619 , \8620 , \8621 , \8622 , \8623 , \8624 , \8625 , \8626 , \8627 ,
         \8628 , \8629 , \8630 , \8631 , \8632 , \8633 , \8634 , \8635 , \8636 , \8637 ,
         \8638 , \8639 , \8640 , \8641 , \8642 , \8643 , \8644 , \8645 , \8646 , \8647 ,
         \8648 , \8649 , \8650 , \8651 , \8652 , \8653 , \8654 , \8655 , \8656 , \8657_nG2e7a ,
         \8658 , \8659 , \8660 , \8661 , \8662 , \8663 , \8664 , \8665 , \8666 , \8667 ,
         \8668 , \8669 , \8670 , \8671 , \8672 , \8673 , \8674 , \8675 , \8676 , \8677 ,
         \8678 , \8679 , \8680 , \8681 , \8682 , \8683 , \8684 , \8685 , \8686 , \8687 ,
         \8688 , \8689 , \8690 , \8691 , \8692 , \8693 , \8694 , \8695 , \8696 , \8697 ,
         \8698 , \8699 , \8700 , \8701 , \8702 , \8703 , \8704 , \8705 , \8706 , \8707 ,
         \8708 , \8709 , \8710 , \8711 , \8712 , \8713 , \8714 , \8715 , \8716 , \8717 ,
         \8718 , \8719 , \8720 , \8721 , \8722 , \8723 , \8724 , \8725 , \8726 , \8727 ,
         \8728 , \8729_nG2d90 , \8730 , \8731 , \8732 , \8733 , \8734 , \8735 , \8736 , \8737 ,
         \8738 , \8739 , \8740 , \8741 , \8742 , \8743 , \8744 , \8745 , \8746 , \8747 ,
         \8748 , \8749 , \8750 , \8751 , \8752 , \8753 , \8754 , \8755 , \8756 , \8757 ,
         \8758 , \8759 , \8760 , \8761 , \8762_nG2c8f , \8763 , \8764 , \8765 , \8766 , \8767 ,
         \8768 , \8769 , \8770 , \8771 , \8772 , \8773 , \8774 , \8775 , \8776 , \8777 ,
         \8778 , \8779 , \8780 , \8781 , \8782 , \8783 , \8784 , \8785 , \8786 , \8787 ,
         \8788 , \8789 , \8790 , \8791 , \8792 , \8793 , \8794 , \8795 , \8796 , \8797 ,
         \8798 , \8799 , \8800 , \8801 , \8802 , \8803 , \8804 , \8805 , \8806 , \8807 ,
         \8808 , \8809 , \8810 , \8811 , \8812 , \8813 , \8814 , \8815 , \8816 , \8817 ,
         \8818 , \8819 , \8820 , \8821 , \8822 , \8823 , \8824 , \8825 , \8826 , \8827 ,
         \8828 , \8829 , \8830 , \8831 , \8832 , \8833 , \8834 , \8835 , \8836 , \8837 ,
         \8838 , \8839 , \8840 , \8841 , \8842 , \8843 , \8844 , \8845 , \8846 , \8847 ,
         \8848 , \8849 , \8850 , \8851 , \8852 , \8853 , \8854 , \8855 , \8856 , \8857 ,
         \8858 , \8859 , \8860 , \8861 , \8862 , \8863 , \8864 , \8865 , \8866 , \8867 ,
         \8868_nG2b9c , \8869 , \8870 , \8871 , \8872 , \8873 , \8874 , \8875 , \8876 , \8877 ,
         \8878 , \8879 , \8880 , \8881 , \8882 , \8883 , \8884 , \8885 , \8886 , \8887 ,
         \8888 , \8889 , \8890 , \8891 , \8892 , \8893 , \8894 , \8895 , \8896 , \8897 ,
         \8898 , \8899 , \8900 , \8901 , \8902 , \8903 , \8904 , \8905 , \8906 , \8907 ,
         \8908 , \8909 , \8910 , \8911 , \8912 , \8913 , \8914 , \8915 , \8916 , \8917 ,
         \8918 , \8919 , \8920 , \8921 , \8922 , \8923 , \8924 , \8925 , \8926 , \8927 ,
         \8928 , \8929 , \8930 , \8931 , \8932 , \8933 , \8934 , \8935 , \8936 , \8937 ,
         \8938 , \8939 , \8940 , \8941 , \8942 , \8943 , \8944 , \8945 , \8946 , \8947_nG2a93 ,
         \8948 , \8949 , \8950 , \8951 , \8952 , \8953 , \8954 , \8955 , \8956 , \8957 ,
         \8958 , \8959 , \8960 , \8961 , \8962 , \8963 , \8964 , \8965 , \8966 , \8967 ,
         \8968 , \8969 , \8970 , \8971 , \8972 , \8973 , \8974 , \8975 , \8976 , \8977 ,
         \8978 , \8979 , \8980 , \8981 , \8982 , \8983 , \8984 , \8985 , \8986 , \8987 ,
         \8988 , \8989 , \8990 , \8991 , \8992 , \8993 , \8994 , \8995 , \8996 , \8997 ,
         \8998 , \8999 , \9000 , \9001 , \9002 , \9003 , \9004 , \9005 , \9006 , \9007 ,
         \9008 , \9009 , \9010 , \9011 , \9012 , \9013 , \9014 , \9015 , \9016 , \9017 ,
         \9018_nG29b3 , \9019 , \9020 , \9021 , \9022 , \9023 , \9024 , \9025 , \9026 , \9027 ,
         \9028 , \9029 , \9030 , \9031 , \9032 , \9033 , \9034 , \9035 , \9036 , \9037 ,
         \9038 , \9039 , \9040 , \9041 , \9042 , \9043 , \9044 , \9045 , \9046 , \9047 ,
         \9048 , \9049 , \9050 , \9051 , \9052 , \9053 , \9054 , \9055 , \9056 , \9057 ,
         \9058 , \9059 , \9060 , \9061 , \9062 , \9063 , \9064 , \9065 , \9066 , \9067 ,
         \9068 , \9069 , \9070 , \9071 , \9072 , \9073 , \9074 , \9075 , \9076 , \9077 ,
         \9078 , \9079 , \9080 , \9081 , \9082 , \9083 , \9084 , \9085 , \9086 , \9087 ,
         \9088 , \9089 , \9090 , \9091 , \9092 , \9093 , \9094 , \9095 , \9096 , \9097 ,
         \9098 , \9099 , \9100 , \9101 , \9102 , \9103 , \9104 , \9105 , \9106 , \9107 ,
         \9108 , \9109 , \9110 , \9111 , \9112 , \9113 , \9114 , \9115 , \9116 , \9117 ,
         \9118 , \9119 , \9120 , \9121 , \9122 , \9123 , \9124 , \9125 , \9126 , \9127 ,
         \9128 , \9129 , \9130 , \9131 , \9132 , \9133 , \9134 , \9135 , \9136 , \9137 ,
         \9138 , \9139 , \9140 , \9141 , \9142 , \9143 , \9144 , \9145 , \9146 , \9147 ,
         \9148 , \9149 , \9150 , \9151 , \9152 , \9153 , \9154 , \9155 , \9156 , \9157 ,
         \9158 , \9159 , \9160 , \9161 , \9162 , \9163 , \9164 , \9165 , \9166 , \9167 ,
         \9168 , \9169 , \9170 , \9171 , \9172 , \9173 , \9174 , \9175 , \9176 , \9177 ,
         \9178 , \9179 , \9180 , \9181 , \9182 , \9183 , \9184 , \9185 , \9186 , \9187 ,
         \9188 , \9189 , \9190 , \9191 , \9192 , \9193 , \9194 , \9195 , \9196 , \9197 ,
         \9198 , \9199 , \9200 , \9201 , \9202 , \9203 , \9204 , \9205 , \9206 , \9207 ,
         \9208 , \9209 , \9210 , \9211 , \9212 , \9213 , \9214 , \9215 , \9216 , \9217 ,
         \9218 , \9219 , \9220 , \9221 , \9222 , \9223 , \9224 , \9225 , \9226 , \9227 ,
         \9228 , \9229 , \9230 , \9231 , \9232 , \9233 , \9234 , \9235 , \9236 , \9237 ,
         \9238 , \9239 , \9240 , \9241 , \9242 , \9243 , \9244 , \9245 , \9246 , \9247 ,
         \9248 , \9249 , \9250 , \9251 , \9252 , \9253 , \9254 , \9255 , \9256 , \9257 ,
         \9258 , \9259 , \9260_nG28b3 , \9261 , \9262 , \9263 , \9264 , \9265 , \9266 , \9267 ,
         \9268 , \9269 , \9270 , \9271 , \9272 , \9273 , \9274 , \9275 , \9276 , \9277 ,
         \9278 , \9279 , \9280 , \9281 , \9282 , \9283 , \9284 , \9285 , \9286 , \9287 ,
         \9288 , \9289 , \9290 , \9291 , \9292 , \9293 , \9294 , \9295 , \9296 , \9297 ,
         \9298 , \9299 , \9300 , \9301 , \9302 , \9303 , \9304 , \9305 , \9306 , \9307 ,
         \9308 , \9309 , \9310 , \9311 , \9312 , \9313 , \9314 , \9315 , \9316 , \9317_nG27da ,
         \9318 , \9319 , \9320 , \9321 , \9322 , \9323 , \9324 , \9325 , \9326 , \9327 ,
         \9328 , \9329 , \9330 , \9331 , \9332 , \9333 , \9334 , \9335 , \9336 , \9337 ,
         \9338 , \9339 , \9340 , \9341 , \9342 , \9343 , \9344 , \9345 , \9346 , \9347 ,
         \9348 , \9349 , \9350 , \9351 , \9352 , \9353 , \9354 , \9355 , \9356 , \9357 ,
         \9358 , \9359 , \9360 , \9361 , \9362 , \9363 , \9364 , \9365 , \9366 , \9367 ,
         \9368 , \9369 , \9370 , \9371 , \9372 , \9373 , \9374 , \9375 , \9376 , \9377 ,
         \9378 , \9379 , \9380 , \9381 , \9382 , \9383 , \9384 , \9385 , \9386 , \9387 ,
         \9388 , \9389 , \9390 , \9391 , \9392 , \9393 , \9394 , \9395 , \9396 , \9397 ,
         \9398 , \9399 , \9400 , \9401 , \9402 , \9403 , \9404 , \9405 , \9406 , \9407 ,
         \9408 , \9409 , \9410 , \9411 , \9412 , \9413 , \9414 , \9415 , \9416 , \9417 ,
         \9418 , \9419 , \9420 , \9421 , \9422 , \9423 , \9424 , \9425 , \9426 , \9427 ,
         \9428 , \9429 , \9430 , \9431 , \9432 , \9433 , \9434 , \9435 , \9436 , \9437 ,
         \9438 , \9439 , \9440 , \9441 , \9442 , \9443 , \9444 , \9445 , \9446 , \9447 ,
         \9448 , \9449 , \9450 , \9451 , \9452 , \9453 , \9454 , \9455 , \9456 , \9457 ,
         \9458 , \9459 , \9460 , \9461 , \9462 , \9463 , \9464 , \9465 , \9466 , \9467 ,
         \9468 , \9469 , \9470 , \9471 , \9472 , \9473 , \9474 , \9475 , \9476 , \9477 ,
         \9478 , \9479 , \9480 , \9481_nG2706 , \9482 , \9483 , \9484 , \9485 , \9486 , \9487 ,
         \9488 , \9489 , \9490 , \9491 , \9492 , \9493 , \9494 , \9495 , \9496 , \9497 ,
         \9498 , \9499 , \9500 , \9501 , \9502 , \9503 , \9504 , \9505 , \9506 , \9507 ,
         \9508 , \9509 , \9510 , \9511 , \9512 , \9513 , \9514 , \9515 , \9516 , \9517 ,
         \9518 , \9519 , \9520 , \9521 , \9522 , \9523 , \9524 , \9525 , \9526 , \9527 ,
         \9528 , \9529 , \9530 , \9531 , \9532 , \9533 , \9534 , \9535 , \9536 , \9537 ,
         \9538 , \9539 , \9540 , \9541 , \9542 , \9543 , \9544 , \9545 , \9546 , \9547 ,
         \9548 , \9549 , \9550 , \9551 , \9552 , \9553 , \9554 , \9555 , \9556 , \9557 ,
         \9558 , \9559 , \9560 , \9561 , \9562 , \9563_nG23ac , \9564 , \9565 , \9566 , \9567 ,
         \9568 , \9569 , \9570 , \9571 , \9572 , \9573 , \9574 , \9575 , \9576 , \9577 ,
         \9578 , \9579 , \9580 , \9581 , \9582 , \9583 , \9584 , \9585 , \9586 , \9587 ,
         \9588 , \9589 , \9590 , \9591 , \9592 , \9593 , \9594 , \9595 , \9596 , \9597 ,
         \9598 , \9599 , \9600 , \9601 , \9602 , \9603 , \9604 , \9605 , \9606 , \9607 ,
         \9608 , \9609 , \9610 , \9611 , \9612 , \9613 , \9614 , \9615 , \9616 , \9617 ,
         \9618 , \9619 , \9620 , \9621 , \9622 , \9623 , \9624 , \9625 , \9626 , \9627 ,
         \9628 , \9629 , \9630 , \9631 , \9632 , \9633 , \9634 , \9635 , \9636 , \9637 ,
         \9638 , \9639 , \9640 , \9641 , \9642 , \9643 , \9644 , \9645 , \9646 , \9647 ,
         \9648 , \9649 , \9650 , \9651 , \9652 , \9653 , \9654 , \9655 , \9656 , \9657 ,
         \9658 , \9659 , \9660_nG2373 , \9661 , \9662 , \9663 , \9664 , \9665 , \9666 , \9667 ,
         \9668 , \9669 , \9670 , \9671 , \9672 , \9673 , \9674 , \9675 , \9676 , \9677 ,
         \9678 , \9679 , \9680 , \9681 , \9682 , \9683 , \9684 , \9685 , \9686 , \9687 ,
         \9688 , \9689 , \9690 , \9691 , \9692 , \9693 , \9694 , \9695 , \9696 , \9697 ,
         \9698 , \9699 , \9700 , \9701 , \9702 , \9703 , \9704 , \9705 , \9706 , \9707 ,
         \9708 , \9709 , \9710 , \9711 , \9712 , \9713 , \9714 , \9715 , \9716 , \9717 ,
         \9718 , \9719 , \9720 , \9721 , \9722 , \9723 , \9724 , \9725 , \9726 , \9727 ,
         \9728 , \9729 , \9730 , \9731 , \9732 , \9733 , \9734 , \9735 , \9736 , \9737 ,
         \9738 , \9739 , \9740 , \9741 , \9742 , \9743 , \9744 , \9745 , \9746 , \9747 ,
         \9748 , \9749 , \9750 , \9751 , \9752 , \9753 , \9754 , \9755 , \9756 , \9757 ,
         \9758 , \9759 , \9760 , \9761 , \9762 , \9763 , \9764 , \9765 , \9766 , \9767 ,
         \9768 , \9769 , \9770 , \9771 , \9772 , \9773 , \9774 , \9775 , \9776 , \9777 ,
         \9778 , \9779 , \9780 , \9781 , \9782 , \9783 , \9784 , \9785 , \9786 , \9787 ,
         \9788 , \9789 , \9790 , \9791 , \9792 , \9793 , \9794 , \9795 , \9796 , \9797 ,
         \9798 , \9799 , \9800 , \9801 , \9802 , \9803 , \9804 , \9805 , \9806 , \9807 ,
         \9808 , \9809 , \9810 , \9811 , \9812 , \9813 , \9814 , \9815 , \9816 , \9817 ,
         \9818 , \9819 , \9820 , \9821 , \9822 , \9823 , \9824 , \9825 , \9826 , \9827 ,
         \9828 , \9829 , \9830 , \9831 , \9832 , \9833 , \9834 , \9835 , \9836 , \9837 ,
         \9838 , \9839 , \9840 , \9841 , \9842 , \9843 , \9844 , \9845 , \9846 , \9847 ,
         \9848 , \9849 , \9850 , \9851 , \9852 , \9853 , \9854 , \9855 , \9856 , \9857 ,
         \9858 , \9859 , \9860 , \9861 , \9862 , \9863 , \9864 , \9865 , \9866 , \9867 ,
         \9868_nG2303 , \9869 , \9870 , \9871 , \9872 , \9873 , \9874 , \9875 , \9876 , \9877 ,
         \9878 , \9879 , \9880 , \9881 , \9882 , \9883 , \9884 , \9885 , \9886 , \9887 ,
         \9888 , \9889 , \9890 , \9891 , \9892 , \9893 , \9894 , \9895 , \9896 , \9897 ,
         \9898_nG233b , \9899 , \9900 , \9901 , \9902 , \9903 , \9904 , \9905 , \9906 , \9907 ,
         \9908 , \9909 , \9910 , \9911 , \9912 , \9913 , \9914 , \9915 , \9916 , \9917 ,
         \9918 , \9919 , \9920 , \9921 , \9922 , \9923 , \9924 , \9925 , \9926 , \9927 ,
         \9928 , \9929 , \9930 , \9931 , \9932 , \9933 , \9934 , \9935 , \9936 , \9937 ,
         \9938 , \9939 , \9940 , \9941 , \9942 , \9943 , \9944 , \9945 , \9946 , \9947 ,
         \9948 , \9949 , \9950 , \9951 , \9952 , \9953 , \9954 , \9955 , \9956 , \9957 ,
         \9958 , \9959 , \9960 , \9961 , \9962 , \9963 , \9964 , \9965 , \9966 , \9967 ,
         \9968 , \9969 , \9970 , \9971 , \9972 , \9973 , \9974 , \9975 , \9976 , \9977 ,
         \9978 , \9979 , \9980 , \9981 , \9982 , \9983 , \9984 , \9985 , \9986 , \9987 ,
         \9988 , \9989 , \9990 , \9991 , \9992 , \9993 , \9994 , \9995 , \9996 , \9997 ,
         \9998 , \9999 , \10000 , \10001 , \10002 , \10003 , \10004 , \10005 , \10006 , \10007 ,
         \10008 , \10009 , \10010 , \10011 , \10012 , \10013 , \10014 , \10015 , \10016 , \10017 ,
         \10018 , \10019 , \10020 , \10021 , \10022 , \10023 , \10024 , \10025 , \10026 , \10027 ,
         \10028 , \10029 , \10030 , \10031 , \10032 , \10033 , \10034 , \10035 , \10036 , \10037 ,
         \10038 , \10039 , \10040 , \10041 , \10042 , \10043 , \10044 , \10045 , \10046 , \10047 ,
         \10048 , \10049 , \10050 , \10051 , \10052 , \10053 , \10054 , \10055 , \10056 , \10057 ,
         \10058 , \10059 , \10060 , \10061 , \10062 , \10063 , \10064 , \10065 , \10066 , \10067 ,
         \10068 , \10069 , \10070 , \10071 , \10072 , \10073 , \10074 , \10075 , \10076 , \10077 ,
         \10078 , \10079 , \10080 , \10081 , \10082 , \10083 , \10084 , \10085 , \10086 , \10087 ,
         \10088 , \10089 , \10090 , \10091 , \10092 , \10093 , \10094 , \10095 , \10096 , \10097 ,
         \10098 , \10099 , \10100 , \10101 , \10102 , \10103 , \10104 , \10105 , \10106 , \10107 ,
         \10108 , \10109 , \10110 , \10111 , \10112 , \10113 , \10114 , \10115 , \10116 , \10117 ,
         \10118 , \10119_nG22ca , \10120 , \10121 , \10122 , \10123 , \10124 , \10125 , \10126 , \10127 ,
         \10128 , \10129 , \10130 , \10131 , \10132 , \10133 , \10134 , \10135 , \10136 , \10137 ,
         \10138 , \10139 , \10140 , \10141 , \10142 , \10143 , \10144 , \10145 , \10146 , \10147 ,
         \10148 , \10149 , \10150 , \10151 , \10152 , \10153 , \10154 , \10155 , \10156 , \10157 ,
         \10158 , \10159 , \10160 , \10161 , \10162 , \10163 , \10164 , \10165 , \10166 , \10167 ,
         \10168 , \10169 , \10170 , \10171 , \10172 , \10173 , \10174 , \10175 , \10176 , \10177 ,
         \10178 , \10179 , \10180 , \10181 , \10182 , \10183 , \10184 , \10185 , \10186 , \10187 ,
         \10188 , \10189 , \10190 , \10191 , \10192 , \10193 , \10194 , \10195 , \10196 , \10197 ,
         \10198 , \10199 , \10200 , \10201 , \10202 , \10203 , \10204 , \10205 , \10206 , \10207 ,
         \10208 , \10209 , \10210 , \10211 , \10212 , \10213 , \10214 , \10215 , \10216 , \10217 ,
         \10218 , \10219 , \10220 , \10221 , \10222 , \10223 , \10224 , \10225 , \10226 , \10227 ,
         \10228 , \10229 , \10230 , \10231 , \10232 , \10233 , \10234 , \10235_nG228e , \10236 , \10237 ,
         \10238 , \10239 , \10240 , \10241 , \10242 , \10243 , \10244 , \10245 , \10246 , \10247 ,
         \10248 , \10249 , \10250 , \10251 , \10252 , \10253 , \10254 , \10255 , \10256 , \10257 ,
         \10258 , \10259 , \10260 , \10261 , \10262 , \10263 , \10264 , \10265 , \10266 , \10267 ,
         \10268 , \10269 , \10270 , \10271 , \10272 , \10273 , \10274 , \10275 , \10276 , \10277 ,
         \10278 , \10279 , \10280 , \10281 , \10282 , \10283 , \10284 , \10285 , \10286 , \10287 ,
         \10288 , \10289 , \10290 , \10291 , \10292 , \10293 , \10294 , \10295 , \10296 , \10297 ,
         \10298 , \10299 , \10300 , \10301 , \10302 , \10303 , \10304 , \10305 , \10306 , \10307 ,
         \10308 , \10309 , \10310 , \10311 , \10312 , \10313 , \10314 , \10315 , \10316 , \10317 ,
         \10318 , \10319 , \10320 , \10321 , \10322 , \10323 , \10324 , \10325 , \10326 , \10327 ,
         \10328 , \10329 , \10330 , \10331 , \10332 , \10333 , \10334 , \10335 , \10336 , \10337 ,
         \10338 , \10339 , \10340 , \10341 , \10342 , \10343 , \10344 , \10345 , \10346 , \10347 ,
         \10348 , \10349 , \10350 , \10351 , \10352 , \10353 , \10354 , \10355 , \10356 , \10357 ,
         \10358 , \10359 , \10360 , \10361 , \10362 , \10363 , \10364 , \10365 , \10366 , \10367 ,
         \10368 , \10369 , \10370 , \10371 , \10372 , \10373 , \10374 , \10375 , \10376 , \10377 ,
         \10378 , \10379 , \10380 , \10381 , \10382 , \10383 , \10384 , \10385 , \10386 , \10387 ,
         \10388 , \10389 , \10390 , \10391 , \10392 , \10393 , \10394 , \10395 , \10396 , \10397 ,
         \10398 , \10399 , \10400 , \10401 , \10402 , \10403 , \10404 , \10405 , \10406 , \10407 ,
         \10408 , \10409_nG225a , \10410 , \10411 , \10412 , \10413 , \10414 , \10415 , \10416 , \10417 ,
         \10418 , \10419 , \10420 , \10421 , \10422 , \10423 , \10424 , \10425 , \10426 , \10427 ,
         \10428 , \10429 , \10430 , \10431 , \10432 , \10433 , \10434 , \10435 , \10436 , \10437 ,
         \10438 , \10439 , \10440 , \10441 , \10442 , \10443 , \10444 , \10445 , \10446 , \10447 ,
         \10448 , \10449 , \10450 , \10451 , \10452 , \10453 , \10454 , \10455 , \10456 , \10457 ,
         \10458 , \10459 , \10460 , \10461 , \10462 , \10463 , \10464 , \10465 , \10466 , \10467 ,
         \10468 , \10469 , \10470 , \10471 , \10472 , \10473 , \10474 , \10475 , \10476 , \10477 ,
         \10478 , \10479 , \10480 , \10481 , \10482 , \10483 , \10484 , \10485 , \10486 , \10487 ,
         \10488 , \10489 , \10490 , \10491 , \10492 , \10493 , \10494 , \10495 , \10496 , \10497 ,
         \10498 , \10499 , \10500 , \10501 , \10502 , \10503 , \10504 , \10505 , \10506_nG221a , \10507 ,
         \10508 , \10509 , \10510 , \10511 , \10512 , \10513 , \10514 , \10515 , \10516 , \10517 ,
         \10518 , \10519 , \10520 , \10521 , \10522 , \10523 , \10524 , \10525 , \10526 , \10527 ,
         \10528 , \10529 , \10530 , \10531 , \10532 , \10533 , \10534 , \10535 , \10536 , \10537 ,
         \10538 , \10539 , \10540 , \10541 , \10542 , \10543 , \10544 , \10545 , \10546 , \10547 ,
         \10548 , \10549 , \10550 , \10551 , \10552 , \10553 , \10554 , \10555 , \10556 , \10557 ,
         \10558 , \10559 , \10560 , \10561 , \10562 , \10563 , \10564 , \10565 , \10566 , \10567 ,
         \10568 , \10569 , \10570 , \10571 , \10572 , \10573 , \10574 , \10575 , \10576 , \10577 ,
         \10578 , \10579 , \10580 , \10581 , \10582 , \10583 , \10584 , \10585 , \10586 , \10587 ,
         \10588 , \10589 , \10590 , \10591 , \10592 , \10593 , \10594 , \10595 , \10596 , \10597 ,
         \10598 , \10599 , \10600 , \10601 , \10602 , \10603 , \10604 , \10605 , \10606 , \10607 ,
         \10608 , \10609 , \10610 , \10611 , \10612 , \10613 , \10614 , \10615 , \10616 , \10617 ,
         \10618 , \10619 , \10620 , \10621 , \10622 , \10623 , \10624 , \10625 , \10626 , \10627 ,
         \10628 , \10629 , \10630 , \10631 , \10632 , \10633 , \10634 , \10635 , \10636 , \10637 ,
         \10638 , \10639 , \10640 , \10641 , \10642 , \10643 , \10644 , \10645 , \10646 , \10647 ,
         \10648 , \10649 , \10650 , \10651 , \10652 , \10653 , \10654 , \10655 , \10656 , \10657 ,
         \10658 , \10659 , \10660 , \10661 , \10662 , \10663 , \10664 , \10665 , \10666 , \10667 ,
         \10668 , \10669 , \10670 , \10671 , \10672 , \10673 , \10674 , \10675 , \10676 , \10677 ,
         \10678 , \10679 , \10680 , \10681 , \10682 , \10683 , \10684 , \10685 , \10686 , \10687 ,
         \10688 , \10689 , \10690 , \10691 , \10692 , \10693 , \10694 , \10695 , \10696 , \10697 ,
         \10698 , \10699 , \10700 , \10701 , \10702 , \10703 , \10704 , \10705 , \10706 , \10707 ,
         \10708 , \10709 , \10710 , \10711 , \10712 , \10713 , \10714 , \10715 , \10716 , \10717 ,
         \10718 , \10719 , \10720 , \10721 , \10722 , \10723 , \10724 , \10725 , \10726 , \10727 ,
         \10728 , \10729 , \10730 , \10731 , \10732 , \10733 , \10734 , \10735 , \10736 , \10737 ,
         \10738 , \10739 , \10740 , \10741 , \10742 , \10743 , \10744 , \10745 , \10746 , \10747 ,
         \10748 , \10749 , \10750 , \10751 , \10752 , \10753 , \10754 , \10755 , \10756 , \10757 ,
         \10758 , \10759 , \10760 , \10761 , \10762 , \10763 , \10764 , \10765 , \10766 , \10767 ,
         \10768 , \10769 , \10770 , \10771 , \10772 , \10773 , \10774 , \10775 , \10776 , \10777 ,
         \10778 , \10779 , \10780 , \10781 , \10782 , \10783 , \10784 , \10785 , \10786 , \10787 ,
         \10788 , \10789 , \10790 , \10791 , \10792 , \10793 , \10794 , \10795 , \10796 , \10797 ,
         \10798 , \10799 , \10800 , \10801 , \10802 , \10803 , \10804 , \10805 , \10806 , \10807 ,
         \10808 , \10809 , \10810 , \10811 , \10812 , \10813 , \10814 , \10815 , \10816 , \10817 ,
         \10818 , \10819 , \10820 , \10821 , \10822 , \10823 , \10824 , \10825 , \10826 , \10827 ,
         \10828 , \10829 , \10830 , \10831 , \10832 , \10833 , \10834 , \10835 , \10836 , \10837 ,
         \10838 , \10839 , \10840 , \10841 , \10842 , \10843 , \10844 , \10845 , \10846 , \10847 ,
         \10848 , \10849 , \10850 , \10851 , \10852 , \10853 , \10854 , \10855 , \10856 , \10857 ,
         \10858 , \10859 , \10860 , \10861 , \10862 , \10863 , \10864 , \10865 , \10866 , \10867 ,
         \10868 , \10869 , \10870 , \10871 , \10872 , \10873 , \10874 , \10875 , \10876 , \10877 ,
         \10878 , \10879 , \10880 , \10881 , \10882 , \10883 , \10884 , \10885 , \10886 , \10887 ,
         \10888 , \10889 , \10890 , \10891 , \10892 , \10893 , \10894 , \10895 , \10896 , \10897 ,
         \10898 , \10899 , \10900 , \10901 , \10902 , \10903 , \10904 , \10905 , \10906 , \10907 ,
         \10908 , \10909 , \10910 , \10911 , \10912 , \10913 , \10914 , \10915 , \10916 , \10917 ,
         \10918 , \10919 , \10920 , \10921 , \10922 , \10923 , \10924 , \10925 , \10926 , \10927 ,
         \10928 , \10929 , \10930 , \10931 , \10932 , \10933 , \10934 , \10935 , \10936 , \10937 ,
         \10938 , \10939 , \10940 , \10941 , \10942 , \10943 , \10944 , \10945 , \10946 , \10947 ,
         \10948 , \10949 , \10950 , \10951 , \10952 , \10953 , \10954 , \10955 , \10956 , \10957 ,
         \10958 , \10959 , \10960 , \10961 , \10962 , \10963 , \10964 , \10965 , \10966 , \10967 ,
         \10968 , \10969 , \10970 , \10971 , \10972 , \10973 , \10974 , \10975 , \10976 , \10977 ,
         \10978 , \10979 , \10980 , \10981 , \10982 , \10983 , \10984 , \10985 , \10986 , \10987 ,
         \10988 , \10989 , \10990 , \10991 , \10992 , \10993 , \10994 , \10995 , \10996 , \10997 ,
         \10998 , \10999 , \11000 , \11001 , \11002 , \11003 , \11004 , \11005 , \11006 , \11007 ,
         \11008 , \11009 , \11010 , \11011 , \11012 , \11013 , \11014 , \11015 , \11016 , \11017 ,
         \11018 , \11019 , \11020 , \11021 , \11022 , \11023 , \11024 , \11025 , \11026 , \11027 ,
         \11028 , \11029 , \11030 , \11031 , \11032 , \11033 , \11034 , \11035 , \11036 , \11037 ,
         \11038 , \11039 , \11040 , \11041 , \11042 , \11043 , \11044 , \11045 , \11046 , \11047 ,
         \11048 , \11049 , \11050 , \11051 , \11052 , \11053 , \11054 , \11055 , \11056 , \11057 ,
         \11058 , \11059 , \11060 , \11061 , \11062 , \11063 , \11064 , \11065 , \11066 , \11067 ,
         \11068 , \11069 , \11070 , \11071 , \11072 , \11073 , \11074 , \11075 , \11076 , \11077 ,
         \11078 , \11079 , \11080 , \11081 , \11082 , \11083 , \11084 , \11085 , \11086 , \11087 ,
         \11088 , \11089 , \11090 , \11091 , \11092 , \11093 , \11094 , \11095 , \11096 , \11097 ,
         \11098 , \11099 , \11100 , \11101 , \11102 , \11103 , \11104 , \11105 , \11106 , \11107 ,
         \11108 , \11109 , \11110 , \11111 , \11112 , \11113 , \11114 , \11115 , \11116 , \11117 ,
         \11118 , \11119 , \11120 , \11121 , \11122 , \11123 , \11124 , \11125 , \11126 , \11127 ,
         \11128 , \11129 , \11130 , \11131 , \11132 , \11133 , \11134 , \11135 , \11136 , \11137 ,
         \11138 , \11139 , \11140 , \11141 , \11142 , \11143 , \11144 , \11145 , \11146 , \11147 ,
         \11148 , \11149 , \11150 , \11151 , \11152 , \11153 , \11154 , \11155 , \11156 , \11157 ,
         \11158 , \11159 , \11160 , \11161 , \11162 , \11163 , \11164 , \11165 , \11166 , \11167 ,
         \11168 , \11169 , \11170 , \11171 , \11172 , \11173 , \11174 , \11175 , \11176 , \11177 ,
         \11178 , \11179 , \11180 , \11181 , \11182 , \11183 , \11184 , \11185 , \11186 , \11187 ,
         \11188 , \11189 , \11190 , \11191 , \11192 , \11193 , \11194 , \11195 , \11196 , \11197 ,
         \11198 , \11199 , \11200 , \11201 , \11202 , \11203 , \11204 , \11205 , \11206 , \11207 ,
         \11208 , \11209 , \11210 , \11211 , \11212 , \11213 , \11214 , \11215 , \11216 , \11217 ,
         \11218 , \11219 , \11220 , \11221 , \11222 , \11223 , \11224 , \11225 , \11226 , \11227 ,
         \11228 , \11229 , \11230 , \11231 , \11232 , \11233 , \11234 , \11235 , \11236 , \11237 ,
         \11238 , \11239 , \11240 , \11241 , \11242 , \11243 , \11244 , \11245 , \11246 , \11247 ,
         \11248 , \11249 , \11250 , \11251 , \11252 , \11253 , \11254 , \11255 , \11256 , \11257 ,
         \11258 , \11259 , \11260 , \11261 , \11262 , \11263 , \11264 , \11265 , \11266 , \11267 ,
         \11268 , \11269 , \11270 , \11271 , \11272 , \11273 , \11274 , \11275 , \11276 , \11277 ,
         \11278 , \11279 , \11280 , \11281 , \11282 , \11283 , \11284 , \11285 , \11286 , \11287 ,
         \11288 , \11289 , \11290 , \11291 , \11292 , \11293 , \11294 , \11295 , \11296 , \11297 ,
         \11298 , \11299 , \11300 , \11301 , \11302 , \11303 , \11304 , \11305 , \11306 , \11307 ,
         \11308 , \11309 , \11310 , \11311 , \11312 , \11313 , \11314 , \11315 , \11316 , \11317 ,
         \11318 , \11319 , \11320 , \11321 , \11322 , \11323 , \11324 , \11325 , \11326 , \11327 ,
         \11328 , \11329 , \11330 , \11331 , \11332 , \11333 , \11334 , \11335 , \11336 , \11337 ,
         \11338 , \11339 , \11340 , \11341 , \11342 , \11343 , \11344 , \11345 , \11346 , \11347 ,
         \11348 , \11349 , \11350 , \11351 , \11352 , \11353 , \11354 , \11355 , \11356 , \11357 ,
         \11358 , \11359 , \11360 , \11361 , \11362 , \11363 , \11364 , \11365 , \11366 , \11367 ,
         \11368 , \11369 , \11370 , \11371 , \11372_nG2a95 , \11373 , \11374 , \11375 , \11376 , \11377 ,
         \11378 , \11379 , \11380 , \11381 , \11382 , \11383 , \11384 , \11385 , \11386 , \11387 ,
         \11388 , \11389 , \11390 , \11391 , \11392 , \11393 , \11394 , \11395 , \11396 , \11397 ,
         \11398 , \11399 , \11400 , \11401_nG28b7 , \11402 , \11403 , \11404 , \11405 , \11406 , \11407 ,
         \11408 , \11409 , \11410 , \11411 , \11412 , \11413 , \11414 , \11415 , \11416 , \11417 ,
         \11418 , \11419 , \11420 , \11421 , \11422 , \11423 , \11424 , \11425 , \11426 , \11427 ,
         \11428 , \11429_nG28b5 , \11430 , \11431 , \11432 , \11433 , \11434 , \11435 , \11436 , \11437 ,
         \11438 , \11439 , \11440 , \11441 , \11442 , \11443 , \11444 , \11445 , \11446 , \11447 ,
         \11448 , \11449 , \11450 , \11451 , \11452 , \11453 , \11454 , \11455 , \11456 , \11457 ,
         \11458_nG270a , \11459 , \11460 , \11461 , \11462 , \11463 , \11464 , \11465 , \11466 , \11467 ,
         \11468 , \11469 , \11470 , \11471 , \11472 , \11473 , \11474 , \11475 , \11476 , \11477 ,
         \11478 , \11479 , \11480 , \11481 , \11482 , \11483 , \11484 , \11485 , \11486 , \11487_nG2708 ,
         \11488 , \11489 , \11490 , \11491 , \11492 , \11493 , \11494 , \11495 , \11496 , \11497 ,
         \11498 , \11499 , \11500 , \11501 , \11502 , \11503 , \11504 , \11505 , \11506 , \11507 ,
         \11508 , \11509 , \11510 , \11511 , \11512 , \11513 , \11514 , \11515 , \11516_nG2377 , \11517 ,
         \11518 , \11519 , \11520 , \11521 , \11522 , \11523 , \11524 , \11525 , \11526 , \11527 ,
         \11528 , \11529 , \11530 , \11531 , \11532 , \11533 , \11534 , \11535 , \11536 , \11537 ,
         \11538 , \11539 , \11540 , \11541 , \11542 , \11543 , \11544 , \11545_nG2375 , \11546 , \11547 ,
         \11548 , \11549 , \11550 , \11551 , \11552 , \11553 , \11554 , \11555 , \11556 , \11557 ,
         \11558 , \11559 , \11560 , \11561 , \11562 , \11563 , \11564 , \11565 , \11566 , \11567 ,
         \11568 , \11569 , \11570 , \11571 , \11572 , \11573_nG2307 , \11574 , \11575 , \11576 , \11577 ,
         \11578 , \11579 , \11580 , \11581 , \11582 , \11583 , \11584 , \11585 , \11586 , \11587 ,
         \11588 , \11589 , \11590 , \11591 , \11592 , \11593 , \11594 , \11595 , \11596 , \11597 ,
         \11598 , \11599 , \11600 , \11601 , \11602_nG2305 , \11603 , \11604 , \11605 , \11606 , \11607 ,
         \11608 , \11609 , \11610 , \11611 , \11612 , \11613 , \11614 , \11615 , \11616 , \11617 ,
         \11618 , \11619 , \11620 , \11621 , \11622 , \11623 , \11624 , \11625 , \11626 , \11627 ,
         \11628 , \11629 , \11630_nG22ad , \11631 , \11632 , \11633 , \11634 , \11635 , \11636 , \11637 ,
         \11638 , \11639 , \11640 , \11641 , \11642 , \11643 , \11644 , \11645 , \11646 , \11647 ,
         \11648 , \11649 , \11650 , \11651 , \11652 , \11653 , \11654 , \11655 , \11656 , \11657 ,
         \11658_nG22af , \11659 , \11660 , \11661 , \11662 , \11663 , \11664 , \11665 , \11666 , \11667 ,
         \11668 , \11669 , \11670 , \11671 , \11672 , \11673 , \11674 , \11675 , \11676 , \11677 ,
         \11678 , \11679 , \11680 , \11681 , \11682 , \11683 , \11684 , \11685 , \11686 , \11687_nG223f ,
         \11688 , \11689 , \11690 , \11691 , \11692 , \11693 , \11694 , \11695 , \11696 , \11697 ,
         \11698 , \11699 , \11700 , \11701 , \11702 , \11703 , \11704 , \11705 , \11706 , \11707 ,
         \11708 , \11709 , \11710 , \11711 , \11712 , \11713 , \11714 , \11715_nG223d , \11716 , \11717 ,
         \11718 , \11719 , \11720 , \11721 , \11722 , \11723 , \11724 , \11725 , \11726 , \11727 ,
         \11728 , \11729 , \11730 , \11731 , \11732 , \11733 , \11734 , \11735 , \11736 , \11737 ,
         \11738 , \11739 , \11740 , \11741 , \11742 , \11743 , \11744 , \11745 , \11746 , \11747 ,
         \11748 , \11749 , \11750 , \11751 , \11752 , \11753 , \11754 , \11755 , \11756 , \11757 ,
         \11758 , \11759 , \11760 , \11761 , \11762 , \11763 , \11764 , \11765 , \11766 , \11767 ,
         \11768 , \11769 , \11770 , \11771 , \11772 , \11773 , \11774 , \11775 , \11776 , \11777 ,
         \11778 , \11779 , \11780 , \11781 , \11782_nG30bb , \11783 , \11784 , \11785 , \11786 , \11787 ,
         \11788 , \11789 , \11790 , \11791 , \11792 , \11793 , \11794 , \11795 , \11796 , \11797 ,
         \11798 , \11799 , \11800 , \11801 , \11802 , \11803 , \11804 , \11805 , \11806 , \11807 ,
         \11808 , \11809 , \11810 , \11811 , \11812 , \11813 , \11814 , \11815 , \11816 , \11817 ,
         \11818 , \11819 , \11820 , \11821_nG31ca , \11822 , \11823 , \11824 , \11825 , \11826 , \11827 ,
         \11828 , \11829 , \11830 , \11831 , \11832 , \11833 , \11834 , \11835 , \11836 , \11837 ,
         \11838 , \11839 , \11840 , \11841 , \11842 , \11843 , \11844 , \11845 , \11846 , \11847 ,
         \11848 , \11849 , \11850 , \11851 , \11852 , \11853 , \11854 , \11855 , \11856 , \11857 ,
         \11858 , \11859 , \11860 , \11861 , \11862 , \11863 , \11864 , \11865 , \11866 , \11867 ,
         \11868 , \11869 , \11870 , \11871 , \11872 , \11873 , \11874_nG2fb5 , \11875 , \11876 , \11877 ,
         \11878 , \11879 , \11880 , \11881 , \11882 , \11883 , \11884 , \11885 , \11886 , \11887 ,
         \11888 , \11889 , \11890 , \11891 , \11892 , \11893 , \11894 , \11895 , \11896 , \11897 ,
         \11898 , \11899 , \11900 , \11901 , \11902 , \11903 , \11904 , \11905 , \11906 , \11907 ,
         \11908 , \11909 , \11910 , \11911 , \11912 , \11913 , \11914 , \11915 , \11916 , \11917 ,
         \11918 , \11919 , \11920 , \11921 , \11922 , \11923 , \11924 , \11925 , \11926 , \11927 ,
         \11928 , \11929 , \11930 , \11931 , \11932 , \11933 , \11934 , \11935 , \11936 , \11937 ,
         \11938 , \11939 , \11940 , \11941 , \11942 , \11943 , \11944 , \11945 , \11946 , \11947 ,
         \11948 , \11949 , \11950 , \11951_nG2e94 , \11952 , \11953 , \11954 , \11955 , \11956 , \11957 ,
         \11958 , \11959 , \11960 , \11961 , \11962 , \11963 , \11964 , \11965 , \11966 , \11967 ,
         \11968 , \11969 , \11970 , \11971 , \11972 , \11973 , \11974 , \11975 , \11976 , \11977 ,
         \11978 , \11979 , \11980 , \11981 , \11982 , \11983 , \11984 , \11985 , \11986 , \11987 ,
         \11988 , \11989 , \11990 , \11991 , \11992 , \11993 , \11994 , \11995 , \11996 , \11997 ,
         \11998 , \11999 , \12000 , \12001 , \12002 , \12003 , \12004 , \12005 , \12006 , \12007 ,
         \12008 , \12009 , \12010 , \12011 , \12012 , \12013 , \12014 , \12015 , \12016 , \12017 ,
         \12018 , \12019 , \12020 , \12021 , \12022 , \12023 , \12024 , \12025 , \12026 , \12027 ,
         \12028 , \12029 , \12030 , \12031 , \12032 , \12033 , \12034 , \12035 , \12036 , \12037 ,
         \12038 , \12039 , \12040 , \12041 , \12042 , \12043 , \12044 , \12045 , \12046 , \12047 ,
         \12048_nG2ca8 , \12049 , \12050 , \12051 , \12052 , \12053 , \12054 , \12055 , \12056 , \12057 ,
         \12058 , \12059 , \12060 , \12061 , \12062 , \12063 , \12064 , \12065 , \12066 , \12067 ,
         \12068 , \12069 , \12070 , \12071 , \12072 , \12073 , \12074 , \12075 , \12076_nG2daa , \12077 ,
         \12078 , \12079 , \12080 , \12081 , \12082 , \12083 , \12084 , \12085 , \12086 , \12087 ,
         \12088 , \12089 , \12090 , \12091 , \12092 , \12093 , \12094 , \12095 , \12096 , \12097 ,
         \12098 , \12099 , \12100 , \12101 , \12102 , \12103 , \12104 , \12105 , \12106 , \12107 ,
         \12108 , \12109 , \12110 , \12111 , \12112 , \12113 , \12114 , \12115 , \12116 , \12117 ,
         \12118 , \12119 , \12120 , \12121 , \12122 , \12123 , \12124 , \12125 , \12126 , \12127 ,
         \12128 , \12129 , \12130 , \12131 , \12132 , \12133 , \12134 , \12135 , \12136 , \12137 ,
         \12138 , \12139 , \12140 , \12141 , \12142 , \12143 , \12144 , \12145 , \12146 , \12147 ,
         \12148 , \12149 , \12150 , \12151 , \12152 , \12153 , \12154 , \12155 , \12156 , \12157 ,
         \12158 , \12159 , \12160_nG2bb5 , \12161 , \12162 , \12163 , \12164 , \12165 , \12166 , \12167 ,
         \12168 , \12169 , \12170 , \12171 , \12172 , \12173 , \12174 , \12175 , \12176 , \12177 ,
         \12178 , \12179 , \12180 , \12181 , \12182 , \12183 , \12184 , \12185 , \12186 , \12187 ,
         \12188 , \12189 , \12190 , \12191 , \12192 , \12193 , \12194 , \12195 , \12196 , \12197 ,
         \12198 , \12199 , \12200 , \12201 , \12202 , \12203 , \12204 , \12205 , \12206 , \12207 ,
         \12208 , \12209 , \12210 , \12211 , \12212 , \12213 , \12214 , \12215 , \12216 , \12217 ,
         \12218 , \12219 , \12220 , \12221 , \12222 , \12223 , \12224 , \12225 , \12226 , \12227 ,
         \12228 , \12229 , \12230 , \12231 , \12232 , \12233 , \12234 , \12235 , \12236 , \12237_nG2aae ,
         \12238 , \12239 , \12240 , \12241 , \12242 , \12243 , \12244 , \12245 , \12246 , \12247 ,
         \12248 , \12249 , \12250 , \12251 , \12252 , \12253 , \12254 , \12255 , \12256 , \12257 ,
         \12258 , \12259 , \12260 , \12261 , \12262 , \12263 , \12264 , \12265 , \12266 , \12267 ,
         \12268 , \12269 , \12270 , \12271 , \12272 , \12273 , \12274 , \12275 , \12276 , \12277 ,
         \12278 , \12279 , \12280 , \12281 , \12282 , \12283 , \12284 , \12285 , \12286 , \12287 ,
         \12288 , \12289 , \12290 , \12291 , \12292 , \12293 , \12294 , \12295 , \12296 , \12297 ,
         \12298 , \12299 , \12300 , \12301 , \12302 , \12303 , \12304 , \12305 , \12306 , \12307_nG29cd ,
         \12308 , \12309 , \12310 , \12311 , \12312 , \12313 , \12314 , \12315 , \12316 , \12317 ,
         \12318 , \12319 , \12320 , \12321 , \12322 , \12323 , \12324 , \12325 , \12326 , \12327 ,
         \12328 , \12329 , \12330 , \12331 , \12332 , \12333 , \12334 , \12335 , \12336 , \12337 ,
         \12338 , \12339 , \12340 , \12341 , \12342 , \12343 , \12344 , \12345 , \12346 , \12347 ,
         \12348 , \12349 , \12350 , \12351 , \12352 , \12353 , \12354 , \12355 , \12356 , \12357 ,
         \12358 , \12359 , \12360 , \12361 , \12362 , \12363 , \12364 , \12365 , \12366 , \12367 ,
         \12368 , \12369 , \12370 , \12371 , \12372 , \12373 , \12374 , \12375 , \12376 , \12377 ,
         \12378 , \12379 , \12380 , \12381 , \12382 , \12383 , \12384 , \12385 , \12386 , \12387 ,
         \12388 , \12389 , \12390 , \12391 , \12392 , \12393 , \12394 , \12395 , \12396 , \12397 ,
         \12398 , \12399 , \12400 , \12401 , \12402 , \12403 , \12404 , \12405 , \12406 , \12407 ,
         \12408 , \12409 , \12410 , \12411 , \12412 , \12413 , \12414 , \12415 , \12416 , \12417 ,
         \12418 , \12419 , \12420 , \12421 , \12422 , \12423 , \12424 , \12425 , \12426 , \12427 ,
         \12428 , \12429 , \12430 , \12431 , \12432 , \12433 , \12434 , \12435 , \12436 , \12437 ,
         \12438 , \12439 , \12440 , \12441 , \12442 , \12443 , \12444 , \12445 , \12446 , \12447 ,
         \12448 , \12449 , \12450 , \12451 , \12452 , \12453 , \12454 , \12455 , \12456 , \12457 ,
         \12458 , \12459 , \12460 , \12461 , \12462 , \12463 , \12464 , \12465 , \12466 , \12467 ,
         \12468 , \12469 , \12470 , \12471 , \12472 , \12473 , \12474 , \12475 , \12476 , \12477 ,
         \12478 , \12479 , \12480 , \12481 , \12482 , \12483 , \12484 , \12485 , \12486 , \12487 ,
         \12488 , \12489 , \12490 , \12491 , \12492 , \12493 , \12494 , \12495 , \12496 , \12497 ,
         \12498 , \12499 , \12500 , \12501 , \12502 , \12503 , \12504 , \12505 , \12506 , \12507 ,
         \12508 , \12509 , \12510 , \12511 , \12512 , \12513 , \12514 , \12515_nG28d0 , \12516 , \12517 ,
         \12518 , \12519 , \12520 , \12521 , \12522 , \12523 , \12524 , \12525 , \12526 , \12527 ,
         \12528 , \12529 , \12530 , \12531 , \12532 , \12533 , \12534 , \12535 , \12536 , \12537 ,
         \12538 , \12539 , \12540 , \12541 , \12542 , \12543 , \12544 , \12545 , \12546 , \12547 ,
         \12548 , \12549 , \12550 , \12551 , \12552 , \12553 , \12554 , \12555 , \12556 , \12557 ,
         \12558 , \12559 , \12560 , \12561 , \12562 , \12563 , \12564 , \12565 , \12566 , \12567 ,
         \12568 , \12569 , \12570 , \12571 , \12572 , \12573 , \12574 , \12575 , \12576 , \12577 ,
         \12578 , \12579 , \12580 , \12581 , \12582 , \12583 , \12584 , \12585 , \12586 , \12587 ,
         \12588 , \12589 , \12590 , \12591 , \12592 , \12593 , \12594 , \12595 , \12596 , \12597 ,
         \12598 , \12599 , \12600 , \12601 , \12602 , \12603 , \12604 , \12605 , \12606 , \12607 ,
         \12608 , \12609 , \12610 , \12611 , \12612 , \12613 , \12614 , \12615 , \12616 , \12617 ,
         \12618 , \12619 , \12620 , \12621 , \12622 , \12623 , \12624 , \12625 , \12626 , \12627 ,
         \12628 , \12629 , \12630 , \12631 , \12632 , \12633 , \12634 , \12635 , \12636 , \12637 ,
         \12638 , \12639 , \12640 , \12641 , \12642 , \12643 , \12644 , \12645 , \12646 , \12647 ,
         \12648 , \12649 , \12650 , \12651 , \12652 , \12653 , \12654 , \12655 , \12656 , \12657 ,
         \12658 , \12659 , \12660 , \12661 , \12662_nG27f3 , \12663 , \12664 , \12665 , \12666 , \12667 ,
         \12668 , \12669 , \12670 , \12671 , \12672 , \12673 , \12674 , \12675 , \12676 , \12677 ,
         \12678 , \12679 , \12680 , \12681 , \12682 , \12683 , \12684 , \12685 , \12686 , \12687 ,
         \12688 , \12689 , \12690 , \12691 , \12692 , \12693 , \12694 , \12695 , \12696 , \12697 ,
         \12698 , \12699 , \12700 , \12701 , \12702 , \12703 , \12704 , \12705 , \12706_nG2723 , \12707 ,
         \12708 , \12709 , \12710 , \12711 , \12712 , \12713 , \12714 , \12715 , \12716 , \12717 ,
         \12718 , \12719 , \12720 , \12721 , \12722 , \12723 , \12724 , \12725 , \12726 , \12727 ,
         \12728 , \12729 , \12730 , \12731 , \12732 , \12733 , \12734 , \12735 , \12736 , \12737 ,
         \12738 , \12739 , \12740 , \12741 , \12742 , \12743 , \12744 , \12745 , \12746 , \12747 ,
         \12748 , \12749 , \12750 , \12751 , \12752 , \12753 , \12754 , \12755 , \12756 , \12757 ,
         \12758 , \12759 , \12760 , \12761 , \12762 , \12763 , \12764 , \12765 , \12766 , \12767 ,
         \12768 , \12769 , \12770 , \12771 , \12772 , \12773 , \12774 , \12775 , \12776 , \12777 ,
         \12778 , \12779 , \12780 , \12781 , \12782 , \12783 , \12784 , \12785 , \12786 , \12787 ,
         \12788 , \12789 , \12790 , \12791 , \12792 , \12793 , \12794 , \12795 , \12796 , \12797 ,
         \12798 , \12799 , \12800 , \12801 , \12802 , \12803 , \12804 , \12805 , \12806 , \12807 ,
         \12808 , \12809 , \12810 , \12811 , \12812 , \12813 , \12814 , \12815 , \12816 , \12817 ,
         \12818 , \12819 , \12820 , \12821 , \12822 , \12823 , \12824 , \12825 , \12826 , \12827 ,
         \12828 , \12829 , \12830 , \12831 , \12832 , \12833 , \12834 , \12835 , \12836 , \12837 ,
         \12838 , \12839 , \12840 , \12841 , \12842 , \12843 , \12844 , \12845 , \12846 , \12847 ,
         \12848 , \12849 , \12850 , \12851 , \12852 , \12853 , \12854 , \12855 , \12856 , \12857 ,
         \12858 , \12859 , \12860 , \12861 , \12862 , \12863 , \12864 , \12865 , \12866 , \12867 ,
         \12868 , \12869 , \12870 , \12871 , \12872 , \12873 , \12874 , \12875 , \12876 , \12877 ,
         \12878 , \12879 , \12880 , \12881_nG23c5 , \12882 , \12883 , \12884 , \12885 , \12886 , \12887 ,
         \12888 , \12889 , \12890 , \12891 , \12892 , \12893 , \12894 , \12895 , \12896 , \12897 ,
         \12898 , \12899 , \12900 , \12901 , \12902 , \12903 , \12904 , \12905 , \12906 , \12907 ,
         \12908 , \12909 , \12910 , \12911 , \12912 , \12913 , \12914 , \12915 , \12916 , \12917 ,
         \12918 , \12919 , \12920 , \12921 , \12922_nG2391 , \12923 , \12924 , \12925 , \12926 , \12927 ,
         \12928 , \12929 , \12930 , \12931 , \12932 , \12933 , \12934 , \12935 , \12936 , \12937 ,
         \12938 , \12939 , \12940 , \12941 , \12942 , \12943 , \12944 , \12945 , \12946 , \12947 ,
         \12948 , \12949 , \12950 , \12951 , \12952 , \12953 , \12954 , \12955 , \12956 , \12957 ,
         \12958 , \12959 , \12960 , \12961 , \12962 , \12963 , \12964 , \12965 , \12966 , \12967 ,
         \12968 , \12969 , \12970 , \12971 , \12972 , \12973 , \12974 , \12975 , \12976 , \12977 ,
         \12978 , \12979 , \12980 , \12981 , \12982 , \12983 , \12984 , \12985 , \12986 , \12987 ,
         \12988 , \12989 , \12990 , \12991 , \12992 , \12993 , \12994 , \12995 , \12996 , \12997 ,
         \12998 , \12999 , \13000 , \13001 , \13002 , \13003 , \13004 , \13005 , \13006 , \13007 ,
         \13008 , \13009 , \13010 , \13011 , \13012 , \13013 , \13014 , \13015 , \13016 , \13017 ,
         \13018 , \13019 , \13020 , \13021 , \13022 , \13023 , \13024 , \13025 , \13026 , \13027 ,
         \13028 , \13029 , \13030 , \13031 , \13032 , \13033 , \13034 , \13035 , \13036 , \13037 ,
         \13038 , \13039 , \13040 , \13041 , \13042 , \13043 , \13044 , \13045 , \13046 , \13047 ,
         \13048 , \13049 , \13050 , \13051 , \13052 , \13053 , \13054 , \13055 , \13056 , \13057 ,
         \13058 , \13059 , \13060 , \13061 , \13062 , \13063 , \13064 , \13065 , \13066 , \13067 ,
         \13068 , \13069 , \13070 , \13071 , \13072 , \13073 , \13074 , \13075 , \13076 , \13077 ,
         \13078 , \13079 , \13080 , \13081 , \13082 , \13083 , \13084 , \13085 , \13086 , \13087 ,
         \13088 , \13089 , \13090 , \13091 , \13092 , \13093 , \13094 , \13095 , \13096 , \13097 ,
         \13098 , \13099 , \13100 , \13101 , \13102 , \13103 , \13104 , \13105 , \13106 , \13107 ,
         \13108 , \13109 , \13110 , \13111 , \13112 , \13113 , \13114 , \13115 , \13116 , \13117 ,
         \13118 , \13119 , \13120 , \13121 , \13122_nG2354 , \13123 , \13124 , \13125 , \13126 , \13127 ,
         \13128 , \13129 , \13130 , \13131 , \13132 , \13133 , \13134 , \13135 , \13136 , \13137 ,
         \13138 , \13139 , \13140 , \13141 , \13142 , \13143 , \13144 , \13145 , \13146 , \13147 ,
         \13148 , \13149 , \13150 , \13151 , \13152 , \13153 , \13154 , \13155 , \13156 , \13157 ,
         \13158 , \13159 , \13160 , \13161 , \13162_nG2320 , \13163 , \13164 , \13165 , \13166 , \13167 ,
         \13168 , \13169 , \13170 , \13171 , \13172 , \13173 , \13174 , \13175 , \13176 , \13177 ,
         \13178 , \13179 , \13180 , \13181 , \13182 , \13183 , \13184 , \13185 , \13186 , \13187 ,
         \13188 , \13189 , \13190 , \13191 , \13192 , \13193 , \13194 , \13195 , \13196 , \13197 ,
         \13198 , \13199 , \13200 , \13201 , \13202 , \13203 , \13204 , \13205 , \13206 , \13207 ,
         \13208 , \13209 , \13210 , \13211 , \13212 , \13213 , \13214 , \13215 , \13216 , \13217 ,
         \13218 , \13219 , \13220 , \13221 , \13222 , \13223 , \13224 , \13225 , \13226 , \13227 ,
         \13228 , \13229 , \13230 , \13231 , \13232 , \13233 , \13234 , \13235 , \13236 , \13237 ,
         \13238 , \13239 , \13240 , \13241 , \13242 , \13243 , \13244 , \13245 , \13246 , \13247 ,
         \13248 , \13249 , \13250 , \13251 , \13252 , \13253 , \13254 , \13255 , \13256 , \13257 ,
         \13258 , \13259 , \13260 , \13261 , \13262 , \13263 , \13264 , \13265 , \13266 , \13267 ,
         \13268 , \13269 , \13270 , \13271 , \13272 , \13273 , \13274 , \13275 , \13276 , \13277 ,
         \13278 , \13279 , \13280 , \13281 , \13282 , \13283 , \13284 , \13285 , \13286 , \13287 ,
         \13288 , \13289 , \13290 , \13291 , \13292 , \13293 , \13294 , \13295 , \13296 , \13297 ,
         \13298 , \13299 , \13300 , \13301 , \13302 , \13303 , \13304 , \13305 , \13306 , \13307 ,
         \13308 , \13309 , \13310 , \13311 , \13312 , \13313 , \13314 , \13315 , \13316 , \13317 ,
         \13318 , \13319 , \13320 , \13321 , \13322 , \13323 , \13324 , \13325 , \13326 , \13327 ,
         \13328 , \13329 , \13330 , \13331 , \13332 , \13333 , \13334 , \13335 , \13336 , \13337 ,
         \13338 , \13339 , \13340 , \13341 , \13342 , \13343 , \13344 , \13345 , \13346 , \13347 ,
         \13348 , \13349 , \13350 , \13351 , \13352 , \13353 , \13354 , \13355 , \13356 , \13357 ,
         \13358 , \13359 , \13360 , \13361 , \13362 , \13363 , \13364_nG22e4 , \13365 , \13366 , \13367 ,
         \13368 , \13369 , \13370 , \13371 , \13372 , \13373 , \13374 , \13375 , \13376 , \13377 ,
         \13378 , \13379 , \13380 , \13381 , \13382 , \13383 , \13384 , \13385 , \13386 , \13387 ,
         \13388 , \13389 , \13390 , \13391 , \13392 , \13393 , \13394 , \13395 , \13396 , \13397 ,
         \13398 , \13399 , \13400 , \13401 , \13402 , \13403 , \13404 , \13405 , \13406 , \13407 ,
         \13408 , \13409 , \13410 , \13411 , \13412 , \13413 , \13414 , \13415 , \13416 , \13417 ,
         \13418 , \13419 , \13420 , \13421 , \13422 , \13423 , \13424 , \13425 , \13426 , \13427 ,
         \13428 , \13429 , \13430 , \13431 , \13432 , \13433 , \13434 , \13435 , \13436 , \13437 ,
         \13438 , \13439 , \13440 , \13441 , \13442 , \13443 , \13444 , \13445 , \13446 , \13447 ,
         \13448 , \13449 , \13450 , \13451 , \13452 , \13453 , \13454 , \13455 , \13456 , \13457 ,
         \13458 , \13459 , \13460 , \13461 , \13462 , \13463 , \13464 , \13465 , \13466 , \13467 ,
         \13468 , \13469 , \13470 , \13471 , \13472 , \13473 , \13474 , \13475 , \13476 , \13477 ,
         \13478 , \13479 , \13480 , \13481_nG22ab , \13482 , \13483 , \13484 , \13485 , \13486 , \13487 ,
         \13488 , \13489 , \13490 , \13491 , \13492 , \13493 , \13494 , \13495 , \13496 , \13497 ,
         \13498 , \13499 , \13500 , \13501 , \13502 , \13503 , \13504 , \13505 , \13506 , \13507 ,
         \13508 , \13509 , \13510 , \13511 , \13512 , \13513 , \13514 , \13515 , \13516 , \13517 ,
         \13518 , \13519 , \13520 , \13521 , \13522 , \13523 , \13524 , \13525 , \13526 , \13527 ,
         \13528 , \13529 , \13530 , \13531 , \13532 , \13533 , \13534 , \13535 , \13536 , \13537 ,
         \13538 , \13539 , \13540 , \13541 , \13542 , \13543 , \13544 , \13545 , \13546 , \13547 ,
         \13548 , \13549 , \13550 , \13551 , \13552 , \13553 , \13554 , \13555 , \13556 , \13557 ,
         \13558 , \13559 , \13560 , \13561 , \13562 , \13563 , \13564 , \13565 , \13566 , \13567 ,
         \13568 , \13569 , \13570 , \13571 , \13572 , \13573 , \13574 , \13575 , \13576 , \13577 ,
         \13578 , \13579 , \13580 , \13581 , \13582 , \13583 , \13584 , \13585 , \13586 , \13587 ,
         \13588 , \13589 , \13590 , \13591 , \13592 , \13593 , \13594 , \13595 , \13596 , \13597 ,
         \13598 , \13599 , \13600 , \13601 , \13602 , \13603 , \13604 , \13605 , \13606 , \13607 ,
         \13608 , \13609 , \13610 , \13611 , \13612 , \13613 , \13614 , \13615 , \13616 , \13617 ,
         \13618 , \13619 , \13620 , \13621 , \13622 , \13623 , \13624 , \13625 , \13626 , \13627 ,
         \13628 , \13629 , \13630 , \13631 , \13632 , \13633 , \13634 , \13635 , \13636 , \13637_nG2273 ,
         \13638 , \13639 , \13640 , \13641 , \13642 , \13643 , \13644 , \13645 , \13646 , \13647 ,
         \13648 , \13649 , \13650 , \13651 , \13652 , \13653 , \13654 , \13655 , \13656 , \13657 ,
         \13658 , \13659 , \13660 , \13661 , \13662 , \13663 , \13664 , \13665 , \13666 , \13667 ,
         \13668 , \13669 , \13670 , \13671 , \13672 , \13673 , \13674 , \13675 , \13676 , \13677 ,
         \13678 , \13679 , \13680 , \13681 , \13682 , \13683 , \13684 , \13685 , \13686 , \13687 ,
         \13688 , \13689 , \13690 , \13691 , \13692 , \13693 , \13694 , \13695 , \13696 , \13697 ,
         \13698 , \13699 , \13700 , \13701 , \13702 , \13703 , \13704 , \13705 , \13706 , \13707 ,
         \13708 , \13709 , \13710 , \13711 , \13712 , \13713 , \13714 , \13715 , \13716 , \13717 ,
         \13718 , \13719 , \13720 , \13721 , \13722 , \13723 , \13724 , \13725 , \13726_nG223a , \13727 ,
         \13728 , \13729 , \13730 , \13731 , \13732 , \13733 , \13734 , \13735 , \13736 , \13737 ,
         \13738 , \13739 , \13740 , \13741 , \13742 , \13743 , \13744 , \13745 , \13746 , \13747 ,
         \13748 , \13749 , \13750 , \13751 , \13752 , \13753 , \13754 , \13755 , \13756 , \13757 ,
         \13758 , \13759 , \13760 , \13761 , \13762 , \13763 , \13764 , \13765 , \13766 , \13767 ,
         \13768 , \13769 , \13770 , \13771 , \13772 , \13773 , \13774 , \13775 , \13776 , \13777 ,
         \13778 , \13779 , \13780 , \13781 , \13782 , \13783 , \13784 , \13785 , \13786 , \13787 ,
         \13788 , \13789 , \13790 , \13791 , \13792 , \13793 , \13794 , \13795 , \13796 , \13797 ,
         \13798 , \13799 , \13800 , \13801 , \13802 , \13803 , \13804 , \13805 , \13806 , \13807 ,
         \13808 , \13809 , \13810 , \13811 , \13812 , \13813 , \13814 , \13815 , \13816 , \13817 ,
         \13818 , \13819 , \13820 , \13821 , \13822 , \13823 , \13824 , \13825 , \13826 , \13827 ,
         \13828 , \13829 , \13830 , \13831 , \13832 , \13833 , \13834 , \13835 , \13836 , \13837 ,
         \13838 , \13839 , \13840 , \13841 , \13842 , \13843 , \13844 , \13845 , \13846 , \13847 ,
         \13848 , \13849 , \13850 , \13851 , \13852 , \13853 , \13854 , \13855 , \13856 , \13857 ,
         \13858 , \13859 , \13860 , \13861 , \13862 , \13863 , \13864 , \13865 , \13866 , \13867 ,
         \13868 , \13869 , \13870 , \13871 , \13872 , \13873 , \13874 , \13875 , \13876 , \13877 ,
         \13878 , \13879 , \13880 , \13881 , \13882 , \13883 , \13884 , \13885 , \13886 , \13887 ,
         \13888 , \13889 , \13890 , \13891 , \13892 , \13893 , \13894 , \13895 , \13896 , \13897 ,
         \13898 , \13899 , \13900 , \13901 , \13902 , \13903 , \13904 , \13905 , \13906 , \13907 ,
         \13908 , \13909 , \13910 , \13911 , \13912 , \13913 , \13914 , \13915 , \13916 , \13917 ,
         \13918 , \13919 , \13920 , \13921 , \13922 , \13923 , \13924 , \13925 , \13926 , \13927 ,
         \13928 , \13929 , \13930 , \13931 , \13932 , \13933 , \13934 , \13935 , \13936 , \13937 ,
         \13938 , \13939 , \13940 , \13941 , \13942 , \13943 , \13944 , \13945 , \13946 , \13947 ,
         \13948 , \13949 , \13950 , \13951 , \13952 , \13953 , \13954 , \13955 , \13956 , \13957 ,
         \13958 , \13959 , \13960 , \13961 , \13962 , \13963 , \13964 , \13965 , \13966 , \13967 ,
         \13968 , \13969 , \13970 , \13971 , \13972 , \13973 , \13974 , \13975 , \13976 , \13977 ,
         \13978 , \13979 , \13980 , \13981 , \13982 , \13983 , \13984 , \13985 , \13986 , \13987 ,
         \13988 , \13989 , \13990 , \13991 , \13992 , \13993 , \13994 , \13995 , \13996 , \13997 ,
         \13998 , \13999 , \14000 , \14001 , \14002 , \14003 , \14004 , \14005 , \14006 , \14007 ,
         \14008 , \14009 , \14010 , \14011 , \14012 , \14013 , \14014 , \14015 , \14016 , \14017 ,
         \14018 , \14019 , \14020 , \14021 , \14022 , \14023 , \14024 , \14025 , \14026 , \14027 ,
         \14028 , \14029 , \14030 , \14031 , \14032 , \14033 , \14034 , \14035 , \14036 , \14037 ,
         \14038 , \14039 , \14040 , \14041 , \14042 , \14043 , \14044 , \14045 , \14046 , \14047 ,
         \14048 , \14049 , \14050 , \14051 , \14052 , \14053 , \14054 , \14055 , \14056 , \14057 ,
         \14058 , \14059 , \14060 , \14061 , \14062 , \14063 , \14064 , \14065 , \14066 , \14067 ,
         \14068 , \14069 , \14070 , \14071 , \14072 , \14073 , \14074 , \14075 , \14076 , \14077 ,
         \14078 , \14079 , \14080 , \14081 , \14082 , \14083 , \14084 , \14085 , \14086 , \14087 ,
         \14088 , \14089 , \14090 , \14091 , \14092 , \14093 , \14094 , \14095 , \14096 , \14097 ,
         \14098 , \14099 , \14100 , \14101 , \14102 , \14103 , \14104 , \14105 , \14106 , \14107 ,
         \14108 , \14109 , \14110 , \14111 , \14112 , \14113 , \14114 , \14115 , \14116 , \14117 ,
         \14118 , \14119 , \14120 , \14121 , \14122 , \14123 , \14124 , \14125 , \14126 , \14127 ,
         \14128 , \14129 , \14130 , \14131 , \14132 , \14133 , \14134 , \14135 , \14136 , \14137 ,
         \14138 , \14139 , \14140 , \14141 , \14142 , \14143 , \14144 , \14145 , \14146 , \14147 ,
         \14148 , \14149 , \14150 , \14151 , \14152 , \14153 , \14154 , \14155 , \14156 , \14157 ,
         \14158 , \14159 , \14160 , \14161 , \14162 , \14163 , \14164 , \14165 , \14166 , \14167 ,
         \14168 , \14169 , \14170 , \14171 , \14172 , \14173 , \14174 , \14175 , \14176 , \14177 ,
         \14178 , \14179 , \14180 , \14181 , \14182 , \14183 , \14184 , \14185 , \14186 , \14187 ,
         \14188 , \14189 , \14190 , \14191 , \14192 , \14193 , \14194 , \14195 , \14196 , \14197 ,
         \14198 , \14199 , \14200 , \14201 , \14202 , \14203 , \14204 , \14205 , \14206 , \14207 ,
         \14208 , \14209 , \14210 , \14211 , \14212 , \14213 , \14214 , \14215 , \14216 , \14217 ,
         \14218 , \14219 , \14220 , \14221 , \14222 , \14223 , \14224 , \14225 , \14226 , \14227 ,
         \14228 , \14229 , \14230 , \14231 , \14232 , \14233 , \14234 , \14235 , \14236 , \14237 ,
         \14238 , \14239 , \14240 , \14241 , \14242 , \14243 , \14244 , \14245 , \14246 , \14247 ,
         \14248 , \14249 , \14250 , \14251 , \14252 , \14253 , \14254 , \14255 , \14256 , \14257 ,
         \14258 , \14259 , \14260 , \14261 , \14262 , \14263 , \14264 , \14265 , \14266 , \14267 ,
         \14268 , \14269 , \14270 , \14271 , \14272 , \14273 , \14274 , \14275 , \14276 , \14277 ,
         \14278 , \14279 , \14280 , \14281 , \14282 , \14283 , \14284 , \14285 , \14286 , \14287 ,
         \14288 , \14289 , \14290 , \14291 , \14292 , \14293 , \14294 , \14295 , \14296 , \14297 ,
         \14298 , \14299 , \14300 , \14301 , \14302 , \14303 , \14304 , \14305 , \14306 , \14307 ,
         \14308 , \14309 , \14310 , \14311 , \14312 , \14313 , \14314 , \14315 , \14316 , \14317 ,
         \14318 , \14319 , \14320 , \14321 , \14322 , \14323 , \14324 , \14325 , \14326 , \14327 ,
         \14328 , \14329 , \14330 , \14331 , \14332 , \14333 , \14334 , \14335 , \14336 , \14337 ,
         \14338 , \14339 , \14340 , \14341 , \14342 , \14343 , \14344 , \14345 , \14346 , \14347 ,
         \14348 , \14349 , \14350 , \14351 , \14352 , \14353 , \14354 , \14355 , \14356 , \14357 ,
         \14358 , \14359 , \14360 , \14361 , \14362 , \14363 , \14364 , \14365 , \14366 , \14367 ,
         \14368 , \14369 , \14370 , \14371 , \14372 , \14373 , \14374 , \14375 , \14376 , \14377 ,
         \14378 , \14379 , \14380 , \14381 , \14382 , \14383 , \14384 , \14385 , \14386 , \14387 ,
         \14388 , \14389 , \14390 , \14391 , \14392 , \14393 , \14394 , \14395 , \14396 , \14397 ,
         \14398 , \14399 , \14400 , \14401 , \14402 , \14403 , \14404 , \14405 , \14406 , \14407 ,
         \14408 , \14409 , \14410 , \14411 , \14412 , \14413 , \14414 , \14415 , \14416 , \14417 ,
         \14418 , \14419 , \14420 , \14421 , \14422 , \14423 , \14424 , \14425 , \14426 , \14427 ,
         \14428 , \14429 , \14430 , \14431 , \14432 , \14433 , \14434 , \14435 , \14436 , \14437 ,
         \14438 , \14439 , \14440 , \14441 , \14442 , \14443 , \14444 , \14445 , \14446 , \14447 ,
         \14448 , \14449 , \14450 , \14451 , \14452 , \14453 , \14454 , \14455 , \14456 , \14457 ,
         \14458 , \14459 , \14460 , \14461 , \14462 , \14463 , \14464 , \14465 , \14466 , \14467 ,
         \14468 , \14469 , \14470 , \14471 , \14472 , \14473 , \14474 , \14475 , \14476 , \14477 ,
         \14478 , \14479 , \14480 , \14481 , \14482 , \14483 , \14484 , \14485 , \14486 , \14487 ,
         \14488 , \14489 , \14490 , \14491 , \14492 , \14493 , \14494 , \14495 , \14496 , \14497 ,
         \14498 , \14499 , \14500 , \14501 , \14502 , \14503 , \14504 , \14505 , \14506 , \14507 ,
         \14508 , \14509 , \14510 , \14511 , \14512 , \14513 , \14514 , \14515 , \14516 , \14517 ,
         \14518 , \14519 , \14520 , \14521 , \14522 , \14523 , \14524 , \14525 , \14526 , \14527 ,
         \14528 , \14529 , \14530 , \14531 , \14532 , \14533 , \14534 , \14535 , \14536 , \14537 ,
         \14538 , \14539 , \14540 , \14541 , \14542 , \14543 , \14544 , \14545 , \14546 , \14547 ,
         \14548 , \14549 , \14550 , \14551 , \14552 , \14553 , \14554 , \14555 , \14556 , \14557 ,
         \14558 , \14559 , \14560 , \14561 , \14562 , \14563 , \14564 , \14565 , \14566 , \14567_nG7eb ,
         \14568 , \14569 , \14570_nG80c , \14571 , \14572 , \14573 , \14574_nG906 , \14575 , \14576 , \14577 ,
         \14578_nG908 , \14579 , \14580 , \14581 , \14582_nG925 , \14583 , \14584 , \14585_nG927 , \14586 , \14587 ,
         \14588 , \14589 , \14590_nG8e5 , \14591 , \14592 , \14593 , \14594 , \14595 , \14596_nG8e7 , \14597 ,
         \14598 , \14599 , \14600_nG8c8 , \14601 , \14602 , \14603 , \14604 , \14605 , \14606_nG8c6 , \14607 ,
         \14608 , \14609 , \14610_nG8a9 , \14611 , \14612 , \14613_nG8a7 , \14614 , \14615 , \14616 , \14617 ,
         \14618 , \14619_nG88a , \14620 , \14621 , \14622 , \14623 , \14624 , \14625_nG888 , \14626 , \14627 ,
         \14628 , \14629_nG86b , \14630 , \14631 , \14632_nG869 , \14633 , \14634 , \14635 , \14636 , \14637 ,
         \14638_nG84c , \14639 , \14640 , \14641 , \14642 , \14643 , \14644_nG84a , \14645 , \14646 , \14647 ,
         \14648_nG829 , \14649 , \14650 , \14651 , \14652 , \14653 , \14654_nG82b , \14655 , \14656 , \14657 ,
         \14658 , \14659 , \14660 , \14661_nG80a , \14662 , \14663 , \14664 , \14665 , \14666 , \14667 ,
         \14668_nG7e9 , \14669 , \14670 , \14671 , \14672_nG7ca , \14673 , \14674 , \14675 , \14676 , \14677 ,
         \14678_nG7c8 , \14679 , \14680 , \14681 , \14682_nG7a9 , \14683 , \14684 , \14685_nG7a6 , \14686 , \14687 ,
         \14688 , \14689 , \14690 , \14691 , \14692_nG62d , \14693 , \14694 , \14695 , \14696 , \14697 ,
         \14698 , \14699 , \14700 , \14701 , \14702 , \14703 , \14704 , \14705 , \14706 , \14707 ,
         \14708 , \14709 , \14710 , \14711 , \14712 , \14713 , \14714 , \14715 , \14716 , \14717 ,
         \14718 , \14719_nG64a , \14720 , \14721 , \14722 , \14723 , \14724_nG683 , \14725 , \14726 , \14727 ,
         \14728 , \14729 , \14730 , \14731 , \14732 , \14733 , \14734 , \14735 , \14736 , \14737_nG6a0 ,
         \14738 , \14739 , \14740_nG6bd , \14741 , \14742 , \14743 , \14744 , \14745 , \14746 , \14747 ,
         \14748 , \14749 , \14750 , \14751_nG6da , \14752 , \14753 , \14754 , \14755 , \14756 , \14757 ,
         \14758 , \14759_nG713 , \14760 , \14761 , \14762 , \14763 , \14764 , \14765 , \14766 , \14767 ,
         \14768 , \14769 , \14770 , \14771_nG784 , \14772 , \14773 , \14774 , \14775 , \14776 , \14777 ,
         \14778_nG768 , \14779 , \14780 , \14781 , \14782_nG74b , \14783 , \14784 , \14785 , \14786 , \14787 ,
         \14788 , \14789 , \14790 , \14791 , \14792_nG72f , \14793 , \14794 , \14795 , \14796 , \14797 ,
         \14798 , \14799 , \14800 , \14801_nG6f6 , \14802 , \14803 , \14804 , \14805 , \14806 , \14807 ,
         \14808 , \14809 , \14810 , \14811 , \14812 , \14813 , \14814 , \14815 , \14816 , \14817 ,
         \14818 , \14819_nG666 , \14820 , \14821 , \14822 , \14823 , \14824 , \14825 , \14826 , \14827_nG3a8a ,
         \14828 , \14829 , \14830 , \14831 , \14832 , \14833_nG3a4f , \14834 , \14835 , \14836 , \14837 ,
         \14838 , \14839_nG3a1e , \14840 , \14841 , \14842 , \14843 , \14844 , \14845_nG39d7 , \14846 , \14847 ,
         \14848 , \14849 , \14850 , \14851_nG397e , \14852 , \14853 , \14854 , \14855 , \14856 , \14857_nG3917 ,
         \14858 , \14859 , \14860 , \14861 , \14862 , \14863_nG38a0 , \14864 , \14865 , \14866 , \14867 ,
         \14868 , \14869_nG3823 , \14870 , \14871 , \14872 , \14873 , \14874 , \14875 , \14876_nG378d , \14877 ,
         \14878 , \14879 , \14880 , \14881 , \14882 , \14883 , \14884 , \14885_nG36d5 , \14886 , \14887 ,
         \14888 , \14889 , \14890 , \14891 , \14892 , \14893 , \14894 , \14895 , \14896_nG3621 , \14897 ,
         \14898 , \14899 , \14900 , \14901 , \14902_nG3562 , \14903 , \14904 , \14905 , \14906 , \14907 ,
         \14908 , \14909_nG347c , \14910 , \14911 , \14912 , \14913 , \14914 , \14915 , \14916 , \14917 ,
         \14918 , \14919 , \14920_nG33a1 , \14921 , \14922 , \14923 , \14924 , \14925 , \14926_nG32a4 , \14927 ,
         \14928 , \14929 , \14930 , \14931 , \14932_nG3195 , \14933 , \14934 , \14935 , \14936 , \14937 ,
         \14938 , \14939_nG3087 , \14940 , \14941 , \14942 , \14943 , \14944 , \14945 , \14946 , \14947 ,
         \14948 , \14949_nG2f81 , \14950 , \14951 , \14952 , \14953 , \14954 , \14955 , \14956 , \14957 ,
         \14958 , \14959 , \14960 , \14961_nG2e5f , \14962 , \14963 , \14964 , \14965 , \14966 , \14967 ,
         \14968 , \14969 , \14970 , \14971 , \14972 , \14973 , \14974 , \14975 , \14976 , \14977_nG2d75 ,
         \14978 , \14979 , \14980 , \14981 , \14982 , \14983_nG2c74 , \14984 , \14985 , \14986 , \14987 ,
         \14988 , \14989_nG2b81 , \14990 , \14991 , \14992 , \14993 , \14994 , \14995_nG2a76 , \14996 , \14997 ,
         \14998 , \14999 , \15000 , \15001_nG2998 , \15002 , \15003 , \15004 , \15005 , \15006 , \15007_nG2894 ,
         \15008 , \15009 , \15010 , \15011 , \15012 , \15013_nG27bf , \15014 , \15015 , \15016 , \15017 ,
         \15018 , \15019_nG26e7 , \15020 ;
buf \U$labajz1574 ( R_267_b0ecd58, \7666 );
buf \U$labajz1575 ( R_268_b0ece00, \7671 );
buf \U$labajz1576 ( R_269_b0ecea8, \7677 );
buf \U$labajz1577 ( R_26a_b0ecf50, \7683 );
buf \U$labajz1578 ( R_26b_b0ecff8, \7689 );
buf \U$labajz1579 ( R_26c_b0ed0a0, \7695 );
buf \U$labajz1580 ( R_26d_b0ed148, \7701 );
buf \U$labajz1581 ( R_26e_b0ed1f0, \7708 );
buf \U$labajz1582 ( R_26f_b0ed298, \7717 );
buf \U$labajz1583 ( R_270_b0ed340, \7727 );
buf \U$labajz1584 ( R_271_b0ed3e8, \7743 );
buf \U$labajz1585 ( R_272_b0ed490, \7749 );
buf \U$labajz1586 ( R_273_b0ed538, \7757 );
buf \U$labajz1587 ( R_274_b0ed5e0, \7773 );
buf \U$labajz1588 ( R_275_b0ed688, \7779 );
buf \U$labajz1589 ( R_276_b0ed730, \7785 );
buf \U$labajz1590 ( R_277_b0ed7d8, \7792 );
buf \U$labajz1591 ( R_278_b0ed880, \7804 );
buf \U$labajz1592 ( R_279_b0ed928, \7816 );
buf \U$labajz1593 ( R_27a_b0ed9d0, \7832 );
buf \U$labajz1594 ( R_27b_b0eda78, \7838 );
buf \U$labajz1595 ( R_27c_b0edb20, \7844 );
buf \U$labajz1596 ( R_27d_b0edbc8, \7850 );
buf \U$labajz1597 ( R_27e_b0edc70, \7856 );
buf \U$labajz1598 ( R_27f_b0edd18, \7862 );
buf \U$labajz1599 ( R_280_b0eddc0, \7868 );
buf \U$labajz1600 ( R_281_b0ede68, \7874 );
buf \U$labajz1601 ( R_282_b0edf10, \14828 );
buf \U$labajz1602 ( R_283_b0edfb8, \14834 );
buf \U$labajz1603 ( R_284_b0ee060, \14840 );
buf \U$labajz1604 ( R_285_b0ee108, \14846 );
buf \U$labajz1605 ( R_286_b0ee1b0, \14852 );
buf \U$labajz1606 ( R_287_b0ee258, \14858 );
buf \U$labajz1607 ( R_288_b0ee300, \14864 );
buf \U$labajz1608 ( R_289_b0ee3a8, \14870 );
buf \U$labajz1609 ( R_28a_b0ee450, \14877 );
buf \U$labajz1610 ( R_28b_b0ee4f8, \14886 );
buf \U$labajz1611 ( R_28c_b0ee5a0, \14897 );
buf \U$labajz1612 ( R_28d_b0ee648, \14903 );
buf \U$labajz1613 ( R_28e_b0ee6f0, \14910 );
buf \U$labajz1614 ( R_28f_b0ee798, \14921 );
buf \U$labajz1615 ( R_290_b0ee840, \14927 );
buf \U$labajz1616 ( R_291_b0ee8e8, \14933 );
buf \U$labajz1617 ( R_292_b0ee990, \14940 );
buf \U$labajz1618 ( R_293_b0eea38, \14950 );
buf \U$labajz1619 ( R_294_b0eeae0, \14962 );
buf \U$labajz1620 ( R_295_b0eeb88, \14978 );
buf \U$labajz1621 ( R_296_b0eec30, \14984 );
buf \U$labajz1622 ( R_297_b0eecd8, \14990 );
buf \U$labajz1623 ( R_298_b0eed80, \14996 );
buf \U$labajz1624 ( R_299_b0eee28, \15002 );
buf \U$labajz1625 ( R_29a_b0eeed0, \15008 );
buf \U$labajz1626 ( R_29b_b0eef78, \15014 );
buf \U$labajz1627 ( R_29c_b0ef020, \15020 );
and \U$1 ( \651 , RIaa97770_3, RIaa977e8_4);
nand \U$2 ( \652 , RIaa976f8_2, \651 );
not \U$3 ( \653 , \652 );
nand \U$4 ( \654 , \653 , RIaa97860_5);
not \U$5 ( \655 , \654 );
nand \U$6 ( \656 , \655 , RIaa978d8_6);
not \U$7 ( \657 , \656 );
nand \U$8 ( \658 , \657 , RIaa97950_7);
not \U$9 ( \659 , \658 );
nand \U$10 ( \660 , \659 , RIaa979c8_8);
not \U$11 ( \661 , \660 );
nand \U$12 ( \662 , \661 , RIaa97ba8_12);
not \U$13 ( \663 , \662 );
nand \U$14 ( \664 , \663 , RIaa97b30_11);
not \U$15 ( \665 , \664 );
nand \U$16 ( \666 , \665 , RIaa97ab8_10);
not \U$17 ( \667 , \666 );
nand \U$18 ( \668 , \667 , RIaa97a40_9);
not \U$19 ( \669 , \668 );
not \U$20 ( \670 , RIaa97680_1);
and \U$21 ( \671 , \669 , \670 );
and \U$22 ( \672 , \668 , RIaa97680_1);
nor \U$23 ( \673 , \671 , \672 );
nor \U$24 ( \674 , RIaa9e958_246, RIaa9e8e0_245, RIaa9e700_241, RIaa9e7f0_243);
nor \U$25 ( \675 , RIaa9e688_240, RIaa9e778_242, RIaa9e868_244, RIaa9e9d0_247);
nand \U$26 ( \676 , \674 , \675 );
nor \U$27 ( \677 , \676 , RIaa97d88_16);
nand \U$28 ( \678 , RIaa97c20_13, \677 );
nor \U$29 ( \679 , \678 , RIaa97e00_17);
not \U$30 ( \680 , RIaa97d10_15);
nor \U$31 ( \681 , \680 , RIaa97c98_14);
and \U$32 ( \682 , \679 , \681 );
and \U$33 ( \683 , \682 , RIaa983a0_29);
not \U$34 ( \684 , RIaa97c98_14);
nor \U$35 ( \685 , \684 , RIaa97d10_15);
and \U$36 ( \686 , \679 , \685 );
and \U$37 ( \687 , \686 , RIaa982b0_27);
not \U$38 ( \688 , RIaa97e00_17);
nor \U$39 ( \689 , \678 , \688 );
and \U$40 ( \690 , \689 , \681 );
and \U$41 ( \691 , RIaa98418_30, \690 );
nor \U$42 ( \692 , \687 , \691 );
not \U$43 ( \693 , RIaa97c20_13);
nand \U$44 ( \694 , \693 , \677 );
nor \U$45 ( \695 , \694 , RIaa97e00_17);
and \U$46 ( \696 , \695 , \685 );
and \U$47 ( \697 , \696 , RIaa98580_33);
nor \U$48 ( \698 , \694 , \688 );
and \U$49 ( \699 , \698 , \681 );
and \U$50 ( \700 , RIaa98058_22, \699 );
nor \U$51 ( \701 , \697 , \700 );
and \U$52 ( \702 , \695 , \681 );
and \U$53 ( \703 , \702 , RIaa97fe0_21);
nor \U$54 ( \704 , RIaa97d10_15, RIaa97c98_14);
not \U$55 ( \705 , \704 );
nor \U$56 ( \706 , \705 , RIaa97e00_17, RIaa97c20_13);
not \U$57 ( \707 , \676 );
and \U$58 ( \708 , \706 , \707 , RIaa97d88_16);
nand \U$59 ( \709 , RIaa97f68_20, \708 );
not \U$60 ( \710 , \709 );
nor \U$61 ( \711 , \703 , \710 );
and \U$62 ( \712 , \689 , \685 );
and \U$63 ( \713 , \712 , RIaa98328_28);
not \U$64 ( \714 , \677 );
and \U$65 ( \715 , RIaa97d10_15, RIaa97c98_14);
nand \U$66 ( \716 , RIaa97e00_17, \715 , RIaa97c20_13);
nor \U$67 ( \717 , \714 , \716 );
and \U$68 ( \718 , RIaa98148_24, \717 );
nor \U$69 ( \719 , \713 , \718 );
nand \U$70 ( \720 , \692 , \701 , \711 , \719 );
and \U$71 ( \721 , \698 , \704 );
and \U$72 ( \722 , \721 , RIaa97ef0_19);
and \U$73 ( \723 , \679 , \704 );
and \U$74 ( \724 , RIaa981c0_25, \723 );
nor \U$75 ( \725 , \722 , \724 );
not \U$76 ( \726 , \725 );
nor \U$77 ( \727 , \683 , \720 , \726 );
and \U$78 ( \728 , \689 , \704 );
and \U$79 ( \729 , \728 , RIaa98238_26);
and \U$80 ( \730 , \698 , \715 );
and \U$81 ( \731 , RIaa985f8_34, \730 );
nor \U$82 ( \732 , \729 , \731 );
and \U$83 ( \733 , \695 , \715 );
and \U$84 ( \734 , \733 , RIaa98490_31);
and \U$85 ( \735 , \698 , \685 );
and \U$86 ( \736 , RIaa98508_32, \735 );
nor \U$87 ( \737 , \734 , \736 );
and \U$88 ( \738 , \677 , \706 );
and \U$89 ( \739 , \738 , RIaa97e78_18);
not \U$90 ( \740 , \715 );
nor \U$91 ( \741 , \740 , \678 );
and \U$92 ( \742 , \741 , \688 );
and \U$93 ( \743 , RIaa980d0_23, \742 );
nor \U$94 ( \744 , \739 , \743 );
nand \U$95 ( \745 , \727 , \732 , \737 , \744 );
buf \U$96 ( \746 , \745 );
not \U$97 ( \747 , RIaa97d88_16);
nor \U$98 ( \748 , \747 , \706 );
or \U$99 ( \749 , \748 , \676 );
buf \U$100 ( \750 , \749 );
_DC g11a6 ( \751_nG11a6 , \746 , \750 );
xor \U$101 ( \752 , \673 , \751_nG11a6 );
not \U$102 ( \753 , \666 );
not \U$103 ( \754 , RIaa97a40_9);
and \U$104 ( \755 , \753 , \754 );
and \U$105 ( \756 , \666 , RIaa97a40_9);
nor \U$106 ( \757 , \755 , \756 );
and \U$107 ( \758 , RIaa98b98_46, \682 );
and \U$108 ( \759 , RIaa986e8_36, \738 );
and \U$109 ( \760 , \742 , RIaa987d8_38);
and \U$110 ( \761 , RIaa98c10_47, \690 );
nor \U$111 ( \762 , \760 , \761 );
and \U$112 ( \763 , \728 , RIaa98a30_43);
and \U$113 ( \764 , RIaa98850_39, \717 );
nor \U$114 ( \765 , \763 , \764 );
and \U$115 ( \766 , \696 , RIaa98b20_45);
and \U$116 ( \767 , RIaa98670_35, \721 );
nor \U$117 ( \768 , \766 , \767 );
and \U$118 ( \769 , \686 , RIaa98c88_48);
and \U$119 ( \770 , RIaa98aa8_44, \712 );
nor \U$120 ( \771 , \769 , \770 );
nand \U$121 ( \772 , \762 , \765 , \768 , \771 );
nor \U$122 ( \773 , \758 , \759 , \772 );
and \U$123 ( \774 , \702 , RIaa988c8_40);
and \U$124 ( \775 , RIaa98940_41, \699 );
nor \U$125 ( \776 , \774 , \775 );
nand \U$126 ( \777 , RIaa98760_37, \708 );
and \U$127 ( \778 , RIaa989b8_42, \723 );
and \U$128 ( \779 , RIaa98d00_49, \730 );
and \U$129 ( \780 , \733 , RIaa98d78_50);
and \U$130 ( \781 , RIaa98df0_51, \735 );
nor \U$131 ( \782 , \780 , \781 );
not \U$132 ( \783 , \782 );
nor \U$133 ( \784 , \778 , \779 , \783 );
nand \U$134 ( \785 , \773 , \776 , \777 , \784 );
buf \U$135 ( \786 , \785 );
_DC gfc6 ( \787_nGfc6 , \786 , \750 );
xor \U$136 ( \788 , \757 , \787_nGfc6 );
not \U$137 ( \789 , \664 );
not \U$138 ( \790 , RIaa97ab8_10);
and \U$139 ( \791 , \789 , \790 );
and \U$140 ( \792 , \664 , RIaa97ab8_10);
nor \U$141 ( \793 , \791 , \792 );
and \U$142 ( \794 , RIaa9e160_229, \717 );
and \U$143 ( \795 , RIaa9de90_223, \721 );
and \U$144 ( \796 , \686 , RIaa9e2c8_232);
and \U$145 ( \797 , RIaa9e430_235, \690 );
nor \U$146 ( \798 , \796 , \797 );
and \U$147 ( \799 , \723 , RIaa9e1d8_230);
and \U$148 ( \800 , RIaa9e4a8_236, \733 );
nor \U$149 ( \801 , \799 , \800 );
and \U$150 ( \802 , \738 , RIaa9df08_224);
and \U$151 ( \803 , RIaa9e598_238, \696 );
nor \U$152 ( \804 , \802 , \803 );
and \U$153 ( \805 , \682 , RIaa9e3b8_234);
and \U$154 ( \806 , RIaa9e250_231, \728 );
nor \U$155 ( \807 , \805 , \806 );
nand \U$156 ( \808 , \798 , \801 , \804 , \807 );
nor \U$157 ( \809 , \794 , \795 , \808 );
and \U$158 ( \810 , \702 , RIaa9dff8_226);
and \U$159 ( \811 , RIaa9e070_227, \699 );
nor \U$160 ( \812 , \810 , \811 );
nand \U$161 ( \813 , RIaa9df80_225, \708 );
and \U$162 ( \814 , RIaa9e0e8_228, \742 );
and \U$163 ( \815 , RIaa9e340_233, \712 );
and \U$164 ( \816 , \735 , RIaa9e520_237);
and \U$165 ( \817 , RIaa9e610_239, \730 );
nor \U$166 ( \818 , \816 , \817 );
not \U$167 ( \819 , \818 );
nor \U$168 ( \820 , \814 , \815 , \819 );
nand \U$169 ( \821 , \809 , \812 , \813 , \820 );
buf \U$170 ( \822 , \821 );
_DC gfc4 ( \823_nGfc4 , \822 , \750 );
xor \U$171 ( \824 , \793 , \823_nGfc4 );
and \U$172 ( \825 , \662 , RIaa97b30_11);
not \U$173 ( \826 , \662 );
not \U$174 ( \827 , RIaa97b30_11);
and \U$175 ( \828 , \826 , \827 );
nor \U$176 ( \829 , \825 , \828 );
and \U$177 ( \830 , \682 , RIaa9d878_210);
and \U$178 ( \831 , \686 , RIaa9d698_206);
and \U$179 ( \832 , RIaa9d8f0_211, \690 );
nor \U$180 ( \833 , \831 , \832 );
and \U$181 ( \834 , \733 , RIaa9d968_212);
and \U$182 ( \835 , RIaa9d9e0_213, \735 );
nor \U$183 ( \836 , \834 , \835 );
and \U$184 ( \837 , \696 , RIaa9d788_208);
nand \U$185 ( \838 , RIaa9db48_216, \708 );
not \U$186 ( \839 , \838 );
nor \U$187 ( \840 , \837 , \839 );
and \U$188 ( \841 , \712 , RIaa9d710_207);
and \U$189 ( \842 , RIaa9de18_222, \717 );
nor \U$190 ( \843 , \841 , \842 );
nand \U$191 ( \844 , \833 , \836 , \840 , \843 );
and \U$192 ( \845 , \723 , RIaa9dcb0_219);
and \U$193 ( \846 , RIaa9dc38_218, \699 );
nor \U$194 ( \847 , \845 , \846 );
not \U$195 ( \848 , \847 );
nor \U$196 ( \849 , \830 , \844 , \848 );
and \U$197 ( \850 , \728 , RIaa9dd28_220);
and \U$198 ( \851 , RIaa9d800_209, \730 );
nor \U$199 ( \852 , \850 , \851 );
and \U$200 ( \853 , \702 , RIaa9dbc0_217);
and \U$201 ( \854 , RIaa9da58_214, \721 );
nor \U$202 ( \855 , \853 , \854 );
and \U$203 ( \856 , \738 , RIaa9dad0_215);
and \U$204 ( \857 , RIaa9dda0_221, \742 );
nor \U$205 ( \858 , \856 , \857 );
nand \U$206 ( \859 , \849 , \852 , \855 , \858 );
buf \U$207 ( \860 , \859 );
_DC ge1a ( \861_nGe1a , \860 , \750 );
xor \U$208 ( \862 , \829 , \861_nGe1a );
not \U$209 ( \863 , \660 );
not \U$210 ( \864 , RIaa97ba8_12);
and \U$211 ( \865 , \863 , \864 );
and \U$212 ( \866 , \660 , RIaa97ba8_12);
nor \U$213 ( \867 , \865 , \866 );
and \U$214 ( \868 , \742 , RIaa98fd0_55);
and \U$215 ( \869 , \723 , RIaa99390_63);
and \U$216 ( \870 , RIaa99408_64, \728 );
nor \U$217 ( \871 , \869 , \870 );
and \U$218 ( \872 , \702 , RIaa99318_62);
and \U$219 ( \873 , RIaa992a0_61, \699 );
nor \U$220 ( \874 , \872 , \873 );
and \U$221 ( \875 , \721 , RIaa98e68_52);
nand \U$222 ( \876 , RIaa98f58_54, \708 );
not \U$223 ( \877 , \876 );
nor \U$224 ( \878 , \875 , \877 );
and \U$225 ( \879 , \682 , RIaa991b0_59);
and \U$226 ( \880 , RIaa99048_56, \717 );
nor \U$227 ( \881 , \879 , \880 );
nand \U$228 ( \882 , \871 , \874 , \878 , \881 );
and \U$229 ( \883 , \686 , RIaa99480_65);
and \U$230 ( \884 , RIaa994f8_66, \730 );
nor \U$231 ( \885 , \883 , \884 );
not \U$232 ( \886 , \885 );
nor \U$233 ( \887 , \868 , \882 , \886 );
and \U$234 ( \888 , \738 , RIaa98ee0_53);
and \U$235 ( \889 , RIaa990c0_57, \712 );
nor \U$236 ( \890 , \888 , \889 );
and \U$237 ( \891 , \696 , RIaa99138_58);
and \U$238 ( \892 , RIaa99570_67, \735 );
nor \U$239 ( \893 , \891 , \892 );
and \U$240 ( \894 , \733 , RIaa995e8_68);
and \U$241 ( \895 , RIaa99228_60, \690 );
nor \U$242 ( \896 , \894 , \895 );
nand \U$243 ( \897 , \887 , \890 , \893 , \896 );
buf \U$244 ( \898 , \897 );
_DC ge18 ( \899_nGe18 , \898 , \750 );
xor \U$245 ( \900 , \867 , \899_nGe18 );
not \U$246 ( \901 , \658 );
not \U$247 ( \902 , RIaa979c8_8);
and \U$248 ( \903 , \901 , \902 );
and \U$249 ( \904 , \658 , RIaa979c8_8);
nor \U$250 ( \905 , \903 , \904 );
and \U$251 ( \906 , \742 , RIaa999a8_76);
and \U$252 ( \907 , \686 , RIaa99cf0_83);
and \U$253 ( \908 , RIaa997c8_72, \690 );
nor \U$254 ( \909 , \907 , \908 );
and \U$255 ( \910 , \702 , RIaa99b10_79);
and \U$256 ( \911 , RIaa99a98_78, \699 );
nor \U$257 ( \912 , \910 , \911 );
and \U$258 ( \913 , \721 , RIaa99840_73);
nand \U$259 ( \914 , RIaa99930_75, \708 );
not \U$260 ( \915 , \914 );
nor \U$261 ( \916 , \913 , \915 );
and \U$262 ( \917 , \712 , RIaa99c78_82);
and \U$263 ( \918 , RIaa99a20_77, \717 );
nor \U$264 ( \919 , \917 , \918 );
nand \U$265 ( \920 , \909 , \912 , \916 , \919 );
and \U$266 ( \921 , \723 , RIaa99b88_80);
and \U$267 ( \922 , RIaa99750_71, \682 );
nor \U$268 ( \923 , \921 , \922 );
not \U$269 ( \924 , \923 );
nor \U$270 ( \925 , \906 , \920 , \924 );
and \U$271 ( \926 , \696 , RIaa99d68_84);
and \U$272 ( \927 , RIaa99660_69, \735 );
nor \U$273 ( \928 , \926 , \927 );
and \U$274 ( \929 , \733 , RIaa996d8_70);
and \U$275 ( \930 , RIaa99de0_85, \730 );
nor \U$276 ( \931 , \929 , \930 );
and \U$277 ( \932 , \738 , RIaa998b8_74);
and \U$278 ( \933 , RIaa99c00_81, \728 );
nor \U$279 ( \934 , \932 , \933 );
nand \U$280 ( \935 , \925 , \928 , \931 , \934 );
buf \U$281 ( \936 , \935 );
_DC ga83 ( \937_nGa83 , \936 , \750 );
xor \U$282 ( \938 , \905 , \937_nGa83 );
not \U$283 ( \939 , \656 );
not \U$284 ( \940 , RIaa97950_7);
and \U$285 ( \941 , \939 , \940 );
and \U$286 ( \942 , \656 , RIaa97950_7);
nor \U$287 ( \943 , \941 , \942 );
and \U$288 ( \944 , \686 , RIaa9a470_99);
and \U$289 ( \945 , \733 , RIaa9a3f8_98);
and \U$290 ( \946 , RIaa9a380_97, \735 );
nor \U$291 ( \947 , \945 , \946 );
and \U$292 ( \948 , \699 , RIaa9a128_92);
and \U$293 ( \949 , RIaa9a038_90, \717 );
nor \U$294 ( \950 , \948 , \949 );
and \U$295 ( \951 , \696 , RIaa9a290_95);
nand \U$296 ( \952 , RIaa99ed0_87, \708 );
not \U$297 ( \953 , \952 );
nor \U$298 ( \954 , \951 , \953 );
and \U$299 ( \955 , \702 , RIaa9a1a0_93);
and \U$300 ( \956 , RIaa99e58_86, \721 );
nor \U$301 ( \957 , \955 , \956 );
nand \U$302 ( \958 , \947 , \950 , \954 , \957 );
and \U$303 ( \959 , \723 , RIaa9a0b0_91);
and \U$304 ( \960 , RIaa9a4e8_100, \682 );
nor \U$305 ( \961 , \959 , \960 );
not \U$306 ( \962 , \961 );
nor \U$307 ( \963 , \944 , \958 , \962 );
and \U$308 ( \964 , \690 , RIaa9a560_101);
and \U$309 ( \965 , RIaa9a308_96, \712 );
nor \U$310 ( \966 , \964 , \965 );
and \U$311 ( \967 , \728 , RIaa9a218_94);
and \U$312 ( \968 , RIaa9a5d8_102, \730 );
nor \U$313 ( \969 , \967 , \968 );
and \U$314 ( \970 , \738 , RIaa99fc0_89);
and \U$315 ( \971 , RIaa99f48_88, \742 );
nor \U$316 ( \972 , \970 , \971 );
nand \U$317 ( \973 , \963 , \966 , \969 , \972 );
buf \U$318 ( \974 , \973 );
_DC ga81 ( \975_nGa81 , \974 , \750 );
xor \U$319 ( \976 , \943 , \975_nGa81 );
not \U$320 ( \977 , \654 );
not \U$321 ( \978 , RIaa978d8_6);
and \U$322 ( \979 , \977 , \978 );
and \U$323 ( \980 , \654 , RIaa978d8_6);
nor \U$324 ( \981 , \979 , \980 );
and \U$325 ( \982 , \717 , RIaa9a830_107);
and \U$326 ( \983 , RIaa9ab78_114, \682 );
and \U$327 ( \984 , \686 , RIaa9aa88_112);
and \U$328 ( \985 , RIaa9a8a8_108, \696 );
nor \U$329 ( \986 , \983 , \984 , \985 );
and \U$330 ( \987 , \728 , RIaa9add0_119);
and \U$331 ( \988 , RIaa9ab00_113, \690 );
nor \U$332 ( \989 , \987 , \988 );
and \U$333 ( \990 , \738 , RIaa9a6c8_104);
and \U$334 ( \991 , RIaa9a998_110, \735 );
nor \U$335 ( \992 , \990 , \991 );
and \U$336 ( \993 , \742 , RIaa9a7b8_106);
and \U$337 ( \994 , RIaa9a920_109, \712 );
nor \U$338 ( \995 , \993 , \994 );
nand \U$339 ( \996 , \986 , \989 , \992 , \995 );
and \U$340 ( \997 , \723 , RIaa9ad58_118);
and \U$341 ( \998 , RIaa9abf0_115, \730 );
nor \U$342 ( \999 , \997 , \998 );
not \U$343 ( \1000 , \999 );
nor \U$344 ( \1001 , \982 , \996 , \1000 );
and \U$345 ( \1002 , \702 , RIaa9ac68_116);
and \U$346 ( \1003 , RIaa9a650_103, \721 );
nor \U$347 ( \1004 , \1002 , \1003 );
nand \U$348 ( \1005 , RIaa9a740_105, \708 );
and \U$349 ( \1006 , \733 , RIaa9aa10_111);
and \U$350 ( \1007 , RIaa9ace0_117, \699 );
nor \U$351 ( \1008 , \1006 , \1007 );
nand \U$352 ( \1009 , \1001 , \1004 , \1005 , \1008 );
buf \U$353 ( \1010 , \1009 );
_DC ga12 ( \1011_nGa12 , \1010 , \750 );
xor \U$354 ( \1012 , \981 , \1011_nGa12 );
not \U$355 ( \1013 , \652 );
not \U$356 ( \1014 , RIaa97860_5);
and \U$357 ( \1015 , \1013 , \1014 );
and \U$358 ( \1016 , \652 , RIaa97860_5);
nor \U$359 ( \1017 , \1015 , \1016 );
and \U$360 ( \1018 , \686 , RIaa9d2d8_198);
and \U$361 ( \1019 , \728 , RIaa9d620_205);
and \U$362 ( \1020 , RIaa9d350_199, \690 );
nor \U$363 ( \1021 , \1019 , \1020 );
and \U$364 ( \1022 , \699 , RIaa9d4b8_202);
and \U$365 ( \1023 , RIaa9cf90_191, \717 );
nor \U$366 ( \1024 , \1022 , \1023 );
and \U$367 ( \1025 , \730 , RIaa9d440_201);
nand \U$368 ( \1026 , RIaa9cea0_189, \708 );
not \U$369 ( \1027 , \1026 );
nor \U$370 ( \1028 , \1025 , \1027 );
and \U$371 ( \1029 , \702 , RIaa9d530_203);
and \U$372 ( \1030 , RIaa9d008_192, \721 );
nor \U$373 ( \1031 , \1029 , \1030 );
nand \U$374 ( \1032 , \1021 , \1024 , \1028 , \1031 );
and \U$375 ( \1033 , \723 , RIaa9d5a8_204);
and \U$376 ( \1034 , RIaa9d3c8_200, \682 );
nor \U$377 ( \1035 , \1033 , \1034 );
not \U$378 ( \1036 , \1035 );
nor \U$379 ( \1037 , \1018 , \1032 , \1036 );
and \U$380 ( \1038 , \733 , RIaa9d260_197);
and \U$381 ( \1039 , RIaa9d0f8_194, \712 );
nor \U$382 ( \1040 , \1038 , \1039 );
and \U$383 ( \1041 , \696 , RIaa9d170_195);
and \U$384 ( \1042 , RIaa9d1e8_196, \735 );
nor \U$385 ( \1043 , \1041 , \1042 );
and \U$386 ( \1044 , \738 , RIaa9d080_193);
and \U$387 ( \1045 , RIaa9cf18_190, \742 );
nor \U$388 ( \1046 , \1044 , \1045 );
nand \U$389 ( \1047 , \1037 , \1040 , \1043 , \1046 );
buf \U$390 ( \1048 , \1047 );
_DC ga10 ( \1049_nGa10 , \1048 , \750 );
xor \U$391 ( \1050 , \1017 , \1049_nGa10 );
xnor \U$392 ( \1051 , RIaa976f8_2, \651 );
and \U$393 ( \1052 , \717 , RIaa9b028_124);
and \U$394 ( \1053 , RIaa9b370_131, \682 );
and \U$395 ( \1054 , \686 , RIaa9b280_129);
and \U$396 ( \1055 , RIaa9b0a0_125, \696 );
nor \U$397 ( \1056 , \1053 , \1054 , \1055 );
and \U$398 ( \1057 , \738 , RIaa9aec0_121);
and \U$399 ( \1058 , RIaa9b460_133, \723 );
nor \U$400 ( \1059 , \1057 , \1058 );
and \U$401 ( \1060 , \733 , RIaa9b208_128);
and \U$402 ( \1061 , RIaa9b190_127, \735 );
nor \U$403 ( \1062 , \1060 , \1061 );
and \U$404 ( \1063 , \742 , RIaa9afb0_123);
and \U$405 ( \1064 , RIaa9b118_126, \712 );
nor \U$406 ( \1065 , \1063 , \1064 );
nand \U$407 ( \1066 , \1056 , \1059 , \1062 , \1065 );
nand \U$408 ( \1067 , RIaa9af38_122, \708 );
not \U$409 ( \1068 , \1067 );
nor \U$410 ( \1069 , \1052 , \1066 , \1068 );
and \U$411 ( \1070 , \721 , RIaa9ae48_120);
and \U$412 ( \1071 , RIaa9b2f8_130, \690 );
nor \U$413 ( \1072 , \1070 , \1071 );
and \U$414 ( \1073 , \702 , RIaa9b5c8_136);
and \U$415 ( \1074 , RIaa9b550_135, \699 );
nor \U$416 ( \1075 , \1073 , \1074 );
and \U$417 ( \1076 , \728 , RIaa9b4d8_134);
and \U$418 ( \1077 , RIaa9b3e8_132, \730 );
nor \U$419 ( \1078 , \1076 , \1077 );
nand \U$420 ( \1079 , \1069 , \1072 , \1075 , \1078 );
buf \U$421 ( \1080 , \1079 );
_DC g9bb ( \1081_nG9bb , \1080 , \750 );
xor \U$422 ( \1082 , \1051 , \1081_nG9bb );
not \U$423 ( \1083 , RIaa977e8_4);
and \U$424 ( \1084 , RIaa97770_3, \1083 );
not \U$425 ( \1085 , RIaa97770_3);
and \U$426 ( \1086 , \1085 , RIaa977e8_4);
nor \U$427 ( \1087 , \1084 , \1086 );
and \U$428 ( \1088 , \717 , RIaa9ba00_145);
and \U$429 ( \1089 , RIaa9bb68_148, \682 );
and \U$430 ( \1090 , \686 , RIaa9ba78_146);
and \U$431 ( \1091 , RIaa9b6b8_138, \696 );
nor \U$432 ( \1092 , \1089 , \1090 , \1091 );
and \U$433 ( \1093 , \738 , RIaa9b898_142);
and \U$434 ( \1094 , RIaa9bd48_152, \723 );
nor \U$435 ( \1095 , \1093 , \1094 );
and \U$436 ( \1096 , \733 , RIaa9b7a8_140);
and \U$437 ( \1097 , RIaa9b730_139, \735 );
nor \U$438 ( \1098 , \1096 , \1097 );
and \U$439 ( \1099 , \742 , RIaa9b988_144);
and \U$440 ( \1100 , RIaa9b640_137, \712 );
nor \U$441 ( \1101 , \1099 , \1100 );
nand \U$442 ( \1102 , \1092 , \1095 , \1098 , \1101 );
nand \U$443 ( \1103 , RIaa9b910_143, \708 );
not \U$444 ( \1104 , \1103 );
nor \U$445 ( \1105 , \1088 , \1102 , \1104 );
and \U$446 ( \1106 , \721 , RIaa9b820_141);
and \U$447 ( \1107 , RIaa9baf0_147, \690 );
nor \U$448 ( \1108 , \1106 , \1107 );
and \U$449 ( \1109 , \702 , RIaa9bcd0_151);
and \U$450 ( \1110 , RIaa9bc58_150, \699 );
nor \U$451 ( \1111 , \1109 , \1110 );
and \U$452 ( \1112 , \728 , RIaa9bdc0_153);
and \U$453 ( \1113 , RIaa9bbe0_149, \730 );
nor \U$454 ( \1114 , \1112 , \1113 );
nand \U$455 ( \1115 , \1105 , \1108 , \1111 , \1114 );
buf \U$456 ( \1116 , \1115 );
_DC g9bd ( \1117_nG9bd , \1116 , \750 );
xor \U$457 ( \1118 , \1087 , \1117_nG9bd );
and \U$458 ( \1119 , RIaa9c180_161, \717 );
and \U$459 ( \1120 , RIaa9c540_169, \733 );
and \U$460 ( \1121 , \723 , RIaa9c450_167);
and \U$461 ( \1122 , RIaa9c360_165, \682 );
nor \U$462 ( \1123 , \1121 , \1122 );
and \U$463 ( \1124 , \702 , RIaa9bf28_156);
and \U$464 ( \1125 , RIaa9bfa0_157, \699 );
nor \U$465 ( \1126 , \1124 , \1125 );
and \U$466 ( \1127 , \738 , RIaa9c090_159);
and \U$467 ( \1128 , RIaa9c018_158, \721 );
nor \U$468 ( \1129 , \1127 , \1128 );
and \U$469 ( \1130 , \696 , RIaa9c2e8_164);
and \U$470 ( \1131 , RIaa9c270_163, \735 );
nor \U$471 ( \1132 , \1130 , \1131 );
nand \U$472 ( \1133 , \1123 , \1126 , \1129 , \1132 );
nor \U$473 ( \1134 , \1119 , \1120 , \1133 );
and \U$474 ( \1135 , \728 , RIaa9c4c8_168);
and \U$475 ( \1136 , RIaa9beb0_155, \730 );
nor \U$476 ( \1137 , \1135 , \1136 );
nand \U$477 ( \1138 , RIaa9c108_160, \708 );
and \U$478 ( \1139 , RIaa9be38_154, \686 );
and \U$479 ( \1140 , RIaa9c3d8_166, \690 );
and \U$480 ( \1141 , \742 , RIaa9c1f8_162);
and \U$481 ( \1142 , RIaa9c5b8_170, \712 );
nor \U$482 ( \1143 , \1141 , \1142 );
not \U$483 ( \1144 , \1143 );
nor \U$484 ( \1145 , \1139 , \1140 , \1144 );
nand \U$485 ( \1146 , \1134 , \1137 , \1138 , \1145 );
buf \U$486 ( \1147 , \1146 );
_DC g949 ( \1148_nG949 , \1147 , \750 );
xor \U$487 ( \1149 , RIaa977e8_4, \1148_nG949 );
and \U$488 ( \1150 , \686 , RIaa9cd38_186);
and \U$489 ( \1151 , \728 , RIaa9cb58_182);
and \U$490 ( \1152 , RIaa9cbd0_183, \690 );
nor \U$491 ( \1153 , \1151 , \1152 );
and \U$492 ( \1154 , \699 , RIaa9c978_178);
and \U$493 ( \1155 , RIaa9c810_175, \717 );
nor \U$494 ( \1156 , \1154 , \1155 );
and \U$495 ( \1157 , \730 , RIaa9cdb0_187);
nand \U$496 ( \1158 , RIaa9c720_173, \708 );
not \U$497 ( \1159 , \1158 );
nor \U$498 ( \1160 , \1157 , \1159 );
and \U$499 ( \1161 , \702 , RIaa9cae0_181);
and \U$500 ( \1162 , RIaa9c6a8_172, \721 );
nor \U$501 ( \1163 , \1161 , \1162 );
nand \U$502 ( \1164 , \1153 , \1156 , \1160 , \1163 );
and \U$503 ( \1165 , \723 , RIaa9ca68_180);
and \U$504 ( \1166 , RIaa9c9f0_179, \682 );
nor \U$505 ( \1167 , \1165 , \1166 );
not \U$506 ( \1168 , \1167 );
nor \U$507 ( \1169 , \1150 , \1164 , \1168 );
and \U$508 ( \1170 , \733 , RIaa9c900_177);
and \U$509 ( \1171 , RIaa9c888_176, \712 );
nor \U$510 ( \1172 , \1170 , \1171 );
and \U$511 ( \1173 , \696 , RIaa9ccc0_185);
and \U$512 ( \1174 , RIaa9cc48_184, \735 );
nor \U$513 ( \1175 , \1173 , \1174 );
and \U$514 ( \1176 , \738 , RIaa9c798_174);
and \U$515 ( \1177 , RIaa9c630_171, \742 );
nor \U$516 ( \1178 , \1176 , \1177 );
nand \U$517 ( \1179 , \1169 , \1172 , \1175 , \1178 );
buf \U$518 ( \1180 , \1179 );
_DC g947 ( \1181_nG947 , \1180 , \750 );
not \U$519 ( \1182 , RIaa9ce28_188);
nand \U$520 ( \1183 , \1181_nG947 , \1182 );
not \U$521 ( \1184 , \1183 );
and \U$522 ( \1185 , \1149 , \1184 );
and \U$523 ( \1186 , RIaa977e8_4, \1148_nG949 );
or \U$524 ( \1187 , \1185 , \1186 );
and \U$525 ( \1188 , \1118 , \1187 );
and \U$526 ( \1189 , \1087 , \1117_nG9bd );
or \U$527 ( \1190 , \1188 , \1189 );
and \U$528 ( \1191 , \1082 , \1190 );
and \U$529 ( \1192 , \1051 , \1081_nG9bb );
or \U$530 ( \1193 , \1191 , \1192 );
and \U$531 ( \1194 , \1050 , \1193 );
and \U$532 ( \1195 , \1017 , \1049_nGa10 );
or \U$533 ( \1196 , \1194 , \1195 );
and \U$534 ( \1197 , \1012 , \1196 );
and \U$535 ( \1198 , \981 , \1011_nGa12 );
or \U$536 ( \1199 , \1197 , \1198 );
and \U$537 ( \1200 , \976 , \1199 );
and \U$538 ( \1201 , \943 , \975_nGa81 );
or \U$539 ( \1202 , \1200 , \1201 );
and \U$540 ( \1203 , \938 , \1202 );
and \U$541 ( \1204 , \905 , \937_nGa83 );
or \U$542 ( \1205 , \1203 , \1204 );
and \U$543 ( \1206 , \900 , \1205 );
and \U$544 ( \1207 , \867 , \899_nGe18 );
or \U$545 ( \1208 , \1206 , \1207 );
and \U$546 ( \1209 , \862 , \1208 );
and \U$547 ( \1210 , \829 , \861_nGe1a );
or \U$548 ( \1211 , \1209 , \1210 );
and \U$549 ( \1212 , \824 , \1211 );
and \U$550 ( \1213 , \793 , \823_nGfc4 );
or \U$551 ( \1214 , \1212 , \1213 );
and \U$552 ( \1215 , \788 , \1214 );
and \U$553 ( \1216 , \757 , \787_nGfc6 );
or \U$554 ( \1217 , \1215 , \1216 );
and \U$555 ( \1218 , \752 , \1217 );
and \U$556 ( \1219 , \673 , \751_nG11a6 );
or \U$557 ( \1220 , \1218 , \1219 );
not \U$558 ( \1221 , \668 );
nand \U$559 ( \1222 , \1221 , RIaa97680_1);
nor \U$560 ( \1223 , \1220 , \1222 );
not \U$561 ( \1224 , \1223 );
and \U$562 ( \1225 , RIaa9f768_276, \730 );
and \U$563 ( \1226 , RIaa9f9c0_281, \712 );
and \U$564 ( \1227 , \721 , RIaa9f330_267);
and \U$565 ( \1228 , RIaa9f600_273, \742 );
nor \U$566 ( \1229 , \1227 , \1228 );
and \U$567 ( \1230 , \738 , RIaa9f510_271);
and \U$568 ( \1231 , RIaa9f3a8_268, \723 );
nor \U$569 ( \1232 , \1230 , \1231 );
and \U$570 ( \1233 , \702 , RIaa9f420_269);
and \U$571 ( \1234 , RIaa9f858_278, \699 );
nor \U$572 ( \1235 , \1233 , \1234 );
and \U$573 ( \1236 , \682 , RIaa9f6f0_275);
and \U$574 ( \1237 , RIaa9f678_274, \728 );
nor \U$575 ( \1238 , \1236 , \1237 );
nand \U$576 ( \1239 , \1229 , \1232 , \1235 , \1238 );
nor \U$577 ( \1240 , \1225 , \1226 , \1239 );
or \U$578 ( \1241 , \708 , \717 );
and \U$579 ( \1242 , \1241 , RIaa9f588_272);
and \U$580 ( \1243 , RIaa9f7e0_277, \690 );
nor \U$581 ( \1244 , \1242 , \1243 );
and \U$582 ( \1245 , \733 , RIaa9f2b8_266);
and \U$583 ( \1246 , RIaa9f948_280, \735 );
nor \U$584 ( \1247 , \1245 , \1246 );
and \U$585 ( \1248 , \696 , RIaa9f498_270);
and \U$586 ( \1249 , RIaa9f8d0_279, \686 );
nor \U$587 ( \1250 , \1248 , \1249 );
nand \U$588 ( \1251 , \1240 , \1244 , \1247 , \1250 );
buf \U$589 ( \1252 , \749 );
_DC g17dd ( \1253_nG17dd , \1251 , \1252 );
not \U$590 ( \1254 , \1253_nG17dd );
nor \U$591 ( \1255 , \1224 , \1254 );
xor \U$592 ( \1256 , \673 , \751_nG11a6 );
xor \U$593 ( \1257 , \1256 , \1217 );
not \U$594 ( \1258 , \1257 );
xor \U$595 ( \1259 , \757 , \787_nGfc6 );
xor \U$596 ( \1260 , \1259 , \1214 );
not \U$597 ( \1261 , \1260 );
and \U$598 ( \1262 , \1258 , \1261 );
and \U$599 ( \1263 , \1220 , \1222 );
nor \U$600 ( \1264 , \1263 , \1223 );
nor \U$601 ( \1265 , \1262 , \1264 );
not \U$602 ( \1266 , \1265 );
and \U$603 ( \1267 , RIaa9f1c8_264, \686 );
and \U$604 ( \1268 , RIaa9efe8_260, \712 );
and \U$605 ( \1269 , \733 , RIaa9ec28_252);
and \U$606 ( \1270 , RIaa9eb38_250, \742 );
nor \U$607 ( \1271 , \1269 , \1270 );
and \U$608 ( \1272 , \723 , RIaa9ed18_254);
and \U$609 ( \1273 , RIaa9f0d8_262, \730 );
nor \U$610 ( \1274 , \1272 , \1273 );
and \U$611 ( \1275 , \738 , RIaa9eac0_249);
and \U$612 ( \1276 , RIaa9ef70_259, \735 );
nor \U$613 ( \1277 , \1275 , \1276 );
and \U$614 ( \1278 , \682 , RIaa9eef8_258);
and \U$615 ( \1279 , RIaa9ee80_257, \728 );
nor \U$616 ( \1280 , \1278 , \1279 );
nand \U$617 ( \1281 , \1271 , \1274 , \1277 , \1280 );
nor \U$618 ( \1282 , \1267 , \1268 , \1281 );
and \U$619 ( \1283 , \696 , RIaa9ed90_255);
and \U$620 ( \1284 , RIaa9eca0_253, \721 );
nor \U$621 ( \1285 , \1283 , \1284 );
and \U$622 ( \1286 , \1241 , RIaa9ebb0_251);
and \U$623 ( \1287 , RIaa9f150_263, \699 );
nor \U$624 ( \1288 , \1286 , \1287 );
and \U$625 ( \1289 , \702 , RIaa9ee08_256);
and \U$626 ( \1290 , RIaa9f060_261, \690 );
nor \U$627 ( \1291 , \1289 , \1290 );
nand \U$628 ( \1292 , \1282 , \1285 , \1288 , \1291 );
_DC g18eb ( \1293_nG18eb , \1292 , \1252 );
or \U$629 ( \1294 , \1266 , \1293_nG18eb );
not \U$630 ( \1295 , \1293_nG18eb );
and \U$631 ( \1296 , \1264 , \1257 );
nor \U$632 ( \1297 , \1264 , \1257 );
xnor \U$633 ( \1298 , \1260 , \1257 );
not \U$634 ( \1299 , \1298 );
nor \U$635 ( \1300 , \1296 , \1297 , \1299 );
nand \U$636 ( \1301 , \1266 , \1300 );
or \U$637 ( \1302 , \1295 , \1301 );
or \U$638 ( \1303 , \1300 , \1266 );
nand \U$639 ( \1304 , \1294 , \1302 , \1303 );
xnor \U$640 ( \1305 , \1255 , \1304 );
nor \U$641 ( \1306 , \1265 , \1298 );
not \U$642 ( \1307 , \1306 );
or \U$643 ( \1308 , \1307 , \1295 );
or \U$644 ( \1309 , \1254 , \1301 );
or \U$645 ( \1310 , \1298 , \1295 );
or \U$646 ( \1311 , \1266 , \1253_nG17dd );
nand \U$647 ( \1312 , \1311 , \1303 );
nand \U$648 ( \1313 , \1310 , \1312 );
nand \U$649 ( \1314 , \1308 , \1309 , \1313 );
xor \U$650 ( \1315 , \793 , \823_nGfc4 );
xor \U$651 ( \1316 , \1315 , \1211 );
xor \U$652 ( \1317 , \829 , \861_nGe1a );
xor \U$653 ( \1318 , \1317 , \1208 );
nor \U$654 ( \1319 , \1316 , \1318 );
or \U$655 ( \1320 , \1260 , \1319 );
and \U$656 ( \1321 , \1314 , \1320 );
and \U$657 ( \1322 , RIaa9fee8_292, \690 );
and \U$658 ( \1323 , RIaa9fd08_288, \735 );
and \U$659 ( \1324 , \742 , RIaa9fc90_287);
and \U$660 ( \1325 , RIaa9fd80_289, \712 );
nor \U$661 ( \1326 , \1324 , \1325 );
and \U$662 ( \1327 , \702 , RIaa9fdf8_290);
and \U$663 ( \1328 , RIaaa0050_295, \723 );
nor \U$664 ( \1329 , \1327 , \1328 );
and \U$665 ( \1330 , \738 , RIaa9fba0_285);
and \U$666 ( \1331 , RIaaa0140_297, \721 );
nor \U$667 ( \1332 , \1330 , \1331 );
and \U$668 ( \1333 , \682 , RIaa9ffd8_294);
and \U$669 ( \1334 , RIaa9fab0_283, \686 );
nor \U$670 ( \1335 , \1333 , \1334 );
nand \U$671 ( \1336 , \1326 , \1329 , \1332 , \1335 );
nor \U$672 ( \1337 , \1322 , \1323 , \1336 );
and \U$673 ( \1338 , \1241 , RIaa9fc18_286);
and \U$674 ( \1339 , RIaa9fa38_282, \699 );
nor \U$675 ( \1340 , \1338 , \1339 );
and \U$676 ( \1341 , \696 , RIaaa00c8_296);
and \U$677 ( \1342 , RIaaa01b8_298, \733 );
nor \U$678 ( \1343 , \1341 , \1342 );
and \U$679 ( \1344 , \728 , RIaa9ff60_293);
and \U$680 ( \1345 , RIaa9fe70_291, \730 );
nor \U$681 ( \1346 , \1344 , \1345 );
nand \U$682 ( \1347 , \1337 , \1340 , \1343 , \1346 );
_DC g16d6 ( \1348_nG16d6 , \1347 , \1252 );
not \U$683 ( \1349 , \1348_nG16d6 );
nor \U$684 ( \1350 , \1224 , \1349 );
nor \U$685 ( \1351 , \1321 , \1350 );
xor \U$686 ( \1352 , \1305 , \1351 );
not \U$687 ( \1353 , \1352 );
not \U$688 ( \1354 , \1316 );
not \U$689 ( \1355 , \1260 );
or \U$690 ( \1356 , \1354 , \1355 );
or \U$691 ( \1357 , \1260 , \1316 );
nand \U$692 ( \1358 , \1356 , \1357 );
xor \U$693 ( \1359 , \1318 , \1316 );
nor \U$694 ( \1360 , \1358 , \1359 );
not \U$695 ( \1361 , \1360 );
not \U$696 ( \1362 , \1320 );
nor \U$697 ( \1363 , \1361 , \1362 );
not \U$698 ( \1364 , \1363 );
or \U$699 ( \1365 , \1364 , \1295 );
or \U$700 ( \1366 , \1361 , \1295 );
nand \U$701 ( \1367 , \1366 , \1362 );
nand \U$702 ( \1368 , \1365 , \1367 );
or \U$703 ( \1369 , \1307 , \1254 );
or \U$704 ( \1370 , \1349 , \1301 );
or \U$705 ( \1371 , \1298 , \1254 );
or \U$706 ( \1372 , \1266 , \1348_nG16d6 );
nand \U$707 ( \1373 , \1372 , \1303 );
nand \U$708 ( \1374 , \1371 , \1373 );
nand \U$709 ( \1375 , \1369 , \1370 , \1374 );
and \U$710 ( \1376 , \1368 , \1375 );
and \U$711 ( \1377 , \1314 , \1320 );
not \U$712 ( \1378 , \1314 );
and \U$713 ( \1379 , \1378 , \1362 );
nor \U$714 ( \1380 , \1377 , \1379 );
xor \U$715 ( \1381 , \1350 , \1380 );
and \U$716 ( \1382 , \1376 , \1381 );
and \U$717 ( \1383 , \1353 , \1382 );
or \U$718 ( \1384 , \1383 , \1265 );
and \U$719 ( \1385 , \1304 , \1255 );
and \U$720 ( \1386 , \1265 , \1383 );
nor \U$721 ( \1387 , \1385 , \1386 );
nand \U$722 ( \1388 , \1384 , \1387 );
not \U$723 ( \1389 , \1388 );
and \U$724 ( \1390 , \1223 , \1293_nG18eb );
and \U$725 ( \1391 , \1305 , \1351 );
nor \U$726 ( \1392 , \1390 , \1391 );
not \U$727 ( \1393 , \1392 );
and \U$728 ( \1394 , \1389 , \1393 );
and \U$729 ( \1395 , \1388 , \1392 );
nor \U$730 ( \1396 , \1394 , \1395 );
not \U$731 ( \1397 , \1396 );
xor \U$732 ( \1398 , \1353 , \1382 );
and \U$733 ( \1399 , \1253_nG17dd , \1363 );
and \U$734 ( \1400 , \1320 , \1359 );
and \U$735 ( \1401 , \1400 , \1293_nG18eb );
nand \U$736 ( \1402 , \1253_nG17dd , \1360 );
or \U$737 ( \1403 , \1320 , \1293_nG18eb );
or \U$738 ( \1404 , \1320 , \1359 );
nand \U$739 ( \1405 , \1403 , \1404 );
and \U$740 ( \1406 , \1402 , \1405 );
nor \U$741 ( \1407 , \1399 , \1401 , \1406 );
and \U$742 ( \1408 , \1348_nG16d6 , \1306 );
and \U$743 ( \1409 , RIaaa07d0_311, \1241 );
and \U$744 ( \1410 , RIaaa06e0_309, \733 );
and \U$745 ( \1411 , \742 , RIaaa0848_312);
and \U$746 ( \1412 , RIaaa0398_302, \712 );
nor \U$747 ( \1413 , \1411 , \1412 );
and \U$748 ( \1414 , \738 , RIaaa0758_310);
and \U$749 ( \1415 , RIaaa0488_304, \723 );
nor \U$750 ( \1416 , \1414 , \1415 );
and \U$751 ( \1417 , \702 , RIaaa0410_303);
and \U$752 ( \1418 , RIaaa0668_308, \721 );
nor \U$753 ( \1419 , \1417 , \1418 );
and \U$754 ( \1420 , \682 , RIaaa05f0_307);
and \U$755 ( \1421 , RIaaa08c0_313, \686 );
nor \U$756 ( \1422 , \1420 , \1421 );
nand \U$757 ( \1423 , \1413 , \1416 , \1419 , \1422 );
nor \U$758 ( \1424 , \1409 , \1410 , \1423 );
and \U$759 ( \1425 , \699 , RIaaa0938_314);
and \U$760 ( \1426 , RIaaa02a8_300, \690 );
nor \U$761 ( \1427 , \1425 , \1426 );
and \U$762 ( \1428 , \696 , RIaaa0500_305);
and \U$763 ( \1429 , RIaaa0320_301, \735 );
nor \U$764 ( \1430 , \1428 , \1429 );
and \U$765 ( \1431 , \728 , RIaaa0578_306);
and \U$766 ( \1432 , RIaaa0230_299, \730 );
nor \U$767 ( \1433 , \1431 , \1432 );
nand \U$768 ( \1434 , \1424 , \1427 , \1430 , \1433 );
_DC g15b1 ( \1435_nG15b1 , \1434 , \1252 );
or \U$769 ( \1436 , \1266 , \1435_nG15b1 );
nand \U$770 ( \1437 , \1436 , \1303 );
nand \U$771 ( \1438 , \1348_nG16d6 , \1299 );
and \U$772 ( \1439 , \1437 , \1438 );
not \U$773 ( \1440 , \1301 );
and \U$774 ( \1441 , \1435_nG15b1 , \1440 );
nor \U$775 ( \1442 , \1408 , \1439 , \1441 );
nand \U$776 ( \1443 , \1407 , \1442 );
xor \U$777 ( \1444 , \867 , \899_nGe18 );
xor \U$778 ( \1445 , \1444 , \1205 );
xor \U$779 ( \1446 , \905 , \937_nGa83 );
xor \U$780 ( \1447 , \1446 , \1202 );
nor \U$781 ( \1448 , \1445 , \1447 );
or \U$782 ( \1449 , \1318 , \1448 );
and \U$783 ( \1450 , \1443 , \1449 );
nor \U$784 ( \1451 , \1442 , \1407 );
nor \U$785 ( \1452 , \1450 , \1451 );
xor \U$786 ( \1453 , \1368 , \1375 );
not \U$787 ( \1454 , \1453 );
nand \U$788 ( \1455 , \1435_nG15b1 , \1223 );
not \U$789 ( \1456 , \1455 );
and \U$790 ( \1457 , \1454 , \1456 );
and \U$791 ( \1458 , \1453 , \1455 );
nor \U$792 ( \1459 , \1457 , \1458 );
nand \U$793 ( \1460 , \1452 , \1459 );
xor \U$794 ( \1461 , \1376 , \1381 );
and \U$795 ( \1462 , \1460 , \1461 );
and \U$796 ( \1463 , \1398 , \1462 );
not \U$797 ( \1464 , \1463 );
and \U$798 ( \1465 , \1397 , \1464 );
and \U$799 ( \1466 , \1396 , \1463 );
nor \U$800 ( \1467 , \1465 , \1466 );
not \U$801 ( \1468 , \1467 );
xor \U$802 ( \1469 , \1460 , \1461 );
not \U$803 ( \1470 , \1453 );
nor \U$804 ( \1471 , \1470 , \1455 );
xor \U$805 ( \1472 , \1469 , \1471 );
or \U$806 ( \1473 , \1459 , \1452 );
nand \U$807 ( \1474 , \1473 , \1460 );
not \U$808 ( \1475 , \1474 );
and \U$809 ( \1476 , RIaaa0a28_316, \723 );
and \U$810 ( \1477 , RIaaa0e60_325, \712 );
and \U$811 ( \1478 , \728 , RIaaa0b18_318);
and \U$812 ( \1479 , RIaaa1040_329, \742 );
nor \U$813 ( \1480 , \1478 , \1479 );
and \U$814 ( \1481 , \733 , RIaaa0c80_321);
and \U$815 ( \1482 , RIaaa0cf8_322, \730 );
nor \U$816 ( \1483 , \1481 , \1482 );
and \U$817 ( \1484 , \1241 , RIaaa0fc8_328);
and \U$818 ( \1485 , RIaaa0de8_324, \735 );
nor \U$819 ( \1486 , \1484 , \1485 );
and \U$820 ( \1487 , \696 , RIaaa0aa0_317);
and \U$821 ( \1488 , RIaaa1130_331, \699 );
nor \U$822 ( \1489 , \1487 , \1488 );
nand \U$823 ( \1490 , \1480 , \1483 , \1486 , \1489 );
nor \U$824 ( \1491 , \1476 , \1477 , \1490 );
and \U$825 ( \1492 , \721 , RIaaa0c08_320);
and \U$826 ( \1493 , RIaaa0b90_319, \682 );
nor \U$827 ( \1494 , \1492 , \1493 );
and \U$828 ( \1495 , \738 , RIaaa0f50_327);
and \U$829 ( \1496 , RIaaa0ed8_326, \702 );
nor \U$830 ( \1497 , \1495 , \1496 );
and \U$831 ( \1498 , \686 , RIaaa10b8_330);
and \U$832 ( \1499 , RIaaa0d70_323, \690 );
nor \U$833 ( \1500 , \1498 , \1499 );
nand \U$834 ( \1501 , \1491 , \1494 , \1497 , \1500 );
_DC g14c8 ( \1502_nG14c8 , \1501 , \1252 );
not \U$835 ( \1503 , \1502_nG14c8 );
nor \U$836 ( \1504 , \1224 , \1503 );
not \U$837 ( \1505 , \1449 );
not \U$838 ( \1506 , \1451 );
nand \U$839 ( \1507 , \1506 , \1443 );
not \U$840 ( \1508 , \1507 );
or \U$841 ( \1509 , \1505 , \1508 );
or \U$842 ( \1510 , \1507 , \1449 );
nand \U$843 ( \1511 , \1509 , \1510 );
xnor \U$844 ( \1512 , \1504 , \1511 );
not \U$845 ( \1513 , \1512 );
and \U$846 ( \1514 , \1348_nG16d6 , \1363 );
and \U$847 ( \1515 , \1400 , \1253_nG17dd );
nand \U$848 ( \1516 , \1348_nG16d6 , \1360 );
or \U$849 ( \1517 , \1320 , \1253_nG17dd );
nand \U$850 ( \1518 , \1517 , \1404 );
and \U$851 ( \1519 , \1516 , \1518 );
nor \U$852 ( \1520 , \1514 , \1515 , \1519 );
and \U$853 ( \1521 , \1318 , \1445 );
nor \U$854 ( \1522 , \1318 , \1445 );
xor \U$855 ( \1523 , \1445 , \1447 );
nor \U$856 ( \1524 , \1521 , \1522 , \1523 );
and \U$857 ( \1525 , \1524 , \1449 );
and \U$858 ( \1526 , \1293_nG18eb , \1525 );
not \U$859 ( \1527 , \1449 );
and \U$860 ( \1528 , \1295 , \1527 );
or \U$861 ( \1529 , \1524 , \1449 );
not \U$862 ( \1530 , \1529 );
nor \U$863 ( \1531 , \1526 , \1528 , \1530 );
or \U$864 ( \1532 , \1520 , \1531 );
and \U$865 ( \1533 , RIaaa20a8_364, \690 );
and \U$866 ( \1534 , RIaaa1f40_361, \735 );
and \U$867 ( \1535 , \742 , RIaaa1b80_353);
and \U$868 ( \1536 , RIaaa1fb8_362, \712 );
nor \U$869 ( \1537 , \1535 , \1536 );
and \U$870 ( \1538 , \738 , RIaaa1a90_351);
and \U$871 ( \1539 , RIaaa2198_366, \686 );
nor \U$872 ( \1540 , \1538 , \1539 );
and \U$873 ( \1541 , \702 , RIaaa1d60_357);
and \U$874 ( \1542 , RIaaa1c70_355, \721 );
nor \U$875 ( \1543 , \1541 , \1542 );
and \U$876 ( \1544 , \723 , RIaaa1ce8_356);
and \U$877 ( \1545 , RIaaa1ec8_360, \682 );
nor \U$878 ( \1546 , \1544 , \1545 );
nand \U$879 ( \1547 , \1537 , \1540 , \1543 , \1546 );
nor \U$880 ( \1548 , \1533 , \1534 , \1547 );
and \U$881 ( \1549 , \1241 , RIaaa1b08_352);
and \U$882 ( \1550 , RIaaa2120_365, \699 );
nor \U$883 ( \1551 , \1549 , \1550 );
and \U$884 ( \1552 , \696 , RIaaa1dd8_358);
and \U$885 ( \1553 , RIaaa1bf8_354, \733 );
nor \U$886 ( \1554 , \1552 , \1553 );
and \U$887 ( \1555 , \728 , RIaaa1e50_359);
and \U$888 ( \1556 , RIaaa2030_363, \730 );
nor \U$889 ( \1557 , \1555 , \1556 );
nand \U$890 ( \1558 , \1548 , \1551 , \1554 , \1557 );
_DC g13c8 ( \1559_nG13c8 , \1558 , \1252 );
nand \U$891 ( \1560 , \1559_nG13c8 , \1223 );
and \U$892 ( \1561 , \1435_nG15b1 , \1306 );
or \U$893 ( \1562 , \1266 , \1502_nG14c8 );
nand \U$894 ( \1563 , \1562 , \1303 );
nand \U$895 ( \1564 , \1435_nG15b1 , \1299 );
and \U$896 ( \1565 , \1563 , \1564 );
and \U$897 ( \1566 , \1502_nG14c8 , \1440 );
nor \U$898 ( \1567 , \1561 , \1565 , \1566 );
or \U$899 ( \1568 , \1560 , \1567 );
nand \U$900 ( \1569 , \1532 , \1568 );
nand \U$901 ( \1570 , \1513 , \1569 );
nor \U$902 ( \1571 , \1475 , \1570 );
xor \U$903 ( \1572 , \1472 , \1571 );
and \U$904 ( \1573 , \1511 , \1504 );
xor \U$905 ( \1574 , \943 , \975_nGa81 );
xor \U$906 ( \1575 , \1574 , \1199 );
xor \U$907 ( \1576 , \981 , \1011_nGa12 );
xor \U$908 ( \1577 , \1576 , \1196 );
nor \U$909 ( \1578 , \1575 , \1577 );
or \U$910 ( \1579 , \1447 , \1578 );
not \U$911 ( \1580 , \1579 );
and \U$912 ( \1581 , \1435_nG15b1 , \1363 );
and \U$913 ( \1582 , \1400 , \1348_nG16d6 );
nand \U$914 ( \1583 , \1435_nG15b1 , \1360 );
or \U$915 ( \1584 , \1320 , \1348_nG16d6 );
nand \U$916 ( \1585 , \1584 , \1404 );
and \U$917 ( \1586 , \1583 , \1585 );
nor \U$918 ( \1587 , \1581 , \1582 , \1586 );
nand \U$919 ( \1588 , \1293_nG18eb , \1523 );
or \U$920 ( \1589 , \1449 , \1253_nG17dd );
nand \U$921 ( \1590 , \1589 , \1529 );
and \U$922 ( \1591 , \1588 , \1590 );
and \U$923 ( \1592 , \1525 , \1253_nG17dd );
not \U$924 ( \1593 , \1523 );
nor \U$925 ( \1594 , \1527 , \1593 );
and \U$926 ( \1595 , \1293_nG18eb , \1594 );
nor \U$927 ( \1596 , \1591 , \1592 , \1595 );
nor \U$928 ( \1597 , \1587 , \1596 );
not \U$929 ( \1598 , \1597 );
nand \U$930 ( \1599 , \1596 , \1587 );
nand \U$931 ( \1600 , \1598 , \1599 );
not \U$932 ( \1601 , \1600 );
or \U$933 ( \1602 , \1580 , \1601 );
or \U$934 ( \1603 , \1600 , \1579 );
nand \U$935 ( \1604 , \1602 , \1603 );
and \U$936 ( \1605 , RIaaa1310_335, \1241 );
and \U$937 ( \1606 , RIaaa17c0_345, \712 );
and \U$938 ( \1607 , \682 , RIaaa16d0_343);
and \U$939 ( \1608 , RIaaa19a0_349, \686 );
nor \U$940 ( \1609 , \1607 , \1608 );
and \U$941 ( \1610 , \702 , RIaaa1568_340);
and \U$942 ( \1611 , RIaaa1478_338, \721 );
nor \U$943 ( \1612 , \1610 , \1611 );
and \U$944 ( \1613 , \738 , RIaaa1298_334);
and \U$945 ( \1614 , RIaaa1400_337, \733 );
nor \U$946 ( \1615 , \1613 , \1614 );
and \U$947 ( \1616 , \723 , RIaaa14f0_339);
and \U$948 ( \1617 , RIaaa1838_346, \730 );
nor \U$949 ( \1618 , \1616 , \1617 );
nand \U$950 ( \1619 , \1609 , \1612 , \1615 , \1618 );
nor \U$951 ( \1620 , \1605 , \1606 , \1619 );
and \U$952 ( \1621 , \699 , RIaaa1928_348);
and \U$953 ( \1622 , RIaaa18b0_347, \690 );
nor \U$954 ( \1623 , \1621 , \1622 );
and \U$955 ( \1624 , \696 , RIaaa15e0_341);
and \U$956 ( \1625 , RIaaa1748_344, \735 );
nor \U$957 ( \1626 , \1624 , \1625 );
and \U$958 ( \1627 , \728 , RIaaa1658_342);
and \U$959 ( \1628 , RIaaa1388_336, \742 );
nor \U$960 ( \1629 , \1627 , \1628 );
nand \U$961 ( \1630 , \1620 , \1623 , \1626 , \1629 );
_DC g12c9 ( \1631_nG12c9 , \1630 , \1252 );
not \U$962 ( \1632 , \1631_nG12c9 );
nor \U$963 ( \1633 , \1224 , \1632 );
or \U$964 ( \1634 , \1307 , \1503 );
not \U$965 ( \1635 , \1559_nG13c8 );
or \U$966 ( \1636 , \1635 , \1301 );
or \U$967 ( \1637 , \1298 , \1503 );
or \U$968 ( \1638 , \1266 , \1559_nG13c8 );
nand \U$969 ( \1639 , \1638 , \1303 );
nand \U$970 ( \1640 , \1637 , \1639 );
nand \U$971 ( \1641 , \1634 , \1636 , \1640 );
xor \U$972 ( \1642 , \1633 , \1641 );
and \U$973 ( \1643 , \1604 , \1642 );
not \U$974 ( \1644 , \1575 );
not \U$975 ( \1645 , \1447 );
or \U$976 ( \1646 , \1644 , \1645 );
or \U$977 ( \1647 , \1447 , \1575 );
nand \U$978 ( \1648 , \1646 , \1647 );
xor \U$979 ( \1649 , \1577 , \1575 );
nor \U$980 ( \1650 , \1648 , \1649 );
not \U$981 ( \1651 , \1650 );
not \U$982 ( \1652 , \1579 );
nor \U$983 ( \1653 , \1651 , \1652 );
not \U$984 ( \1654 , \1653 );
or \U$985 ( \1655 , \1654 , \1295 );
or \U$986 ( \1656 , \1651 , \1295 );
nand \U$987 ( \1657 , \1656 , \1652 );
nand \U$988 ( \1658 , \1655 , \1657 );
not \U$989 ( \1659 , \1594 );
or \U$990 ( \1660 , \1659 , \1254 );
not \U$991 ( \1661 , \1525 );
or \U$992 ( \1662 , \1349 , \1661 );
or \U$993 ( \1663 , \1593 , \1254 );
or \U$994 ( \1664 , \1449 , \1348_nG16d6 );
nand \U$995 ( \1665 , \1664 , \1529 );
nand \U$996 ( \1666 , \1663 , \1665 );
nand \U$997 ( \1667 , \1660 , \1662 , \1666 );
and \U$998 ( \1668 , \1658 , \1667 );
and \U$999 ( \1669 , \1559_nG13c8 , \1306 );
or \U$1000 ( \1670 , \1266 , \1631_nG12c9 );
nand \U$1001 ( \1671 , \1670 , \1303 );
nand \U$1002 ( \1672 , \1559_nG13c8 , \1299 );
and \U$1003 ( \1673 , \1671 , \1672 );
and \U$1004 ( \1674 , \1631_nG12c9 , \1440 );
nor \U$1005 ( \1675 , \1669 , \1673 , \1674 );
and \U$1006 ( \1676 , \1502_nG14c8 , \1363 );
and \U$1007 ( \1677 , \1400 , \1435_nG15b1 );
nand \U$1008 ( \1678 , \1502_nG14c8 , \1360 );
or \U$1009 ( \1679 , \1320 , \1435_nG15b1 );
nand \U$1010 ( \1680 , \1679 , \1404 );
and \U$1011 ( \1681 , \1678 , \1680 );
nor \U$1012 ( \1682 , \1676 , \1677 , \1681 );
and \U$1013 ( \1683 , \1675 , \1682 );
and \U$1014 ( \1684 , RIaaa3098_398, \742 );
and \U$1015 ( \1685 , RIaaa2e40_393, \735 );
and \U$1016 ( \1686 , \682 , RIaaa2a08_384);
and \U$1017 ( \1687 , RIaaa2f30_395, \686 );
nor \U$1018 ( \1688 , \1686 , \1687 );
and \U$1019 ( \1689 , \702 , RIaaa2eb8_394);
and \U$1020 ( \1690 , RIaaa2c60_389, \721 );
nor \U$1021 ( \1691 , \1689 , \1690 );
and \U$1022 ( \1692 , \733 , RIaaa2be8_388);
and \U$1023 ( \1693 , RIaaa2d50_391, \730 );
nor \U$1024 ( \1694 , \1692 , \1693 );
and \U$1025 ( \1695 , \738 , RIaaa3020_397);
and \U$1026 ( \1696 , RIaaa2b70_387, \723 );
nor \U$1027 ( \1697 , \1695 , \1696 );
nand \U$1028 ( \1698 , \1688 , \1691 , \1694 , \1697 );
nor \U$1029 ( \1699 , \1684 , \1685 , \1698 );
and \U$1030 ( \1700 , \696 , RIaaa2af8_386);
and \U$1031 ( \1701 , RIaaa2a80_385, \728 );
nor \U$1032 ( \1702 , \1700 , \1701 );
and \U$1033 ( \1703 , \1241 , RIaaa3110_399);
and \U$1034 ( \1704 , RIaaa2fa8_396, \699 );
nor \U$1035 ( \1705 , \1703 , \1704 );
and \U$1036 ( \1706 , \690 , RIaaa2cd8_390);
and \U$1037 ( \1707 , RIaaa2dc8_392, \712 );
nor \U$1038 ( \1708 , \1706 , \1707 );
nand \U$1039 ( \1709 , \1699 , \1702 , \1705 , \1708 );
_DC g11c1 ( \1710_nG11c1 , \1709 , \1252 );
nand \U$1040 ( \1711 , \1710_nG11c1 , \1223 );
or \U$1041 ( \1712 , \1683 , \1711 );
or \U$1042 ( \1713 , \1675 , \1682 );
nand \U$1043 ( \1714 , \1712 , \1713 );
and \U$1044 ( \1715 , \1668 , \1714 );
and \U$1045 ( \1716 , \1643 , \1715 );
and \U$1046 ( \1717 , \1599 , \1579 );
and \U$1047 ( \1718 , \1633 , \1641 );
nor \U$1048 ( \1719 , \1717 , \1718 , \1597 );
xor \U$1049 ( \1720 , \1560 , \1567 );
not \U$1050 ( \1721 , \1720 );
xnor \U$1051 ( \1722 , \1531 , \1520 );
not \U$1052 ( \1723 , \1722 );
and \U$1053 ( \1724 , \1721 , \1723 );
and \U$1054 ( \1725 , \1720 , \1722 );
nor \U$1055 ( \1726 , \1724 , \1725 );
nand \U$1056 ( \1727 , \1719 , \1726 );
xor \U$1057 ( \1728 , \1716 , \1727 );
not \U$1058 ( \1729 , \1569 );
not \U$1059 ( \1730 , \1512 );
or \U$1060 ( \1731 , \1729 , \1730 );
or \U$1061 ( \1732 , \1512 , \1569 );
nand \U$1062 ( \1733 , \1731 , \1732 );
and \U$1063 ( \1734 , \1728 , \1733 );
and \U$1064 ( \1735 , \1716 , \1727 );
or \U$1065 ( \1736 , \1734 , \1735 );
nor \U$1066 ( \1737 , \1573 , \1736 );
not \U$1067 ( \1738 , \1474 );
not \U$1068 ( \1739 , \1570 );
and \U$1069 ( \1740 , \1738 , \1739 );
and \U$1070 ( \1741 , \1474 , \1570 );
nor \U$1071 ( \1742 , \1740 , \1741 );
nor \U$1072 ( \1743 , \1737 , \1742 );
xor \U$1073 ( \1744 , \1572 , \1743 );
and \U$1074 ( \1745 , \1631_nG12c9 , \1306 );
or \U$1075 ( \1746 , \1266 , \1710_nG11c1 );
nand \U$1076 ( \1747 , \1746 , \1303 );
nand \U$1077 ( \1748 , \1631_nG12c9 , \1299 );
and \U$1078 ( \1749 , \1747 , \1748 );
and \U$1079 ( \1750 , \1710_nG11c1 , \1440 );
nor \U$1080 ( \1751 , \1745 , \1749 , \1750 );
and \U$1081 ( \1752 , \1559_nG13c8 , \1363 );
and \U$1082 ( \1753 , \1400 , \1502_nG14c8 );
nand \U$1083 ( \1754 , \1559_nG13c8 , \1360 );
or \U$1084 ( \1755 , \1320 , \1502_nG14c8 );
nand \U$1085 ( \1756 , \1755 , \1404 );
and \U$1086 ( \1757 , \1754 , \1756 );
nor \U$1087 ( \1758 , \1752 , \1753 , \1757 );
and \U$1088 ( \1759 , \1751 , \1758 );
not \U$1089 ( \1760 , \1759 );
and \U$1090 ( \1761 , RIaaa2648_376, \721 );
and \U$1091 ( \1762 , RIaaa27b0_379, \686 );
and \U$1092 ( \1763 , \742 , RIaaa2918_382);
and \U$1093 ( \1764 , RIaaa2210_367, \712 );
nor \U$1094 ( \1765 , \1763 , \1764 );
and \U$1095 ( \1766 , \696 , RIaaa25d0_375);
and \U$1096 ( \1767 , RIaaa2738_378, \699 );
nor \U$1097 ( \1768 , \1766 , \1767 );
and \U$1098 ( \1769 , \1241 , RIaaa28a0_381);
and \U$1099 ( \1770 , RIaaa2288_368, \735 );
nor \U$1100 ( \1771 , \1769 , \1770 );
and \U$1101 ( \1772 , \728 , RIaaa2468_372);
and \U$1102 ( \1773 , RIaaa2378_370, \690 );
nor \U$1103 ( \1774 , \1772 , \1773 );
nand \U$1104 ( \1775 , \1765 , \1768 , \1771 , \1774 );
nor \U$1105 ( \1776 , \1761 , \1762 , \1775 );
and \U$1106 ( \1777 , \738 , RIaaa2828_380);
and \U$1107 ( \1778 , RIaaa2300_369, \730 );
nor \U$1108 ( \1779 , \1777 , \1778 );
and \U$1109 ( \1780 , \702 , RIaaa23f0_371);
and \U$1110 ( \1781 , RIaaa26c0_377, \733 );
nor \U$1111 ( \1782 , \1780 , \1781 );
and \U$1112 ( \1783 , \723 , RIaaa2558_374);
and \U$1113 ( \1784 , RIaaa24e0_373, \682 );
nor \U$1114 ( \1785 , \1783 , \1784 );
nand \U$1115 ( \1786 , \1776 , \1779 , \1782 , \1785 );
_DC g10e2 ( \1787_nG10e2 , \1786 , \1252 );
nand \U$1116 ( \1788 , \1787_nG10e2 , \1223 );
not \U$1117 ( \1789 , \1788 );
and \U$1118 ( \1790 , \1760 , \1789 );
nor \U$1119 ( \1791 , \1751 , \1758 );
nor \U$1120 ( \1792 , \1790 , \1791 );
or \U$1121 ( \1793 , \1654 , \1254 );
and \U$1122 ( \1794 , \1579 , \1649 );
not \U$1123 ( \1795 , \1794 );
or \U$1124 ( \1796 , \1295 , \1795 );
or \U$1125 ( \1797 , \1651 , \1254 );
or \U$1126 ( \1798 , \1579 , \1293_nG18eb );
or \U$1127 ( \1799 , \1579 , \1649 );
nand \U$1128 ( \1800 , \1798 , \1799 );
nand \U$1129 ( \1801 , \1797 , \1800 );
nand \U$1130 ( \1802 , \1793 , \1796 , \1801 );
xor \U$1131 ( \1803 , \1051 , \1081_nG9bb );
xor \U$1132 ( \1804 , \1803 , \1190 );
not \U$1133 ( \1805 , \1804 );
xor \U$1134 ( \1806 , \1017 , \1049_nGa10 );
xor \U$1135 ( \1807 , \1806 , \1193 );
not \U$1136 ( \1808 , \1807 );
and \U$1137 ( \1809 , \1805 , \1808 );
or \U$1138 ( \1810 , \1577 , \1809 );
and \U$1139 ( \1811 , \1802 , \1810 );
not \U$1140 ( \1812 , \1802 );
not \U$1141 ( \1813 , \1810 );
and \U$1142 ( \1814 , \1812 , \1813 );
nand \U$1143 ( \1815 , \1348_nG16d6 , \1523 );
or \U$1144 ( \1816 , \1449 , \1435_nG15b1 );
nand \U$1145 ( \1817 , \1816 , \1529 );
and \U$1146 ( \1818 , \1815 , \1817 );
and \U$1147 ( \1819 , \1525 , \1435_nG15b1 );
and \U$1148 ( \1820 , \1348_nG16d6 , \1594 );
nor \U$1149 ( \1821 , \1818 , \1819 , \1820 );
nor \U$1150 ( \1822 , \1814 , \1821 );
nor \U$1151 ( \1823 , \1811 , \1822 );
nor \U$1152 ( \1824 , \1792 , \1823 );
xor \U$1153 ( \1825 , \1658 , \1667 );
not \U$1154 ( \1826 , \1825 );
not \U$1155 ( \1827 , \1713 );
nor \U$1156 ( \1828 , \1827 , \1683 );
not \U$1157 ( \1829 , \1828 );
not \U$1158 ( \1830 , \1711 );
and \U$1159 ( \1831 , \1829 , \1830 );
and \U$1160 ( \1832 , \1828 , \1711 );
nor \U$1161 ( \1833 , \1831 , \1832 );
nor \U$1162 ( \1834 , \1826 , \1833 );
and \U$1163 ( \1835 , \1824 , \1834 );
xor \U$1164 ( \1836 , \1668 , \1714 );
xor \U$1165 ( \1837 , \1604 , \1642 );
and \U$1166 ( \1838 , \1836 , \1837 );
xor \U$1167 ( \1839 , \1835 , \1838 );
or \U$1168 ( \1840 , \1726 , \1719 );
nand \U$1169 ( \1841 , \1840 , \1727 );
and \U$1170 ( \1842 , \1839 , \1841 );
and \U$1171 ( \1843 , \1835 , \1838 );
or \U$1172 ( \1844 , \1842 , \1843 );
not \U$1173 ( \1845 , \1720 );
nor \U$1174 ( \1846 , \1845 , \1722 );
xor \U$1175 ( \1847 , \1844 , \1846 );
xor \U$1176 ( \1848 , \1716 , \1727 );
xor \U$1177 ( \1849 , \1848 , \1733 );
and \U$1178 ( \1850 , \1847 , \1849 );
and \U$1179 ( \1851 , \1844 , \1846 );
or \U$1180 ( \1852 , \1850 , \1851 );
and \U$1181 ( \1853 , \1737 , \1742 );
nor \U$1182 ( \1854 , \1853 , \1743 );
xor \U$1183 ( \1855 , \1852 , \1854 );
xor \U$1184 ( \1856 , \1844 , \1846 );
xor \U$1185 ( \1857 , \1856 , \1849 );
xor \U$1186 ( \1858 , \1836 , \1837 );
not \U$1187 ( \1859 , \1807 );
not \U$1188 ( \1860 , \1577 );
or \U$1189 ( \1861 , \1859 , \1860 );
or \U$1190 ( \1862 , \1577 , \1807 );
nand \U$1191 ( \1863 , \1861 , \1862 );
xor \U$1192 ( \1864 , \1805 , \1808 );
nor \U$1193 ( \1865 , \1863 , \1864 );
not \U$1194 ( \1866 , \1865 );
not \U$1195 ( \1867 , \1810 );
nor \U$1196 ( \1868 , \1866 , \1867 );
not \U$1197 ( \1869 , \1868 );
or \U$1198 ( \1870 , \1869 , \1295 );
or \U$1199 ( \1871 , \1866 , \1295 );
nand \U$1200 ( \1872 , \1871 , \1867 );
nand \U$1201 ( \1873 , \1870 , \1872 );
or \U$1202 ( \1874 , \1654 , \1349 );
or \U$1203 ( \1875 , \1254 , \1795 );
or \U$1204 ( \1876 , \1651 , \1349 );
or \U$1205 ( \1877 , \1579 , \1253_nG17dd );
nand \U$1206 ( \1878 , \1877 , \1799 );
nand \U$1207 ( \1879 , \1876 , \1878 );
nand \U$1208 ( \1880 , \1874 , \1875 , \1879 );
and \U$1209 ( \1881 , \1873 , \1880 );
not \U$1210 ( \1882 , \1881 );
and \U$1211 ( \1883 , \1631_nG12c9 , \1363 );
and \U$1212 ( \1884 , \1400 , \1559_nG13c8 );
nand \U$1213 ( \1885 , \1631_nG12c9 , \1360 );
or \U$1214 ( \1886 , \1320 , \1559_nG13c8 );
nand \U$1215 ( \1887 , \1886 , \1404 );
and \U$1216 ( \1888 , \1885 , \1887 );
nor \U$1217 ( \1889 , \1883 , \1884 , \1888 );
nand \U$1218 ( \1890 , \1435_nG15b1 , \1523 );
or \U$1219 ( \1891 , \1449 , \1502_nG14c8 );
nand \U$1220 ( \1892 , \1891 , \1529 );
and \U$1221 ( \1893 , \1890 , \1892 );
and \U$1222 ( \1894 , \1525 , \1502_nG14c8 );
and \U$1223 ( \1895 , \1435_nG15b1 , \1594 );
nor \U$1224 ( \1896 , \1893 , \1894 , \1895 );
xor \U$1225 ( \1897 , \1889 , \1896 );
and \U$1226 ( \1898 , \1710_nG11c1 , \1306 );
or \U$1227 ( \1899 , \1266 , \1787_nG10e2 );
nand \U$1228 ( \1900 , \1899 , \1303 );
nand \U$1229 ( \1901 , \1710_nG11c1 , \1299 );
and \U$1230 ( \1902 , \1900 , \1901 );
and \U$1231 ( \1903 , \1787_nG10e2 , \1440 );
nor \U$1232 ( \1904 , \1898 , \1902 , \1903 );
and \U$1233 ( \1905 , \1897 , \1904 );
and \U$1234 ( \1906 , \1889 , \1896 );
or \U$1235 ( \1907 , \1905 , \1906 );
nor \U$1236 ( \1908 , \1882 , \1907 );
and \U$1237 ( \1909 , \1802 , \1810 );
not \U$1238 ( \1910 , \1802 );
and \U$1239 ( \1911 , \1910 , \1867 );
nor \U$1240 ( \1912 , \1909 , \1911 );
not \U$1241 ( \1913 , \1912 );
not \U$1242 ( \1914 , \1821 );
or \U$1243 ( \1915 , \1913 , \1914 );
or \U$1244 ( \1916 , \1821 , \1912 );
nand \U$1245 ( \1917 , \1915 , \1916 );
not \U$1246 ( \1918 , \1788 );
nor \U$1247 ( \1919 , \1759 , \1791 );
not \U$1248 ( \1920 , \1919 );
or \U$1249 ( \1921 , \1918 , \1920 );
or \U$1250 ( \1922 , \1919 , \1788 );
nand \U$1251 ( \1923 , \1921 , \1922 );
and \U$1252 ( \1924 , \1917 , \1923 );
and \U$1253 ( \1925 , \1908 , \1924 );
xor \U$1254 ( \1926 , \1858 , \1925 );
xnor \U$1255 ( \1927 , \1823 , \1792 );
not \U$1256 ( \1928 , \1833 );
not \U$1257 ( \1929 , \1825 );
and \U$1258 ( \1930 , \1928 , \1929 );
and \U$1259 ( \1931 , \1833 , \1825 );
nor \U$1260 ( \1932 , \1930 , \1931 );
nand \U$1261 ( \1933 , \1927 , \1932 );
and \U$1262 ( \1934 , \1926 , \1933 );
and \U$1263 ( \1935 , \1858 , \1925 );
or \U$1264 ( \1936 , \1934 , \1935 );
xor \U$1265 ( \1937 , \1643 , \1715 );
xor \U$1266 ( \1938 , \1936 , \1937 );
xor \U$1267 ( \1939 , \1835 , \1838 );
xor \U$1268 ( \1940 , \1939 , \1841 );
and \U$1269 ( \1941 , \1938 , \1940 );
and \U$1270 ( \1942 , \1936 , \1937 );
or \U$1271 ( \1943 , \1941 , \1942 );
xor \U$1272 ( \1944 , \1857 , \1943 );
xor \U$1273 ( \1945 , \1824 , \1834 );
xor \U$1274 ( \1946 , \1858 , \1925 );
xor \U$1275 ( \1947 , \1946 , \1933 );
and \U$1276 ( \1948 , \1945 , \1947 );
xor \U$1277 ( \1949 , \1917 , \1923 );
not \U$1278 ( \1950 , \1949 );
not \U$1279 ( \1951 , \1907 );
not \U$1280 ( \1952 , \1881 );
and \U$1281 ( \1953 , \1951 , \1952 );
and \U$1282 ( \1954 , \1907 , \1881 );
nor \U$1283 ( \1955 , \1953 , \1954 );
nor \U$1284 ( \1956 , \1950 , \1955 );
xor \U$1285 ( \1957 , \1873 , \1880 );
xor \U$1286 ( \1958 , \1889 , \1896 );
xor \U$1287 ( \1959 , \1958 , \1904 );
not \U$1288 ( \1960 , \1959 );
and \U$1289 ( \1961 , \1957 , \1960 );
xor \U$1290 ( \1962 , RIaa977e8_4, \1148_nG949 );
xor \U$1291 ( \1963 , \1962 , \1184 );
not \U$1292 ( \1964 , \1963 );
xor \U$1293 ( \1965 , \1087 , \1117_nG9bd );
xor \U$1294 ( \1966 , \1965 , \1187 );
not \U$1295 ( \1967 , \1966 );
and \U$1296 ( \1968 , \1964 , \1967 );
or \U$1297 ( \1969 , \1804 , \1968 );
not \U$1298 ( \1970 , \1969 );
nand \U$1299 ( \1971 , \1253_nG17dd , \1865 );
or \U$1300 ( \1972 , \1810 , \1293_nG18eb );
or \U$1301 ( \1973 , \1810 , \1864 );
nand \U$1302 ( \1974 , \1972 , \1973 );
and \U$1303 ( \1975 , \1971 , \1974 );
and \U$1304 ( \1976 , \1810 , \1864 );
and \U$1305 ( \1977 , \1976 , \1293_nG18eb );
and \U$1306 ( \1978 , \1253_nG17dd , \1868 );
nor \U$1307 ( \1979 , \1975 , \1977 , \1978 );
and \U$1308 ( \1980 , \1435_nG15b1 , \1653 );
or \U$1309 ( \1981 , \1579 , \1348_nG16d6 );
nand \U$1310 ( \1982 , \1981 , \1799 );
nand \U$1311 ( \1983 , \1435_nG15b1 , \1650 );
and \U$1312 ( \1984 , \1982 , \1983 );
and \U$1313 ( \1985 , \1348_nG16d6 , \1794 );
nor \U$1314 ( \1986 , \1980 , \1984 , \1985 );
nand \U$1315 ( \1987 , \1979 , \1986 );
not \U$1316 ( \1988 , \1987 );
or \U$1317 ( \1989 , \1970 , \1988 );
or \U$1318 ( \1990 , \1986 , \1979 );
nand \U$1319 ( \1991 , \1989 , \1990 );
and \U$1320 ( \1992 , \1710_nG11c1 , \1363 );
and \U$1321 ( \1993 , \1400 , \1631_nG12c9 );
nand \U$1322 ( \1994 , \1710_nG11c1 , \1360 );
or \U$1323 ( \1995 , \1320 , \1631_nG12c9 );
nand \U$1324 ( \1996 , \1995 , \1404 );
and \U$1325 ( \1997 , \1994 , \1996 );
nor \U$1326 ( \1998 , \1992 , \1993 , \1997 );
nand \U$1327 ( \1999 , \1502_nG14c8 , \1523 );
or \U$1328 ( \2000 , \1449 , \1559_nG13c8 );
nand \U$1329 ( \2001 , \2000 , \1529 );
and \U$1330 ( \2002 , \1999 , \2001 );
and \U$1331 ( \2003 , \1525 , \1559_nG13c8 );
and \U$1332 ( \2004 , \1502_nG14c8 , \1594 );
nor \U$1333 ( \2005 , \2002 , \2003 , \2004 );
xor \U$1334 ( \2006 , \1998 , \2005 );
and \U$1335 ( \2007 , \1787_nG10e2 , \1306 );
and \U$1336 ( \2008 , RIaaa3ea8_428, \723 );
and \U$1337 ( \2009 , RIaaa3a70_419, \682 );
and \U$1338 ( \2010 , \742 , RIaaa4178_434);
and \U$1339 ( \2011 , RIaaa3d40_425, \712 );
nor \U$1340 ( \2012 , \2010 , \2011 );
and \U$1341 ( \2013 , \696 , RIaaa4010_431);
and \U$1342 ( \2014 , RIaaa3bd8_422, \699 );
nor \U$1343 ( \2015 , \2013 , \2014 );
and \U$1344 ( \2016 , \1241 , RIaaa4100_433);
and \U$1345 ( \2017 , RIaaa3cc8_424, \735 );
nor \U$1346 ( \2018 , \2016 , \2017 );
and \U$1347 ( \2019 , \728 , RIaaa39f8_418);
and \U$1348 ( \2020 , RIaaa3b60_421, \690 );
nor \U$1349 ( \2021 , \2019 , \2020 );
nand \U$1350 ( \2022 , \2012 , \2015 , \2018 , \2021 );
nor \U$1351 ( \2023 , \2008 , \2009 , \2022 );
and \U$1352 ( \2024 , \702 , RIaaa3f98_430);
and \U$1353 ( \2025 , RIaaa3f20_429, \721 );
nor \U$1354 ( \2026 , \2024 , \2025 );
and \U$1355 ( \2027 , \738 , RIaaa4088_432);
and \U$1356 ( \2028 , RIaaa3ae8_420, \730 );
nor \U$1357 ( \2029 , \2027 , \2028 );
and \U$1358 ( \2030 , \733 , RIaaa3e30_427);
and \U$1359 ( \2031 , RIaaa3c50_423, \686 );
nor \U$1360 ( \2032 , \2030 , \2031 );
nand \U$1361 ( \2033 , \2023 , \2026 , \2029 , \2032 );
_DC gfe1 ( \2034_nGfe1 , \2033 , \1252 );
or \U$1362 ( \2035 , \1266 , \2034_nGfe1 );
nand \U$1363 ( \2036 , \2035 , \1303 );
nand \U$1364 ( \2037 , \1787_nG10e2 , \1299 );
and \U$1365 ( \2038 , \2036 , \2037 );
and \U$1366 ( \2039 , \2034_nGfe1 , \1440 );
nor \U$1367 ( \2040 , \2007 , \2038 , \2039 );
and \U$1368 ( \2041 , \2006 , \2040 );
and \U$1369 ( \2042 , \1998 , \2005 );
or \U$1370 ( \2043 , \2041 , \2042 );
not \U$1371 ( \2044 , \2043 );
and \U$1372 ( \2045 , \1991 , \2044 );
and \U$1373 ( \2046 , \1961 , \2045 );
xor \U$1374 ( \2047 , \1956 , \2046 );
or \U$1375 ( \2048 , \1932 , \1927 );
nand \U$1376 ( \2049 , \2048 , \1933 );
and \U$1377 ( \2050 , \2047 , \2049 );
and \U$1378 ( \2051 , \1956 , \2046 );
or \U$1379 ( \2052 , \2050 , \2051 );
xor \U$1380 ( \2053 , \1858 , \1925 );
xor \U$1381 ( \2054 , \2053 , \1933 );
and \U$1382 ( \2055 , \2052 , \2054 );
and \U$1383 ( \2056 , \1945 , \2052 );
or \U$1384 ( \2057 , \1948 , \2055 , \2056 );
xor \U$1385 ( \2058 , \1936 , \1937 );
xor \U$1386 ( \2059 , \2058 , \1940 );
xor \U$1387 ( \2060 , \2057 , \2059 );
xor \U$1388 ( \2061 , \1908 , \1924 );
xor \U$1389 ( \2062 , \1956 , \2046 );
xor \U$1390 ( \2063 , \2062 , \2049 );
nand \U$1391 ( \2064 , \2061 , \2063 );
not \U$1392 ( \2065 , \1949 );
not \U$1393 ( \2066 , \1955 );
and \U$1394 ( \2067 , \2065 , \2066 );
and \U$1395 ( \2068 , \1949 , \1955 );
nor \U$1396 ( \2069 , \2067 , \2068 );
nand \U$1397 ( \2070 , \1559_nG13c8 , \1523 );
or \U$1398 ( \2071 , \1449 , \1631_nG12c9 );
nand \U$1399 ( \2072 , \2071 , \1529 );
and \U$1400 ( \2073 , \2070 , \2072 );
and \U$1401 ( \2074 , \1525 , \1631_nG12c9 );
and \U$1402 ( \2075 , \1559_nG13c8 , \1594 );
nor \U$1403 ( \2076 , \2073 , \2074 , \2075 );
and \U$1404 ( \2077 , \1502_nG14c8 , \1653 );
or \U$1405 ( \2078 , \1579 , \1435_nG15b1 );
nand \U$1406 ( \2079 , \2078 , \1799 );
nand \U$1407 ( \2080 , \1502_nG14c8 , \1650 );
and \U$1408 ( \2081 , \2079 , \2080 );
and \U$1409 ( \2082 , \1435_nG15b1 , \1794 );
nor \U$1410 ( \2083 , \2077 , \2081 , \2082 );
xor \U$1411 ( \2084 , \2076 , \2083 );
and \U$1412 ( \2085 , \1787_nG10e2 , \1363 );
and \U$1413 ( \2086 , \1400 , \1710_nG11c1 );
nand \U$1414 ( \2087 , \1787_nG10e2 , \1360 );
or \U$1415 ( \2088 , \1320 , \1710_nG11c1 );
nand \U$1416 ( \2089 , \2088 , \1404 );
and \U$1417 ( \2090 , \2087 , \2089 );
nor \U$1418 ( \2091 , \2085 , \2086 , \2090 );
and \U$1419 ( \2092 , \2084 , \2091 );
and \U$1420 ( \2093 , \2076 , \2083 );
or \U$1421 ( \2094 , \2092 , \2093 );
not \U$1422 ( \2095 , \2094 );
or \U$1423 ( \2096 , \1804 , \1966 );
nand \U$1424 ( \2097 , \1966 , \1804 );
nand \U$1425 ( \2098 , \2096 , \2097 );
xor \U$1426 ( \2099 , \1964 , \1967 );
nor \U$1427 ( \2100 , \2098 , \2099 );
not \U$1428 ( \2101 , \2100 );
not \U$1429 ( \2102 , \1969 );
nor \U$1430 ( \2103 , \2101 , \2102 );
not \U$1431 ( \2104 , \2103 );
or \U$1432 ( \2105 , \2104 , \1295 );
or \U$1433 ( \2106 , \2101 , \1295 );
nand \U$1434 ( \2107 , \2106 , \2102 );
nand \U$1435 ( \2108 , \2105 , \2107 );
not \U$1436 ( \2109 , \2108 );
nand \U$1437 ( \2110 , \1348_nG16d6 , \1865 );
or \U$1438 ( \2111 , \1810 , \1253_nG17dd );
nand \U$1439 ( \2112 , \2111 , \1973 );
and \U$1440 ( \2113 , \2110 , \2112 );
and \U$1441 ( \2114 , \1976 , \1253_nG17dd );
and \U$1442 ( \2115 , \1348_nG16d6 , \1868 );
nor \U$1443 ( \2116 , \2113 , \2114 , \2115 );
nor \U$1444 ( \2117 , \2109 , \2116 );
nand \U$1445 ( \2118 , \2095 , \2117 );
not \U$1446 ( \2119 , \2118 );
xor \U$1447 ( \2120 , \1998 , \2005 );
xor \U$1448 ( \2121 , \2120 , \2040 );
nand \U$1449 ( \2122 , \1987 , \1990 );
not \U$1450 ( \2123 , \2122 );
not \U$1451 ( \2124 , \1969 );
and \U$1452 ( \2125 , \2123 , \2124 );
and \U$1453 ( \2126 , \2122 , \1969 );
nor \U$1454 ( \2127 , \2125 , \2126 );
nor \U$1455 ( \2128 , \2121 , \2127 );
not \U$1456 ( \2129 , \2128 );
and \U$1457 ( \2130 , RIaaa32f0_403, \723 );
and \U$1458 ( \2131 , RIaaa3818_414, \728 );
and \U$1459 ( \2132 , \742 , RIaaa35c0_409);
and \U$1460 ( \2133 , RIaaa3728_412, \730 );
nor \U$1461 ( \2134 , \2132 , \2133 );
and \U$1462 ( \2135 , \1241 , RIaaa3548_408);
and \U$1463 ( \2136 , RIaaa3980_417, \712 );
nor \U$1464 ( \2137 , \2135 , \2136 );
and \U$1465 ( \2138 , \733 , RIaaa3278_402);
and \U$1466 ( \2139 , RIaaa3908_416, \735 );
nor \U$1467 ( \2140 , \2138 , \2139 );
and \U$1468 ( \2141 , \686 , RIaaa36b0_411);
and \U$1469 ( \2142 , RIaaa37a0_413, \690 );
nor \U$1470 ( \2143 , \2141 , \2142 );
nand \U$1471 ( \2144 , \2134 , \2137 , \2140 , \2143 );
nor \U$1472 ( \2145 , \2130 , \2131 , \2144 );
and \U$1473 ( \2146 , \696 , RIaaa3458_406);
and \U$1474 ( \2147 , RIaaa3638_410, \699 );
nor \U$1475 ( \2148 , \2146 , \2147 );
and \U$1476 ( \2149 , \738 , RIaaa34d0_407);
and \U$1477 ( \2150 , RIaaa33e0_405, \702 );
nor \U$1478 ( \2151 , \2149 , \2150 );
and \U$1479 ( \2152 , \721 , RIaaa3368_404);
and \U$1480 ( \2153 , RIaaa3890_415, \682 );
nor \U$1481 ( \2154 , \2152 , \2153 );
nand \U$1482 ( \2155 , \2145 , \2148 , \2151 , \2154 );
_DC gf08 ( \2156_nGf08 , \2155 , \1252 );
nand \U$1483 ( \2157 , \2156_nGf08 , \1223 );
nand \U$1484 ( \2158 , \2129 , \2157 );
nand \U$1485 ( \2159 , \2119 , \2158 );
xor \U$1486 ( \2160 , \2069 , \2159 );
xor \U$1487 ( \2161 , \1957 , \1960 );
nand \U$1488 ( \2162 , \2034_nGfe1 , \1223 );
and \U$1489 ( \2163 , \2161 , \2162 );
xor \U$1490 ( \2164 , \1991 , \2044 );
nor \U$1491 ( \2165 , \2163 , \2164 );
and \U$1492 ( \2166 , \2160 , \2165 );
and \U$1493 ( \2167 , \2069 , \2159 );
or \U$1494 ( \2168 , \2166 , \2167 );
and \U$1495 ( \2169 , \2064 , \2168 );
nor \U$1496 ( \2170 , \2063 , \2061 );
nor \U$1497 ( \2171 , \2169 , \2170 );
xor \U$1498 ( \2172 , \1858 , \1925 );
xor \U$1499 ( \2173 , \2172 , \1933 );
xor \U$1500 ( \2174 , \1945 , \2052 );
xor \U$1501 ( \2175 , \2173 , \2174 );
xor \U$1502 ( \2176 , \2171 , \2175 );
not \U$1503 ( \2177 , \2168 );
not \U$1504 ( \2178 , \2170 );
nand \U$1505 ( \2179 , \2178 , \2064 );
not \U$1506 ( \2180 , \2179 );
or \U$1507 ( \2181 , \2177 , \2180 );
or \U$1508 ( \2182 , \2179 , \2168 );
nand \U$1509 ( \2183 , \2181 , \2182 );
xor \U$1510 ( \2184 , \2069 , \2159 );
xor \U$1511 ( \2185 , \2184 , \2165 );
not \U$1512 ( \2186 , \1961 );
not \U$1513 ( \2187 , \2162 );
nor \U$1514 ( \2188 , \2187 , \2045 );
not \U$1515 ( \2189 , \2188 );
and \U$1516 ( \2190 , \2186 , \2189 );
and \U$1517 ( \2191 , \1961 , \2188 );
nor \U$1518 ( \2192 , \2190 , \2191 );
xor \U$1519 ( \2193 , \2185 , \2192 );
and \U$1520 ( \2194 , \2121 , \2127 );
nor \U$1521 ( \2195 , \2194 , \2128 );
not \U$1522 ( \2196 , \2195 );
not \U$1523 ( \2197 , \2157 );
and \U$1524 ( \2198 , \2196 , \2197 );
and \U$1525 ( \2199 , \2195 , \2157 );
nor \U$1526 ( \2200 , \2198 , \2199 );
not \U$1527 ( \2201 , \2200 );
or \U$1528 ( \2202 , \2094 , \2117 );
and \U$1529 ( \2203 , RIaaa42e0_437, \1241 );
and \U$1530 ( \2204 , RIaaa4448_440, \721 );
and \U$1531 ( \2205 , \742 , RIaaa4358_438);
and \U$1532 ( \2206 , RIaaa4790_447, \712 );
nor \U$1533 ( \2207 , \2205 , \2206 );
and \U$1534 ( \2208 , \738 , RIaaa4268_436);
and \U$1535 ( \2209 , RIaaa4718_446, \735 );
nor \U$1536 ( \2210 , \2208 , \2209 );
and \U$1537 ( \2211 , \733 , RIaaa43d0_439);
and \U$1538 ( \2212 , RIaaa4808_448, \730 );
nor \U$1539 ( \2213 , \2211 , \2212 );
and \U$1540 ( \2214 , \686 , RIaaa4970_451);
and \U$1541 ( \2215 , RIaaa4880_449, \690 );
nor \U$1542 ( \2216 , \2214 , \2215 );
nand \U$1543 ( \2217 , \2207 , \2210 , \2213 , \2216 );
nor \U$1544 ( \2218 , \2203 , \2204 , \2217 );
and \U$1545 ( \2219 , \696 , RIaaa45b0_443);
and \U$1546 ( \2220 , RIaaa46a0_445, \682 );
nor \U$1547 ( \2221 , \2219 , \2220 );
and \U$1548 ( \2222 , \702 , RIaaa4538_442);
and \U$1549 ( \2223 , RIaaa44c0_441, \723 );
nor \U$1550 ( \2224 , \2222 , \2223 );
and \U$1551 ( \2225 , \699 , RIaaa48f8_450);
and \U$1552 ( \2226 , RIaaa4628_444, \728 );
nor \U$1553 ( \2227 , \2225 , \2226 );
nand \U$1554 ( \2228 , \2218 , \2221 , \2224 , \2227 );
_DC ge35 ( \2229_nGe35 , \2228 , \1252 );
nand \U$1555 ( \2230 , \2229_nGe35 , \1223 );
and \U$1556 ( \2231 , \2034_nGfe1 , \1306 );
or \U$1557 ( \2232 , \1266 , \2156_nGf08 );
nand \U$1558 ( \2233 , \2232 , \1303 );
nand \U$1559 ( \2234 , \2034_nGfe1 , \1299 );
and \U$1560 ( \2235 , \2233 , \2234 );
and \U$1561 ( \2236 , \2156_nGf08 , \1440 );
nor \U$1562 ( \2237 , \2231 , \2235 , \2236 );
or \U$1563 ( \2238 , \2230 , \2237 );
nand \U$1564 ( \2239 , \2117 , \2094 );
nand \U$1565 ( \2240 , \2202 , \2238 , \2239 );
nand \U$1566 ( \2241 , \2201 , \2240 );
not \U$1567 ( \2242 , \2116 );
not \U$1568 ( \2243 , \2108 );
and \U$1569 ( \2244 , \2242 , \2243 );
and \U$1570 ( \2245 , \2116 , \2108 );
nor \U$1571 ( \2246 , \2244 , \2245 );
xor \U$1572 ( \2247 , \2076 , \2083 );
xor \U$1573 ( \2248 , \2247 , \2091 );
and \U$1574 ( \2249 , \2246 , \2248 );
xnor \U$1575 ( \2250 , \2230 , \2237 );
xor \U$1576 ( \2251 , \2076 , \2083 );
xor \U$1577 ( \2252 , \2251 , \2091 );
and \U$1578 ( \2253 , \2250 , \2252 );
and \U$1579 ( \2254 , \2246 , \2250 );
or \U$1580 ( \2255 , \2249 , \2253 , \2254 );
not \U$1581 ( \2256 , \2255 );
not \U$1582 ( \2257 , \2034_nGfe1 );
or \U$1583 ( \2258 , \1364 , \2257 );
and \U$1584 ( \2259 , \1400 , \1787_nG10e2 );
nand \U$1585 ( \2260 , \2034_nGfe1 , \1360 );
or \U$1586 ( \2261 , \1320 , \1787_nG10e2 );
nand \U$1587 ( \2262 , \2261 , \1404 );
and \U$1588 ( \2263 , \2260 , \2262 );
nor \U$1589 ( \2264 , \2259 , \2263 );
nand \U$1590 ( \2265 , \2258 , \2264 );
and \U$1591 ( \2266 , \1559_nG13c8 , \1653 );
or \U$1592 ( \2267 , \1579 , \1502_nG14c8 );
nand \U$1593 ( \2268 , \2267 , \1799 );
nand \U$1594 ( \2269 , \1559_nG13c8 , \1650 );
and \U$1595 ( \2270 , \2268 , \2269 );
and \U$1596 ( \2271 , \1502_nG14c8 , \1794 );
nor \U$1597 ( \2272 , \2266 , \2270 , \2271 );
nand \U$1598 ( \2273 , \1631_nG12c9 , \1523 );
or \U$1599 ( \2274 , \1449 , \1710_nG11c1 );
nand \U$1600 ( \2275 , \2274 , \1529 );
and \U$1601 ( \2276 , \2273 , \2275 );
and \U$1602 ( \2277 , \1525 , \1710_nG11c1 );
and \U$1603 ( \2278 , \1631_nG12c9 , \1594 );
nor \U$1604 ( \2279 , \2276 , \2277 , \2278 );
nand \U$1605 ( \2280 , \2272 , \2279 );
and \U$1606 ( \2281 , \2265 , \2280 );
nor \U$1607 ( \2282 , \2279 , \2272 );
nor \U$1608 ( \2283 , \2281 , \2282 );
nand \U$1609 ( \2284 , \1253_nG17dd , \2100 );
or \U$1610 ( \2285 , \1969 , \1293_nG18eb );
or \U$1611 ( \2286 , \1969 , \2099 );
nand \U$1612 ( \2287 , \2285 , \2286 );
and \U$1613 ( \2288 , \2284 , \2287 );
and \U$1614 ( \2289 , \1969 , \2099 );
and \U$1615 ( \2290 , \2289 , \1293_nG18eb );
and \U$1616 ( \2291 , \1253_nG17dd , \2103 );
nor \U$1617 ( \2292 , \2288 , \2290 , \2291 );
xor \U$1618 ( \2293 , \2292 , \1964 );
nand \U$1619 ( \2294 , \1435_nG15b1 , \1865 );
or \U$1620 ( \2295 , \1810 , \1348_nG16d6 );
nand \U$1621 ( \2296 , \2295 , \1973 );
and \U$1622 ( \2297 , \2294 , \2296 );
and \U$1623 ( \2298 , \1976 , \1348_nG16d6 );
and \U$1624 ( \2299 , \1435_nG15b1 , \1868 );
nor \U$1625 ( \2300 , \2297 , \2298 , \2299 );
and \U$1626 ( \2301 , \2293 , \2300 );
and \U$1627 ( \2302 , \2292 , \1964 );
or \U$1628 ( \2303 , \2301 , \2302 );
nor \U$1629 ( \2304 , \2283 , \2303 );
nand \U$1630 ( \2305 , \2256 , \2304 );
xor \U$1631 ( \2306 , \2241 , \2305 );
not \U$1632 ( \2307 , \2164 );
not \U$1633 ( \2308 , \2161 );
or \U$1634 ( \2309 , \2307 , \2308 );
or \U$1635 ( \2310 , \2161 , \2164 );
nand \U$1636 ( \2311 , \2309 , \2310 );
not \U$1637 ( \2312 , \2311 );
not \U$1638 ( \2313 , \2162 );
and \U$1639 ( \2314 , \2312 , \2313 );
and \U$1640 ( \2315 , \2311 , \2162 );
nor \U$1641 ( \2316 , \2314 , \2315 );
and \U$1642 ( \2317 , \2306 , \2316 );
and \U$1643 ( \2318 , \2241 , \2305 );
or \U$1644 ( \2319 , \2317 , \2318 );
and \U$1645 ( \2320 , \2193 , \2319 );
and \U$1646 ( \2321 , \2185 , \2192 );
or \U$1647 ( \2322 , \2320 , \2321 );
xor \U$1648 ( \2323 , \2183 , \2322 );
not \U$1649 ( \2324 , \2200 );
not \U$1650 ( \2325 , \2240 );
and \U$1651 ( \2326 , \2324 , \2325 );
and \U$1652 ( \2327 , \2200 , \2240 );
nor \U$1653 ( \2328 , \2326 , \2327 );
not \U$1654 ( \2329 , \2255 );
not \U$1655 ( \2330 , \2304 );
and \U$1656 ( \2331 , \2329 , \2330 );
and \U$1657 ( \2332 , \2255 , \2304 );
nor \U$1658 ( \2333 , \2331 , \2332 );
xor \U$1659 ( \2334 , \2328 , \2333 );
and \U$1660 ( \2335 , \1631_nG12c9 , \1653 );
or \U$1661 ( \2336 , \1579 , \1559_nG13c8 );
nand \U$1662 ( \2337 , \2336 , \1799 );
nand \U$1663 ( \2338 , \1631_nG12c9 , \1650 );
and \U$1664 ( \2339 , \2337 , \2338 );
and \U$1665 ( \2340 , \1559_nG13c8 , \1794 );
nor \U$1666 ( \2341 , \2335 , \2339 , \2340 );
nand \U$1667 ( \2342 , \1502_nG14c8 , \1865 );
or \U$1668 ( \2343 , \1810 , \1435_nG15b1 );
nand \U$1669 ( \2344 , \2343 , \1973 );
and \U$1670 ( \2345 , \2342 , \2344 );
and \U$1671 ( \2346 , \1976 , \1435_nG15b1 );
and \U$1672 ( \2347 , \1502_nG14c8 , \1868 );
nor \U$1673 ( \2348 , \2345 , \2346 , \2347 );
xor \U$1674 ( \2349 , \2341 , \2348 );
nand \U$1675 ( \2350 , \1710_nG11c1 , \1523 );
or \U$1676 ( \2351 , \1449 , \1787_nG10e2 );
nand \U$1677 ( \2352 , \2351 , \1529 );
and \U$1678 ( \2353 , \2350 , \2352 );
and \U$1679 ( \2354 , \1525 , \1787_nG10e2 );
and \U$1680 ( \2355 , \1710_nG11c1 , \1594 );
nor \U$1681 ( \2356 , \2353 , \2354 , \2355 );
and \U$1682 ( \2357 , \2349 , \2356 );
and \U$1683 ( \2358 , \2341 , \2348 );
or \U$1684 ( \2359 , \2357 , \2358 );
nand \U$1685 ( \2360 , \1348_nG16d6 , \2100 );
or \U$1686 ( \2361 , \1969 , \1253_nG17dd );
nand \U$1687 ( \2362 , \2361 , \2286 );
and \U$1688 ( \2363 , \2360 , \2362 );
and \U$1689 ( \2364 , \2289 , \1253_nG17dd );
and \U$1690 ( \2365 , \1348_nG16d6 , \2103 );
nor \U$1691 ( \2366 , \2363 , \2364 , \2365 );
not \U$1692 ( \2367 , \2366 );
or \U$1693 ( \2368 , \1963 , \1293_nG18eb );
or \U$1694 ( \2369 , \1182 , \1181_nG947 );
nand \U$1695 ( \2370 , \2369 , \1183 );
nor \U$1696 ( \2371 , \1963 , \2370 );
not \U$1697 ( \2372 , \2371 );
nand \U$1698 ( \2373 , \1964 , \2372 );
nand \U$1699 ( \2374 , \2368 , \2373 );
nand \U$1700 ( \2375 , \2367 , \2374 );
xor \U$1701 ( \2376 , \2359 , \2375 );
and \U$1702 ( \2377 , \2229_nGe35 , \1306 );
and \U$1703 ( \2378 , RIaaa62c0_505, \1241 );
and \U$1704 ( \2379 , RIaaa6428_508, \721 );
and \U$1705 ( \2380 , \742 , RIaaa6338_506);
and \U$1706 ( \2381 , RIaaa6680_513, \730 );
nor \U$1707 ( \2382 , \2380 , \2381 );
and \U$1708 ( \2383 , \723 , RIaaa64a0_509);
and \U$1709 ( \2384 , RIaaa63b0_507, \733 );
nor \U$1710 ( \2385 , \2383 , \2384 );
and \U$1711 ( \2386 , \738 , RIaaa6248_504);
and \U$1712 ( \2387 , RIaaa68d8_518, \735 );
nor \U$1713 ( \2388 , \2386 , \2387 );
and \U$1714 ( \2389 , \682 , RIaaa67e8_516);
and \U$1715 ( \2390 , RIaaa6860_517, \728 );
nor \U$1716 ( \2391 , \2389 , \2390 );
nand \U$1717 ( \2392 , \2382 , \2385 , \2388 , \2391 );
nor \U$1718 ( \2393 , \2378 , \2379 , \2392 );
and \U$1719 ( \2394 , \696 , RIaaa6518_510);
and \U$1720 ( \2395 , RIaaa6608_512, \690 );
nor \U$1721 ( \2396 , \2394 , \2395 );
and \U$1722 ( \2397 , \702 , RIaaa6590_511);
and \U$1723 ( \2398 , RIaaa66f8_514, \699 );
nor \U$1724 ( \2399 , \2397 , \2398 );
and \U$1725 ( \2400 , \686 , RIaaa6770_515);
and \U$1726 ( \2401 , RIaaa6950_519, \712 );
nor \U$1727 ( \2402 , \2400 , \2401 );
nand \U$1728 ( \2403 , \2393 , \2396 , \2399 , \2402 );
_DC gad6 ( \2404_nGad6 , \2403 , \1252 );
or \U$1729 ( \2405 , \1266 , \2404_nGad6 );
nand \U$1730 ( \2406 , \2405 , \1303 );
nand \U$1731 ( \2407 , \2229_nGe35 , \1299 );
and \U$1732 ( \2408 , \2406 , \2407 );
and \U$1733 ( \2409 , \2404_nGad6 , \1440 );
nor \U$1734 ( \2410 , \2377 , \2408 , \2409 );
and \U$1735 ( \2411 , \2156_nGf08 , \1363 );
and \U$1736 ( \2412 , \1400 , \2034_nGfe1 );
nand \U$1737 ( \2413 , \2156_nGf08 , \1360 );
or \U$1738 ( \2414 , \1320 , \2034_nGfe1 );
nand \U$1739 ( \2415 , \2414 , \1404 );
and \U$1740 ( \2416 , \2413 , \2415 );
nor \U$1741 ( \2417 , \2411 , \2412 , \2416 );
and \U$1742 ( \2418 , \2410 , \2417 );
not \U$1743 ( \2419 , \2418 );
and \U$1744 ( \2420 , RIaaa5708_480, \730 );
and \U$1745 ( \2421 , RIaaa58e8_484, \712 );
and \U$1746 ( \2422 , \682 , RIaaa5690_479);
and \U$1747 ( \2423 , RIaaa5780_481, \690 );
nor \U$1748 ( \2424 , \2422 , \2423 );
and \U$1749 ( \2425 , \702 , RIaaa53c0_473);
and \U$1750 ( \2426 , RIaaa5348_472, \721 );
nor \U$1751 ( \2427 , \2425 , \2426 );
and \U$1752 ( \2428 , \696 , RIaaa5438_474);
and \U$1753 ( \2429 , RIaaa57f8_482, \699 );
nor \U$1754 ( \2430 , \2428 , \2429 );
and \U$1755 ( \2431 , \1241 , RIaaa55a0_477);
and \U$1756 ( \2432 , RIaaa5870_483, \686 );
nor \U$1757 ( \2433 , \2431 , \2432 );
nand \U$1758 ( \2434 , \2424 , \2427 , \2430 , \2433 );
nor \U$1759 ( \2435 , \2420 , \2421 , \2434 );
and \U$1760 ( \2436 , \738 , RIaaa54b0_475);
and \U$1761 ( \2437 , RIaaa5618_478, \728 );
nor \U$1762 ( \2438 , \2436 , \2437 );
and \U$1763 ( \2439 , \733 , RIaaa5258_470);
and \U$1764 ( \2440 , RIaaa5960_485, \735 );
nor \U$1765 ( \2441 , \2439 , \2440 );
and \U$1766 ( \2442 , \723 , RIaaa52d0_471);
and \U$1767 ( \2443 , RIaaa5528_476, \742 );
nor \U$1768 ( \2444 , \2442 , \2443 );
nand \U$1769 ( \2445 , \2435 , \2438 , \2441 , \2444 );
_DC ga9e ( \2446_nGa9e , \2445 , \1252 );
nand \U$1770 ( \2447 , \2446_nGa9e , \1223 );
not \U$1771 ( \2448 , \2447 );
and \U$1772 ( \2449 , \2419 , \2448 );
nor \U$1773 ( \2450 , \2410 , \2417 );
nor \U$1774 ( \2451 , \2449 , \2450 );
and \U$1775 ( \2452 , \2376 , \2451 );
and \U$1776 ( \2453 , \2359 , \2375 );
or \U$1777 ( \2454 , \2452 , \2453 );
nand \U$1778 ( \2455 , \2404_nGad6 , \1223 );
and \U$1779 ( \2456 , \2156_nGf08 , \1306 );
or \U$1780 ( \2457 , \1266 , \2229_nGe35 );
nand \U$1781 ( \2458 , \2457 , \1303 );
nand \U$1782 ( \2459 , \2156_nGf08 , \1299 );
and \U$1783 ( \2460 , \2458 , \2459 );
and \U$1784 ( \2461 , \2229_nGe35 , \1440 );
nor \U$1785 ( \2462 , \2456 , \2460 , \2461 );
xnor \U$1786 ( \2463 , \2455 , \2462 );
xor \U$1787 ( \2464 , \2454 , \2463 );
xor \U$1788 ( \2465 , \2076 , \2083 );
xor \U$1789 ( \2466 , \2465 , \2091 );
xor \U$1790 ( \2467 , \2246 , \2250 );
xor \U$1791 ( \2468 , \2466 , \2467 );
and \U$1792 ( \2469 , \2464 , \2468 );
and \U$1793 ( \2470 , \2454 , \2463 );
or \U$1794 ( \2471 , \2469 , \2470 );
and \U$1795 ( \2472 , \2334 , \2471 );
and \U$1796 ( \2473 , \2328 , \2333 );
or \U$1797 ( \2474 , \2472 , \2473 );
not \U$1798 ( \2475 , \2158 );
not \U$1799 ( \2476 , \2118 );
and \U$1800 ( \2477 , \2475 , \2476 );
and \U$1801 ( \2478 , \2158 , \2118 );
nor \U$1802 ( \2479 , \2477 , \2478 );
xor \U$1803 ( \2480 , \2474 , \2479 );
xor \U$1804 ( \2481 , \2241 , \2305 );
xor \U$1805 ( \2482 , \2481 , \2316 );
and \U$1806 ( \2483 , \2480 , \2482 );
and \U$1807 ( \2484 , \2474 , \2479 );
or \U$1808 ( \2485 , \2483 , \2484 );
xor \U$1809 ( \2486 , \2185 , \2192 );
xor \U$1810 ( \2487 , \2486 , \2319 );
and \U$1811 ( \2488 , \2485 , \2487 );
xor \U$1812 ( \2489 , \2454 , \2463 );
xor \U$1813 ( \2490 , \2489 , \2468 );
not \U$1814 ( \2491 , \2490 );
or \U$1815 ( \2492 , \2462 , \2455 );
not \U$1816 ( \2493 , \2303 );
or \U$1817 ( \2494 , \2493 , \2283 );
not \U$1818 ( \2495 , \2283 );
or \U$1819 ( \2496 , \2303 , \2495 );
nand \U$1820 ( \2497 , \2492 , \2494 , \2496 );
nand \U$1821 ( \2498 , \2491 , \2497 );
not \U$1822 ( \2499 , \2463 );
xor \U$1823 ( \2500 , \2292 , \1964 );
xor \U$1824 ( \2501 , \2500 , \2300 );
xor \U$1825 ( \2502 , \2499 , \2501 );
xor \U$1826 ( \2503 , \2359 , \2375 );
xor \U$1827 ( \2504 , \2503 , \2451 );
and \U$1828 ( \2505 , \2502 , \2504 );
and \U$1829 ( \2506 , \2499 , \2501 );
or \U$1830 ( \2507 , \2505 , \2506 );
not \U$1831 ( \2508 , \2507 );
nand \U$1832 ( \2509 , \1787_nG10e2 , \1523 );
or \U$1833 ( \2510 , \1449 , \2034_nGfe1 );
nand \U$1834 ( \2511 , \2510 , \1529 );
and \U$1835 ( \2512 , \2509 , \2511 );
and \U$1836 ( \2513 , \1525 , \2034_nGfe1 );
and \U$1837 ( \2514 , \1787_nG10e2 , \1594 );
nor \U$1838 ( \2515 , \2512 , \2513 , \2514 );
and \U$1839 ( \2516 , \1710_nG11c1 , \1653 );
or \U$1840 ( \2517 , \1579 , \1631_nG12c9 );
nand \U$1841 ( \2518 , \2517 , \1799 );
nand \U$1842 ( \2519 , \1710_nG11c1 , \1650 );
and \U$1843 ( \2520 , \2518 , \2519 );
and \U$1844 ( \2521 , \1631_nG12c9 , \1794 );
nor \U$1845 ( \2522 , \2516 , \2520 , \2521 );
xor \U$1846 ( \2523 , \2515 , \2522 );
and \U$1847 ( \2524 , \2229_nGe35 , \1363 );
and \U$1848 ( \2525 , \1400 , \2156_nGf08 );
nand \U$1849 ( \2526 , \2229_nGe35 , \1360 );
or \U$1850 ( \2527 , \1320 , \2156_nGf08 );
nand \U$1851 ( \2528 , \2527 , \1404 );
and \U$1852 ( \2529 , \2526 , \2528 );
nor \U$1853 ( \2530 , \2524 , \2525 , \2529 );
and \U$1854 ( \2531 , \2523 , \2530 );
and \U$1855 ( \2532 , \2515 , \2522 );
or \U$1856 ( \2533 , \2531 , \2532 );
nand \U$1857 ( \2534 , \1435_nG15b1 , \2100 );
or \U$1858 ( \2535 , \1969 , \1348_nG16d6 );
nand \U$1859 ( \2536 , \2535 , \2286 );
and \U$1860 ( \2537 , \2534 , \2536 );
and \U$1861 ( \2538 , \2289 , \1348_nG16d6 );
and \U$1862 ( \2539 , \1435_nG15b1 , \2103 );
nor \U$1863 ( \2540 , \2537 , \2538 , \2539 );
not \U$1864 ( \2541 , \2373 );
and \U$1865 ( \2542 , \1295 , \2541 );
and \U$1866 ( \2543 , \2371 , \1254 );
nand \U$1867 ( \2544 , \2370 , \1963 );
not \U$1868 ( \2545 , \2544 );
and \U$1869 ( \2546 , \1293_nG18eb , \2545 );
nor \U$1870 ( \2547 , \2542 , \2543 , \2546 );
xor \U$1871 ( \2548 , \2540 , \2547 );
nand \U$1872 ( \2549 , \1559_nG13c8 , \1865 );
or \U$1873 ( \2550 , \1810 , \1502_nG14c8 );
nand \U$1874 ( \2551 , \2550 , \1973 );
and \U$1875 ( \2552 , \2549 , \2551 );
and \U$1876 ( \2553 , \1976 , \1502_nG14c8 );
and \U$1877 ( \2554 , \1559_nG13c8 , \1868 );
nor \U$1878 ( \2555 , \2552 , \2553 , \2554 );
and \U$1879 ( \2556 , \2548 , \2555 );
and \U$1880 ( \2557 , \2540 , \2547 );
or \U$1881 ( \2558 , \2556 , \2557 );
nor \U$1882 ( \2559 , \2533 , \2558 );
not \U$1883 ( \2560 , \2282 );
nand \U$1884 ( \2561 , \2560 , \2280 );
not \U$1885 ( \2562 , \2561 );
not \U$1886 ( \2563 , \2265 );
or \U$1887 ( \2564 , \2562 , \2563 );
or \U$1888 ( \2565 , \2265 , \2561 );
nand \U$1889 ( \2566 , \2564 , \2565 );
xor \U$1890 ( \2567 , \2559 , \2566 );
not \U$1891 ( \2568 , \2447 );
nor \U$1892 ( \2569 , \2418 , \2450 );
not \U$1893 ( \2570 , \2569 );
or \U$1894 ( \2571 , \2568 , \2570 );
or \U$1895 ( \2572 , \2569 , \2447 );
nand \U$1896 ( \2573 , \2571 , \2572 );
not \U$1897 ( \2574 , \2573 );
xor \U$1898 ( \2575 , \2341 , \2348 );
xor \U$1899 ( \2576 , \2575 , \2356 );
nor \U$1900 ( \2577 , \2574 , \2576 );
and \U$1901 ( \2578 , \2567 , \2577 );
and \U$1902 ( \2579 , \2559 , \2566 );
or \U$1903 ( \2580 , \2578 , \2579 );
nor \U$1904 ( \2581 , \2508 , \2580 );
xor \U$1905 ( \2582 , \2498 , \2581 );
xor \U$1906 ( \2583 , \2328 , \2333 );
xor \U$1907 ( \2584 , \2583 , \2471 );
and \U$1908 ( \2585 , \2582 , \2584 );
and \U$1909 ( \2586 , \2498 , \2581 );
or \U$1910 ( \2587 , \2585 , \2586 );
xor \U$1911 ( \2588 , \2474 , \2479 );
xor \U$1912 ( \2589 , \2588 , \2482 );
and \U$1913 ( \2590 , \2587 , \2589 );
not \U$1914 ( \2591 , \2490 );
not \U$1915 ( \2592 , \2497 );
and \U$1916 ( \2593 , \2591 , \2592 );
and \U$1917 ( \2594 , \2490 , \2497 );
nor \U$1918 ( \2595 , \2593 , \2594 );
not \U$1919 ( \2596 , \2366 );
not \U$1920 ( \2597 , \2374 );
and \U$1921 ( \2598 , \2596 , \2597 );
and \U$1922 ( \2599 , \2366 , \2374 );
nor \U$1923 ( \2600 , \2598 , \2599 );
and \U$1924 ( \2601 , \1787_nG10e2 , \1653 );
or \U$1925 ( \2602 , \1579 , \1710_nG11c1 );
nand \U$1926 ( \2603 , \2602 , \1799 );
nand \U$1927 ( \2604 , \1787_nG10e2 , \1650 );
and \U$1928 ( \2605 , \2603 , \2604 );
and \U$1929 ( \2606 , \1710_nG11c1 , \1794 );
nor \U$1930 ( \2607 , \2601 , \2605 , \2606 );
nand \U$1931 ( \2608 , \1631_nG12c9 , \1865 );
or \U$1932 ( \2609 , \1810 , \1559_nG13c8 );
nand \U$1933 ( \2610 , \2609 , \1973 );
and \U$1934 ( \2611 , \2608 , \2610 );
and \U$1935 ( \2612 , \1976 , \1559_nG13c8 );
and \U$1936 ( \2613 , \1631_nG12c9 , \1868 );
nor \U$1937 ( \2614 , \2611 , \2612 , \2613 );
xor \U$1938 ( \2615 , \2607 , \2614 );
nand \U$1939 ( \2616 , \2034_nGfe1 , \1523 );
or \U$1940 ( \2617 , \1449 , \2156_nGf08 );
nand \U$1941 ( \2618 , \2617 , \1529 );
and \U$1942 ( \2619 , \2616 , \2618 );
and \U$1943 ( \2620 , \1525 , \2156_nGf08 );
and \U$1944 ( \2621 , \2034_nGfe1 , \1594 );
nor \U$1945 ( \2622 , \2619 , \2620 , \2621 );
and \U$1946 ( \2623 , \2615 , \2622 );
and \U$1947 ( \2624 , \2607 , \2614 );
or \U$1948 ( \2625 , \2623 , \2624 );
and \U$1949 ( \2626 , \2446_nGa9e , \1306 );
and \U$1950 ( \2627 , RIaaa4bc8_456, \1241 );
and \U$1951 ( \2628 , RIaaa5168_468, \690 );
and \U$1952 ( \2629 , \721 , RIaaa5078_466);
and \U$1953 ( \2630 , RIaaa4c40_457, \742 );
nor \U$1954 ( \2631 , \2629 , \2630 );
and \U$1955 ( \2632 , \723 , RIaaa4f88_464);
and \U$1956 ( \2633 , RIaaa50f0_467, \730 );
nor \U$1957 ( \2634 , \2632 , \2633 );
and \U$1958 ( \2635 , \738 , RIaaa4b50_455);
and \U$1959 ( \2636 , RIaaa5000_465, \733 );
nor \U$1960 ( \2637 , \2635 , \2636 );
and \U$1961 ( \2638 , \682 , RIaaa4e20_461);
and \U$1962 ( \2639 , RIaaa4e98_462, \728 );
nor \U$1963 ( \2640 , \2638 , \2639 );
nand \U$1964 ( \2641 , \2631 , \2634 , \2637 , \2640 );
nor \U$1965 ( \2642 , \2627 , \2628 , \2641 );
and \U$1966 ( \2643 , \702 , RIaaa4da8_460);
and \U$1967 ( \2644 , RIaaa4a60_453, \686 );
nor \U$1968 ( \2645 , \2643 , \2644 );
and \U$1969 ( \2646 , \696 , RIaaa4f10_463);
and \U$1970 ( \2647 , RIaaa49e8_452, \699 );
nor \U$1971 ( \2648 , \2646 , \2647 );
and \U$1972 ( \2649 , \735 , RIaaa4d30_459);
and \U$1973 ( \2650 , RIaaa4cb8_458, \712 );
nor \U$1974 ( \2651 , \2649 , \2650 );
nand \U$1975 ( \2652 , \2642 , \2645 , \2648 , \2651 );
_DC ga66 ( \2653_nGa66 , \2652 , \1252 );
or \U$1976 ( \2654 , \1266 , \2653_nGa66 );
nand \U$1977 ( \2655 , \2654 , \1303 );
nand \U$1978 ( \2656 , \2446_nGa9e , \1299 );
and \U$1979 ( \2657 , \2655 , \2656 );
and \U$1980 ( \2658 , \2653_nGa66 , \1440 );
nor \U$1981 ( \2659 , \2626 , \2657 , \2658 );
and \U$1982 ( \2660 , \2404_nGad6 , \1363 );
and \U$1983 ( \2661 , \1400 , \2229_nGe35 );
nand \U$1984 ( \2662 , \2404_nGad6 , \1360 );
or \U$1985 ( \2663 , \1320 , \2229_nGe35 );
nand \U$1986 ( \2664 , \2663 , \1404 );
and \U$1987 ( \2665 , \2662 , \2664 );
nor \U$1988 ( \2666 , \2660 , \2661 , \2665 );
and \U$1989 ( \2667 , \2659 , \2666 );
not \U$1990 ( \2668 , \2667 );
and \U$1991 ( \2669 , RIaaa5e88_496, \1241 );
and \U$1992 ( \2670 , RIaaa5ca8_492, \699 );
and \U$1993 ( \2671 , \742 , RIaaa5f00_497);
and \U$1994 ( \2672 , RIaaa60e0_501, \730 );
nor \U$1995 ( \2673 , \2671 , \2672 );
and \U$1996 ( \2674 , \723 , RIaaa5b40_489);
and \U$1997 ( \2675 , RIaaa5bb8_490, \733 );
nor \U$1998 ( \2676 , \2674 , \2675 );
and \U$1999 ( \2677 , \738 , RIaaa5e10_495);
and \U$2000 ( \2678 , RIaaa5ff0_499, \735 );
nor \U$2001 ( \2679 , \2677 , \2678 );
and \U$2002 ( \2680 , \682 , RIaaa5a50_487);
and \U$2003 ( \2681 , RIaaa59d8_486, \728 );
nor \U$2004 ( \2682 , \2680 , \2681 );
nand \U$2005 ( \2683 , \2673 , \2676 , \2679 , \2682 );
nor \U$2006 ( \2684 , \2669 , \2670 , \2683 );
and \U$2007 ( \2685 , \702 , RIaaa6068_500);
and \U$2008 ( \2686 , RIaaa5f78_498, \712 );
nor \U$2009 ( \2687 , \2685 , \2686 );
and \U$2010 ( \2688 , \696 , RIaaa5ac8_488);
and \U$2011 ( \2689 , RIaaa6158_502, \690 );
nor \U$2012 ( \2690 , \2688 , \2689 );
and \U$2013 ( \2691 , \721 , RIaaa5c30_491);
and \U$2014 ( \2692 , RIaaa5d20_493, \686 );
nor \U$2015 ( \2693 , \2691 , \2692 );
nand \U$2016 ( \2694 , \2684 , \2687 , \2690 , \2693 );
_DC ga2d ( \2695_nGa2d , \2694 , \1252 );
nand \U$2017 ( \2696 , \2695_nGa2d , \1223 );
not \U$2018 ( \2697 , \2696 );
and \U$2019 ( \2698 , \2668 , \2697 );
nor \U$2020 ( \2699 , \2659 , \2666 );
nor \U$2021 ( \2700 , \2698 , \2699 );
nand \U$2022 ( \2701 , \2625 , \2700 );
or \U$2023 ( \2702 , \2544 , \1254 );
or \U$2024 ( \2703 , \1253_nG17dd , \2373 );
or \U$2025 ( \2704 , \1348_nG16d6 , \2372 );
nand \U$2026 ( \2705 , \2702 , \2703 , \2704 );
or \U$2027 ( \2706 , \2104 , \1503 );
or \U$2028 ( \2707 , \1969 , \1435_nG15b1 );
nand \U$2029 ( \2708 , \2707 , \2286 );
nand \U$2030 ( \2709 , \1502_nG14c8 , \2100 );
and \U$2031 ( \2710 , \2708 , \2709 );
and \U$2032 ( \2711 , \1435_nG15b1 , \2289 );
nor \U$2033 ( \2712 , \2710 , \2711 );
nand \U$2034 ( \2713 , \2706 , \2712 );
and \U$2035 ( \2714 , \2705 , \2713 );
and \U$2036 ( \2715 , \2701 , \2714 );
nor \U$2037 ( \2716 , \2700 , \2625 );
nor \U$2038 ( \2717 , \2715 , \2716 );
nand \U$2039 ( \2718 , \2600 , \2717 );
xor \U$2040 ( \2719 , \2515 , \2522 );
xor \U$2041 ( \2720 , \2719 , \2530 );
not \U$2042 ( \2721 , \2720 );
nand \U$2043 ( \2722 , \2653_nGa66 , \1223 );
and \U$2044 ( \2723 , \2404_nGad6 , \1306 );
or \U$2045 ( \2724 , \1266 , \2446_nGa9e );
nand \U$2046 ( \2725 , \2724 , \1303 );
nand \U$2047 ( \2726 , \2404_nGad6 , \1299 );
and \U$2048 ( \2727 , \2725 , \2726 );
and \U$2049 ( \2728 , \2446_nGa9e , \1440 );
nor \U$2050 ( \2729 , \2723 , \2727 , \2728 );
xor \U$2051 ( \2730 , \2722 , \2729 );
and \U$2052 ( \2731 , \2721 , \2730 );
and \U$2053 ( \2732 , \2718 , \2731 );
nor \U$2054 ( \2733 , \2717 , \2600 );
nor \U$2055 ( \2734 , \2732 , \2733 );
not \U$2056 ( \2735 , \2573 );
not \U$2057 ( \2736 , \2576 );
and \U$2058 ( \2737 , \2735 , \2736 );
and \U$2059 ( \2738 , \2573 , \2576 );
nor \U$2060 ( \2739 , \2737 , \2738 );
not \U$2061 ( \2740 , \2739 );
not \U$2062 ( \2741 , \2558 );
or \U$2063 ( \2742 , \2533 , \2741 );
not \U$2064 ( \2743 , \2533 );
or \U$2065 ( \2744 , \2558 , \2743 );
or \U$2066 ( \2745 , \2722 , \2729 );
nand \U$2067 ( \2746 , \2742 , \2744 , \2745 );
nand \U$2068 ( \2747 , \2740 , \2746 );
xor \U$2069 ( \2748 , \2734 , \2747 );
xor \U$2070 ( \2749 , \2499 , \2501 );
xor \U$2071 ( \2750 , \2749 , \2504 );
and \U$2072 ( \2751 , \2748 , \2750 );
and \U$2073 ( \2752 , \2734 , \2747 );
or \U$2074 ( \2753 , \2751 , \2752 );
nand \U$2075 ( \2754 , \2595 , \2753 );
not \U$2076 ( \2755 , \2754 );
nor \U$2077 ( \2756 , \2753 , \2595 );
nor \U$2078 ( \2757 , \2755 , \2756 );
not \U$2079 ( \2758 , \2757 );
not \U$2080 ( \2759 , \2507 );
not \U$2081 ( \2760 , \2580 );
and \U$2082 ( \2761 , \2759 , \2760 );
and \U$2083 ( \2762 , \2507 , \2580 );
nor \U$2084 ( \2763 , \2761 , \2762 );
not \U$2085 ( \2764 , \2763 );
and \U$2086 ( \2765 , \2758 , \2764 );
and \U$2087 ( \2766 , \2757 , \2763 );
nor \U$2088 ( \2767 , \2765 , \2766 );
xor \U$2089 ( \2768 , \2734 , \2747 );
xor \U$2090 ( \2769 , \2768 , \2750 );
not \U$2091 ( \2770 , \2746 );
not \U$2092 ( \2771 , \2739 );
or \U$2093 ( \2772 , \2770 , \2771 );
or \U$2094 ( \2773 , \2739 , \2746 );
nand \U$2095 ( \2774 , \2772 , \2773 );
not \U$2096 ( \2775 , \2774 );
xor \U$2097 ( \2776 , \2540 , \2547 );
xor \U$2098 ( \2777 , \2776 , \2555 );
not \U$2099 ( \2778 , \2777 );
nand \U$2100 ( \2779 , \2156_nGf08 , \1523 );
or \U$2101 ( \2780 , \1449 , \2229_nGe35 );
nand \U$2102 ( \2781 , \2780 , \1529 );
and \U$2103 ( \2782 , \2779 , \2781 );
and \U$2104 ( \2783 , \1525 , \2229_nGe35 );
and \U$2105 ( \2784 , \2156_nGf08 , \1594 );
nor \U$2106 ( \2785 , \2782 , \2783 , \2784 );
and \U$2107 ( \2786 , \2034_nGfe1 , \1653 );
or \U$2108 ( \2787 , \1579 , \1787_nG10e2 );
nand \U$2109 ( \2788 , \2787 , \1799 );
nand \U$2110 ( \2789 , \2034_nGfe1 , \1650 );
and \U$2111 ( \2790 , \2788 , \2789 );
and \U$2112 ( \2791 , \1787_nG10e2 , \1794 );
nor \U$2113 ( \2792 , \2786 , \2790 , \2791 );
xor \U$2114 ( \2793 , \2785 , \2792 );
and \U$2115 ( \2794 , \2446_nGa9e , \1363 );
and \U$2116 ( \2795 , \1400 , \2404_nGad6 );
nand \U$2117 ( \2796 , \2446_nGa9e , \1360 );
or \U$2118 ( \2797 , \1320 , \2404_nGad6 );
nand \U$2119 ( \2798 , \2797 , \1404 );
and \U$2120 ( \2799 , \2796 , \2798 );
nor \U$2121 ( \2800 , \2794 , \2795 , \2799 );
and \U$2122 ( \2801 , \2793 , \2800 );
and \U$2123 ( \2802 , \2785 , \2792 );
or \U$2124 ( \2803 , \2801 , \2802 );
nand \U$2125 ( \2804 , \1559_nG13c8 , \2100 );
or \U$2126 ( \2805 , \1969 , \1502_nG14c8 );
nand \U$2127 ( \2806 , \2805 , \2286 );
and \U$2128 ( \2807 , \2804 , \2806 );
and \U$2129 ( \2808 , \2289 , \1502_nG14c8 );
and \U$2130 ( \2809 , \1559_nG13c8 , \2103 );
nor \U$2131 ( \2810 , \2807 , \2808 , \2809 );
and \U$2132 ( \2811 , \1349 , \2541 );
not \U$2133 ( \2812 , \1435_nG15b1 );
and \U$2134 ( \2813 , \2371 , \2812 );
and \U$2135 ( \2814 , \1348_nG16d6 , \2545 );
nor \U$2136 ( \2815 , \2811 , \2813 , \2814 );
xor \U$2137 ( \2816 , \2810 , \2815 );
nand \U$2138 ( \2817 , \1710_nG11c1 , \1865 );
or \U$2139 ( \2818 , \1810 , \1631_nG12c9 );
nand \U$2140 ( \2819 , \2818 , \1973 );
and \U$2141 ( \2820 , \2817 , \2819 );
and \U$2142 ( \2821 , \1976 , \1631_nG12c9 );
and \U$2143 ( \2822 , \1710_nG11c1 , \1868 );
nor \U$2144 ( \2823 , \2820 , \2821 , \2822 );
and \U$2145 ( \2824 , \2816 , \2823 );
and \U$2146 ( \2825 , \2810 , \2815 );
or \U$2147 ( \2826 , \2824 , \2825 );
nor \U$2148 ( \2827 , \2803 , \2826 );
nand \U$2149 ( \2828 , \2778 , \2827 );
or \U$2150 ( \2829 , \2775 , \2828 );
not \U$2151 ( \2830 , \2828 );
not \U$2152 ( \2831 , \2775 );
or \U$2153 ( \2832 , \2830 , \2831 );
not \U$2154 ( \2833 , \2731 );
not \U$2155 ( \2834 , \2733 );
nand \U$2156 ( \2835 , \2834 , \2718 );
not \U$2157 ( \2836 , \2835 );
or \U$2158 ( \2837 , \2833 , \2836 );
or \U$2159 ( \2838 , \2835 , \2731 );
nand \U$2160 ( \2839 , \2837 , \2838 );
nand \U$2161 ( \2840 , \2832 , \2839 );
nand \U$2162 ( \2841 , \2829 , \2840 );
xor \U$2163 ( \2842 , \2559 , \2566 );
xor \U$2164 ( \2843 , \2842 , \2577 );
nor \U$2165 ( \2844 , \2841 , \2843 );
or \U$2166 ( \2845 , \2769 , \2844 );
nand \U$2167 ( \2846 , \2843 , \2841 );
nand \U$2168 ( \2847 , \2845 , \2846 );
xor \U$2169 ( \2848 , \2767 , \2847 );
not \U$2170 ( \2849 , \2844 );
nand \U$2171 ( \2850 , \2849 , \2846 );
not \U$2172 ( \2851 , \2850 );
not \U$2173 ( \2852 , \2769 );
or \U$2174 ( \2853 , \2851 , \2852 );
or \U$2175 ( \2854 , \2769 , \2850 );
nand \U$2176 ( \2855 , \2853 , \2854 );
not \U$2177 ( \2856 , \2826 );
or \U$2178 ( \2857 , \2803 , \2856 );
not \U$2179 ( \2858 , \2803 );
or \U$2180 ( \2859 , \2826 , \2858 );
and \U$2181 ( \2860 , RIaaa6d88_528, \730 );
and \U$2182 ( \2861 , RIaaa6ab8_522, \682 );
and \U$2183 ( \2862 , \686 , RIaaa6f68_532);
and \U$2184 ( \2863 , RIaaa6e00_529, \690 );
nor \U$2185 ( \2864 , \2862 , \2863 );
and \U$2186 ( \2865 , \702 , RIaaa6e78_530);
and \U$2187 ( \2866 , RIaaa6ba8_524, \721 );
nor \U$2188 ( \2867 , \2865 , \2866 );
and \U$2189 ( \2868 , \696 , RIaaa6a40_521);
and \U$2190 ( \2869 , RIaaa6ef0_531, \699 );
nor \U$2191 ( \2870 , \2868 , \2869 );
and \U$2192 ( \2871 , \1241 , RIaaa7058_534);
and \U$2193 ( \2872 , RIaaa6d10_527, \712 );
nor \U$2194 ( \2873 , \2871 , \2872 );
nand \U$2195 ( \2874 , \2864 , \2867 , \2870 , \2873 );
nor \U$2196 ( \2875 , \2860 , \2861 , \2874 );
and \U$2197 ( \2876 , \723 , RIaaa69c8_520);
and \U$2198 ( \2877 , RIaaa6b30_523, \728 );
nor \U$2199 ( \2878 , \2876 , \2877 );
and \U$2200 ( \2879 , \738 , RIaaa6fe0_533);
and \U$2201 ( \2880 , RIaaa6c20_525, \733 );
nor \U$2202 ( \2881 , \2879 , \2880 );
and \U$2203 ( \2882 , \735 , RIaaa6c98_526);
and \U$2204 ( \2883 , RIaaa70d0_535, \742 );
nor \U$2205 ( \2884 , \2882 , \2883 );
nand \U$2206 ( \2885 , \2875 , \2878 , \2881 , \2884 );
_DC g9f5 ( \2886_nG9f5 , \2885 , \1252 );
nand \U$2207 ( \2887 , \2886_nG9f5 , \1223 );
and \U$2208 ( \2888 , \2653_nGa66 , \1306 );
or \U$2209 ( \2889 , \1266 , \2695_nGa2d );
nand \U$2210 ( \2890 , \2889 , \1303 );
nand \U$2211 ( \2891 , \2653_nGa66 , \1299 );
and \U$2212 ( \2892 , \2890 , \2891 );
and \U$2213 ( \2893 , \2695_nGa2d , \1440 );
nor \U$2214 ( \2894 , \2888 , \2892 , \2893 );
or \U$2215 ( \2895 , \2887 , \2894 );
nand \U$2216 ( \2896 , \2857 , \2859 , \2895 );
xor \U$2217 ( \2897 , \2705 , \2713 );
xor \U$2218 ( \2898 , \2896 , \2897 );
not \U$2219 ( \2899 , \2696 );
nor \U$2220 ( \2900 , \2667 , \2699 );
not \U$2221 ( \2901 , \2900 );
or \U$2222 ( \2902 , \2899 , \2901 );
or \U$2223 ( \2903 , \2900 , \2696 );
nand \U$2224 ( \2904 , \2902 , \2903 );
and \U$2225 ( \2905 , \2898 , \2904 );
and \U$2226 ( \2906 , \2896 , \2897 );
or \U$2227 ( \2907 , \2905 , \2906 );
xor \U$2228 ( \2908 , \2721 , \2730 );
and \U$2229 ( \2909 , \2907 , \2908 );
not \U$2230 ( \2910 , \2907 );
not \U$2231 ( \2911 , \2908 );
and \U$2232 ( \2912 , \2910 , \2911 );
xnor \U$2233 ( \2913 , \2887 , \2894 );
xor \U$2234 ( \2914 , \2785 , \2792 );
xor \U$2235 ( \2915 , \2914 , \2800 );
and \U$2236 ( \2916 , \2913 , \2915 );
not \U$2237 ( \2917 , \2916 );
xor \U$2238 ( \2918 , \2810 , \2815 );
xor \U$2239 ( \2919 , \2918 , \2823 );
not \U$2240 ( \2920 , \2919 );
and \U$2241 ( \2921 , \2917 , \2920 );
nor \U$2242 ( \2922 , \2913 , \2915 );
nor \U$2243 ( \2923 , \2921 , \2922 );
xor \U$2244 ( \2924 , \2607 , \2614 );
xor \U$2245 ( \2925 , \2924 , \2622 );
xor \U$2246 ( \2926 , \2923 , \2925 );
and \U$2247 ( \2927 , \2156_nGf08 , \1653 );
or \U$2248 ( \2928 , \1579 , \2034_nGfe1 );
nand \U$2249 ( \2929 , \2928 , \1799 );
nand \U$2250 ( \2930 , \2156_nGf08 , \1650 );
and \U$2251 ( \2931 , \2929 , \2930 );
and \U$2252 ( \2932 , \2034_nGfe1 , \1794 );
nor \U$2253 ( \2933 , \2927 , \2931 , \2932 );
nand \U$2254 ( \2934 , \1787_nG10e2 , \1865 );
or \U$2255 ( \2935 , \1810 , \1710_nG11c1 );
nand \U$2256 ( \2936 , \2935 , \1973 );
and \U$2257 ( \2937 , \2934 , \2936 );
and \U$2258 ( \2938 , \1976 , \1710_nG11c1 );
and \U$2259 ( \2939 , \1787_nG10e2 , \1868 );
nor \U$2260 ( \2940 , \2937 , \2938 , \2939 );
xor \U$2261 ( \2941 , \2933 , \2940 );
nand \U$2262 ( \2942 , \2229_nGe35 , \1523 );
or \U$2263 ( \2943 , \1449 , \2404_nGad6 );
nand \U$2264 ( \2944 , \2943 , \1529 );
and \U$2265 ( \2945 , \2942 , \2944 );
and \U$2266 ( \2946 , \1525 , \2404_nGad6 );
and \U$2267 ( \2947 , \2229_nGe35 , \1594 );
nor \U$2268 ( \2948 , \2945 , \2946 , \2947 );
and \U$2269 ( \2949 , \2941 , \2948 );
and \U$2270 ( \2950 , \2933 , \2940 );
or \U$2271 ( \2951 , \2949 , \2950 );
nand \U$2272 ( \2952 , \1631_nG12c9 , \2100 );
or \U$2273 ( \2953 , \1969 , \1559_nG13c8 );
nand \U$2274 ( \2954 , \2953 , \2286 );
and \U$2275 ( \2955 , \2952 , \2954 );
and \U$2276 ( \2956 , \2289 , \1559_nG13c8 );
and \U$2277 ( \2957 , \1631_nG12c9 , \2103 );
nor \U$2278 ( \2958 , \2955 , \2956 , \2957 );
not \U$2279 ( \2959 , \2958 );
or \U$2280 ( \2960 , \2544 , \2812 );
or \U$2281 ( \2961 , \1435_nG15b1 , \2373 );
or \U$2282 ( \2962 , \1502_nG14c8 , \2372 );
nand \U$2283 ( \2963 , \2960 , \2961 , \2962 );
nand \U$2284 ( \2964 , \2959 , \2963 );
xor \U$2285 ( \2965 , \2951 , \2964 );
and \U$2286 ( \2966 , \2695_nGa2d , \1306 );
or \U$2287 ( \2967 , \1266 , \2886_nG9f5 );
nand \U$2288 ( \2968 , \2967 , \1303 );
nand \U$2289 ( \2969 , \2695_nGa2d , \1299 );
and \U$2290 ( \2970 , \2968 , \2969 );
and \U$2291 ( \2971 , \2886_nG9f5 , \1440 );
nor \U$2292 ( \2972 , \2966 , \2970 , \2971 );
and \U$2293 ( \2973 , \2653_nGa66 , \1363 );
and \U$2294 ( \2974 , \1400 , \2446_nGa9e );
nand \U$2295 ( \2975 , \2653_nGa66 , \1360 );
or \U$2296 ( \2976 , \1320 , \2446_nGa9e );
nand \U$2297 ( \2977 , \2976 , \1404 );
and \U$2298 ( \2978 , \2975 , \2977 );
nor \U$2299 ( \2979 , \2973 , \2974 , \2978 );
and \U$2300 ( \2980 , \2972 , \2979 );
not \U$2301 ( \2981 , \2980 );
and \U$2302 ( \2982 , RIaaa7418_542, \721 );
and \U$2303 ( \2983 , RIaaa7940_553, \686 );
and \U$2304 ( \2984 , \742 , RIaaa7328_540);
and \U$2305 ( \2985 , RIaaa77d8_550, \730 );
nor \U$2306 ( \2986 , \2984 , \2985 );
and \U$2307 ( \2987 , \723 , RIaaa7490_543);
and \U$2308 ( \2988 , RIaaa73a0_541, \733 );
nor \U$2309 ( \2989 , \2987 , \2988 );
and \U$2310 ( \2990 , \738 , RIaaa7238_538);
and \U$2311 ( \2991 , RIaaa76e8_548, \735 );
nor \U$2312 ( \2992 , \2990 , \2991 );
and \U$2313 ( \2993 , \682 , RIaaa7670_547);
and \U$2314 ( \2994 , RIaaa75f8_546, \728 );
nor \U$2315 ( \2995 , \2993 , \2994 );
nand \U$2316 ( \2996 , \2986 , \2989 , \2992 , \2995 );
nor \U$2317 ( \2997 , \2982 , \2983 , \2996 );
and \U$2318 ( \2998 , \702 , RIaaa7508_544);
and \U$2319 ( \2999 , RIaaa7760_549, \712 );
nor \U$2320 ( \3000 , \2998 , \2999 );
and \U$2321 ( \3001 , \1241 , RIaaa72b0_539);
and \U$2322 ( \3002 , RIaaa78c8_552, \699 );
nor \U$2323 ( \3003 , \3001 , \3002 );
and \U$2324 ( \3004 , \696 , RIaaa7580_545);
and \U$2325 ( \3005 , RIaaa7850_551, \690 );
nor \U$2326 ( \3006 , \3004 , \3005 );
nand \U$2327 ( \3007 , \2997 , \3000 , \3003 , \3006 );
_DC g9b9 ( \3008_nG9b9 , \3007 , \1252 );
nand \U$2328 ( \3009 , \3008_nG9b9 , \1223 );
not \U$2329 ( \3010 , \3009 );
and \U$2330 ( \3011 , \2981 , \3010 );
nor \U$2331 ( \3012 , \2972 , \2979 );
nor \U$2332 ( \3013 , \3011 , \3012 );
and \U$2333 ( \3014 , \2965 , \3013 );
and \U$2334 ( \3015 , \2951 , \2964 );
or \U$2335 ( \3016 , \3014 , \3015 );
and \U$2336 ( \3017 , \2926 , \3016 );
and \U$2337 ( \3018 , \2923 , \2925 );
or \U$2338 ( \3019 , \3017 , \3018 );
nor \U$2339 ( \3020 , \2912 , \3019 );
nor \U$2340 ( \3021 , \2909 , \3020 );
not \U$2341 ( \3022 , \2827 );
not \U$2342 ( \3023 , \2777 );
and \U$2343 ( \3024 , \3022 , \3023 );
and \U$2344 ( \3025 , \2827 , \2777 );
nor \U$2345 ( \3026 , \3024 , \3025 );
not \U$2346 ( \3027 , \3026 );
not \U$2347 ( \3028 , \2714 );
not \U$2348 ( \3029 , \2716 );
nand \U$2349 ( \3030 , \3029 , \2701 );
not \U$2350 ( \3031 , \3030 );
or \U$2351 ( \3032 , \3028 , \3031 );
or \U$2352 ( \3033 , \3030 , \2714 );
nand \U$2353 ( \3034 , \3032 , \3033 );
nand \U$2354 ( \3035 , \3027 , \3034 );
xor \U$2355 ( \3036 , \3021 , \3035 );
not \U$2356 ( \3037 , \2839 );
not \U$2357 ( \3038 , \2828 );
and \U$2358 ( \3039 , \3037 , \3038 );
and \U$2359 ( \3040 , \2839 , \2828 );
nor \U$2360 ( \3041 , \3039 , \3040 );
not \U$2361 ( \3042 , \3041 );
not \U$2362 ( \3043 , \2774 );
and \U$2363 ( \3044 , \3042 , \3043 );
and \U$2364 ( \3045 , \3041 , \2774 );
nor \U$2365 ( \3046 , \3044 , \3045 );
and \U$2366 ( \3047 , \3036 , \3046 );
and \U$2367 ( \3048 , \3021 , \3035 );
or \U$2368 ( \3049 , \3047 , \3048 );
xor \U$2369 ( \3050 , \2855 , \3049 );
xor \U$2370 ( \3051 , \2923 , \2925 );
xor \U$2371 ( \3052 , \3051 , \3016 );
not \U$2372 ( \3053 , \3009 );
nor \U$2373 ( \3054 , \2980 , \3012 );
not \U$2374 ( \3055 , \3054 );
or \U$2375 ( \3056 , \3053 , \3055 );
or \U$2376 ( \3057 , \3054 , \3009 );
nand \U$2377 ( \3058 , \3056 , \3057 );
not \U$2378 ( \3059 , \3058 );
xor \U$2379 ( \3060 , \2933 , \2940 );
xor \U$2380 ( \3061 , \3060 , \2948 );
nor \U$2381 ( \3062 , \3059 , \3061 );
nand \U$2382 ( \3063 , \2404_nGad6 , \1523 );
or \U$2383 ( \3064 , \1449 , \2446_nGa9e );
nand \U$2384 ( \3065 , \3064 , \1529 );
and \U$2385 ( \3066 , \3063 , \3065 );
and \U$2386 ( \3067 , \1525 , \2446_nGa9e );
and \U$2387 ( \3068 , \2404_nGad6 , \1594 );
nor \U$2388 ( \3069 , \3066 , \3067 , \3068 );
and \U$2389 ( \3070 , \2229_nGe35 , \1653 );
or \U$2390 ( \3071 , \1579 , \2156_nGf08 );
nand \U$2391 ( \3072 , \3071 , \1799 );
nand \U$2392 ( \3073 , \2229_nGe35 , \1650 );
and \U$2393 ( \3074 , \3072 , \3073 );
and \U$2394 ( \3075 , \2156_nGf08 , \1794 );
nor \U$2395 ( \3076 , \3070 , \3074 , \3075 );
xor \U$2396 ( \3077 , \3069 , \3076 );
and \U$2397 ( \3078 , \2695_nGa2d , \1363 );
and \U$2398 ( \3079 , \1400 , \2653_nGa66 );
nand \U$2399 ( \3080 , \2695_nGa2d , \1360 );
or \U$2400 ( \3081 , \1320 , \2653_nGa66 );
nand \U$2401 ( \3082 , \3081 , \1404 );
and \U$2402 ( \3083 , \3080 , \3082 );
nor \U$2403 ( \3084 , \3078 , \3079 , \3083 );
and \U$2404 ( \3085 , \3077 , \3084 );
and \U$2405 ( \3086 , \3069 , \3076 );
or \U$2406 ( \3087 , \3085 , \3086 );
nand \U$2407 ( \3088 , \1710_nG11c1 , \2100 );
or \U$2408 ( \3089 , \1969 , \1631_nG12c9 );
nand \U$2409 ( \3090 , \3089 , \2286 );
and \U$2410 ( \3091 , \3088 , \3090 );
and \U$2411 ( \3092 , \2289 , \1631_nG12c9 );
and \U$2412 ( \3093 , \1710_nG11c1 , \2103 );
nor \U$2413 ( \3094 , \3091 , \3092 , \3093 );
and \U$2414 ( \3095 , \1503 , \2541 );
and \U$2415 ( \3096 , \2371 , \1635 );
and \U$2416 ( \3097 , \1502_nG14c8 , \2545 );
nor \U$2417 ( \3098 , \3095 , \3096 , \3097 );
xor \U$2418 ( \3099 , \3094 , \3098 );
nand \U$2419 ( \3100 , \2034_nGfe1 , \1865 );
or \U$2420 ( \3101 , \1810 , \1787_nG10e2 );
nand \U$2421 ( \3102 , \3101 , \1973 );
and \U$2422 ( \3103 , \3100 , \3102 );
and \U$2423 ( \3104 , \1976 , \1787_nG10e2 );
and \U$2424 ( \3105 , \2034_nGfe1 , \1868 );
nor \U$2425 ( \3106 , \3103 , \3104 , \3105 );
and \U$2426 ( \3107 , \3099 , \3106 );
and \U$2427 ( \3108 , \3094 , \3098 );
or \U$2428 ( \3109 , \3107 , \3108 );
nor \U$2429 ( \3110 , \3087 , \3109 );
xor \U$2430 ( \3111 , \3062 , \3110 );
not \U$2431 ( \3112 , \2919 );
nor \U$2432 ( \3113 , \2922 , \2916 );
not \U$2433 ( \3114 , \3113 );
or \U$2434 ( \3115 , \3112 , \3114 );
or \U$2435 ( \3116 , \3113 , \2919 );
nand \U$2436 ( \3117 , \3115 , \3116 );
and \U$2437 ( \3118 , \3111 , \3117 );
and \U$2438 ( \3119 , \3062 , \3110 );
or \U$2439 ( \3120 , \3118 , \3119 );
xor \U$2440 ( \3121 , \2896 , \2897 );
xor \U$2441 ( \3122 , \3121 , \2904 );
nor \U$2442 ( \3123 , \3120 , \3122 );
or \U$2443 ( \3124 , \3052 , \3123 );
nand \U$2444 ( \3125 , \3122 , \3120 );
nand \U$2445 ( \3126 , \3124 , \3125 );
not \U$2446 ( \3127 , \3026 );
not \U$2447 ( \3128 , \3034 );
or \U$2448 ( \3129 , \3127 , \3128 );
or \U$2449 ( \3130 , \3034 , \3026 );
nand \U$2450 ( \3131 , \3129 , \3130 );
xor \U$2451 ( \3132 , \3126 , \3131 );
not \U$2452 ( \3133 , \2907 );
not \U$2453 ( \3134 , \3019 );
not \U$2454 ( \3135 , \2908 );
and \U$2455 ( \3136 , \3134 , \3135 );
and \U$2456 ( \3137 , \3019 , \2908 );
nor \U$2457 ( \3138 , \3136 , \3137 );
not \U$2458 ( \3139 , \3138 );
or \U$2459 ( \3140 , \3133 , \3139 );
or \U$2460 ( \3141 , \3138 , \2907 );
nand \U$2461 ( \3142 , \3140 , \3141 );
xor \U$2462 ( \3143 , \3132 , \3142 );
not \U$2463 ( \3144 , \3125 );
nor \U$2464 ( \3145 , \3144 , \3123 );
not \U$2465 ( \3146 , \3145 );
not \U$2466 ( \3147 , \3052 );
and \U$2467 ( \3148 , \3146 , \3147 );
and \U$2468 ( \3149 , \3145 , \3052 );
nor \U$2469 ( \3150 , \3148 , \3149 );
xor \U$2470 ( \3151 , \3069 , \3076 );
xor \U$2471 ( \3152 , \3151 , \3084 );
xor \U$2472 ( \3153 , \3094 , \3098 );
xor \U$2473 ( \3154 , \3153 , \3106 );
xor \U$2474 ( \3155 , \3152 , \3154 );
and \U$2475 ( \3156 , RIaaa87c8_584, \730 );
and \U$2476 ( \3157 , RIaaa8660_581, \682 );
and \U$2477 ( \3158 , \686 , RIaaa8930_587);
and \U$2478 ( \3159 , RIaaa8840_585, \690 );
nor \U$2479 ( \3160 , \3158 , \3159 );
and \U$2480 ( \3161 , \702 , RIaaa84f8_578);
and \U$2481 ( \3162 , RIaaa8480_577, \721 );
nor \U$2482 ( \3163 , \3161 , \3162 );
and \U$2483 ( \3164 , \696 , RIaaa8570_579);
and \U$2484 ( \3165 , RIaaa88b8_586, \699 );
nor \U$2485 ( \3166 , \3164 , \3165 );
and \U$2486 ( \3167 , \1241 , RIaaa82a0_573);
and \U$2487 ( \3168 , RIaaa8750_583, \712 );
nor \U$2488 ( \3169 , \3167 , \3168 );
nand \U$2489 ( \3170 , \3160 , \3163 , \3166 , \3169 );
nor \U$2490 ( \3171 , \3156 , \3157 , \3170 );
and \U$2491 ( \3172 , \723 , RIaaa8408_576);
and \U$2492 ( \3173 , RIaaa85e8_580, \728 );
nor \U$2493 ( \3174 , \3172 , \3173 );
and \U$2494 ( \3175 , \738 , RIaaa8228_572);
and \U$2495 ( \3176 , RIaaa8390_575, \733 );
nor \U$2496 ( \3177 , \3175 , \3176 );
and \U$2497 ( \3178 , \735 , RIaaa86d8_582);
and \U$2498 ( \3179 , RIaaa8318_574, \742 );
nor \U$2499 ( \3180 , \3178 , \3179 );
nand \U$2500 ( \3181 , \3171 , \3174 , \3177 , \3180 );
_DC g984 ( \3182_nG984 , \3181 , \1252 );
nand \U$2501 ( \3183 , \3182_nG984 , \1223 );
and \U$2502 ( \3184 , \2886_nG9f5 , \1306 );
or \U$2503 ( \3185 , \1266 , \3008_nG9b9 );
nand \U$2504 ( \3186 , \3185 , \1303 );
nand \U$2505 ( \3187 , \2886_nG9f5 , \1299 );
and \U$2506 ( \3188 , \3186 , \3187 );
and \U$2507 ( \3189 , \3008_nG9b9 , \1440 );
nor \U$2508 ( \3190 , \3184 , \3188 , \3189 );
xnor \U$2509 ( \3191 , \3183 , \3190 );
and \U$2510 ( \3192 , \3155 , \3191 );
and \U$2511 ( \3193 , \3152 , \3154 );
or \U$2512 ( \3194 , \3192 , \3193 );
not \U$2513 ( \3195 , \2958 );
not \U$2514 ( \3196 , \2963 );
and \U$2515 ( \3197 , \3195 , \3196 );
and \U$2516 ( \3198 , \2958 , \2963 );
nor \U$2517 ( \3199 , \3197 , \3198 );
xor \U$2518 ( \3200 , \3194 , \3199 );
and \U$2519 ( \3201 , \2404_nGad6 , \1653 );
or \U$2520 ( \3202 , \1579 , \2229_nGe35 );
nand \U$2521 ( \3203 , \3202 , \1799 );
nand \U$2522 ( \3204 , \2404_nGad6 , \1650 );
and \U$2523 ( \3205 , \3203 , \3204 );
and \U$2524 ( \3206 , \2229_nGe35 , \1794 );
nor \U$2525 ( \3207 , \3201 , \3205 , \3206 );
nand \U$2526 ( \3208 , \2156_nGf08 , \1865 );
or \U$2527 ( \3209 , \1810 , \2034_nGfe1 );
nand \U$2528 ( \3210 , \3209 , \1973 );
and \U$2529 ( \3211 , \3208 , \3210 );
and \U$2530 ( \3212 , \1976 , \2034_nGfe1 );
and \U$2531 ( \3213 , \2156_nGf08 , \1868 );
nor \U$2532 ( \3214 , \3211 , \3212 , \3213 );
xor \U$2533 ( \3215 , \3207 , \3214 );
nand \U$2534 ( \3216 , \2446_nGa9e , \1523 );
or \U$2535 ( \3217 , \1449 , \2653_nGa66 );
nand \U$2536 ( \3218 , \3217 , \1529 );
and \U$2537 ( \3219 , \3216 , \3218 );
and \U$2538 ( \3220 , \1525 , \2653_nGa66 );
and \U$2539 ( \3221 , \2446_nGa9e , \1594 );
nor \U$2540 ( \3222 , \3219 , \3220 , \3221 );
and \U$2541 ( \3223 , \3215 , \3222 );
and \U$2542 ( \3224 , \3207 , \3214 );
or \U$2543 ( \3225 , \3223 , \3224 );
nand \U$2544 ( \3226 , \1787_nG10e2 , \2100 );
or \U$2545 ( \3227 , \1969 , \1710_nG11c1 );
nand \U$2546 ( \3228 , \3227 , \2286 );
and \U$2547 ( \3229 , \3226 , \3228 );
and \U$2548 ( \3230 , \2289 , \1710_nG11c1 );
and \U$2549 ( \3231 , \1787_nG10e2 , \2103 );
nor \U$2550 ( \3232 , \3229 , \3230 , \3231 );
not \U$2551 ( \3233 , \3232 );
or \U$2552 ( \3234 , \2544 , \1635 );
or \U$2553 ( \3235 , \1559_nG13c8 , \2373 );
or \U$2554 ( \3236 , \1631_nG12c9 , \2372 );
nand \U$2555 ( \3237 , \3234 , \3235 , \3236 );
nand \U$2556 ( \3238 , \3233 , \3237 );
xor \U$2557 ( \3239 , \3225 , \3238 );
and \U$2558 ( \3240 , \2886_nG9f5 , \1363 );
and \U$2559 ( \3241 , \1400 , \2695_nGa2d );
nand \U$2560 ( \3242 , \2886_nG9f5 , \1360 );
or \U$2561 ( \3243 , \1320 , \2695_nGa2d );
nand \U$2562 ( \3244 , \3243 , \1404 );
and \U$2563 ( \3245 , \3242 , \3244 );
nor \U$2564 ( \3246 , \3240 , \3241 , \3245 );
and \U$2565 ( \3247 , RIaaa7aa8_556, \723 );
and \U$2566 ( \3248 , RIaaa80c0_569, \730 );
and \U$2567 ( \3249 , \686 , RIaaa7c88_560);
and \U$2568 ( \3250 , RIaaa8138_570, \690 );
nor \U$2569 ( \3251 , \3249 , \3250 );
and \U$2570 ( \3252 , \702 , RIaaa8048_568);
and \U$2571 ( \3253 , RIaaa7c10_559, \721 );
nor \U$2572 ( \3254 , \3252 , \3253 );
and \U$2573 ( \3255 , \696 , RIaaa7b20_557);
and \U$2574 ( \3256 , RIaaa7d00_561, \699 );
nor \U$2575 ( \3257 , \3255 , \3256 );
and \U$2576 ( \3258 , \1241 , RIaaa7e68_564);
and \U$2577 ( \3259 , RIaaa7fd0_567, \712 );
nor \U$2578 ( \3260 , \3258 , \3259 );
nand \U$2579 ( \3261 , \3251 , \3254 , \3257 , \3260 );
nor \U$2580 ( \3262 , \3247 , \3248 , \3261 );
and \U$2581 ( \3263 , \738 , RIaaa7d78_562);
and \U$2582 ( \3264 , RIaaa7a30_555, \682 );
nor \U$2583 ( \3265 , \3263 , \3264 );
and \U$2584 ( \3266 , \733 , RIaaa7b98_558);
and \U$2585 ( \3267 , RIaaa7f58_566, \735 );
nor \U$2586 ( \3268 , \3266 , \3267 );
and \U$2587 ( \3269 , \728 , RIaaa79b8_554);
and \U$2588 ( \3270 , RIaaa7df0_563, \742 );
nor \U$2589 ( \3271 , \3269 , \3270 );
nand \U$2590 ( \3272 , \3262 , \3265 , \3268 , \3271 );
_DC g944 ( \3273_nG944 , \3272 , \1252 );
nand \U$2591 ( \3274 , \3273_nG944 , \1223 );
xor \U$2592 ( \3275 , \3246 , \3274 );
and \U$2593 ( \3276 , \3008_nG9b9 , \1306 );
or \U$2594 ( \3277 , \1266 , \3182_nG984 );
nand \U$2595 ( \3278 , \3277 , \1303 );
nand \U$2596 ( \3279 , \3008_nG9b9 , \1299 );
and \U$2597 ( \3280 , \3278 , \3279 );
and \U$2598 ( \3281 , \3182_nG984 , \1440 );
nor \U$2599 ( \3282 , \3276 , \3280 , \3281 );
and \U$2600 ( \3283 , \3275 , \3282 );
and \U$2601 ( \3284 , \3246 , \3274 );
or \U$2602 ( \3285 , \3283 , \3284 );
and \U$2603 ( \3286 , \3239 , \3285 );
and \U$2604 ( \3287 , \3225 , \3238 );
or \U$2605 ( \3288 , \3286 , \3287 );
and \U$2606 ( \3289 , \3200 , \3288 );
and \U$2607 ( \3290 , \3194 , \3199 );
or \U$2608 ( \3291 , \3289 , \3290 );
xor \U$2609 ( \3292 , \2951 , \2964 );
xor \U$2610 ( \3293 , \3292 , \3013 );
and \U$2611 ( \3294 , \3291 , \3293 );
not \U$2612 ( \3295 , \3294 );
not \U$2613 ( \3296 , \3058 );
not \U$2614 ( \3297 , \3061 );
and \U$2615 ( \3298 , \3296 , \3297 );
and \U$2616 ( \3299 , \3058 , \3061 );
nor \U$2617 ( \3300 , \3298 , \3299 );
not \U$2618 ( \3301 , \3300 );
not \U$2619 ( \3302 , \3109 );
or \U$2620 ( \3303 , \3087 , \3302 );
not \U$2621 ( \3304 , \3087 );
or \U$2622 ( \3305 , \3109 , \3304 );
or \U$2623 ( \3306 , \3183 , \3190 );
nand \U$2624 ( \3307 , \3303 , \3305 , \3306 );
nand \U$2625 ( \3308 , \3301 , \3307 );
not \U$2626 ( \3309 , \3308 );
and \U$2627 ( \3310 , \3295 , \3309 );
nor \U$2628 ( \3311 , \3291 , \3293 );
nor \U$2629 ( \3312 , \3310 , \3311 );
nor \U$2630 ( \3313 , \3150 , \3312 );
xor \U$2631 ( \3314 , \3143 , \3313 );
and \U$2632 ( \3315 , \3150 , \3312 );
nor \U$2633 ( \3316 , \3315 , \3313 );
xor \U$2634 ( \3317 , \3062 , \3110 );
xor \U$2635 ( \3318 , \3317 , \3117 );
not \U$2636 ( \3319 , \3308 );
nor \U$2637 ( \3320 , \3311 , \3294 );
not \U$2638 ( \3321 , \3320 );
or \U$2639 ( \3322 , \3319 , \3321 );
or \U$2640 ( \3323 , \3320 , \3308 );
nand \U$2641 ( \3324 , \3322 , \3323 );
nand \U$2642 ( \3325 , \3318 , \3324 );
not \U$2643 ( \3326 , \3325 );
xor \U$2644 ( \3327 , \3316 , \3326 );
or \U$2645 ( \3328 , \3324 , \3318 );
nand \U$2646 ( \3329 , \3328 , \3325 );
xor \U$2647 ( \3330 , \3194 , \3199 );
xor \U$2648 ( \3331 , \3330 , \3288 );
not \U$2649 ( \3332 , \3300 );
not \U$2650 ( \3333 , \3307 );
and \U$2651 ( \3334 , \3332 , \3333 );
and \U$2652 ( \3335 , \3300 , \3307 );
nor \U$2653 ( \3336 , \3334 , \3335 );
xor \U$2654 ( \3337 , \3331 , \3336 );
xor \U$2655 ( \3338 , \3207 , \3214 );
xor \U$2656 ( \3339 , \3338 , \3222 );
not \U$2657 ( \3340 , \3339 );
not \U$2658 ( \3341 , \3237 );
not \U$2659 ( \3342 , \3232 );
or \U$2660 ( \3343 , \3341 , \3342 );
or \U$2661 ( \3344 , \3232 , \3237 );
nand \U$2662 ( \3345 , \3343 , \3344 );
nand \U$2663 ( \3346 , \3340 , \3345 );
xor \U$2664 ( \3347 , \3152 , \3154 );
xor \U$2665 ( \3348 , \3347 , \3191 );
and \U$2666 ( \3349 , \3346 , \3348 );
nand \U$2667 ( \3350 , \2653_nGa66 , \1523 );
or \U$2668 ( \3351 , \1449 , \2695_nGa2d );
nand \U$2669 ( \3352 , \3351 , \1529 );
and \U$2670 ( \3353 , \3350 , \3352 );
and \U$2671 ( \3354 , \1525 , \2695_nGa2d );
and \U$2672 ( \3355 , \2653_nGa66 , \1594 );
nor \U$2673 ( \3356 , \3353 , \3354 , \3355 );
and \U$2674 ( \3357 , \2446_nGa9e , \1653 );
or \U$2675 ( \3358 , \1579 , \2404_nGad6 );
nand \U$2676 ( \3359 , \3358 , \1799 );
nand \U$2677 ( \3360 , \2446_nGa9e , \1650 );
and \U$2678 ( \3361 , \3359 , \3360 );
and \U$2679 ( \3362 , \2404_nGad6 , \1794 );
nor \U$2680 ( \3363 , \3357 , \3361 , \3362 );
xor \U$2681 ( \3364 , \3356 , \3363 );
and \U$2682 ( \3365 , \3008_nG9b9 , \1363 );
and \U$2683 ( \3366 , \1400 , \2886_nG9f5 );
nand \U$2684 ( \3367 , \3008_nG9b9 , \1360 );
or \U$2685 ( \3368 , \1320 , \2886_nG9f5 );
nand \U$2686 ( \3369 , \3368 , \1404 );
and \U$2687 ( \3370 , \3367 , \3369 );
nor \U$2688 ( \3371 , \3365 , \3366 , \3370 );
and \U$2689 ( \3372 , \3364 , \3371 );
and \U$2690 ( \3373 , \3356 , \3363 );
or \U$2691 ( \3374 , \3372 , \3373 );
nand \U$2692 ( \3375 , \2034_nGfe1 , \2100 );
or \U$2693 ( \3376 , \1969 , \1787_nG10e2 );
nand \U$2694 ( \3377 , \3376 , \2286 );
and \U$2695 ( \3378 , \3375 , \3377 );
and \U$2696 ( \3379 , \2289 , \1787_nG10e2 );
and \U$2697 ( \3380 , \2034_nGfe1 , \2103 );
nor \U$2698 ( \3381 , \3378 , \3379 , \3380 );
and \U$2699 ( \3382 , \1632 , \2541 );
not \U$2700 ( \3383 , \1710_nG11c1 );
and \U$2701 ( \3384 , \2371 , \3383 );
and \U$2702 ( \3385 , \1631_nG12c9 , \2545 );
nor \U$2703 ( \3386 , \3382 , \3384 , \3385 );
xor \U$2704 ( \3387 , \3381 , \3386 );
nand \U$2705 ( \3388 , \2229_nGe35 , \1865 );
or \U$2706 ( \3389 , \1810 , \2156_nGf08 );
nand \U$2707 ( \3390 , \3389 , \1973 );
and \U$2708 ( \3391 , \3388 , \3390 );
and \U$2709 ( \3392 , \1976 , \2156_nGf08 );
and \U$2710 ( \3393 , \2229_nGe35 , \1868 );
nor \U$2711 ( \3394 , \3391 , \3392 , \3393 );
and \U$2712 ( \3395 , \3387 , \3394 );
and \U$2713 ( \3396 , \3381 , \3386 );
or \U$2714 ( \3397 , \3395 , \3396 );
xor \U$2715 ( \3398 , \3374 , \3397 );
xor \U$2716 ( \3399 , \3246 , \3274 );
xor \U$2717 ( \3400 , \3399 , \3282 );
and \U$2718 ( \3401 , \3398 , \3400 );
and \U$2719 ( \3402 , \3374 , \3397 );
or \U$2720 ( \3403 , \3401 , \3402 );
xor \U$2721 ( \3404 , \3152 , \3154 );
xor \U$2722 ( \3405 , \3404 , \3191 );
and \U$2723 ( \3406 , \3403 , \3405 );
and \U$2724 ( \3407 , \3346 , \3403 );
or \U$2725 ( \3408 , \3349 , \3406 , \3407 );
and \U$2726 ( \3409 , \3337 , \3408 );
and \U$2727 ( \3410 , \3331 , \3336 );
or \U$2728 ( \3411 , \3409 , \3410 );
xor \U$2729 ( \3412 , \3329 , \3411 );
nand \U$2730 ( \3413 , \2156_nGf08 , \2100 );
or \U$2731 ( \3414 , \1969 , \2034_nGfe1 );
nand \U$2732 ( \3415 , \3414 , \2286 );
and \U$2733 ( \3416 , \3413 , \3415 );
and \U$2734 ( \3417 , \2289 , \2034_nGfe1 );
and \U$2735 ( \3418 , \2156_nGf08 , \2103 );
nor \U$2736 ( \3419 , \3416 , \3417 , \3418 );
and \U$2737 ( \3420 , \3383 , \2541 );
not \U$2738 ( \3421 , \1787_nG10e2 );
and \U$2739 ( \3422 , \2371 , \3421 );
and \U$2740 ( \3423 , \1710_nG11c1 , \2545 );
nor \U$2741 ( \3424 , \3420 , \3422 , \3423 );
xor \U$2742 ( \3425 , \3419 , \3424 );
and \U$2743 ( \3426 , \3425 , \1266 );
and \U$2744 ( \3427 , \3419 , \3424 );
or \U$2745 ( \3428 , \3426 , \3427 );
and \U$2746 ( \3429 , \2653_nGa66 , \1653 );
or \U$2747 ( \3430 , \1579 , \2446_nGa9e );
nand \U$2748 ( \3431 , \3430 , \1799 );
nand \U$2749 ( \3432 , \2653_nGa66 , \1650 );
and \U$2750 ( \3433 , \3431 , \3432 );
and \U$2751 ( \3434 , \2446_nGa9e , \1794 );
nor \U$2752 ( \3435 , \3429 , \3433 , \3434 );
nand \U$2753 ( \3436 , \2404_nGad6 , \1865 );
or \U$2754 ( \3437 , \1810 , \2229_nGe35 );
nand \U$2755 ( \3438 , \3437 , \1973 );
and \U$2756 ( \3439 , \3436 , \3438 );
and \U$2757 ( \3440 , \1976 , \2229_nGe35 );
and \U$2758 ( \3441 , \2404_nGad6 , \1868 );
nor \U$2759 ( \3442 , \3439 , \3440 , \3441 );
xor \U$2760 ( \3443 , \3435 , \3442 );
nand \U$2761 ( \3444 , \2695_nGa2d , \1523 );
or \U$2762 ( \3445 , \1449 , \2886_nG9f5 );
nand \U$2763 ( \3446 , \3445 , \1529 );
and \U$2764 ( \3447 , \3444 , \3446 );
and \U$2765 ( \3448 , \1525 , \2886_nG9f5 );
and \U$2766 ( \3449 , \2695_nGa2d , \1594 );
nor \U$2767 ( \3450 , \3447 , \3448 , \3449 );
and \U$2768 ( \3451 , \3443 , \3450 );
and \U$2769 ( \3452 , \3435 , \3442 );
or \U$2770 ( \3453 , \3451 , \3452 );
xor \U$2771 ( \3454 , \3428 , \3453 );
and \U$2772 ( \3455 , \3182_nG984 , \1306 );
or \U$2773 ( \3456 , \1266 , \3273_nG944 );
nand \U$2774 ( \3457 , \3456 , \1303 );
nand \U$2775 ( \3458 , \3182_nG984 , \1299 );
and \U$2776 ( \3459 , \3457 , \3458 );
and \U$2777 ( \3460 , \3273_nG944 , \1440 );
nor \U$2778 ( \3461 , \3455 , \3459 , \3460 );
and \U$2779 ( \3462 , \3454 , \3461 );
and \U$2780 ( \3463 , \3428 , \3453 );
or \U$2781 ( \3464 , \3462 , \3463 );
not \U$2782 ( \3465 , \3339 );
not \U$2783 ( \3466 , \3345 );
and \U$2784 ( \3467 , \3465 , \3466 );
and \U$2785 ( \3468 , \3339 , \3345 );
nor \U$2786 ( \3469 , \3467 , \3468 );
xor \U$2787 ( \3470 , \3464 , \3469 );
xor \U$2788 ( \3471 , \3374 , \3397 );
xor \U$2789 ( \3472 , \3471 , \3400 );
and \U$2790 ( \3473 , \3470 , \3472 );
and \U$2791 ( \3474 , \3464 , \3469 );
or \U$2792 ( \3475 , \3473 , \3474 );
xor \U$2793 ( \3476 , \3225 , \3238 );
xor \U$2794 ( \3477 , \3476 , \3285 );
xor \U$2795 ( \3478 , \3475 , \3477 );
xor \U$2796 ( \3479 , \3152 , \3154 );
xor \U$2797 ( \3480 , \3479 , \3191 );
xor \U$2798 ( \3481 , \3346 , \3403 );
xor \U$2799 ( \3482 , \3480 , \3481 );
and \U$2800 ( \3483 , \3478 , \3482 );
and \U$2801 ( \3484 , \3475 , \3477 );
or \U$2802 ( \3485 , \3483 , \3484 );
xor \U$2803 ( \3486 , \3331 , \3336 );
xor \U$2804 ( \3487 , \3486 , \3408 );
and \U$2805 ( \3488 , \3485 , \3487 );
xor \U$2806 ( \3489 , \3428 , \3453 );
xor \U$2807 ( \3490 , \3489 , \3461 );
xor \U$2808 ( \3491 , \3381 , \3386 );
xor \U$2809 ( \3492 , \3491 , \3394 );
or \U$2810 ( \3493 , \3490 , \3492 );
and \U$2811 ( \3494 , \3182_nG984 , \1363 );
and \U$2812 ( \3495 , \1400 , \3008_nG9b9 );
nand \U$2813 ( \3496 , \3182_nG984 , \1360 );
or \U$2814 ( \3497 , \1320 , \3008_nG9b9 );
nand \U$2815 ( \3498 , \3497 , \1404 );
and \U$2816 ( \3499 , \3496 , \3498 );
nor \U$2817 ( \3500 , \3494 , \3495 , \3499 );
nand \U$2818 ( \3501 , \2229_nGe35 , \2100 );
or \U$2819 ( \3502 , \1969 , \2156_nGf08 );
nand \U$2820 ( \3503 , \3502 , \2286 );
and \U$2821 ( \3504 , \3501 , \3503 );
and \U$2822 ( \3505 , \2289 , \2156_nGf08 );
and \U$2823 ( \3506 , \2229_nGe35 , \2103 );
nor \U$2824 ( \3507 , \3504 , \3505 , \3506 );
and \U$2825 ( \3508 , \3421 , \2541 );
and \U$2826 ( \3509 , \2371 , \2257 );
and \U$2827 ( \3510 , \1787_nG10e2 , \2545 );
nor \U$2828 ( \3511 , \3508 , \3509 , \3510 );
xor \U$2829 ( \3512 , \3507 , \3511 );
nand \U$2830 ( \3513 , \2446_nGa9e , \1865 );
or \U$2831 ( \3514 , \1810 , \2404_nGad6 );
nand \U$2832 ( \3515 , \3514 , \1973 );
and \U$2833 ( \3516 , \3513 , \3515 );
and \U$2834 ( \3517 , \1976 , \2404_nGad6 );
and \U$2835 ( \3518 , \2446_nGa9e , \1868 );
nor \U$2836 ( \3519 , \3516 , \3517 , \3518 );
and \U$2837 ( \3520 , \3512 , \3519 );
and \U$2838 ( \3521 , \3507 , \3511 );
or \U$2839 ( \3522 , \3520 , \3521 );
xor \U$2840 ( \3523 , \3500 , \3522 );
nand \U$2841 ( \3524 , \2886_nG9f5 , \1523 );
or \U$2842 ( \3525 , \1449 , \3008_nG9b9 );
nand \U$2843 ( \3526 , \3525 , \1529 );
and \U$2844 ( \3527 , \3524 , \3526 );
and \U$2845 ( \3528 , \1525 , \3008_nG9b9 );
and \U$2846 ( \3529 , \2886_nG9f5 , \1594 );
nor \U$2847 ( \3530 , \3527 , \3528 , \3529 );
and \U$2848 ( \3531 , \2695_nGa2d , \1653 );
or \U$2849 ( \3532 , \1579 , \2653_nGa66 );
nand \U$2850 ( \3533 , \3532 , \1799 );
nand \U$2851 ( \3534 , \2695_nGa2d , \1650 );
and \U$2852 ( \3535 , \3533 , \3534 );
and \U$2853 ( \3536 , \2653_nGa66 , \1794 );
nor \U$2854 ( \3537 , \3531 , \3535 , \3536 );
xor \U$2855 ( \3538 , \3530 , \3537 );
and \U$2856 ( \3539 , \3273_nG944 , \1363 );
and \U$2857 ( \3540 , \1400 , \3182_nG984 );
nand \U$2858 ( \3541 , \3273_nG944 , \1360 );
or \U$2859 ( \3542 , \1320 , \3182_nG984 );
nand \U$2860 ( \3543 , \3542 , \1404 );
and \U$2861 ( \3544 , \3541 , \3543 );
nor \U$2862 ( \3545 , \3539 , \3540 , \3544 );
and \U$2863 ( \3546 , \3538 , \3545 );
and \U$2864 ( \3547 , \3530 , \3537 );
or \U$2865 ( \3548 , \3546 , \3547 );
and \U$2866 ( \3549 , \3523 , \3548 );
and \U$2867 ( \3550 , \3500 , \3522 );
or \U$2868 ( \3551 , \3549 , \3550 );
xor \U$2869 ( \3552 , \3356 , \3363 );
xor \U$2870 ( \3553 , \3552 , \3371 );
xor \U$2871 ( \3554 , \3551 , \3553 );
xor \U$2872 ( \3555 , \3435 , \3442 );
xor \U$2873 ( \3556 , \3555 , \3450 );
xor \U$2874 ( \3557 , \3419 , \3424 );
xor \U$2875 ( \3558 , \3557 , \1266 );
and \U$2876 ( \3559 , \3556 , \3558 );
nand \U$2877 ( \3560 , \3273_nG944 , \1299 );
and \U$2878 ( \3561 , \1265 , \3560 );
and \U$2879 ( \3562 , \3273_nG944 , \1306 );
nor \U$2880 ( \3563 , \3561 , \3562 );
xor \U$2881 ( \3564 , \3419 , \3424 );
xor \U$2882 ( \3565 , \3564 , \1266 );
and \U$2883 ( \3566 , \3563 , \3565 );
and \U$2884 ( \3567 , \3556 , \3563 );
or \U$2885 ( \3568 , \3559 , \3566 , \3567 );
and \U$2886 ( \3569 , \3554 , \3568 );
and \U$2887 ( \3570 , \3551 , \3553 );
or \U$2888 ( \3571 , \3569 , \3570 );
xor \U$2889 ( \3572 , \3493 , \3571 );
xor \U$2890 ( \3573 , \3464 , \3469 );
xor \U$2891 ( \3574 , \3573 , \3472 );
and \U$2892 ( \3575 , \3572 , \3574 );
and \U$2893 ( \3576 , \3493 , \3571 );
or \U$2894 ( \3577 , \3575 , \3576 );
xor \U$2895 ( \3578 , \3475 , \3477 );
xor \U$2896 ( \3579 , \3578 , \3482 );
and \U$2897 ( \3580 , \3577 , \3579 );
and \U$2898 ( \3581 , \2886_nG9f5 , \1653 );
or \U$2899 ( \3582 , \1579 , \2695_nGa2d );
nand \U$2900 ( \3583 , \3582 , \1799 );
nand \U$2901 ( \3584 , \2886_nG9f5 , \1650 );
and \U$2902 ( \3585 , \3583 , \3584 );
and \U$2903 ( \3586 , \2695_nGa2d , \1794 );
nor \U$2904 ( \3587 , \3581 , \3585 , \3586 );
nand \U$2905 ( \3588 , \2653_nGa66 , \1865 );
or \U$2906 ( \3589 , \1810 , \2446_nGa9e );
nand \U$2907 ( \3590 , \3589 , \1973 );
and \U$2908 ( \3591 , \3588 , \3590 );
and \U$2909 ( \3592 , \1976 , \2446_nGa9e );
and \U$2910 ( \3593 , \2653_nGa66 , \1868 );
nor \U$2911 ( \3594 , \3591 , \3592 , \3593 );
xor \U$2912 ( \3595 , \3587 , \3594 );
nand \U$2913 ( \3596 , \3008_nG9b9 , \1523 );
or \U$2914 ( \3597 , \1449 , \3182_nG984 );
nand \U$2915 ( \3598 , \3597 , \1529 );
and \U$2916 ( \3599 , \3596 , \3598 );
and \U$2917 ( \3600 , \1525 , \3182_nG984 );
and \U$2918 ( \3601 , \3008_nG9b9 , \1594 );
nor \U$2919 ( \3602 , \3599 , \3600 , \3601 );
and \U$2920 ( \3603 , \3595 , \3602 );
and \U$2921 ( \3604 , \3587 , \3594 );
or \U$2922 ( \3605 , \3603 , \3604 );
nand \U$2923 ( \3606 , \2404_nGad6 , \2100 );
or \U$2924 ( \3607 , \1969 , \2229_nGe35 );
nand \U$2925 ( \3608 , \3607 , \2286 );
and \U$2926 ( \3609 , \3606 , \3608 );
and \U$2927 ( \3610 , \2289 , \2229_nGe35 );
and \U$2928 ( \3611 , \2404_nGad6 , \2103 );
nor \U$2929 ( \3612 , \3609 , \3610 , \3611 );
and \U$2930 ( \3613 , \2257 , \2541 );
not \U$2931 ( \3614 , \2156_nGf08 );
and \U$2932 ( \3615 , \2371 , \3614 );
and \U$2933 ( \3616 , \2034_nGfe1 , \2545 );
nor \U$2934 ( \3617 , \3613 , \3615 , \3616 );
xor \U$2935 ( \3618 , \3612 , \3617 );
and \U$2936 ( \3619 , \3618 , \1320 );
and \U$2937 ( \3620 , \3612 , \3617 );
or \U$2938 ( \3621 , \3619 , \3620 );
xor \U$2939 ( \3622 , \3605 , \3621 );
xor \U$2940 ( \3623 , \3530 , \3537 );
xor \U$2941 ( \3624 , \3623 , \3545 );
and \U$2942 ( \3625 , \3622 , \3624 );
and \U$2943 ( \3626 , \3605 , \3621 );
or \U$2944 ( \3627 , \3625 , \3626 );
xor \U$2945 ( \3628 , \3500 , \3522 );
xor \U$2946 ( \3629 , \3628 , \3548 );
xor \U$2947 ( \3630 , \3627 , \3629 );
xor \U$2948 ( \3631 , \3419 , \3424 );
xor \U$2949 ( \3632 , \3631 , \1266 );
xor \U$2950 ( \3633 , \3556 , \3563 );
xor \U$2951 ( \3634 , \3632 , \3633 );
and \U$2952 ( \3635 , \3630 , \3634 );
and \U$2953 ( \3636 , \3627 , \3629 );
or \U$2954 ( \3637 , \3635 , \3636 );
xor \U$2955 ( \3638 , \3551 , \3553 );
xor \U$2956 ( \3639 , \3638 , \3568 );
xor \U$2957 ( \3640 , \3637 , \3639 );
xnor \U$2958 ( \3641 , \3492 , \3490 );
xor \U$2959 ( \3642 , \3640 , \3641 );
not \U$2960 ( \3643 , \3642 );
xor \U$2961 ( \3644 , \3627 , \3629 );
xor \U$2962 ( \3645 , \3644 , \3634 );
nand \U$2963 ( \3646 , \2446_nGa9e , \2100 );
or \U$2964 ( \3647 , \1969 , \2404_nGad6 );
nand \U$2965 ( \3648 , \3647 , \2286 );
and \U$2966 ( \3649 , \3646 , \3648 );
and \U$2967 ( \3650 , \2289 , \2404_nGad6 );
and \U$2968 ( \3651 , \2446_nGa9e , \2103 );
nor \U$2969 ( \3652 , \3649 , \3650 , \3651 );
and \U$2970 ( \3653 , \3614 , \2541 );
not \U$2971 ( \3654 , \2229_nGe35 );
and \U$2972 ( \3655 , \2371 , \3654 );
and \U$2973 ( \3656 , \2156_nGf08 , \2545 );
nor \U$2974 ( \3657 , \3653 , \3655 , \3656 );
xor \U$2975 ( \3658 , \3652 , \3657 );
nand \U$2976 ( \3659 , \2695_nGa2d , \1865 );
or \U$2977 ( \3660 , \1810 , \2653_nGa66 );
nand \U$2978 ( \3661 , \3660 , \1973 );
and \U$2979 ( \3662 , \3659 , \3661 );
and \U$2980 ( \3663 , \1976 , \2653_nGa66 );
and \U$2981 ( \3664 , \2695_nGa2d , \1868 );
nor \U$2982 ( \3665 , \3662 , \3663 , \3664 );
and \U$2983 ( \3666 , \3658 , \3665 );
and \U$2984 ( \3667 , \3652 , \3657 );
or \U$2985 ( \3668 , \3666 , \3667 );
xor \U$2986 ( \3669 , \3587 , \3594 );
xor \U$2987 ( \3670 , \3669 , \3602 );
and \U$2988 ( \3671 , \3668 , \3670 );
and \U$2989 ( \3672 , \3273_nG944 , \1400 );
not \U$2990 ( \3673 , \3273_nG944 );
and \U$2991 ( \3674 , \3673 , \1362 );
not \U$2992 ( \3675 , \1404 );
nor \U$2993 ( \3676 , \3672 , \3674 , \3675 );
xor \U$2994 ( \3677 , \3587 , \3594 );
xor \U$2995 ( \3678 , \3677 , \3602 );
and \U$2996 ( \3679 , \3676 , \3678 );
and \U$2997 ( \3680 , \3668 , \3676 );
or \U$2998 ( \3681 , \3671 , \3679 , \3680 );
xor \U$2999 ( \3682 , \3507 , \3511 );
xor \U$3000 ( \3683 , \3682 , \3519 );
xor \U$3001 ( \3684 , \3681 , \3683 );
xor \U$3002 ( \3685 , \3605 , \3621 );
xor \U$3003 ( \3686 , \3685 , \3624 );
and \U$3004 ( \3687 , \3684 , \3686 );
and \U$3005 ( \3688 , \3681 , \3683 );
or \U$3006 ( \3689 , \3687 , \3688 );
nor \U$3007 ( \3690 , \3645 , \3689 );
xor \U$3008 ( \3691 , \3643 , \3690 );
and \U$3009 ( \3692 , \3645 , \3689 );
nor \U$3010 ( \3693 , \3692 , \3690 );
xor \U$3011 ( \3694 , \3681 , \3683 );
xor \U$3012 ( \3695 , \3694 , \3686 );
xor \U$3013 ( \3696 , \3612 , \3617 );
xor \U$3014 ( \3697 , \3696 , \1320 );
nand \U$3015 ( \3698 , \2653_nGa66 , \2100 );
or \U$3016 ( \3699 , \1969 , \2446_nGa9e );
nand \U$3017 ( \3700 , \3699 , \2286 );
and \U$3018 ( \3701 , \3698 , \3700 );
and \U$3019 ( \3702 , \2289 , \2446_nGa9e );
and \U$3020 ( \3703 , \2653_nGa66 , \2103 );
nor \U$3021 ( \3704 , \3701 , \3702 , \3703 );
and \U$3022 ( \3705 , \3654 , \2541 );
not \U$3023 ( \3706 , \2404_nGad6 );
and \U$3024 ( \3707 , \2371 , \3706 );
and \U$3025 ( \3708 , \2229_nGe35 , \2545 );
nor \U$3026 ( \3709 , \3705 , \3707 , \3708 );
xor \U$3027 ( \3710 , \3704 , \3709 );
and \U$3028 ( \3711 , \3710 , \1449 );
and \U$3029 ( \3712 , \3704 , \3709 );
or \U$3030 ( \3713 , \3711 , \3712 );
and \U$3031 ( \3714 , \3008_nG9b9 , \1653 );
or \U$3032 ( \3715 , \1579 , \2886_nG9f5 );
nand \U$3033 ( \3716 , \3715 , \1799 );
nand \U$3034 ( \3717 , \3008_nG9b9 , \1650 );
and \U$3035 ( \3718 , \3716 , \3717 );
and \U$3036 ( \3719 , \2886_nG9f5 , \1794 );
nor \U$3037 ( \3720 , \3714 , \3718 , \3719 );
xor \U$3038 ( \3721 , \3713 , \3720 );
and \U$3039 ( \3722 , \3182_nG984 , \1653 );
or \U$3040 ( \3723 , \1579 , \3008_nG9b9 );
nand \U$3041 ( \3724 , \3723 , \1799 );
nand \U$3042 ( \3725 , \3182_nG984 , \1650 );
and \U$3043 ( \3726 , \3724 , \3725 );
and \U$3044 ( \3727 , \3008_nG9b9 , \1794 );
nor \U$3045 ( \3728 , \3722 , \3726 , \3727 );
nand \U$3046 ( \3729 , \2886_nG9f5 , \1865 );
or \U$3047 ( \3730 , \1810 , \2695_nGa2d );
nand \U$3048 ( \3731 , \3730 , \1973 );
and \U$3049 ( \3732 , \3729 , \3731 );
and \U$3050 ( \3733 , \1976 , \2695_nGa2d );
and \U$3051 ( \3734 , \2886_nG9f5 , \1868 );
nor \U$3052 ( \3735 , \3732 , \3733 , \3734 );
xor \U$3053 ( \3736 , \3728 , \3735 );
and \U$3054 ( \3737 , \1594 , \3273_nG944 );
nand \U$3055 ( \3738 , \3273_nG944 , \1523 );
and \U$3056 ( \3739 , \3738 , \1527 );
nor \U$3057 ( \3740 , \3737 , \3739 );
and \U$3058 ( \3741 , \3736 , \3740 );
and \U$3059 ( \3742 , \3728 , \3735 );
or \U$3060 ( \3743 , \3741 , \3742 );
and \U$3061 ( \3744 , \3721 , \3743 );
and \U$3062 ( \3745 , \3713 , \3720 );
or \U$3063 ( \3746 , \3744 , \3745 );
nand \U$3064 ( \3747 , \3697 , \3746 );
not \U$3065 ( \3748 , \3182_nG984 );
or \U$3066 ( \3749 , \1659 , \3748 );
or \U$3067 ( \3750 , \3673 , \1661 );
or \U$3068 ( \3751 , \1593 , \3748 );
or \U$3069 ( \3752 , \1449 , \3273_nG944 );
nand \U$3070 ( \3753 , \3752 , \1529 );
nand \U$3071 ( \3754 , \3751 , \3753 );
nand \U$3072 ( \3755 , \3749 , \3750 , \3754 );
not \U$3073 ( \3756 , \3755 );
xor \U$3074 ( \3757 , \3652 , \3657 );
xor \U$3075 ( \3758 , \3757 , \3665 );
nor \U$3076 ( \3759 , \3756 , \3758 );
and \U$3077 ( \3760 , \3747 , \3759 );
nor \U$3078 ( \3761 , \3746 , \3697 );
nor \U$3079 ( \3762 , \3760 , \3761 );
nor \U$3080 ( \3763 , \3695 , \3762 );
xor \U$3081 ( \3764 , \3693 , \3763 );
not \U$3082 ( \3765 , \3759 );
not \U$3083 ( \3766 , \3761 );
nand \U$3084 ( \3767 , \3766 , \3747 );
not \U$3085 ( \3768 , \3767 );
or \U$3086 ( \3769 , \3765 , \3768 );
or \U$3087 ( \3770 , \3767 , \3759 );
nand \U$3088 ( \3771 , \3769 , \3770 );
xor \U$3089 ( \3772 , \3587 , \3594 );
xor \U$3090 ( \3773 , \3772 , \3602 );
xor \U$3091 ( \3774 , \3668 , \3676 );
xor \U$3092 ( \3775 , \3773 , \3774 );
not \U$3093 ( \3776 , \3775 );
xor \U$3094 ( \3777 , \3771 , \3776 );
not \U$3095 ( \3778 , \3755 );
not \U$3096 ( \3779 , \3758 );
and \U$3097 ( \3780 , \3778 , \3779 );
and \U$3098 ( \3781 , \3755 , \3758 );
nor \U$3099 ( \3782 , \3780 , \3781 );
not \U$3100 ( \3783 , \3782 );
xor \U$3101 ( \3784 , \3713 , \3720 );
xor \U$3102 ( \3785 , \3784 , \3743 );
nand \U$3103 ( \3786 , \2695_nGa2d , \2100 );
or \U$3104 ( \3787 , \1969 , \2653_nGa66 );
nand \U$3105 ( \3788 , \3787 , \2286 );
and \U$3106 ( \3789 , \3786 , \3788 );
and \U$3107 ( \3790 , \2289 , \2653_nGa66 );
and \U$3108 ( \3791 , \2695_nGa2d , \2103 );
nor \U$3109 ( \3792 , \3789 , \3790 , \3791 );
not \U$3110 ( \3793 , \3792 );
and \U$3111 ( \3794 , \3706 , \2541 );
not \U$3112 ( \3795 , \2446_nGa9e );
and \U$3113 ( \3796 , \2371 , \3795 );
and \U$3114 ( \3797 , \2404_nGad6 , \2545 );
nor \U$3115 ( \3798 , \3794 , \3796 , \3797 );
not \U$3116 ( \3799 , \3798 );
and \U$3117 ( \3800 , \3793 , \3799 );
and \U$3118 ( \3801 , \3792 , \3798 );
nand \U$3119 ( \3802 , \3008_nG9b9 , \1865 );
or \U$3120 ( \3803 , \1810 , \2886_nG9f5 );
nand \U$3121 ( \3804 , \3803 , \1973 );
and \U$3122 ( \3805 , \3802 , \3804 );
and \U$3123 ( \3806 , \1976 , \2886_nG9f5 );
and \U$3124 ( \3807 , \3008_nG9b9 , \1868 );
nor \U$3125 ( \3808 , \3805 , \3806 , \3807 );
nor \U$3126 ( \3809 , \3801 , \3808 );
nor \U$3127 ( \3810 , \3800 , \3809 );
xor \U$3128 ( \3811 , \3704 , \3709 );
xor \U$3129 ( \3812 , \3811 , \1449 );
and \U$3130 ( \3813 , \3810 , \3812 );
xor \U$3131 ( \3814 , \3728 , \3735 );
xor \U$3132 ( \3815 , \3814 , \3740 );
xor \U$3133 ( \3816 , \3704 , \3709 );
xor \U$3134 ( \3817 , \3816 , \1449 );
and \U$3135 ( \3818 , \3815 , \3817 );
and \U$3136 ( \3819 , \3810 , \3815 );
or \U$3137 ( \3820 , \3813 , \3818 , \3819 );
or \U$3138 ( \3821 , \3785 , \3820 );
not \U$3139 ( \3822 , \3821 );
or \U$3140 ( \3823 , \3783 , \3822 );
nand \U$3141 ( \3824 , \3820 , \3785 );
nand \U$3142 ( \3825 , \3823 , \3824 );
not \U$3143 ( \3826 , \3825 );
xor \U$3144 ( \3827 , \3777 , \3826 );
nand \U$3145 ( \3828 , \3821 , \3824 );
not \U$3146 ( \3829 , \3828 );
not \U$3147 ( \3830 , \3782 );
and \U$3148 ( \3831 , \3829 , \3830 );
and \U$3149 ( \3832 , \3828 , \3782 );
nor \U$3150 ( \3833 , \3831 , \3832 );
xor \U$3151 ( \3834 , \3704 , \3709 );
xor \U$3152 ( \3835 , \3834 , \1449 );
xor \U$3153 ( \3836 , \3810 , \3815 );
xor \U$3154 ( \3837 , \3835 , \3836 );
or \U$3155 ( \3838 , \1795 , \3673 );
or \U$3156 ( \3839 , \3273_nG944 , \1579 );
nand \U$3157 ( \3840 , \3838 , \3839 , \1799 );
not \U$3158 ( \3841 , \3840 );
nand \U$3159 ( \3842 , \3182_nG984 , \1865 );
or \U$3160 ( \3843 , \1810 , \3008_nG9b9 );
nand \U$3161 ( \3844 , \3843 , \1973 );
and \U$3162 ( \3845 , \3842 , \3844 );
and \U$3163 ( \3846 , \1976 , \3008_nG9b9 );
and \U$3164 ( \3847 , \3182_nG984 , \1868 );
nor \U$3165 ( \3848 , \3845 , \3846 , \3847 );
nor \U$3166 ( \3849 , \3841 , \3848 );
nand \U$3167 ( \3850 , \2886_nG9f5 , \2100 );
or \U$3168 ( \3851 , \1969 , \2695_nGa2d );
nand \U$3169 ( \3852 , \3851 , \2286 );
and \U$3170 ( \3853 , \3850 , \3852 );
and \U$3171 ( \3854 , \2289 , \2695_nGa2d );
and \U$3172 ( \3855 , \2886_nG9f5 , \2103 );
nor \U$3173 ( \3856 , \3853 , \3854 , \3855 );
and \U$3174 ( \3857 , \3795 , \2541 );
not \U$3175 ( \3858 , \2653_nGa66 );
and \U$3176 ( \3859 , \2371 , \3858 );
and \U$3177 ( \3860 , \2446_nGa9e , \2545 );
nor \U$3178 ( \3861 , \3857 , \3859 , \3860 );
xor \U$3179 ( \3862 , \3856 , \3861 );
and \U$3180 ( \3863 , \3862 , \1579 );
and \U$3181 ( \3864 , \3856 , \3861 );
or \U$3182 ( \3865 , \3863 , \3864 );
and \U$3183 ( \3866 , \3273_nG944 , \1653 );
or \U$3184 ( \3867 , \1579 , \3182_nG984 );
nand \U$3185 ( \3868 , \3867 , \1799 );
nand \U$3186 ( \3869 , \3273_nG944 , \1650 );
and \U$3187 ( \3870 , \3868 , \3869 );
and \U$3188 ( \3871 , \3182_nG984 , \1794 );
nor \U$3189 ( \3872 , \3866 , \3870 , \3871 );
nand \U$3190 ( \3873 , \3865 , \3872 );
and \U$3191 ( \3874 , \3849 , \3873 );
nor \U$3192 ( \3875 , \3872 , \3865 );
nor \U$3193 ( \3876 , \3874 , \3875 );
nor \U$3194 ( \3877 , \3837 , \3876 );
xor \U$3195 ( \3878 , \3833 , \3877 );
not \U$3196 ( \3879 , \3792 );
xor \U$3197 ( \3880 , \3798 , \3808 );
not \U$3198 ( \3881 , \3880 );
or \U$3199 ( \3882 , \3879 , \3881 );
or \U$3200 ( \3883 , \3880 , \3792 );
nand \U$3201 ( \3884 , \3882 , \3883 );
not \U$3202 ( \3885 , \3849 );
not \U$3203 ( \3886 , \3875 );
nand \U$3204 ( \3887 , \3886 , \3873 );
not \U$3205 ( \3888 , \3887 );
or \U$3206 ( \3889 , \3885 , \3888 );
or \U$3207 ( \3890 , \3887 , \3849 );
nand \U$3208 ( \3891 , \3889 , \3890 );
xor \U$3209 ( \3892 , \3884 , \3891 );
not \U$3210 ( \3893 , \3840 );
not \U$3211 ( \3894 , \3848 );
and \U$3212 ( \3895 , \3893 , \3894 );
and \U$3213 ( \3896 , \3840 , \3848 );
nor \U$3214 ( \3897 , \3895 , \3896 );
xor \U$3215 ( \3898 , \3856 , \3861 );
xor \U$3216 ( \3899 , \3898 , \1579 );
nand \U$3217 ( \3900 , \3008_nG9b9 , \2100 );
or \U$3218 ( \3901 , \1969 , \2886_nG9f5 );
nand \U$3219 ( \3902 , \3901 , \2286 );
and \U$3220 ( \3903 , \3900 , \3902 );
and \U$3221 ( \3904 , \2289 , \2886_nG9f5 );
and \U$3222 ( \3905 , \3008_nG9b9 , \2103 );
nor \U$3223 ( \3906 , \3903 , \3904 , \3905 );
not \U$3224 ( \3907 , \3906 );
and \U$3225 ( \3908 , \3858 , \2541 );
not \U$3226 ( \3909 , \2695_nGa2d );
and \U$3227 ( \3910 , \2371 , \3909 );
and \U$3228 ( \3911 , \2653_nGa66 , \2545 );
nor \U$3229 ( \3912 , \3908 , \3910 , \3911 );
not \U$3230 ( \3913 , \3912 );
and \U$3231 ( \3914 , \3907 , \3913 );
and \U$3232 ( \3915 , \3906 , \3912 );
nand \U$3233 ( \3916 , \3273_nG944 , \1865 );
or \U$3234 ( \3917 , \1810 , \3182_nG984 );
nand \U$3235 ( \3918 , \3917 , \1973 );
and \U$3236 ( \3919 , \3916 , \3918 );
and \U$3237 ( \3920 , \1976 , \3182_nG984 );
and \U$3238 ( \3921 , \3273_nG944 , \1868 );
nor \U$3239 ( \3922 , \3919 , \3920 , \3921 );
nor \U$3240 ( \3923 , \3915 , \3922 );
nor \U$3241 ( \3924 , \3914 , \3923 );
or \U$3242 ( \3925 , \3899 , \3924 );
and \U$3243 ( \3926 , \3897 , \3925 );
and \U$3244 ( \3927 , \3924 , \3899 );
nor \U$3245 ( \3928 , \3926 , \3927 );
xor \U$3246 ( \3929 , \3892 , \3928 );
xor \U$3247 ( \3930 , \3899 , \3924 );
and \U$3248 ( \3931 , \3897 , \3930 );
nor \U$3249 ( \3932 , \3897 , \3930 );
or \U$3250 ( \3933 , \2544 , \3909 );
or \U$3251 ( \3934 , \2695_nGa2d , \2373 );
or \U$3252 ( \3935 , \2886_nG9f5 , \2372 );
nand \U$3253 ( \3936 , \3933 , \3934 , \3935 );
nor \U$3254 ( \3937 , \1867 , \3936 );
nand \U$3255 ( \3938 , \3182_nG984 , \2100 );
or \U$3256 ( \3939 , \1969 , \3008_nG9b9 );
nand \U$3257 ( \3940 , \3939 , \2286 );
and \U$3258 ( \3941 , \3938 , \3940 );
and \U$3259 ( \3942 , \2289 , \3008_nG9b9 );
and \U$3260 ( \3943 , \3182_nG984 , \2103 );
nor \U$3261 ( \3944 , \3941 , \3942 , \3943 );
or \U$3262 ( \3945 , \3937 , \3944 );
nand \U$3263 ( \3946 , \3936 , \1867 );
nand \U$3264 ( \3947 , \3945 , \3946 );
not \U$3265 ( \3948 , \3906 );
xor \U$3266 ( \3949 , \3912 , \3922 );
not \U$3267 ( \3950 , \3949 );
or \U$3268 ( \3951 , \3948 , \3950 );
or \U$3269 ( \3952 , \3949 , \3906 );
nand \U$3270 ( \3953 , \3951 , \3952 );
and \U$3271 ( \3954 , \3947 , \3953 );
nor \U$3272 ( \3955 , \3931 , \3932 , \3954 );
xor \U$3273 ( \3956 , \3947 , \3953 );
not \U$3274 ( \3957 , \1976 );
or \U$3275 ( \3958 , \3957 , \3673 );
or \U$3276 ( \3959 , \3273_nG944 , \1810 );
nand \U$3277 ( \3960 , \3958 , \3959 , \1973 );
not \U$3278 ( \3961 , \3960 );
not \U$3279 ( \3962 , \3946 );
nor \U$3280 ( \3963 , \3962 , \3937 );
not \U$3281 ( \3964 , \3963 );
not \U$3282 ( \3965 , \3944 );
and \U$3283 ( \3966 , \3964 , \3965 );
and \U$3284 ( \3967 , \3963 , \3944 );
nor \U$3285 ( \3968 , \3966 , \3967 );
nor \U$3286 ( \3969 , \3961 , \3968 );
and \U$3287 ( \3970 , \3956 , \3969 );
and \U$3288 ( \3971 , \2370 , \3182_nG984 );
nor \U$3289 ( \3972 , \3971 , \1963 , \3273_nG944 );
not \U$3290 ( \3973 , \3972 );
not \U$3291 ( \3974 , \2289 );
or \U$3292 ( \3975 , \3974 , \3673 );
or \U$3293 ( \3976 , \3273_nG944 , \1969 );
nand \U$3294 ( \3977 , \3975 , \3976 , \2286 );
not \U$3295 ( \3978 , \3977 );
or \U$3296 ( \3979 , \3973 , \3978 );
or \U$3297 ( \3980 , \3977 , \3972 );
not \U$3298 ( \3981 , \3008_nG9b9 );
or \U$3299 ( \3982 , \2544 , \3981 );
or \U$3300 ( \3983 , \3008_nG9b9 , \2373 );
or \U$3301 ( \3984 , \3182_nG984 , \2372 );
nand \U$3302 ( \3985 , \3982 , \3983 , \3984 );
xor \U$3303 ( \3986 , \3985 , \2102 );
nand \U$3304 ( \3987 , \3980 , \3986 );
nand \U$3305 ( \3988 , \3979 , \3987 );
and \U$3306 ( \3989 , \3985 , \2102 );
and \U$3307 ( \3990 , \3988 , \3989 );
not \U$3308 ( \3991 , \3960 );
not \U$3309 ( \3992 , \3968 );
and \U$3310 ( \3993 , \3991 , \3992 );
and \U$3311 ( \3994 , \3960 , \3968 );
nor \U$3312 ( \3995 , \3993 , \3994 );
not \U$3313 ( \3996 , \3995 );
nor \U$3314 ( \3997 , \3990 , \3996 );
nand \U$3315 ( \3998 , \3273_nG944 , \2100 );
or \U$3316 ( \3999 , \1969 , \3182_nG984 );
nand \U$3317 ( \4000 , \3999 , \2286 );
and \U$3318 ( \4001 , \3998 , \4000 );
and \U$3319 ( \4002 , \2289 , \3182_nG984 );
and \U$3320 ( \4003 , \3273_nG944 , \2103 );
nor \U$3321 ( \4004 , \4001 , \4002 , \4003 );
not \U$3322 ( \4005 , \2886_nG9f5 );
and \U$3323 ( \4006 , \4005 , \2541 );
and \U$3324 ( \4007 , \2371 , \3981 );
and \U$3325 ( \4008 , \2886_nG9f5 , \2545 );
nor \U$3326 ( \4009 , \4006 , \4007 , \4008 );
or \U$3327 ( \4010 , \3997 , \4004 , \4009 );
nand \U$3328 ( \4011 , \4009 , \4004 );
or \U$3329 ( \4012 , \4011 , \3989 );
and \U$3330 ( \4013 , \4012 , \3988 );
and \U$3331 ( \4014 , \3989 , \4011 );
nor \U$3332 ( \4015 , \4013 , \4014 );
or \U$3333 ( \4016 , \3995 , \4015 );
nand \U$3334 ( \4017 , \4010 , \4016 );
or \U$3335 ( \4018 , \3956 , \3969 );
and \U$3336 ( \4019 , \4017 , \4018 );
nor \U$3337 ( \4020 , \3970 , \4019 );
or \U$3338 ( \4021 , \3955 , \4020 );
or \U$3339 ( \4022 , \3931 , \3932 );
nand \U$3340 ( \4023 , \4022 , \3954 );
nand \U$3341 ( \4024 , \4021 , \4023 );
and \U$3342 ( \4025 , \3929 , \4024 );
and \U$3343 ( \4026 , \3892 , \3928 );
or \U$3344 ( \4027 , \4025 , \4026 );
and \U$3345 ( \4028 , \3884 , \3891 );
xor \U$3346 ( \4029 , \4027 , \4028 );
and \U$3347 ( \4030 , \3837 , \3876 );
nor \U$3348 ( \4031 , \4030 , \3877 );
and \U$3349 ( \4032 , \4029 , \4031 );
and \U$3350 ( \4033 , \4027 , \4028 );
or \U$3351 ( \4034 , \4032 , \4033 );
and \U$3352 ( \4035 , \3878 , \4034 );
and \U$3353 ( \4036 , \3833 , \3877 );
or \U$3354 ( \4037 , \4035 , \4036 );
and \U$3355 ( \4038 , \3827 , \4037 );
and \U$3356 ( \4039 , \3777 , \3826 );
or \U$3357 ( \4040 , \4038 , \4039 );
and \U$3358 ( \4041 , \3771 , \3776 );
xor \U$3359 ( \4042 , \4040 , \4041 );
and \U$3360 ( \4043 , \3695 , \3762 );
nor \U$3361 ( \4044 , \4043 , \3763 );
and \U$3362 ( \4045 , \4042 , \4044 );
and \U$3363 ( \4046 , \4040 , \4041 );
or \U$3364 ( \4047 , \4045 , \4046 );
and \U$3365 ( \4048 , \3764 , \4047 );
and \U$3366 ( \4049 , \3693 , \3763 );
or \U$3367 ( \4050 , \4048 , \4049 );
and \U$3368 ( \4051 , \3691 , \4050 );
and \U$3369 ( \4052 , \3643 , \3690 );
or \U$3370 ( \4053 , \4051 , \4052 );
xor \U$3371 ( \4054 , \3637 , \3639 );
and \U$3372 ( \4055 , \4054 , \3641 );
and \U$3373 ( \4056 , \3637 , \3639 );
or \U$3374 ( \4057 , \4055 , \4056 );
xor \U$3375 ( \4058 , \3493 , \3571 );
xor \U$3376 ( \4059 , \4058 , \3574 );
nand \U$3377 ( \4060 , \4057 , \4059 );
and \U$3378 ( \4061 , \4053 , \4060 );
nor \U$3379 ( \4062 , \4059 , \4057 );
nor \U$3380 ( \4063 , \4061 , \4062 );
xor \U$3381 ( \4064 , \3475 , \3477 );
xor \U$3382 ( \4065 , \4064 , \3482 );
and \U$3383 ( \4066 , \4063 , \4065 );
and \U$3384 ( \4067 , \3577 , \4063 );
or \U$3385 ( \4068 , \3580 , \4066 , \4067 );
xor \U$3386 ( \4069 , \3331 , \3336 );
xor \U$3387 ( \4070 , \4069 , \3408 );
and \U$3388 ( \4071 , \4068 , \4070 );
and \U$3389 ( \4072 , \3485 , \4068 );
or \U$3390 ( \4073 , \3488 , \4071 , \4072 );
and \U$3391 ( \4074 , \3412 , \4073 );
and \U$3392 ( \4075 , \3329 , \3411 );
or \U$3393 ( \4076 , \4074 , \4075 );
not \U$3394 ( \4077 , \4076 );
and \U$3395 ( \4078 , \3327 , \4077 );
and \U$3396 ( \4079 , \3316 , \3326 );
or \U$3397 ( \4080 , \4078 , \4079 );
and \U$3398 ( \4081 , \3314 , \4080 );
and \U$3399 ( \4082 , \3143 , \3313 );
or \U$3400 ( \4083 , \4081 , \4082 );
xor \U$3401 ( \4084 , \3126 , \3131 );
and \U$3402 ( \4085 , \4084 , \3142 );
and \U$3403 ( \4086 , \3126 , \3131 );
or \U$3404 ( \4087 , \4085 , \4086 );
not \U$3405 ( \4088 , \4087 );
xor \U$3406 ( \4089 , \3021 , \3035 );
xor \U$3407 ( \4090 , \4089 , \3046 );
nand \U$3408 ( \4091 , \4088 , \4090 );
and \U$3409 ( \4092 , \4083 , \4091 );
not \U$3410 ( \4093 , \4087 );
nor \U$3411 ( \4094 , \4093 , \4090 );
nor \U$3412 ( \4095 , \4092 , \4094 );
and \U$3413 ( \4096 , \3050 , \4095 );
and \U$3414 ( \4097 , \2855 , \3049 );
or \U$3415 ( \4098 , \4096 , \4097 );
not \U$3416 ( \4099 , \4098 );
and \U$3417 ( \4100 , \2848 , \4099 );
and \U$3418 ( \4101 , \2767 , \2847 );
or \U$3419 ( \4102 , \4100 , \4101 );
xor \U$3420 ( \4103 , \2498 , \2581 );
xor \U$3421 ( \4104 , \4103 , \2584 );
or \U$3422 ( \4105 , \2756 , \2763 );
nand \U$3423 ( \4106 , \4105 , \2754 );
nand \U$3424 ( \4107 , \4104 , \4106 );
and \U$3425 ( \4108 , \4102 , \4107 );
nor \U$3426 ( \4109 , \4106 , \4104 );
nor \U$3427 ( \4110 , \4108 , \4109 );
xor \U$3428 ( \4111 , \2474 , \2479 );
xor \U$3429 ( \4112 , \4111 , \2482 );
and \U$3430 ( \4113 , \4110 , \4112 );
and \U$3431 ( \4114 , \2587 , \4110 );
or \U$3432 ( \4115 , \2590 , \4113 , \4114 );
xor \U$3433 ( \4116 , \2185 , \2192 );
xor \U$3434 ( \4117 , \4116 , \2319 );
and \U$3435 ( \4118 , \4115 , \4117 );
and \U$3436 ( \4119 , \2485 , \4115 );
or \U$3437 ( \4120 , \2488 , \4118 , \4119 );
and \U$3438 ( \4121 , \2323 , \4120 );
and \U$3439 ( \4122 , \2183 , \2322 );
or \U$3440 ( \4123 , \4121 , \4122 );
not \U$3441 ( \4124 , \4123 );
and \U$3442 ( \4125 , \2176 , \4124 );
and \U$3443 ( \4126 , \2171 , \2175 );
or \U$3444 ( \4127 , \4125 , \4126 );
and \U$3445 ( \4128 , \2060 , \4127 );
and \U$3446 ( \4129 , \2057 , \2059 );
or \U$3447 ( \4130 , \4128 , \4129 );
and \U$3448 ( \4131 , \1944 , \4130 );
and \U$3449 ( \4132 , \1857 , \1943 );
or \U$3450 ( \4133 , \4131 , \4132 );
and \U$3451 ( \4134 , \1855 , \4133 );
and \U$3452 ( \4135 , \1852 , \1854 );
or \U$3453 ( \4136 , \4134 , \4135 );
and \U$3454 ( \4137 , \1744 , \4136 );
and \U$3455 ( \4138 , \1572 , \1743 );
or \U$3456 ( \4139 , \4137 , \4138 );
xor \U$3457 ( \4140 , \1469 , \1471 );
and \U$3458 ( \4141 , \4140 , \1571 );
and \U$3459 ( \4142 , \1469 , \1471 );
or \U$3460 ( \4143 , \4141 , \4142 );
or \U$3461 ( \4144 , \4139 , \4143 );
xor \U$3462 ( \4145 , \1398 , \1462 );
and \U$3463 ( \4146 , \4144 , \4145 );
and \U$3464 ( \4147 , \4143 , \4139 );
nor \U$3465 ( \4148 , \4146 , \4147 );
not \U$3466 ( \4149 , \4148 );
or \U$3467 ( \4150 , \1468 , \4149 );
or \U$3468 ( \4151 , \4148 , \1467 );
nand \U$3469 ( \4152 , \4150 , \4151 );
and \U$3470 ( \4153 , RIaa97fe0_21, \721 );
and \U$3471 ( \4154 , RIaa98418_30, \682 );
and \U$3472 ( \4155 , \686 , RIaa98328_28);
and \U$3473 ( \4156 , RIaa983a0_29, \728 );
nor \U$3474 ( \4157 , \4155 , \4156 );
and \U$3475 ( \4158 , RIaa982b0_27, \690 );
and \U$3476 ( \4159 , \712 , RIaa980d0_23);
and \U$3477 ( \4160 , RIaa981c0_25, \730 );
nor \U$3478 ( \4161 , \4158 , \4159 , \4160 );
and \U$3479 ( \4162 , \738 , RIaa97ef0_19);
and \U$3480 ( \4163 , RIaa98148_24, \741 );
nor \U$3481 ( \4164 , \4162 , \4163 );
nand \U$3482 ( \4165 , \4157 , \4161 , \4164 );
nor \U$3483 ( \4166 , \4153 , \4154 , \4165 );
and \U$3484 ( \4167 , \702 , RIaa98058_22);
and \U$3485 ( \4168 , RIaa98580_33, \699 );
nor \U$3486 ( \4169 , \4167 , \4168 );
and \U$3487 ( \4170 , RIaa98238_26, \723 );
and \U$3488 ( \4171 , RIaa985f8_34, \733 );
and \U$3489 ( \4172 , \696 , RIaa98508_32);
and \U$3490 ( \4173 , RIaa98490_31, \735 );
nor \U$3491 ( \4174 , \4172 , \4173 );
not \U$3492 ( \4175 , \4174 );
nor \U$3493 ( \4176 , \4170 , \4171 , \4175 );
nand \U$3494 ( \4177 , \4166 , \4169 , \709 , \4176 );
buf \U$3495 ( \4178 , \4177 );
buf \U$3496 ( \4179 , \749 );
_DC g11c3 ( \4180_nG11c3 , \4178 , \4179 );
xor \U$3497 ( \4181 , \673 , \4180_nG11c3 );
and \U$3498 ( \4182 , \712 , RIaa987d8_38);
and \U$3499 ( \4183 , \682 , RIaa98c10_47);
and \U$3500 ( \4184 , RIaa98aa8_44, \686 );
nor \U$3501 ( \4185 , \4183 , \4184 );
and \U$3502 ( \4186 , \702 , RIaa98940_41);
and \U$3503 ( \4187 , RIaa988c8_40, \721 );
nor \U$3504 ( \4188 , \4186 , \4187 );
and \U$3505 ( \4189 , \733 , RIaa98d00_49);
and \U$3506 ( \4190 , RIaa98850_39, \741 );
nor \U$3507 ( \4191 , \4189 , \4190 );
and \U$3508 ( \4192 , \738 , RIaa98670_35);
and \U$3509 ( \4193 , RIaa98a30_43, \723 );
nor \U$3510 ( \4194 , \4192 , \4193 );
nand \U$3511 ( \4195 , \4185 , \4188 , \4191 , \4194 );
not \U$3512 ( \4196 , \777 );
nor \U$3513 ( \4197 , \4182 , \4195 , \4196 );
and \U$3514 ( \4198 , \735 , RIaa98d78_50);
and \U$3515 ( \4199 , RIaa989b8_42, \730 );
nor \U$3516 ( \4200 , \4198 , \4199 );
and \U$3517 ( \4201 , \696 , RIaa98df0_51);
and \U$3518 ( \4202 , RIaa98b20_45, \699 );
nor \U$3519 ( \4203 , \4201 , \4202 );
and \U$3520 ( \4204 , \728 , RIaa98b98_46);
and \U$3521 ( \4205 , RIaa98c88_48, \690 );
nor \U$3522 ( \4206 , \4204 , \4205 );
nand \U$3523 ( \4207 , \4197 , \4200 , \4203 , \4206 );
buf \U$3524 ( \4208 , \4207 );
_DC gfe5 ( \4209_nGfe5 , \4208 , \4179 );
xor \U$3525 ( \4210 , \757 , \4209_nGfe5 );
and \U$3526 ( \4211 , \712 , RIaa9e0e8_228);
and \U$3527 ( \4212 , \682 , RIaa9e430_235);
and \U$3528 ( \4213 , RIaa9e340_233, \686 );
nor \U$3529 ( \4214 , \4212 , \4213 );
and \U$3530 ( \4215 , \702 , RIaa9e070_227);
and \U$3531 ( \4216 , RIaa9e250_231, \723 );
nor \U$3532 ( \4217 , \4215 , \4216 );
and \U$3533 ( \4218 , \738 , RIaa9de90_223);
and \U$3534 ( \4219 , RIaa9dff8_226, \721 );
nor \U$3535 ( \4220 , \4218 , \4219 );
and \U$3536 ( \4221 , \690 , RIaa9e2c8_232);
and \U$3537 ( \4222 , RIaa9e160_229, \741 );
nor \U$3538 ( \4223 , \4221 , \4222 );
nand \U$3539 ( \4224 , \4214 , \4217 , \4220 , \4223 );
not \U$3540 ( \4225 , \813 );
nor \U$3541 ( \4226 , \4211 , \4224 , \4225 );
and \U$3542 ( \4227 , \696 , RIaa9e520_237);
and \U$3543 ( \4228 , RIaa9e598_238, \699 );
nor \U$3544 ( \4229 , \4227 , \4228 );
and \U$3545 ( \4230 , \733 , RIaa9e610_239);
and \U$3546 ( \4231 , RIaa9e4a8_236, \735 );
nor \U$3547 ( \4232 , \4230 , \4231 );
and \U$3548 ( \4233 , \728 , RIaa9e3b8_234);
and \U$3549 ( \4234 , RIaa9e1d8_230, \730 );
nor \U$3550 ( \4235 , \4233 , \4234 );
nand \U$3551 ( \4236 , \4226 , \4229 , \4232 , \4235 );
buf \U$3552 ( \4237 , \4236 );
_DC gfe3 ( \4238_nGfe3 , \4237 , \4179 );
xor \U$3553 ( \4239 , \793 , \4238_nGfe3 );
and \U$3554 ( \4240 , RIaa9dbc0_217, \721 );
and \U$3555 ( \4241 , RIaa9d8f0_211, \682 );
and \U$3556 ( \4242 , \686 , RIaa9d710_207);
and \U$3557 ( \4243 , RIaa9d878_210, \728 );
nor \U$3558 ( \4244 , \4242 , \4243 );
and \U$3559 ( \4245 , RIaa9d698_206, \690 );
and \U$3560 ( \4246 , \712 , RIaa9dda0_221);
and \U$3561 ( \4247 , RIaa9dcb0_219, \730 );
nor \U$3562 ( \4248 , \4245 , \4246 , \4247 );
and \U$3563 ( \4249 , \738 , RIaa9da58_214);
and \U$3564 ( \4250 , RIaa9de18_222, \741 );
nor \U$3565 ( \4251 , \4249 , \4250 );
nand \U$3566 ( \4252 , \4244 , \4248 , \4251 );
nor \U$3567 ( \4253 , \4240 , \4241 , \4252 );
and \U$3568 ( \4254 , \702 , RIaa9dc38_218);
and \U$3569 ( \4255 , RIaa9d788_208, \699 );
nor \U$3570 ( \4256 , \4254 , \4255 );
and \U$3571 ( \4257 , RIaa9dd28_220, \723 );
and \U$3572 ( \4258 , RIaa9d800_209, \733 );
and \U$3573 ( \4259 , \696 , RIaa9d9e0_213);
and \U$3574 ( \4260 , RIaa9d968_212, \735 );
nor \U$3575 ( \4261 , \4259 , \4260 );
not \U$3576 ( \4262 , \4261 );
nor \U$3577 ( \4263 , \4257 , \4258 , \4262 );
nand \U$3578 ( \4264 , \4253 , \4256 , \838 , \4263 );
buf \U$3579 ( \4265 , \4264 );
_DC ge39 ( \4266_nGe39 , \4265 , \4179 );
xor \U$3580 ( \4267 , \829 , \4266_nGe39 );
and \U$3581 ( \4268 , \741 , RIaa99048_56);
and \U$3582 ( \4269 , \723 , RIaa99408_64);
and \U$3583 ( \4270 , RIaa99228_60, \682 );
nor \U$3584 ( \4271 , \4269 , \4270 );
and \U$3585 ( \4272 , \702 , RIaa992a0_61);
and \U$3586 ( \4273 , RIaa99318_62, \721 );
nor \U$3587 ( \4274 , \4272 , \4273 );
and \U$3588 ( \4275 , \733 , RIaa994f8_66);
and \U$3589 ( \4276 , RIaa995e8_68, \735 );
nor \U$3590 ( \4277 , \4275 , \4276 );
and \U$3591 ( \4278 , \696 , RIaa99570_67);
and \U$3592 ( \4279 , RIaa99138_58, \699 );
nor \U$3593 ( \4280 , \4278 , \4279 );
nand \U$3594 ( \4281 , \4271 , \4274 , \4277 , \4280 );
and \U$3595 ( \4282 , \686 , RIaa990c0_57);
and \U$3596 ( \4283 , RIaa98fd0_55, \712 );
nor \U$3597 ( \4284 , \4282 , \4283 );
not \U$3598 ( \4285 , \4284 );
nor \U$3599 ( \4286 , \4268 , \4281 , \4285 );
and \U$3600 ( \4287 , \738 , RIaa98e68_52);
and \U$3601 ( \4288 , RIaa99390_63, \730 );
nor \U$3602 ( \4289 , \4287 , \4288 );
and \U$3603 ( \4290 , \728 , RIaa991b0_59);
and \U$3604 ( \4291 , RIaa99480_65, \690 );
nor \U$3605 ( \4292 , \4290 , \4291 );
nand \U$3606 ( \4293 , \4286 , \4289 , \876 , \4292 );
buf \U$3607 ( \4294 , \4293 );
_DC ge37 ( \4295_nGe37 , \4294 , \4179 );
xor \U$3608 ( \4296 , \867 , \4295_nGe37 );
and \U$3609 ( \4297 , \741 , RIaa99a20_77);
and \U$3610 ( \4298 , \723 , RIaa99c00_81);
and \U$3611 ( \4299 , RIaa997c8_72, \682 );
nor \U$3612 ( \4300 , \4298 , \4299 );
and \U$3613 ( \4301 , \702 , RIaa99a98_78);
and \U$3614 ( \4302 , RIaa99b10_79, \721 );
nor \U$3615 ( \4303 , \4301 , \4302 );
and \U$3616 ( \4304 , \733 , RIaa99de0_85);
and \U$3617 ( \4305 , RIaa996d8_70, \735 );
nor \U$3618 ( \4306 , \4304 , \4305 );
and \U$3619 ( \4307 , \696 , RIaa99660_69);
and \U$3620 ( \4308 , RIaa99d68_84, \699 );
nor \U$3621 ( \4309 , \4307 , \4308 );
nand \U$3622 ( \4310 , \4300 , \4303 , \4306 , \4309 );
and \U$3623 ( \4311 , \686 , RIaa99c78_82);
and \U$3624 ( \4312 , RIaa999a8_76, \712 );
nor \U$3625 ( \4313 , \4311 , \4312 );
not \U$3626 ( \4314 , \4313 );
nor \U$3627 ( \4315 , \4297 , \4310 , \4314 );
and \U$3628 ( \4316 , \738 , RIaa99840_73);
and \U$3629 ( \4317 , RIaa99b88_80, \730 );
nor \U$3630 ( \4318 , \4316 , \4317 );
and \U$3631 ( \4319 , \728 , RIaa99750_71);
and \U$3632 ( \4320 , RIaa99cf0_83, \690 );
nor \U$3633 ( \4321 , \4319 , \4320 );
nand \U$3634 ( \4322 , \4315 , \4318 , \914 , \4321 );
buf \U$3635 ( \4323 , \4322 );
_DC gaa2 ( \4324_nGaa2 , \4323 , \4179 );
xor \U$3636 ( \4325 , \905 , \4324_nGaa2 );
and \U$3637 ( \4326 , \741 , RIaa9a038_90);
and \U$3638 ( \4327 , \723 , RIaa9a218_94);
and \U$3639 ( \4328 , RIaa9a560_101, \682 );
nor \U$3640 ( \4329 , \4327 , \4328 );
and \U$3641 ( \4330 , \702 , RIaa9a128_92);
and \U$3642 ( \4331 , RIaa9a1a0_93, \721 );
nor \U$3643 ( \4332 , \4330 , \4331 );
and \U$3644 ( \4333 , \733 , RIaa9a5d8_102);
and \U$3645 ( \4334 , RIaa9a3f8_98, \735 );
nor \U$3646 ( \4335 , \4333 , \4334 );
and \U$3647 ( \4336 , \696 , RIaa9a380_97);
and \U$3648 ( \4337 , RIaa9a290_95, \699 );
nor \U$3649 ( \4338 , \4336 , \4337 );
nand \U$3650 ( \4339 , \4329 , \4332 , \4335 , \4338 );
and \U$3651 ( \4340 , \686 , RIaa9a308_96);
and \U$3652 ( \4341 , RIaa99f48_88, \712 );
nor \U$3653 ( \4342 , \4340 , \4341 );
not \U$3654 ( \4343 , \4342 );
nor \U$3655 ( \4344 , \4326 , \4339 , \4343 );
and \U$3656 ( \4345 , \738 , RIaa99e58_86);
and \U$3657 ( \4346 , RIaa9a0b0_91, \730 );
nor \U$3658 ( \4347 , \4345 , \4346 );
and \U$3659 ( \4348 , \728 , RIaa9a4e8_100);
and \U$3660 ( \4349 , RIaa9a470_99, \690 );
nor \U$3661 ( \4350 , \4348 , \4349 );
nand \U$3662 ( \4351 , \4344 , \4347 , \952 , \4350 );
buf \U$3663 ( \4352 , \4351 );
_DC gaa0 ( \4353_nGaa0 , \4352 , \4179 );
xor \U$3664 ( \4354 , \943 , \4353_nGaa0 );
and \U$3665 ( \4355 , RIaa9a830_107, \741 );
and \U$3666 ( \4356 , RIaa9a650_103, \738 );
and \U$3667 ( \4357 , \723 , RIaa9add0_119);
and \U$3668 ( \4358 , RIaa9ab00_113, \682 );
nor \U$3669 ( \4359 , \4357 , \4358 );
and \U$3670 ( \4360 , \696 , RIaa9a998_110);
and \U$3671 ( \4361 , RIaa9a8a8_108, \699 );
nor \U$3672 ( \4362 , \4360 , \4361 );
and \U$3673 ( \4363 , \702 , RIaa9ace0_117);
and \U$3674 ( \4364 , RIaa9ac68_116, \721 );
nor \U$3675 ( \4365 , \4363 , \4364 );
and \U$3676 ( \4366 , \733 , RIaa9abf0_115);
and \U$3677 ( \4367 , RIaa9aa10_111, \735 );
nor \U$3678 ( \4368 , \4366 , \4367 );
nand \U$3679 ( \4369 , \4359 , \4362 , \4365 , \4368 );
nor \U$3680 ( \4370 , \4355 , \4356 , \4369 );
and \U$3681 ( \4371 , \686 , RIaa9a920_109);
and \U$3682 ( \4372 , RIaa9ab78_114, \728 );
nor \U$3683 ( \4373 , \4371 , \4372 );
and \U$3684 ( \4374 , \730 , RIaa9ad58_118);
not \U$3685 ( \4375 , \1005 );
nor \U$3686 ( \4376 , \4374 , \4375 );
and \U$3687 ( \4377 , \690 , RIaa9aa88_112);
and \U$3688 ( \4378 , RIaa9a7b8_106, \712 );
nor \U$3689 ( \4379 , \4377 , \4378 );
nand \U$3690 ( \4380 , \4370 , \4373 , \4376 , \4379 );
buf \U$3691 ( \4381 , \4380 );
_DC ga31 ( \4382_nGa31 , \4381 , \4179 );
xor \U$3692 ( \4383 , \981 , \4382_nGa31 );
and \U$3693 ( \4384 , \741 , RIaa9cf90_191);
and \U$3694 ( \4385 , \723 , RIaa9d620_205);
and \U$3695 ( \4386 , RIaa9d350_199, \682 );
nor \U$3696 ( \4387 , \4385 , \4386 );
and \U$3697 ( \4388 , \702 , RIaa9d4b8_202);
and \U$3698 ( \4389 , RIaa9d530_203, \721 );
nor \U$3699 ( \4390 , \4388 , \4389 );
and \U$3700 ( \4391 , \733 , RIaa9d440_201);
and \U$3701 ( \4392 , RIaa9d260_197, \735 );
nor \U$3702 ( \4393 , \4391 , \4392 );
and \U$3703 ( \4394 , \696 , RIaa9d1e8_196);
and \U$3704 ( \4395 , RIaa9d170_195, \699 );
nor \U$3705 ( \4396 , \4394 , \4395 );
nand \U$3706 ( \4397 , \4387 , \4390 , \4393 , \4396 );
and \U$3707 ( \4398 , \686 , RIaa9d0f8_194);
and \U$3708 ( \4399 , RIaa9cf18_190, \712 );
nor \U$3709 ( \4400 , \4398 , \4399 );
not \U$3710 ( \4401 , \4400 );
nor \U$3711 ( \4402 , \4384 , \4397 , \4401 );
and \U$3712 ( \4403 , \738 , RIaa9d008_192);
and \U$3713 ( \4404 , RIaa9d5a8_204, \730 );
nor \U$3714 ( \4405 , \4403 , \4404 );
and \U$3715 ( \4406 , \728 , RIaa9d3c8_200);
and \U$3716 ( \4407 , RIaa9d2d8_198, \690 );
nor \U$3717 ( \4408 , \4406 , \4407 );
nand \U$3718 ( \4409 , \4402 , \4405 , \1026 , \4408 );
buf \U$3719 ( \4410 , \4409 );
_DC ga2f ( \4411_nGa2f , \4410 , \4179 );
xor \U$3720 ( \4412 , \1017 , \4411_nGa2f );
and \U$3721 ( \4413 , \741 , RIaa9b028_124);
and \U$3722 ( \4414 , \723 , RIaa9b4d8_134);
and \U$3723 ( \4415 , RIaa9b2f8_130, \682 );
nor \U$3724 ( \4416 , \4414 , \4415 );
and \U$3725 ( \4417 , \702 , RIaa9b550_135);
and \U$3726 ( \4418 , RIaa9b5c8_136, \721 );
nor \U$3727 ( \4419 , \4417 , \4418 );
and \U$3728 ( \4420 , \733 , RIaa9b3e8_132);
and \U$3729 ( \4421 , RIaa9b208_128, \735 );
nor \U$3730 ( \4422 , \4420 , \4421 );
and \U$3731 ( \4423 , \696 , RIaa9b190_127);
and \U$3732 ( \4424 , RIaa9b0a0_125, \699 );
nor \U$3733 ( \4425 , \4423 , \4424 );
nand \U$3734 ( \4426 , \4416 , \4419 , \4422 , \4425 );
and \U$3735 ( \4427 , \686 , RIaa9b118_126);
and \U$3736 ( \4428 , RIaa9afb0_123, \712 );
nor \U$3737 ( \4429 , \4427 , \4428 );
not \U$3738 ( \4430 , \4429 );
nor \U$3739 ( \4431 , \4413 , \4426 , \4430 );
and \U$3740 ( \4432 , \738 , RIaa9ae48_120);
and \U$3741 ( \4433 , RIaa9b460_133, \730 );
nor \U$3742 ( \4434 , \4432 , \4433 );
and \U$3743 ( \4435 , \728 , RIaa9b370_131);
and \U$3744 ( \4436 , RIaa9b280_129, \690 );
nor \U$3745 ( \4437 , \4435 , \4436 );
nand \U$3746 ( \4438 , \4431 , \4434 , \1067 , \4437 );
buf \U$3747 ( \4439 , \4438 );
_DC g9d8 ( \4440_nG9d8 , \4439 , \4179 );
xor \U$3748 ( \4441 , \1051 , \4440_nG9d8 );
and \U$3749 ( \4442 , \741 , RIaa9ba00_145);
and \U$3750 ( \4443 , \682 , RIaa9baf0_147);
and \U$3751 ( \4444 , RIaa9ba78_146, \690 );
nor \U$3752 ( \4445 , \4443 , \4444 );
and \U$3753 ( \4446 , \699 , RIaa9b6b8_138);
and \U$3754 ( \4447 , RIaa9bd48_152, \730 );
nor \U$3755 ( \4448 , \4446 , \4447 );
and \U$3756 ( \4449 , \702 , RIaa9bc58_150);
and \U$3757 ( \4450 , RIaa9bcd0_151, \721 );
nor \U$3758 ( \4451 , \4449 , \4450 );
and \U$3759 ( \4452 , \723 , RIaa9bdc0_153);
and \U$3760 ( \4453 , RIaa9bb68_148, \728 );
nor \U$3761 ( \4454 , \4452 , \4453 );
nand \U$3762 ( \4455 , \4445 , \4448 , \4451 , \4454 );
and \U$3763 ( \4456 , \686 , RIaa9b640_137);
and \U$3764 ( \4457 , RIaa9b988_144, \712 );
nor \U$3765 ( \4458 , \4456 , \4457 );
not \U$3766 ( \4459 , \4458 );
nor \U$3767 ( \4460 , \4442 , \4455 , \4459 );
and \U$3768 ( \4461 , \738 , RIaa9b820_141);
and \U$3769 ( \4462 , RIaa9b730_139, \696 );
nor \U$3770 ( \4463 , \4461 , \4462 );
and \U$3771 ( \4464 , \733 , RIaa9bbe0_149);
and \U$3772 ( \4465 , RIaa9b7a8_140, \735 );
nor \U$3773 ( \4466 , \4464 , \4465 );
nand \U$3774 ( \4467 , \4460 , \4463 , \1103 , \4466 );
buf \U$3775 ( \4468 , \4467 );
_DC g9da ( \4469_nG9da , \4468 , \4179 );
xor \U$3776 ( \4470 , \1087 , \4469_nG9da );
and \U$3777 ( \4471 , \712 , RIaa9c1f8_162);
and \U$3778 ( \4472 , \682 , RIaa9c3d8_166);
and \U$3779 ( \4473 , RIaa9c5b8_170, \686 );
nor \U$3780 ( \4474 , \4472 , \4473 );
and \U$3781 ( \4475 , \702 , RIaa9bfa0_157);
and \U$3782 ( \4476 , RIaa9bf28_156, \721 );
nor \U$3783 ( \4477 , \4475 , \4476 );
and \U$3784 ( \4478 , \738 , RIaa9c018_158);
and \U$3785 ( \4479 , RIaa9beb0_155, \733 );
nor \U$3786 ( \4480 , \4478 , \4479 );
and \U$3787 ( \4481 , \723 , RIaa9c4c8_168);
and \U$3788 ( \4482 , RIaa9c180_161, \741 );
nor \U$3789 ( \4483 , \4481 , \4482 );
nand \U$3790 ( \4484 , \4474 , \4477 , \4480 , \4483 );
not \U$3791 ( \4485 , \1138 );
nor \U$3792 ( \4486 , \4471 , \4484 , \4485 );
and \U$3793 ( \4487 , \735 , RIaa9c540_169);
and \U$3794 ( \4488 , RIaa9c450_167, \730 );
nor \U$3795 ( \4489 , \4487 , \4488 );
and \U$3796 ( \4490 , \696 , RIaa9c270_163);
and \U$3797 ( \4491 , RIaa9c2e8_164, \699 );
nor \U$3798 ( \4492 , \4490 , \4491 );
and \U$3799 ( \4493 , \728 , RIaa9c360_165);
and \U$3800 ( \4494 , RIaa9be38_154, \690 );
nor \U$3801 ( \4495 , \4493 , \4494 );
nand \U$3802 ( \4496 , \4486 , \4489 , \4492 , \4495 );
buf \U$3803 ( \4497 , \4496 );
_DC g969 ( \4498_nG969 , \4497 , \4179 );
xor \U$3804 ( \4499 , RIaa977e8_4, \4498_nG969 );
and \U$3805 ( \4500 , RIaa9cae0_181, \721 );
and \U$3806 ( \4501 , RIaa9cbd0_183, \682 );
and \U$3807 ( \4502 , \686 , RIaa9c888_176);
and \U$3808 ( \4503 , RIaa9c9f0_179, \728 );
nor \U$3809 ( \4504 , \4502 , \4503 );
and \U$3810 ( \4505 , RIaa9cd38_186, \690 );
and \U$3811 ( \4506 , \712 , RIaa9c630_171);
and \U$3812 ( \4507 , RIaa9ca68_180, \730 );
nor \U$3813 ( \4508 , \4505 , \4506 , \4507 );
and \U$3814 ( \4509 , \738 , RIaa9c6a8_172);
and \U$3815 ( \4510 , RIaa9c810_175, \741 );
nor \U$3816 ( \4511 , \4509 , \4510 );
nand \U$3817 ( \4512 , \4504 , \4508 , \4511 );
nor \U$3818 ( \4513 , \4500 , \4501 , \4512 );
and \U$3819 ( \4514 , \702 , RIaa9c978_178);
and \U$3820 ( \4515 , RIaa9ccc0_185, \699 );
nor \U$3821 ( \4516 , \4514 , \4515 );
and \U$3822 ( \4517 , RIaa9cb58_182, \723 );
and \U$3823 ( \4518 , RIaa9cdb0_187, \733 );
and \U$3824 ( \4519 , \696 , RIaa9cc48_184);
and \U$3825 ( \4520 , RIaa9c900_177, \735 );
nor \U$3826 ( \4521 , \4519 , \4520 );
not \U$3827 ( \4522 , \4521 );
nor \U$3828 ( \4523 , \4517 , \4518 , \4522 );
nand \U$3829 ( \4524 , \4513 , \4516 , \1158 , \4523 );
buf \U$3830 ( \4525 , \4524 );
_DC g967 ( \4526_nG967 , \4525 , \4179 );
nand \U$3831 ( \4527 , \4526_nG967 , \1182 );
not \U$3832 ( \4528 , \4527 );
and \U$3833 ( \4529 , \4499 , \4528 );
and \U$3834 ( \4530 , RIaa977e8_4, \4498_nG969 );
or \U$3835 ( \4531 , \4529 , \4530 );
and \U$3836 ( \4532 , \4470 , \4531 );
and \U$3837 ( \4533 , \1087 , \4469_nG9da );
or \U$3838 ( \4534 , \4532 , \4533 );
and \U$3839 ( \4535 , \4441 , \4534 );
and \U$3840 ( \4536 , \1051 , \4440_nG9d8 );
or \U$3841 ( \4537 , \4535 , \4536 );
and \U$3842 ( \4538 , \4412 , \4537 );
and \U$3843 ( \4539 , \1017 , \4411_nGa2f );
or \U$3844 ( \4540 , \4538 , \4539 );
and \U$3845 ( \4541 , \4383 , \4540 );
and \U$3846 ( \4542 , \981 , \4382_nGa31 );
or \U$3847 ( \4543 , \4541 , \4542 );
and \U$3848 ( \4544 , \4354 , \4543 );
and \U$3849 ( \4545 , \943 , \4353_nGaa0 );
or \U$3850 ( \4546 , \4544 , \4545 );
and \U$3851 ( \4547 , \4325 , \4546 );
and \U$3852 ( \4548 , \905 , \4324_nGaa2 );
or \U$3853 ( \4549 , \4547 , \4548 );
and \U$3854 ( \4550 , \4296 , \4549 );
and \U$3855 ( \4551 , \867 , \4295_nGe37 );
or \U$3856 ( \4552 , \4550 , \4551 );
and \U$3857 ( \4553 , \4267 , \4552 );
and \U$3858 ( \4554 , \829 , \4266_nGe39 );
or \U$3859 ( \4555 , \4553 , \4554 );
and \U$3860 ( \4556 , \4239 , \4555 );
and \U$3861 ( \4557 , \793 , \4238_nGfe3 );
or \U$3862 ( \4558 , \4556 , \4557 );
and \U$3863 ( \4559 , \4210 , \4558 );
and \U$3864 ( \4560 , \757 , \4209_nGfe5 );
or \U$3865 ( \4561 , \4559 , \4560 );
and \U$3866 ( \4562 , \4181 , \4561 );
and \U$3867 ( \4563 , \673 , \4180_nG11c3 );
or \U$3868 ( \4564 , \4562 , \4563 );
nor \U$3869 ( \4565 , \4564 , \1222 );
not \U$3870 ( \4566 , \4565 );
and \U$3871 ( \4567 , RIaa9f678_274, \723 );
and \U$3872 ( \4568 , RIaa9f420_269, \721 );
and \U$3873 ( \4569 , \728 , RIaa9f6f0_275);
and \U$3874 ( \4570 , RIaa9f8d0_279, \690 );
nor \U$3875 ( \4571 , \4569 , \4570 );
or \U$3876 ( \4572 , \741 , \708 );
and \U$3877 ( \4573 , RIaa9f588_272, \4572 );
and \U$3878 ( \4574 , \712 , RIaa9f600_273);
and \U$3879 ( \4575 , RIaa9f2b8_266, \735 );
nor \U$3880 ( \4576 , \4573 , \4574 , \4575 );
and \U$3881 ( \4577 , \733 , RIaa9f768_276);
and \U$3882 ( \4578 , RIaa9f3a8_268, \730 );
nor \U$3883 ( \4579 , \4577 , \4578 );
nand \U$3884 ( \4580 , \4571 , \4576 , \4579 );
nor \U$3885 ( \4581 , \4567 , \4568 , \4580 );
and \U$3886 ( \4582 , \702 , RIaa9f858_278);
and \U$3887 ( \4583 , RIaa9f7e0_277, \682 );
nor \U$3888 ( \4584 , \4582 , \4583 );
and \U$3889 ( \4585 , \696 , RIaa9f948_280);
and \U$3890 ( \4586 , RIaa9f498_270, \699 );
nor \U$3891 ( \4587 , \4585 , \4586 );
and \U$3892 ( \4588 , \738 , RIaa9f330_267);
and \U$3893 ( \4589 , RIaa9f9c0_281, \686 );
nor \U$3894 ( \4590 , \4588 , \4589 );
nand \U$3895 ( \4591 , \4581 , \4584 , \4587 , \4590 );
buf \U$3896 ( \4592 , \749 );
_DC g17f6 ( \4593_nG17f6 , \4591 , \4592 );
not \U$3897 ( \4594 , \4593_nG17f6 );
nor \U$3898 ( \4595 , \4566 , \4594 );
xor \U$3899 ( \4596 , \673 , \4180_nG11c3 );
xor \U$3900 ( \4597 , \4596 , \4561 );
not \U$3901 ( \4598 , \4597 );
xor \U$3902 ( \4599 , \757 , \4209_nGfe5 );
xor \U$3903 ( \4600 , \4599 , \4558 );
not \U$3904 ( \4601 , \4600 );
and \U$3905 ( \4602 , \4598 , \4601 );
and \U$3906 ( \4603 , \4564 , \1222 );
nor \U$3907 ( \4604 , \4603 , \4565 );
nor \U$3908 ( \4605 , \4602 , \4604 );
not \U$3909 ( \4606 , \4605 );
and \U$3910 ( \4607 , \4572 , RIaa9ebb0_251);
and \U$3911 ( \4608 , \682 , RIaa9f060_261);
and \U$3912 ( \4609 , RIaa9efe8_260, \686 );
nor \U$3913 ( \4610 , \4608 , \4609 );
and \U$3914 ( \4611 , \738 , RIaa9eca0_253);
and \U$3915 ( \4612 , RIaa9ed90_255, \699 );
nor \U$3916 ( \4613 , \4611 , \4612 );
and \U$3917 ( \4614 , \702 , RIaa9f150_263);
and \U$3918 ( \4615 , RIaa9ee08_256, \721 );
nor \U$3919 ( \4616 , \4614 , \4615 );
and \U$3920 ( \4617 , \696 , RIaa9ef70_259);
and \U$3921 ( \4618 , RIaa9ee80_257, \723 );
nor \U$3922 ( \4619 , \4617 , \4618 );
nand \U$3923 ( \4620 , \4610 , \4613 , \4616 , \4619 );
nor \U$3924 ( \4621 , \4607 , \4620 );
and \U$3925 ( \4622 , \730 , RIaa9ed18_254);
and \U$3926 ( \4623 , RIaa9f1c8_264, \690 );
nor \U$3927 ( \4624 , \4622 , \4623 );
and \U$3928 ( \4625 , \733 , RIaa9f0d8_262);
and \U$3929 ( \4626 , RIaa9ec28_252, \735 );
nor \U$3930 ( \4627 , \4625 , \4626 );
and \U$3931 ( \4628 , \728 , RIaa9eef8_258);
and \U$3932 ( \4629 , RIaa9eb38_250, \712 );
nor \U$3933 ( \4630 , \4628 , \4629 );
nand \U$3934 ( \4631 , \4621 , \4624 , \4627 , \4630 );
_DC g1905 ( \4632_nG1905 , \4631 , \4592 );
or \U$3935 ( \4633 , \4606 , \4632_nG1905 );
not \U$3936 ( \4634 , \4632_nG1905 );
and \U$3937 ( \4635 , \4604 , \4597 );
nor \U$3938 ( \4636 , \4604 , \4597 );
xnor \U$3939 ( \4637 , \4600 , \4597 );
not \U$3940 ( \4638 , \4637 );
nor \U$3941 ( \4639 , \4635 , \4636 , \4638 );
nand \U$3942 ( \4640 , \4606 , \4639 );
or \U$3943 ( \4641 , \4634 , \4640 );
or \U$3944 ( \4642 , \4639 , \4606 );
nand \U$3945 ( \4643 , \4633 , \4641 , \4642 );
xnor \U$3946 ( \4644 , \4595 , \4643 );
nor \U$3947 ( \4645 , \4605 , \4637 );
not \U$3948 ( \4646 , \4645 );
or \U$3949 ( \4647 , \4646 , \4634 );
or \U$3950 ( \4648 , \4594 , \4640 );
or \U$3951 ( \4649 , \4637 , \4634 );
or \U$3952 ( \4650 , \4606 , \4593_nG17f6 );
nand \U$3953 ( \4651 , \4650 , \4642 );
nand \U$3954 ( \4652 , \4649 , \4651 );
nand \U$3955 ( \4653 , \4647 , \4648 , \4652 );
xor \U$3956 ( \4654 , \793 , \4238_nGfe3 );
xor \U$3957 ( \4655 , \4654 , \4555 );
xor \U$3958 ( \4656 , \829 , \4266_nGe39 );
xor \U$3959 ( \4657 , \4656 , \4552 );
nor \U$3960 ( \4658 , \4655 , \4657 );
or \U$3961 ( \4659 , \4600 , \4658 );
and \U$3962 ( \4660 , \4653 , \4659 );
and \U$3963 ( \4661 , \690 , RIaa9fab0_283);
and \U$3964 ( \4662 , \721 , RIaa9fdf8_290);
and \U$3965 ( \4663 , RIaa9fd80_289, \686 );
nor \U$3966 ( \4664 , \4662 , \4663 );
and \U$3967 ( \4665 , \738 , RIaaa0140_297);
and \U$3968 ( \4666 , RIaaa00c8_296, \699 );
nor \U$3969 ( \4667 , \4665 , \4666 );
and \U$3970 ( \4668 , \733 , RIaa9fe70_291);
and \U$3971 ( \4669 , RIaaa0050_295, \730 );
nor \U$3972 ( \4670 , \4668 , \4669 );
and \U$3973 ( \4671 , \696 , RIaa9fd08_288);
and \U$3974 ( \4672 , RIaaa01b8_298, \735 );
nor \U$3975 ( \4673 , \4671 , \4672 );
nand \U$3976 ( \4674 , \4664 , \4667 , \4670 , \4673 );
nor \U$3977 ( \4675 , \4661 , \4674 );
and \U$3978 ( \4676 , \682 , RIaa9fee8_292);
and \U$3979 ( \4677 , RIaa9ffd8_294, \728 );
nor \U$3980 ( \4678 , \4676 , \4677 );
and \U$3981 ( \4679 , \702 , RIaa9fa38_282);
and \U$3982 ( \4680 , RIaa9fc90_287, \712 );
nor \U$3983 ( \4681 , \4679 , \4680 );
and \U$3984 ( \4682 , \4572 , RIaa9fc18_286);
and \U$3985 ( \4683 , RIaa9ff60_293, \723 );
nor \U$3986 ( \4684 , \4682 , \4683 );
nand \U$3987 ( \4685 , \4675 , \4678 , \4681 , \4684 );
_DC g16f0 ( \4686_nG16f0 , \4685 , \4592 );
not \U$3988 ( \4687 , \4686_nG16f0 );
nor \U$3989 ( \4688 , \4566 , \4687 );
nor \U$3990 ( \4689 , \4660 , \4688 );
xor \U$3991 ( \4690 , \4644 , \4689 );
not \U$3992 ( \4691 , \4690 );
not \U$3993 ( \4692 , \4655 );
not \U$3994 ( \4693 , \4600 );
or \U$3995 ( \4694 , \4692 , \4693 );
or \U$3996 ( \4695 , \4600 , \4655 );
nand \U$3997 ( \4696 , \4694 , \4695 );
xor \U$3998 ( \4697 , \4657 , \4655 );
nor \U$3999 ( \4698 , \4696 , \4697 );
not \U$4000 ( \4699 , \4698 );
not \U$4001 ( \4700 , \4659 );
nor \U$4002 ( \4701 , \4699 , \4700 );
not \U$4003 ( \4702 , \4701 );
or \U$4004 ( \4703 , \4702 , \4634 );
or \U$4005 ( \4704 , \4699 , \4634 );
nand \U$4006 ( \4705 , \4704 , \4700 );
nand \U$4007 ( \4706 , \4703 , \4705 );
or \U$4008 ( \4707 , \4646 , \4594 );
or \U$4009 ( \4708 , \4687 , \4640 );
or \U$4010 ( \4709 , \4637 , \4594 );
or \U$4011 ( \4710 , \4606 , \4686_nG16f0 );
nand \U$4012 ( \4711 , \4710 , \4642 );
nand \U$4013 ( \4712 , \4709 , \4711 );
nand \U$4014 ( \4713 , \4707 , \4708 , \4712 );
and \U$4015 ( \4714 , \4706 , \4713 );
and \U$4016 ( \4715 , \4653 , \4659 );
not \U$4017 ( \4716 , \4653 );
and \U$4018 ( \4717 , \4716 , \4700 );
nor \U$4019 ( \4718 , \4715 , \4717 );
xor \U$4020 ( \4719 , \4688 , \4718 );
and \U$4021 ( \4720 , \4714 , \4719 );
xor \U$4022 ( \4721 , \4691 , \4720 );
xor \U$4023 ( \4722 , \4714 , \4719 );
nand \U$4024 ( \4723 , \4593_nG17f6 , \4698 );
or \U$4025 ( \4724 , \4659 , \4632_nG1905 );
or \U$4026 ( \4725 , \4659 , \4697 );
nand \U$4027 ( \4726 , \4724 , \4725 );
and \U$4028 ( \4727 , \4723 , \4726 );
and \U$4029 ( \4728 , \4659 , \4697 );
and \U$4030 ( \4729 , \4728 , \4632_nG1905 );
and \U$4031 ( \4730 , \4593_nG17f6 , \4701 );
nor \U$4032 ( \4731 , \4727 , \4729 , \4730 );
and \U$4033 ( \4732 , \4686_nG16f0 , \4645 );
and \U$4034 ( \4733 , RIaaa0578_306, \723 );
and \U$4035 ( \4734 , RIaaa02a8_300, \682 );
and \U$4036 ( \4735 , \728 , RIaaa05f0_307);
and \U$4037 ( \4736 , RIaaa08c0_313, \690 );
nor \U$4038 ( \4737 , \4735 , \4736 );
and \U$4039 ( \4738 , RIaaa07d0_311, \4572 );
and \U$4040 ( \4739 , \712 , RIaaa0848_312);
and \U$4041 ( \4740 , RIaaa06e0_309, \735 );
nor \U$4042 ( \4741 , \4738 , \4739 , \4740 );
and \U$4043 ( \4742 , \733 , RIaaa0230_299);
and \U$4044 ( \4743 , RIaaa0488_304, \730 );
nor \U$4045 ( \4744 , \4742 , \4743 );
nand \U$4046 ( \4745 , \4737 , \4741 , \4744 );
nor \U$4047 ( \4746 , \4733 , \4734 , \4745 );
and \U$4048 ( \4747 , \702 , RIaaa0938_314);
and \U$4049 ( \4748 , RIaaa0410_303, \721 );
nor \U$4050 ( \4749 , \4747 , \4748 );
and \U$4051 ( \4750 , \738 , RIaaa0668_308);
and \U$4052 ( \4751 , RIaaa0320_301, \696 );
nor \U$4053 ( \4752 , \4750 , \4751 );
and \U$4054 ( \4753 , \699 , RIaaa0500_305);
and \U$4055 ( \4754 , RIaaa0398_302, \686 );
nor \U$4056 ( \4755 , \4753 , \4754 );
nand \U$4057 ( \4756 , \4746 , \4749 , \4752 , \4755 );
_DC g15ca ( \4757_nG15ca , \4756 , \4592 );
or \U$4058 ( \4758 , \4606 , \4757_nG15ca );
nand \U$4059 ( \4759 , \4758 , \4642 );
nand \U$4060 ( \4760 , \4686_nG16f0 , \4638 );
and \U$4061 ( \4761 , \4759 , \4760 );
not \U$4062 ( \4762 , \4640 );
and \U$4063 ( \4763 , \4757_nG15ca , \4762 );
nor \U$4064 ( \4764 , \4732 , \4761 , \4763 );
nand \U$4065 ( \4765 , \4731 , \4764 );
xor \U$4066 ( \4766 , \867 , \4295_nGe37 );
xor \U$4067 ( \4767 , \4766 , \4549 );
xor \U$4068 ( \4768 , \905 , \4324_nGaa2 );
xor \U$4069 ( \4769 , \4768 , \4546 );
nor \U$4070 ( \4770 , \4767 , \4769 );
or \U$4071 ( \4771 , \4657 , \4770 );
and \U$4072 ( \4772 , \4765 , \4771 );
nor \U$4073 ( \4773 , \4764 , \4731 );
nor \U$4074 ( \4774 , \4772 , \4773 );
xor \U$4075 ( \4775 , \4706 , \4713 );
not \U$4076 ( \4776 , \4775 );
nand \U$4077 ( \4777 , \4757_nG15ca , \4565 );
not \U$4078 ( \4778 , \4777 );
and \U$4079 ( \4779 , \4776 , \4778 );
and \U$4080 ( \4780 , \4775 , \4777 );
nor \U$4081 ( \4781 , \4779 , \4780 );
nand \U$4082 ( \4782 , \4774 , \4781 );
and \U$4083 ( \4783 , \4722 , \4782 );
and \U$4084 ( \4784 , \4721 , \4783 );
not \U$4085 ( \4785 , \4784 );
and \U$4086 ( \4786 , \4691 , \4720 );
or \U$4087 ( \4787 , \4786 , \4605 );
and \U$4088 ( \4788 , \4643 , \4595 );
and \U$4089 ( \4789 , \4605 , \4786 );
nor \U$4090 ( \4790 , \4788 , \4789 );
nand \U$4091 ( \4791 , \4787 , \4790 );
not \U$4092 ( \4792 , \4791 );
and \U$4093 ( \4793 , \4565 , \4632_nG1905 );
and \U$4094 ( \4794 , \4644 , \4689 );
nor \U$4095 ( \4795 , \4793 , \4794 );
not \U$4096 ( \4796 , \4795 );
and \U$4097 ( \4797 , \4792 , \4796 );
and \U$4098 ( \4798 , \4791 , \4795 );
nor \U$4099 ( \4799 , \4797 , \4798 );
not \U$4100 ( \4800 , \4799 );
or \U$4101 ( \4801 , \4785 , \4800 );
or \U$4102 ( \4802 , \4799 , \4784 );
nand \U$4103 ( \4803 , \4801 , \4802 );
not \U$4104 ( \4804 , \4803 );
xor \U$4105 ( \4805 , \4722 , \4782 );
not \U$4106 ( \4806 , \4775 );
nor \U$4107 ( \4807 , \4806 , \4777 );
xor \U$4108 ( \4808 , \4805 , \4807 );
or \U$4109 ( \4809 , \4781 , \4774 );
nand \U$4110 ( \4810 , \4809 , \4782 );
not \U$4111 ( \4811 , \4810 );
and \U$4112 ( \4812 , RIaaa0b18_318, \723 );
and \U$4113 ( \4813 , RIaaa0ed8_326, \721 );
and \U$4114 ( \4814 , \728 , RIaaa0b90_319);
and \U$4115 ( \4815 , RIaaa10b8_330, \690 );
nor \U$4116 ( \4816 , \4814 , \4815 );
and \U$4117 ( \4817 , RIaaa0fc8_328, \4572 );
and \U$4118 ( \4818 , \712 , RIaaa1040_329);
and \U$4119 ( \4819 , RIaaa0c80_321, \735 );
nor \U$4120 ( \4820 , \4817 , \4818 , \4819 );
and \U$4121 ( \4821 , \733 , RIaaa0cf8_322);
and \U$4122 ( \4822 , RIaaa0a28_316, \730 );
nor \U$4123 ( \4823 , \4821 , \4822 );
nand \U$4124 ( \4824 , \4816 , \4820 , \4823 );
nor \U$4125 ( \4825 , \4812 , \4813 , \4824 );
and \U$4126 ( \4826 , \702 , RIaaa1130_331);
and \U$4127 ( \4827 , RIaaa0d70_323, \682 );
nor \U$4128 ( \4828 , \4826 , \4827 );
and \U$4129 ( \4829 , \696 , RIaaa0de8_324);
and \U$4130 ( \4830 , RIaaa0aa0_317, \699 );
nor \U$4131 ( \4831 , \4829 , \4830 );
and \U$4132 ( \4832 , \738 , RIaaa0c08_320);
and \U$4133 ( \4833 , RIaaa0e60_325, \686 );
nor \U$4134 ( \4834 , \4832 , \4833 );
nand \U$4135 ( \4835 , \4825 , \4828 , \4831 , \4834 );
_DC g14e1 ( \4836_nG14e1 , \4835 , \4592 );
not \U$4136 ( \4837 , \4836_nG14e1 );
nor \U$4137 ( \4838 , \4566 , \4837 );
not \U$4138 ( \4839 , \4771 );
not \U$4139 ( \4840 , \4773 );
nand \U$4140 ( \4841 , \4840 , \4765 );
not \U$4141 ( \4842 , \4841 );
or \U$4142 ( \4843 , \4839 , \4842 );
or \U$4143 ( \4844 , \4841 , \4771 );
nand \U$4144 ( \4845 , \4843 , \4844 );
xnor \U$4145 ( \4846 , \4838 , \4845 );
not \U$4146 ( \4847 , \4846 );
nand \U$4147 ( \4848 , \4686_nG16f0 , \4698 );
or \U$4148 ( \4849 , \4659 , \4593_nG17f6 );
nand \U$4149 ( \4850 , \4849 , \4725 );
and \U$4150 ( \4851 , \4848 , \4850 );
and \U$4151 ( \4852 , \4728 , \4593_nG17f6 );
and \U$4152 ( \4853 , \4686_nG16f0 , \4701 );
nor \U$4153 ( \4854 , \4851 , \4852 , \4853 );
and \U$4154 ( \4855 , \4657 , \4767 );
nor \U$4155 ( \4856 , \4657 , \4767 );
xor \U$4156 ( \4857 , \4767 , \4769 );
nor \U$4157 ( \4858 , \4855 , \4856 , \4857 );
and \U$4158 ( \4859 , \4771 , \4858 );
and \U$4159 ( \4860 , \4632_nG1905 , \4859 );
not \U$4160 ( \4861 , \4771 );
and \U$4161 ( \4862 , \4634 , \4861 );
or \U$4162 ( \4863 , \4858 , \4771 );
not \U$4163 ( \4864 , \4863 );
nor \U$4164 ( \4865 , \4860 , \4862 , \4864 );
or \U$4165 ( \4866 , \4854 , \4865 );
and \U$4166 ( \4867 , RIaaa1fb8_362, \686 );
and \U$4167 ( \4868 , RIaaa1dd8_358, \699 );
and \U$4168 ( \4869 , \728 , RIaaa1ec8_360);
and \U$4169 ( \4870 , RIaaa2198_366, \690 );
nor \U$4170 ( \4871 , \4869 , \4870 );
and \U$4171 ( \4872 , RIaaa1b08_352, \4572 );
and \U$4172 ( \4873 , \712 , RIaaa1b80_353);
and \U$4173 ( \4874 , RIaaa1bf8_354, \735 );
nor \U$4174 ( \4875 , \4872 , \4873 , \4874 );
and \U$4175 ( \4876 , \733 , RIaaa2030_363);
and \U$4176 ( \4877 , RIaaa1ce8_356, \730 );
nor \U$4177 ( \4878 , \4876 , \4877 );
nand \U$4178 ( \4879 , \4871 , \4875 , \4878 );
nor \U$4179 ( \4880 , \4867 , \4868 , \4879 );
and \U$4180 ( \4881 , \702 , RIaaa2120_365);
and \U$4181 ( \4882 , RIaaa20a8_364, \682 );
nor \U$4182 ( \4883 , \4881 , \4882 );
and \U$4183 ( \4884 , \738 , RIaaa1c70_355);
and \U$4184 ( \4885 , RIaaa1f40_361, \696 );
nor \U$4185 ( \4886 , \4884 , \4885 );
and \U$4186 ( \4887 , \721 , RIaaa1d60_357);
and \U$4187 ( \4888 , RIaaa1e50_359, \723 );
nor \U$4188 ( \4889 , \4887 , \4888 );
nand \U$4189 ( \4890 , \4880 , \4883 , \4886 , \4889 );
_DC g13e1 ( \4891_nG13e1 , \4890 , \4592 );
nand \U$4190 ( \4892 , \4891_nG13e1 , \4565 );
and \U$4191 ( \4893 , \4757_nG15ca , \4645 );
or \U$4192 ( \4894 , \4606 , \4836_nG14e1 );
nand \U$4193 ( \4895 , \4894 , \4642 );
nand \U$4194 ( \4896 , \4757_nG15ca , \4638 );
and \U$4195 ( \4897 , \4895 , \4896 );
and \U$4196 ( \4898 , \4836_nG14e1 , \4762 );
nor \U$4197 ( \4899 , \4893 , \4897 , \4898 );
or \U$4198 ( \4900 , \4892 , \4899 );
nand \U$4199 ( \4901 , \4866 , \4900 );
nand \U$4200 ( \4902 , \4847 , \4901 );
nor \U$4201 ( \4903 , \4811 , \4902 );
and \U$4202 ( \4904 , \4808 , \4903 );
and \U$4203 ( \4905 , \4805 , \4807 );
or \U$4204 ( \4906 , \4904 , \4905 );
xor \U$4205 ( \4907 , \4721 , \4783 );
xor \U$4206 ( \4908 , \4906 , \4907 );
xor \U$4207 ( \4909 , \4805 , \4807 );
xor \U$4208 ( \4910 , \4909 , \4903 );
and \U$4209 ( \4911 , \4845 , \4838 );
nand \U$4210 ( \4912 , \4632_nG1905 , \4857 );
or \U$4211 ( \4913 , \4771 , \4593_nG17f6 );
nand \U$4212 ( \4914 , \4913 , \4863 );
and \U$4213 ( \4915 , \4912 , \4914 );
and \U$4214 ( \4916 , \4859 , \4593_nG17f6 );
not \U$4215 ( \4917 , \4857 );
nor \U$4216 ( \4918 , \4861 , \4917 );
and \U$4217 ( \4919 , \4632_nG1905 , \4918 );
nor \U$4218 ( \4920 , \4915 , \4916 , \4919 );
nand \U$4219 ( \4921 , \4757_nG15ca , \4698 );
or \U$4220 ( \4922 , \4659 , \4686_nG16f0 );
nand \U$4221 ( \4923 , \4922 , \4725 );
and \U$4222 ( \4924 , \4921 , \4923 );
and \U$4223 ( \4925 , \4728 , \4686_nG16f0 );
and \U$4224 ( \4926 , \4757_nG15ca , \4701 );
nor \U$4225 ( \4927 , \4924 , \4925 , \4926 );
nand \U$4226 ( \4928 , \4920 , \4927 );
xor \U$4227 ( \4929 , \943 , \4353_nGaa0 );
xor \U$4228 ( \4930 , \4929 , \4543 );
xor \U$4229 ( \4931 , \981 , \4382_nGa31 );
xor \U$4230 ( \4932 , \4931 , \4540 );
nor \U$4231 ( \4933 , \4930 , \4932 );
or \U$4232 ( \4934 , \4769 , \4933 );
and \U$4233 ( \4935 , \4928 , \4934 );
and \U$4234 ( \4936 , RIaaa1568_340, \721 );
and \U$4235 ( \4937 , RIaaa17c0_345, \686 );
and \U$4236 ( \4938 , \728 , RIaaa16d0_343);
and \U$4237 ( \4939 , RIaaa19a0_349, \690 );
nor \U$4238 ( \4940 , \4938 , \4939 );
and \U$4239 ( \4941 , RIaaa1310_335, \4572 );
and \U$4240 ( \4942 , \712 , RIaaa1388_336);
and \U$4241 ( \4943 , RIaaa1400_337, \735 );
nor \U$4242 ( \4944 , \4941 , \4942 , \4943 );
and \U$4243 ( \4945 , \733 , RIaaa1838_346);
and \U$4244 ( \4946 , RIaaa14f0_339, \730 );
nor \U$4245 ( \4947 , \4945 , \4946 );
nand \U$4246 ( \4948 , \4940 , \4944 , \4947 );
nor \U$4247 ( \4949 , \4936 , \4937 , \4948 );
and \U$4248 ( \4950 , \702 , RIaaa1928_348);
and \U$4249 ( \4951 , RIaaa15e0_341, \699 );
nor \U$4250 ( \4952 , \4950 , \4951 );
and \U$4251 ( \4953 , \738 , RIaaa1478_338);
and \U$4252 ( \4954 , RIaaa1748_344, \696 );
nor \U$4253 ( \4955 , \4953 , \4954 );
and \U$4254 ( \4956 , \723 , RIaaa1658_342);
and \U$4255 ( \4957 , RIaaa18b0_347, \682 );
nor \U$4256 ( \4958 , \4956 , \4957 );
nand \U$4257 ( \4959 , \4949 , \4952 , \4955 , \4958 );
_DC g12e2 ( \4960_nG12e2 , \4959 , \4592 );
not \U$4258 ( \4961 , \4960_nG12e2 );
nor \U$4259 ( \4962 , \4566 , \4961 );
or \U$4260 ( \4963 , \4646 , \4837 );
not \U$4261 ( \4964 , \4891_nG13e1 );
or \U$4262 ( \4965 , \4964 , \4640 );
or \U$4263 ( \4966 , \4637 , \4837 );
or \U$4264 ( \4967 , \4606 , \4891_nG13e1 );
nand \U$4265 ( \4968 , \4967 , \4642 );
nand \U$4266 ( \4969 , \4966 , \4968 );
nand \U$4267 ( \4970 , \4963 , \4965 , \4969 );
and \U$4268 ( \4971 , \4962 , \4970 );
nor \U$4269 ( \4972 , \4927 , \4920 );
nor \U$4270 ( \4973 , \4935 , \4971 , \4972 );
xnor \U$4271 ( \4974 , \4892 , \4899 );
not \U$4272 ( \4975 , \4974 );
xor \U$4273 ( \4976 , \4865 , \4854 );
not \U$4274 ( \4977 , \4976 );
and \U$4275 ( \4978 , \4975 , \4977 );
and \U$4276 ( \4979 , \4974 , \4976 );
nor \U$4277 ( \4980 , \4978 , \4979 );
nand \U$4278 ( \4981 , \4973 , \4980 );
not \U$4279 ( \4982 , \4934 );
not \U$4280 ( \4983 , \4972 );
nand \U$4281 ( \4984 , \4983 , \4928 );
not \U$4282 ( \4985 , \4984 );
or \U$4283 ( \4986 , \4982 , \4985 );
or \U$4284 ( \4987 , \4984 , \4934 );
nand \U$4285 ( \4988 , \4986 , \4987 );
xor \U$4286 ( \4989 , \4962 , \4970 );
and \U$4287 ( \4990 , \4988 , \4989 );
not \U$4288 ( \4991 , \4930 );
not \U$4289 ( \4992 , \4769 );
or \U$4290 ( \4993 , \4991 , \4992 );
or \U$4291 ( \4994 , \4769 , \4930 );
nand \U$4292 ( \4995 , \4993 , \4994 );
xor \U$4293 ( \4996 , \4932 , \4930 );
nor \U$4294 ( \4997 , \4995 , \4996 );
not \U$4295 ( \4998 , \4997 );
not \U$4296 ( \4999 , \4934 );
nor \U$4297 ( \5000 , \4998 , \4999 );
not \U$4298 ( \5001 , \5000 );
or \U$4299 ( \5002 , \5001 , \4634 );
or \U$4300 ( \5003 , \4998 , \4634 );
nand \U$4301 ( \5004 , \5003 , \4999 );
nand \U$4302 ( \5005 , \5002 , \5004 );
not \U$4303 ( \5006 , \4918 );
or \U$4304 ( \5007 , \5006 , \4594 );
not \U$4305 ( \5008 , \4859 );
or \U$4306 ( \5009 , \4687 , \5008 );
or \U$4307 ( \5010 , \4917 , \4594 );
or \U$4308 ( \5011 , \4771 , \4686_nG16f0 );
nand \U$4309 ( \5012 , \5011 , \4863 );
nand \U$4310 ( \5013 , \5010 , \5012 );
nand \U$4311 ( \5014 , \5007 , \5009 , \5013 );
and \U$4312 ( \5015 , \5005 , \5014 );
and \U$4313 ( \5016 , \4891_nG13e1 , \4645 );
or \U$4314 ( \5017 , \4606 , \4960_nG12e2 );
nand \U$4315 ( \5018 , \5017 , \4642 );
nand \U$4316 ( \5019 , \4891_nG13e1 , \4638 );
and \U$4317 ( \5020 , \5018 , \5019 );
and \U$4318 ( \5021 , \4960_nG12e2 , \4762 );
nor \U$4319 ( \5022 , \5016 , \5020 , \5021 );
nand \U$4320 ( \5023 , \4836_nG14e1 , \4698 );
or \U$4321 ( \5024 , \4659 , \4757_nG15ca );
nand \U$4322 ( \5025 , \5024 , \4725 );
and \U$4323 ( \5026 , \5023 , \5025 );
and \U$4324 ( \5027 , \4728 , \4757_nG15ca );
and \U$4325 ( \5028 , \4836_nG14e1 , \4701 );
nor \U$4326 ( \5029 , \5026 , \5027 , \5028 );
and \U$4327 ( \5030 , \5022 , \5029 );
and \U$4328 ( \5031 , RIaaa2dc8_392, \686 );
and \U$4329 ( \5032 , RIaaa2af8_386, \699 );
and \U$4330 ( \5033 , \728 , RIaaa2a08_384);
and \U$4331 ( \5034 , RIaaa2f30_395, \690 );
nor \U$4332 ( \5035 , \5033 , \5034 );
and \U$4333 ( \5036 , RIaaa3110_399, \4572 );
and \U$4334 ( \5037 , \712 , RIaaa3098_398);
and \U$4335 ( \5038 , RIaaa2be8_388, \735 );
nor \U$4336 ( \5039 , \5036 , \5037 , \5038 );
and \U$4337 ( \5040 , \733 , RIaaa2d50_391);
and \U$4338 ( \5041 , RIaaa2b70_387, \730 );
nor \U$4339 ( \5042 , \5040 , \5041 );
nand \U$4340 ( \5043 , \5035 , \5039 , \5042 );
nor \U$4341 ( \5044 , \5031 , \5032 , \5043 );
and \U$4342 ( \5045 , \696 , RIaaa2e40_393);
and \U$4343 ( \5046 , RIaaa2eb8_394, \721 );
nor \U$4344 ( \5047 , \5045 , \5046 );
and \U$4345 ( \5048 , \738 , RIaaa2c60_389);
and \U$4346 ( \5049 , RIaaa2fa8_396, \702 );
nor \U$4347 ( \5050 , \5048 , \5049 );
and \U$4348 ( \5051 , \723 , RIaaa2a80_385);
and \U$4349 ( \5052 , RIaaa2cd8_390, \682 );
nor \U$4350 ( \5053 , \5051 , \5052 );
nand \U$4351 ( \5054 , \5044 , \5047 , \5050 , \5053 );
_DC g11dc ( \5055_nG11dc , \5054 , \4592 );
nand \U$4352 ( \5056 , \5055_nG11dc , \4565 );
or \U$4353 ( \5057 , \5030 , \5056 );
or \U$4354 ( \5058 , \5022 , \5029 );
nand \U$4355 ( \5059 , \5057 , \5058 );
and \U$4356 ( \5060 , \5015 , \5059 );
and \U$4357 ( \5061 , \4990 , \5060 );
xor \U$4358 ( \5062 , \4981 , \5061 );
not \U$4359 ( \5063 , \4901 );
not \U$4360 ( \5064 , \4846 );
or \U$4361 ( \5065 , \5063 , \5064 );
or \U$4362 ( \5066 , \4846 , \4901 );
nand \U$4363 ( \5067 , \5065 , \5066 );
and \U$4364 ( \5068 , \5062 , \5067 );
and \U$4365 ( \5069 , \4981 , \5061 );
or \U$4366 ( \5070 , \5068 , \5069 );
nor \U$4367 ( \5071 , \4911 , \5070 );
not \U$4368 ( \5072 , \4810 );
not \U$4369 ( \5073 , \4902 );
and \U$4370 ( \5074 , \5072 , \5073 );
and \U$4371 ( \5075 , \4810 , \4902 );
nor \U$4372 ( \5076 , \5074 , \5075 );
nor \U$4373 ( \5077 , \5071 , \5076 );
xor \U$4374 ( \5078 , \4910 , \5077 );
and \U$4375 ( \5079 , \4960_nG12e2 , \4645 );
or \U$4376 ( \5080 , \4606 , \5055_nG11dc );
nand \U$4377 ( \5081 , \5080 , \4642 );
nand \U$4378 ( \5082 , \4960_nG12e2 , \4638 );
and \U$4379 ( \5083 , \5081 , \5082 );
and \U$4380 ( \5084 , \5055_nG11dc , \4762 );
nor \U$4381 ( \5085 , \5079 , \5083 , \5084 );
nand \U$4382 ( \5086 , \4891_nG13e1 , \4698 );
or \U$4383 ( \5087 , \4659 , \4836_nG14e1 );
nand \U$4384 ( \5088 , \5087 , \4725 );
and \U$4385 ( \5089 , \5086 , \5088 );
and \U$4386 ( \5090 , \4728 , \4836_nG14e1 );
and \U$4387 ( \5091 , \4891_nG13e1 , \4701 );
nor \U$4388 ( \5092 , \5089 , \5090 , \5091 );
and \U$4389 ( \5093 , \5085 , \5092 );
not \U$4390 ( \5094 , \5093 );
and \U$4391 ( \5095 , RIaaa2210_367, \686 );
and \U$4392 ( \5096 , RIaaa2738_378, \702 );
and \U$4393 ( \5097 , \728 , RIaaa24e0_373);
and \U$4394 ( \5098 , RIaaa27b0_379, \690 );
nor \U$4395 ( \5099 , \5097 , \5098 );
and \U$4396 ( \5100 , RIaaa28a0_381, \4572 );
and \U$4397 ( \5101 , \712 , RIaaa2918_382);
and \U$4398 ( \5102 , RIaaa2300_369, \733 );
nor \U$4399 ( \5103 , \5100 , \5101 , \5102 );
and \U$4400 ( \5104 , \723 , RIaaa2468_372);
and \U$4401 ( \5105 , RIaaa2558_374, \730 );
nor \U$4402 ( \5106 , \5104 , \5105 );
nand \U$4403 ( \5107 , \5099 , \5103 , \5106 );
nor \U$4404 ( \5108 , \5095 , \5096 , \5107 );
and \U$4405 ( \5109 , \738 , RIaaa2648_376);
and \U$4406 ( \5110 , RIaaa25d0_375, \699 );
nor \U$4407 ( \5111 , \5109 , \5110 );
and \U$4408 ( \5112 , \696 , RIaaa2288_368);
and \U$4409 ( \5113 , RIaaa23f0_371, \721 );
nor \U$4410 ( \5114 , \5112 , \5113 );
and \U$4411 ( \5115 , \735 , RIaaa26c0_377);
and \U$4412 ( \5116 , RIaaa2378_370, \682 );
nor \U$4413 ( \5117 , \5115 , \5116 );
nand \U$4414 ( \5118 , \5108 , \5111 , \5114 , \5117 );
_DC g10fb ( \5119_nG10fb , \5118 , \4592 );
nand \U$4415 ( \5120 , \5119_nG10fb , \4565 );
not \U$4416 ( \5121 , \5120 );
and \U$4417 ( \5122 , \5094 , \5121 );
nor \U$4418 ( \5123 , \5085 , \5092 );
nor \U$4419 ( \5124 , \5122 , \5123 );
and \U$4420 ( \5125 , \4934 , \4996 );
and \U$4421 ( \5126 , \4632_nG1905 , \5125 );
or \U$4422 ( \5127 , \4934 , \4632_nG1905 );
or \U$4423 ( \5128 , \4934 , \4996 );
nand \U$4424 ( \5129 , \5127 , \5128 );
nand \U$4425 ( \5130 , \4593_nG17f6 , \4997 );
and \U$4426 ( \5131 , \5129 , \5130 );
and \U$4427 ( \5132 , \4593_nG17f6 , \5000 );
nor \U$4428 ( \5133 , \5126 , \5131 , \5132 );
nand \U$4429 ( \5134 , \4686_nG16f0 , \4857 );
or \U$4430 ( \5135 , \4771 , \4757_nG15ca );
nand \U$4431 ( \5136 , \5135 , \4863 );
and \U$4432 ( \5137 , \5134 , \5136 );
and \U$4433 ( \5138 , \4859 , \4757_nG15ca );
and \U$4434 ( \5139 , \4686_nG16f0 , \4918 );
nor \U$4435 ( \5140 , \5137 , \5138 , \5139 );
nand \U$4436 ( \5141 , \5133 , \5140 );
xor \U$4437 ( \5142 , \1051 , \4440_nG9d8 );
xor \U$4438 ( \5143 , \5142 , \4534 );
not \U$4439 ( \5144 , \5143 );
xor \U$4440 ( \5145 , \1017 , \4411_nGa2f );
xor \U$4441 ( \5146 , \5145 , \4537 );
not \U$4442 ( \5147 , \5146 );
and \U$4443 ( \5148 , \5144 , \5147 );
or \U$4444 ( \5149 , \4932 , \5148 );
and \U$4445 ( \5150 , \5141 , \5149 );
nor \U$4446 ( \5151 , \5140 , \5133 );
nor \U$4447 ( \5152 , \5150 , \5151 );
nor \U$4448 ( \5153 , \5124 , \5152 );
xor \U$4449 ( \5154 , \5005 , \5014 );
not \U$4450 ( \5155 , \5154 );
not \U$4451 ( \5156 , \5058 );
nor \U$4452 ( \5157 , \5156 , \5030 );
not \U$4453 ( \5158 , \5157 );
not \U$4454 ( \5159 , \5056 );
and \U$4455 ( \5160 , \5158 , \5159 );
and \U$4456 ( \5161 , \5157 , \5056 );
nor \U$4457 ( \5162 , \5160 , \5161 );
nor \U$4458 ( \5163 , \5155 , \5162 );
and \U$4459 ( \5164 , \5153 , \5163 );
xor \U$4460 ( \5165 , \4988 , \4989 );
xor \U$4461 ( \5166 , \5015 , \5059 );
and \U$4462 ( \5167 , \5165 , \5166 );
xor \U$4463 ( \5168 , \5164 , \5167 );
or \U$4464 ( \5169 , \4980 , \4973 );
nand \U$4465 ( \5170 , \5169 , \4981 );
and \U$4466 ( \5171 , \5168 , \5170 );
and \U$4467 ( \5172 , \5164 , \5167 );
or \U$4468 ( \5173 , \5171 , \5172 );
not \U$4469 ( \5174 , \4976 );
nor \U$4470 ( \5175 , \5174 , \4974 );
xor \U$4471 ( \5176 , \5173 , \5175 );
xor \U$4472 ( \5177 , \4981 , \5061 );
xor \U$4473 ( \5178 , \5177 , \5067 );
and \U$4474 ( \5179 , \5176 , \5178 );
and \U$4475 ( \5180 , \5173 , \5175 );
or \U$4476 ( \5181 , \5179 , \5180 );
and \U$4477 ( \5182 , \5071 , \5076 );
nor \U$4478 ( \5183 , \5182 , \5077 );
xor \U$4479 ( \5184 , \5181 , \5183 );
xor \U$4480 ( \5185 , \5173 , \5175 );
xor \U$4481 ( \5186 , \5185 , \5178 );
xnor \U$4482 ( \5187 , \5152 , \5124 );
not \U$4483 ( \5188 , \5162 );
not \U$4484 ( \5189 , \5154 );
and \U$4485 ( \5190 , \5188 , \5189 );
and \U$4486 ( \5191 , \5162 , \5154 );
nor \U$4487 ( \5192 , \5190 , \5191 );
nand \U$4488 ( \5193 , \5187 , \5192 );
not \U$4489 ( \5194 , \5146 );
not \U$4490 ( \5195 , \4932 );
or \U$4491 ( \5196 , \5194 , \5195 );
or \U$4492 ( \5197 , \4932 , \5146 );
nand \U$4493 ( \5198 , \5196 , \5197 );
xor \U$4494 ( \5199 , \5144 , \5147 );
nor \U$4495 ( \5200 , \5198 , \5199 );
not \U$4496 ( \5201 , \5200 );
not \U$4497 ( \5202 , \5149 );
nor \U$4498 ( \5203 , \5201 , \5202 );
not \U$4499 ( \5204 , \5203 );
or \U$4500 ( \5205 , \5204 , \4634 );
or \U$4501 ( \5206 , \5201 , \4634 );
nand \U$4502 ( \5207 , \5206 , \5202 );
nand \U$4503 ( \5208 , \5205 , \5207 );
not \U$4504 ( \5209 , \5125 );
or \U$4505 ( \5210 , \5209 , \4594 );
or \U$4506 ( \5211 , \4687 , \5001 );
or \U$4507 ( \5212 , \4998 , \4687 );
or \U$4508 ( \5213 , \4934 , \4593_nG17f6 );
nand \U$4509 ( \5214 , \5213 , \5128 );
nand \U$4510 ( \5215 , \5212 , \5214 );
nand \U$4511 ( \5216 , \5210 , \5211 , \5215 );
and \U$4512 ( \5217 , \5208 , \5216 );
nand \U$4513 ( \5218 , \4960_nG12e2 , \4698 );
or \U$4514 ( \5219 , \4659 , \4891_nG13e1 );
nand \U$4515 ( \5220 , \5219 , \4725 );
and \U$4516 ( \5221 , \5218 , \5220 );
and \U$4517 ( \5222 , \4728 , \4891_nG13e1 );
and \U$4518 ( \5223 , \4960_nG12e2 , \4701 );
nor \U$4519 ( \5224 , \5221 , \5222 , \5223 );
nand \U$4520 ( \5225 , \4757_nG15ca , \4857 );
or \U$4521 ( \5226 , \4771 , \4836_nG14e1 );
nand \U$4522 ( \5227 , \5226 , \4863 );
and \U$4523 ( \5228 , \5225 , \5227 );
and \U$4524 ( \5229 , \4859 , \4836_nG14e1 );
and \U$4525 ( \5230 , \4757_nG15ca , \4918 );
nor \U$4526 ( \5231 , \5228 , \5229 , \5230 );
xor \U$4527 ( \5232 , \5224 , \5231 );
and \U$4528 ( \5233 , \5055_nG11dc , \4645 );
or \U$4529 ( \5234 , \4606 , \5119_nG10fb );
nand \U$4530 ( \5235 , \5234 , \4642 );
nand \U$4531 ( \5236 , \5055_nG11dc , \4638 );
and \U$4532 ( \5237 , \5235 , \5236 );
and \U$4533 ( \5238 , \5119_nG10fb , \4762 );
nor \U$4534 ( \5239 , \5233 , \5237 , \5238 );
and \U$4535 ( \5240 , \5232 , \5239 );
and \U$4536 ( \5241 , \5224 , \5231 );
or \U$4537 ( \5242 , \5240 , \5241 );
not \U$4538 ( \5243 , \5242 );
and \U$4539 ( \5244 , \5217 , \5243 );
not \U$4540 ( \5245 , \5149 );
not \U$4541 ( \5246 , \5151 );
nand \U$4542 ( \5247 , \5246 , \5141 );
not \U$4543 ( \5248 , \5247 );
or \U$4544 ( \5249 , \5245 , \5248 );
or \U$4545 ( \5250 , \5247 , \5149 );
nand \U$4546 ( \5251 , \5249 , \5250 );
not \U$4547 ( \5252 , \5120 );
nor \U$4548 ( \5253 , \5093 , \5123 );
not \U$4549 ( \5254 , \5253 );
or \U$4550 ( \5255 , \5252 , \5254 );
or \U$4551 ( \5256 , \5253 , \5120 );
nand \U$4552 ( \5257 , \5255 , \5256 );
and \U$4553 ( \5258 , \5251 , \5257 );
and \U$4554 ( \5259 , \5244 , \5258 );
xor \U$4555 ( \5260 , \5193 , \5259 );
xor \U$4556 ( \5261 , \5165 , \5166 );
and \U$4557 ( \5262 , \5260 , \5261 );
and \U$4558 ( \5263 , \5193 , \5259 );
or \U$4559 ( \5264 , \5262 , \5263 );
xor \U$4560 ( \5265 , \4990 , \5060 );
xor \U$4561 ( \5266 , \5264 , \5265 );
xor \U$4562 ( \5267 , \5164 , \5167 );
xor \U$4563 ( \5268 , \5267 , \5170 );
and \U$4564 ( \5269 , \5266 , \5268 );
and \U$4565 ( \5270 , \5264 , \5265 );
or \U$4566 ( \5271 , \5269 , \5270 );
xor \U$4567 ( \5272 , \5186 , \5271 );
xor \U$4568 ( \5273 , \5217 , \5243 );
xor \U$4569 ( \5274 , \5251 , \5257 );
and \U$4570 ( \5275 , \5273 , \5274 );
xor \U$4571 ( \5276 , \5208 , \5216 );
xor \U$4572 ( \5277 , \5224 , \5231 );
xor \U$4573 ( \5278 , \5277 , \5239 );
not \U$4574 ( \5279 , \5278 );
and \U$4575 ( \5280 , \5276 , \5279 );
xor \U$4576 ( \5281 , RIaa977e8_4, \4498_nG969 );
xor \U$4577 ( \5282 , \5281 , \4528 );
not \U$4578 ( \5283 , \5282 );
xor \U$4579 ( \5284 , \1087 , \4469_nG9da );
xor \U$4580 ( \5285 , \5284 , \4531 );
not \U$4581 ( \5286 , \5285 );
and \U$4582 ( \5287 , \5283 , \5286 );
or \U$4583 ( \5288 , \5143 , \5287 );
not \U$4584 ( \5289 , \5288 );
nand \U$4585 ( \5290 , \4593_nG17f6 , \5200 );
or \U$4586 ( \5291 , \5149 , \4632_nG1905 );
or \U$4587 ( \5292 , \5149 , \5199 );
nand \U$4588 ( \5293 , \5291 , \5292 );
and \U$4589 ( \5294 , \5290 , \5293 );
and \U$4590 ( \5295 , \5149 , \5199 );
and \U$4591 ( \5296 , \5295 , \4632_nG1905 );
and \U$4592 ( \5297 , \4593_nG17f6 , \5203 );
nor \U$4593 ( \5298 , \5294 , \5296 , \5297 );
and \U$4594 ( \5299 , \4686_nG16f0 , \5125 );
or \U$4595 ( \5300 , \4934 , \4686_nG16f0 );
nand \U$4596 ( \5301 , \5300 , \5128 );
nand \U$4597 ( \5302 , \4757_nG15ca , \4997 );
and \U$4598 ( \5303 , \5301 , \5302 );
and \U$4599 ( \5304 , \4757_nG15ca , \5000 );
nor \U$4600 ( \5305 , \5299 , \5303 , \5304 );
nand \U$4601 ( \5306 , \5298 , \5305 );
not \U$4602 ( \5307 , \5306 );
or \U$4603 ( \5308 , \5289 , \5307 );
or \U$4604 ( \5309 , \5305 , \5298 );
nand \U$4605 ( \5310 , \5308 , \5309 );
nand \U$4606 ( \5311 , \5055_nG11dc , \4698 );
or \U$4607 ( \5312 , \4659 , \4960_nG12e2 );
nand \U$4608 ( \5313 , \5312 , \4725 );
and \U$4609 ( \5314 , \5311 , \5313 );
and \U$4610 ( \5315 , \4728 , \4960_nG12e2 );
and \U$4611 ( \5316 , \5055_nG11dc , \4701 );
nor \U$4612 ( \5317 , \5314 , \5315 , \5316 );
nand \U$4613 ( \5318 , \4836_nG14e1 , \4857 );
or \U$4614 ( \5319 , \4771 , \4891_nG13e1 );
nand \U$4615 ( \5320 , \5319 , \4863 );
and \U$4616 ( \5321 , \5318 , \5320 );
and \U$4617 ( \5322 , \4859 , \4891_nG13e1 );
and \U$4618 ( \5323 , \4836_nG14e1 , \4918 );
nor \U$4619 ( \5324 , \5321 , \5322 , \5323 );
xor \U$4620 ( \5325 , \5317 , \5324 );
and \U$4621 ( \5326 , \5119_nG10fb , \4645 );
and \U$4622 ( \5327 , RIaaa3d40_425, \686 );
and \U$4623 ( \5328 , RIaaa3f20_429, \738 );
and \U$4624 ( \5329 , \682 , RIaaa3b60_421);
and \U$4625 ( \5330 , RIaaa3a70_419, \728 );
nor \U$4626 ( \5331 , \5329 , \5330 );
and \U$4627 ( \5332 , RIaaa4100_433, \4572 );
and \U$4628 ( \5333 , \712 , RIaaa4178_434);
and \U$4629 ( \5334 , RIaaa4010_431, \699 );
nor \U$4630 ( \5335 , \5332 , \5333 , \5334 );
and \U$4631 ( \5336 , \702 , RIaaa3bd8_422);
and \U$4632 ( \5337 , RIaaa3c50_423, \690 );
nor \U$4633 ( \5338 , \5336 , \5337 );
nand \U$4634 ( \5339 , \5331 , \5335 , \5338 );
nor \U$4635 ( \5340 , \5327 , \5328 , \5339 );
and \U$4636 ( \5341 , \696 , RIaaa3cc8_424);
and \U$4637 ( \5342 , RIaaa3e30_427, \735 );
nor \U$4638 ( \5343 , \5341 , \5342 );
and \U$4639 ( \5344 , \721 , RIaaa3f98_430);
and \U$4640 ( \5345 , RIaaa3ae8_420, \733 );
nor \U$4641 ( \5346 , \5344 , \5345 );
and \U$4642 ( \5347 , \723 , RIaaa39f8_418);
and \U$4643 ( \5348 , RIaaa3ea8_428, \730 );
nor \U$4644 ( \5349 , \5347 , \5348 );
nand \U$4645 ( \5350 , \5340 , \5343 , \5346 , \5349 );
_DC gffe ( \5351_nGffe , \5350 , \4592 );
or \U$4646 ( \5352 , \4606 , \5351_nGffe );
nand \U$4647 ( \5353 , \5352 , \4642 );
nand \U$4648 ( \5354 , \5119_nG10fb , \4638 );
and \U$4649 ( \5355 , \5353 , \5354 );
and \U$4650 ( \5356 , \5351_nGffe , \4762 );
nor \U$4651 ( \5357 , \5326 , \5355 , \5356 );
and \U$4652 ( \5358 , \5325 , \5357 );
and \U$4653 ( \5359 , \5317 , \5324 );
or \U$4654 ( \5360 , \5358 , \5359 );
not \U$4655 ( \5361 , \5360 );
and \U$4656 ( \5362 , \5310 , \5361 );
and \U$4657 ( \5363 , \5280 , \5362 );
xor \U$4658 ( \5364 , \5275 , \5363 );
or \U$4659 ( \5365 , \5192 , \5187 );
nand \U$4660 ( \5366 , \5365 , \5193 );
and \U$4661 ( \5367 , \5364 , \5366 );
and \U$4662 ( \5368 , \5275 , \5363 );
or \U$4663 ( \5369 , \5367 , \5368 );
xor \U$4664 ( \5370 , \5153 , \5163 );
xor \U$4665 ( \5371 , \5369 , \5370 );
xor \U$4666 ( \5372 , \5193 , \5259 );
xor \U$4667 ( \5373 , \5372 , \5261 );
and \U$4668 ( \5374 , \5371 , \5373 );
and \U$4669 ( \5375 , \5369 , \5370 );
or \U$4670 ( \5376 , \5374 , \5375 );
xor \U$4671 ( \5377 , \5264 , \5265 );
xor \U$4672 ( \5378 , \5377 , \5268 );
xor \U$4673 ( \5379 , \5376 , \5378 );
xor \U$4674 ( \5380 , \5369 , \5370 );
xor \U$4675 ( \5381 , \5380 , \5373 );
xor \U$4676 ( \5382 , \5276 , \5279 );
nand \U$4677 ( \5383 , \5351_nGffe , \4565 );
and \U$4678 ( \5384 , \5382 , \5383 );
xor \U$4679 ( \5385 , \5310 , \5361 );
nor \U$4680 ( \5386 , \5384 , \5385 );
not \U$4681 ( \5387 , \5386 );
or \U$4682 ( \5388 , \5143 , \5285 );
nand \U$4683 ( \5389 , \5285 , \5143 );
nand \U$4684 ( \5390 , \5388 , \5389 );
xor \U$4685 ( \5391 , \5283 , \5286 );
nor \U$4686 ( \5392 , \5390 , \5391 );
not \U$4687 ( \5393 , \5392 );
not \U$4688 ( \5394 , \5288 );
nor \U$4689 ( \5395 , \5393 , \5394 );
not \U$4690 ( \5396 , \5395 );
or \U$4691 ( \5397 , \5396 , \4634 );
or \U$4692 ( \5398 , \5393 , \4634 );
nand \U$4693 ( \5399 , \5398 , \5394 );
nand \U$4694 ( \5400 , \5397 , \5399 );
not \U$4695 ( \5401 , \5400 );
nand \U$4696 ( \5402 , \4686_nG16f0 , \5200 );
or \U$4697 ( \5403 , \5149 , \4593_nG17f6 );
nand \U$4698 ( \5404 , \5403 , \5292 );
and \U$4699 ( \5405 , \5402 , \5404 );
and \U$4700 ( \5406 , \5295 , \4593_nG17f6 );
and \U$4701 ( \5407 , \4686_nG16f0 , \5203 );
nor \U$4702 ( \5408 , \5405 , \5406 , \5407 );
nor \U$4703 ( \5409 , \5401 , \5408 );
not \U$4704 ( \5410 , \5409 );
nand \U$4705 ( \5411 , \4891_nG13e1 , \4857 );
or \U$4706 ( \5412 , \4771 , \4960_nG12e2 );
nand \U$4707 ( \5413 , \5412 , \4863 );
and \U$4708 ( \5414 , \5411 , \5413 );
and \U$4709 ( \5415 , \4859 , \4960_nG12e2 );
and \U$4710 ( \5416 , \4891_nG13e1 , \4918 );
nor \U$4711 ( \5417 , \5414 , \5415 , \5416 );
and \U$4712 ( \5418 , \4757_nG15ca , \5125 );
or \U$4713 ( \5419 , \4934 , \4757_nG15ca );
nand \U$4714 ( \5420 , \5419 , \5128 );
nand \U$4715 ( \5421 , \4836_nG14e1 , \4997 );
and \U$4716 ( \5422 , \5420 , \5421 );
and \U$4717 ( \5423 , \4836_nG14e1 , \5000 );
nor \U$4718 ( \5424 , \5418 , \5422 , \5423 );
xor \U$4719 ( \5425 , \5417 , \5424 );
nand \U$4720 ( \5426 , \5119_nG10fb , \4698 );
or \U$4721 ( \5427 , \4659 , \5055_nG11dc );
nand \U$4722 ( \5428 , \5427 , \4725 );
and \U$4723 ( \5429 , \5426 , \5428 );
and \U$4724 ( \5430 , \4728 , \5055_nG11dc );
and \U$4725 ( \5431 , \5119_nG10fb , \4701 );
nor \U$4726 ( \5432 , \5429 , \5430 , \5431 );
and \U$4727 ( \5433 , \5425 , \5432 );
and \U$4728 ( \5434 , \5417 , \5424 );
or \U$4729 ( \5435 , \5433 , \5434 );
nor \U$4730 ( \5436 , \5410 , \5435 );
xor \U$4731 ( \5437 , \5317 , \5324 );
xor \U$4732 ( \5438 , \5437 , \5357 );
nand \U$4733 ( \5439 , \5306 , \5309 );
not \U$4734 ( \5440 , \5439 );
not \U$4735 ( \5441 , \5288 );
and \U$4736 ( \5442 , \5440 , \5441 );
and \U$4737 ( \5443 , \5439 , \5288 );
nor \U$4738 ( \5444 , \5442 , \5443 );
nor \U$4739 ( \5445 , \5438 , \5444 );
not \U$4740 ( \5446 , \5445 );
and \U$4741 ( \5447 , RIaaa3890_415, \728 );
and \U$4742 ( \5448 , RIaaa3368_404, \738 );
and \U$4743 ( \5449 , \682 , RIaaa37a0_413);
and \U$4744 ( \5450 , RIaaa36b0_411, \690 );
nor \U$4745 ( \5451 , \5449 , \5450 );
and \U$4746 ( \5452 , RIaaa3548_408, \4572 );
and \U$4747 ( \5453 , \712 , RIaaa35c0_409);
and \U$4748 ( \5454 , RIaaa3278_402, \735 );
nor \U$4749 ( \5455 , \5452 , \5453 , \5454 );
and \U$4750 ( \5456 , \696 , RIaaa3908_416);
and \U$4751 ( \5457 , RIaaa3980_417, \686 );
nor \U$4752 ( \5458 , \5456 , \5457 );
nand \U$4753 ( \5459 , \5451 , \5455 , \5458 );
nor \U$4754 ( \5460 , \5447 , \5448 , \5459 );
and \U$4755 ( \5461 , \702 , RIaaa3638_410);
and \U$4756 ( \5462 , RIaaa33e0_405, \721 );
nor \U$4757 ( \5463 , \5461 , \5462 );
and \U$4758 ( \5464 , \733 , RIaaa3728_412);
and \U$4759 ( \5465 , RIaaa3458_406, \699 );
nor \U$4760 ( \5466 , \5464 , \5465 );
and \U$4761 ( \5467 , \723 , RIaaa3818_414);
and \U$4762 ( \5468 , RIaaa32f0_403, \730 );
nor \U$4763 ( \5469 , \5467 , \5468 );
nand \U$4764 ( \5470 , \5460 , \5463 , \5466 , \5469 );
_DC gf21 ( \5471_nGf21 , \5470 , \4592 );
nand \U$4765 ( \5472 , \5471_nGf21 , \4565 );
nand \U$4766 ( \5473 , \5446 , \5472 );
and \U$4767 ( \5474 , \5436 , \5473 );
xor \U$4768 ( \5475 , \5387 , \5474 );
xor \U$4769 ( \5476 , \5273 , \5274 );
and \U$4770 ( \5477 , \5475 , \5476 );
and \U$4771 ( \5478 , \5387 , \5474 );
or \U$4772 ( \5479 , \5477 , \5478 );
xor \U$4773 ( \5480 , \5244 , \5258 );
xor \U$4774 ( \5481 , \5479 , \5480 );
xor \U$4775 ( \5482 , \5275 , \5363 );
xor \U$4776 ( \5483 , \5482 , \5366 );
and \U$4777 ( \5484 , \5481 , \5483 );
and \U$4778 ( \5485 , \5479 , \5480 );
or \U$4779 ( \5486 , \5484 , \5485 );
xor \U$4780 ( \5487 , \5381 , \5486 );
xor \U$4781 ( \5488 , \5479 , \5480 );
xor \U$4782 ( \5489 , \5488 , \5483 );
not \U$4783 ( \5490 , \5280 );
not \U$4784 ( \5491 , \5383 );
nor \U$4785 ( \5492 , \5491 , \5362 );
not \U$4786 ( \5493 , \5492 );
or \U$4787 ( \5494 , \5490 , \5493 );
or \U$4788 ( \5495 , \5280 , \5492 );
nand \U$4789 ( \5496 , \5494 , \5495 );
xor \U$4790 ( \5497 , \5387 , \5474 );
xor \U$4791 ( \5498 , \5497 , \5476 );
and \U$4792 ( \5499 , \5496 , \5498 );
or \U$4793 ( \5500 , \5435 , \5409 );
and \U$4794 ( \5501 , \4572 , RIaaa42e0_437);
and \U$4795 ( \5502 , \735 , RIaaa43d0_439);
and \U$4796 ( \5503 , RIaaa4880_449, \682 );
nor \U$4797 ( \5504 , \5502 , \5503 );
and \U$4798 ( \5505 , \738 , RIaaa4448_440);
and \U$4799 ( \5506 , RIaaa45b0_443, \699 );
nor \U$4800 ( \5507 , \5505 , \5506 );
and \U$4801 ( \5508 , \702 , RIaaa48f8_450);
and \U$4802 ( \5509 , RIaaa4538_442, \721 );
nor \U$4803 ( \5510 , \5508 , \5509 );
and \U$4804 ( \5511 , \696 , RIaaa4718_446);
and \U$4805 ( \5512 , RIaaa4790_447, \686 );
nor \U$4806 ( \5513 , \5511 , \5512 );
nand \U$4807 ( \5514 , \5504 , \5507 , \5510 , \5513 );
nor \U$4808 ( \5515 , \5501 , \5514 );
and \U$4809 ( \5516 , \723 , RIaaa4628_444);
and \U$4810 ( \5517 , RIaaa4970_451, \690 );
nor \U$4811 ( \5518 , \5516 , \5517 );
and \U$4812 ( \5519 , \733 , RIaaa4808_448);
and \U$4813 ( \5520 , RIaaa44c0_441, \730 );
nor \U$4814 ( \5521 , \5519 , \5520 );
and \U$4815 ( \5522 , \728 , RIaaa46a0_445);
and \U$4816 ( \5523 , RIaaa4358_438, \712 );
nor \U$4817 ( \5524 , \5522 , \5523 );
nand \U$4818 ( \5525 , \5515 , \5518 , \5521 , \5524 );
_DC ge53 ( \5526_nGe53 , \5525 , \4592 );
nand \U$4819 ( \5527 , \5526_nGe53 , \4565 );
and \U$4820 ( \5528 , \5351_nGffe , \4645 );
or \U$4821 ( \5529 , \4606 , \5471_nGf21 );
nand \U$4822 ( \5530 , \5529 , \4642 );
nand \U$4823 ( \5531 , \5351_nGffe , \4638 );
and \U$4824 ( \5532 , \5530 , \5531 );
and \U$4825 ( \5533 , \5471_nGf21 , \4762 );
nor \U$4826 ( \5534 , \5528 , \5532 , \5533 );
or \U$4827 ( \5535 , \5527 , \5534 );
nand \U$4828 ( \5536 , \5409 , \5435 );
nand \U$4829 ( \5537 , \5500 , \5535 , \5536 );
not \U$4830 ( \5538 , \5537 );
and \U$4831 ( \5539 , \5438 , \5444 );
nor \U$4832 ( \5540 , \5539 , \5445 );
not \U$4833 ( \5541 , \5540 );
not \U$4834 ( \5542 , \5472 );
and \U$4835 ( \5543 , \5541 , \5542 );
and \U$4836 ( \5544 , \5540 , \5472 );
nor \U$4837 ( \5545 , \5543 , \5544 );
nor \U$4838 ( \5546 , \5538 , \5545 );
nand \U$4839 ( \5547 , \4960_nG12e2 , \4857 );
or \U$4840 ( \5548 , \4771 , \5055_nG11dc );
nand \U$4841 ( \5549 , \5548 , \4863 );
and \U$4842 ( \5550 , \5547 , \5549 );
and \U$4843 ( \5551 , \4859 , \5055_nG11dc );
and \U$4844 ( \5552 , \4960_nG12e2 , \4918 );
nor \U$4845 ( \5553 , \5550 , \5551 , \5552 );
and \U$4846 ( \5554 , \4836_nG14e1 , \5125 );
or \U$4847 ( \5555 , \4934 , \4836_nG14e1 );
nand \U$4848 ( \5556 , \5555 , \5128 );
nand \U$4849 ( \5557 , \4891_nG13e1 , \4997 );
and \U$4850 ( \5558 , \5556 , \5557 );
and \U$4851 ( \5559 , \4891_nG13e1 , \5000 );
nor \U$4852 ( \5560 , \5554 , \5558 , \5559 );
xor \U$4853 ( \5561 , \5553 , \5560 );
nand \U$4854 ( \5562 , \5351_nGffe , \4698 );
or \U$4855 ( \5563 , \4659 , \5119_nG10fb );
nand \U$4856 ( \5564 , \5563 , \4725 );
and \U$4857 ( \5565 , \5562 , \5564 );
and \U$4858 ( \5566 , \4728 , \5119_nG10fb );
and \U$4859 ( \5567 , \5351_nGffe , \4701 );
nor \U$4860 ( \5568 , \5565 , \5566 , \5567 );
and \U$4861 ( \5569 , \5561 , \5568 );
and \U$4862 ( \5570 , \5553 , \5560 );
or \U$4863 ( \5571 , \5569 , \5570 );
nand \U$4864 ( \5572 , \4593_nG17f6 , \5392 );
or \U$4865 ( \5573 , \5288 , \4632_nG1905 );
or \U$4866 ( \5574 , \5288 , \5391 );
nand \U$4867 ( \5575 , \5573 , \5574 );
and \U$4868 ( \5576 , \5572 , \5575 );
and \U$4869 ( \5577 , \5288 , \5391 );
and \U$4870 ( \5578 , \5577 , \4632_nG1905 );
and \U$4871 ( \5579 , \4593_nG17f6 , \5395 );
nor \U$4872 ( \5580 , \5576 , \5578 , \5579 );
xor \U$4873 ( \5581 , \5580 , \5283 );
nand \U$4874 ( \5582 , \4757_nG15ca , \5200 );
or \U$4875 ( \5583 , \5149 , \4686_nG16f0 );
nand \U$4876 ( \5584 , \5583 , \5292 );
and \U$4877 ( \5585 , \5582 , \5584 );
and \U$4878 ( \5586 , \5295 , \4686_nG16f0 );
and \U$4879 ( \5587 , \4757_nG15ca , \5203 );
nor \U$4880 ( \5588 , \5585 , \5586 , \5587 );
and \U$4881 ( \5589 , \5581 , \5588 );
and \U$4882 ( \5590 , \5580 , \5283 );
or \U$4883 ( \5591 , \5589 , \5590 );
nor \U$4884 ( \5592 , \5571 , \5591 );
not \U$4885 ( \5593 , \5592 );
xor \U$4886 ( \5594 , \5417 , \5424 );
xor \U$4887 ( \5595 , \5594 , \5432 );
not \U$4888 ( \5596 , \5408 );
not \U$4889 ( \5597 , \5400 );
and \U$4890 ( \5598 , \5596 , \5597 );
and \U$4891 ( \5599 , \5408 , \5400 );
nor \U$4892 ( \5600 , \5598 , \5599 );
xor \U$4893 ( \5601 , \5595 , \5600 );
xnor \U$4894 ( \5602 , \5527 , \5534 );
and \U$4895 ( \5603 , \5601 , \5602 );
and \U$4896 ( \5604 , \5595 , \5600 );
or \U$4897 ( \5605 , \5603 , \5604 );
nor \U$4898 ( \5606 , \5593 , \5605 );
xor \U$4899 ( \5607 , \5546 , \5606 );
not \U$4900 ( \5608 , \5385 );
xnor \U$4901 ( \5609 , \5383 , \5382 );
not \U$4902 ( \5610 , \5609 );
or \U$4903 ( \5611 , \5608 , \5610 );
or \U$4904 ( \5612 , \5609 , \5385 );
nand \U$4905 ( \5613 , \5611 , \5612 );
and \U$4906 ( \5614 , \5607 , \5613 );
and \U$4907 ( \5615 , \5546 , \5606 );
or \U$4908 ( \5616 , \5614 , \5615 );
xor \U$4909 ( \5617 , \5387 , \5474 );
xor \U$4910 ( \5618 , \5617 , \5476 );
and \U$4911 ( \5619 , \5616 , \5618 );
and \U$4912 ( \5620 , \5496 , \5616 );
or \U$4913 ( \5621 , \5499 , \5619 , \5620 );
xor \U$4914 ( \5622 , \5489 , \5621 );
xor \U$4915 ( \5623 , \5387 , \5474 );
xor \U$4916 ( \5624 , \5623 , \5476 );
xor \U$4917 ( \5625 , \5496 , \5616 );
xor \U$4918 ( \5626 , \5624 , \5625 );
xor \U$4919 ( \5627 , \5436 , \5473 );
xor \U$4920 ( \5628 , \5546 , \5606 );
xor \U$4921 ( \5629 , \5628 , \5613 );
nand \U$4922 ( \5630 , \5627 , \5629 );
and \U$4923 ( \5631 , \690 , RIaaa6770_515);
and \U$4924 ( \5632 , \723 , RIaaa6860_517);
and \U$4925 ( \5633 , RIaaa64a0_509, \730 );
nor \U$4926 ( \5634 , \5632 , \5633 );
and \U$4927 ( \5635 , \696 , RIaaa68d8_518);
and \U$4928 ( \5636 , RIaaa6518_510, \699 );
nor \U$4929 ( \5637 , \5635 , \5636 );
and \U$4930 ( \5638 , \738 , RIaaa6428_508);
and \U$4931 ( \5639 , RIaaa6590_511, \721 );
nor \U$4932 ( \5640 , \5638 , \5639 );
and \U$4933 ( \5641 , \702 , RIaaa66f8_514);
and \U$4934 ( \5642 , RIaaa6950_519, \686 );
nor \U$4935 ( \5643 , \5641 , \5642 );
nand \U$4936 ( \5644 , \5634 , \5637 , \5640 , \5643 );
nor \U$4937 ( \5645 , \5631 , \5644 );
and \U$4938 ( \5646 , \682 , RIaaa6608_512);
and \U$4939 ( \5647 , RIaaa67e8_516, \728 );
nor \U$4940 ( \5648 , \5646 , \5647 );
and \U$4941 ( \5649 , \735 , RIaaa63b0_507);
and \U$4942 ( \5650 , RIaaa6338_506, \712 );
nor \U$4943 ( \5651 , \5649 , \5650 );
and \U$4944 ( \5652 , \4572 , RIaaa62c0_505);
and \U$4945 ( \5653 , RIaaa6680_513, \733 );
nor \U$4946 ( \5654 , \5652 , \5653 );
nand \U$4947 ( \5655 , \5645 , \5648 , \5651 , \5654 );
_DC gaf0 ( \5656_nGaf0 , \5655 , \4592 );
nand \U$4948 ( \5657 , \5656_nGaf0 , \4565 );
and \U$4949 ( \5658 , \5471_nGf21 , \4645 );
or \U$4950 ( \5659 , \4606 , \5526_nGe53 );
nand \U$4951 ( \5660 , \5659 , \4642 );
nand \U$4952 ( \5661 , \5471_nGf21 , \4638 );
and \U$4953 ( \5662 , \5660 , \5661 );
and \U$4954 ( \5663 , \5526_nGe53 , \4762 );
nor \U$4955 ( \5664 , \5658 , \5662 , \5663 );
xnor \U$4956 ( \5665 , \5657 , \5664 );
xor \U$4957 ( \5666 , \5595 , \5600 );
xor \U$4958 ( \5667 , \5666 , \5602 );
and \U$4959 ( \5668 , \5665 , \5667 );
and \U$4960 ( \5669 , \4891_nG13e1 , \5125 );
or \U$4961 ( \5670 , \4934 , \4891_nG13e1 );
nand \U$4962 ( \5671 , \5670 , \5128 );
nand \U$4963 ( \5672 , \4960_nG12e2 , \4997 );
and \U$4964 ( \5673 , \5671 , \5672 );
and \U$4965 ( \5674 , \4960_nG12e2 , \5000 );
nor \U$4966 ( \5675 , \5669 , \5673 , \5674 );
nand \U$4967 ( \5676 , \4836_nG14e1 , \5200 );
or \U$4968 ( \5677 , \5149 , \4757_nG15ca );
nand \U$4969 ( \5678 , \5677 , \5292 );
and \U$4970 ( \5679 , \5676 , \5678 );
and \U$4971 ( \5680 , \5295 , \4757_nG15ca );
and \U$4972 ( \5681 , \4836_nG14e1 , \5203 );
nor \U$4973 ( \5682 , \5679 , \5680 , \5681 );
xor \U$4974 ( \5683 , \5675 , \5682 );
nand \U$4975 ( \5684 , \5055_nG11dc , \4857 );
or \U$4976 ( \5685 , \4771 , \5119_nG10fb );
nand \U$4977 ( \5686 , \5685 , \4863 );
and \U$4978 ( \5687 , \5684 , \5686 );
and \U$4979 ( \5688 , \4859 , \5119_nG10fb );
and \U$4980 ( \5689 , \5055_nG11dc , \4918 );
nor \U$4981 ( \5690 , \5687 , \5688 , \5689 );
and \U$4982 ( \5691 , \5683 , \5690 );
and \U$4983 ( \5692 , \5675 , \5682 );
or \U$4984 ( \5693 , \5691 , \5692 );
nand \U$4985 ( \5694 , \4686_nG16f0 , \5392 );
or \U$4986 ( \5695 , \5288 , \4593_nG17f6 );
nand \U$4987 ( \5696 , \5695 , \5574 );
and \U$4988 ( \5697 , \5694 , \5696 );
and \U$4989 ( \5698 , \5577 , \4593_nG17f6 );
and \U$4990 ( \5699 , \4686_nG16f0 , \5395 );
nor \U$4991 ( \5700 , \5697 , \5698 , \5699 );
not \U$4992 ( \5701 , \5700 );
or \U$4993 ( \5702 , \5282 , \4632_nG1905 );
or \U$4994 ( \5703 , \1182 , \4526_nG967 );
nand \U$4995 ( \5704 , \5703 , \4527 );
nor \U$4996 ( \5705 , \5282 , \5704 );
not \U$4997 ( \5706 , \5705 );
nand \U$4998 ( \5707 , \5283 , \5706 );
nand \U$4999 ( \5708 , \5702 , \5707 );
nand \U$5000 ( \5709 , \5701 , \5708 );
xor \U$5001 ( \5710 , \5693 , \5709 );
and \U$5002 ( \5711 , \5526_nGe53 , \4645 );
or \U$5003 ( \5712 , \4606 , \5656_nGaf0 );
nand \U$5004 ( \5713 , \5712 , \4642 );
nand \U$5005 ( \5714 , \5526_nGe53 , \4638 );
and \U$5006 ( \5715 , \5713 , \5714 );
and \U$5007 ( \5716 , \5656_nGaf0 , \4762 );
nor \U$5008 ( \5717 , \5711 , \5715 , \5716 );
nand \U$5009 ( \5718 , \5471_nGf21 , \4698 );
or \U$5010 ( \5719 , \4659 , \5351_nGffe );
nand \U$5011 ( \5720 , \5719 , \4725 );
and \U$5012 ( \5721 , \5718 , \5720 );
and \U$5013 ( \5722 , \4728 , \5351_nGffe );
and \U$5014 ( \5723 , \5471_nGf21 , \4701 );
nor \U$5015 ( \5724 , \5721 , \5722 , \5723 );
and \U$5016 ( \5725 , \5717 , \5724 );
not \U$5017 ( \5726 , \5725 );
and \U$5018 ( \5727 , RIaaa58e8_484, \686 );
and \U$5019 ( \5728 , RIaaa5438_474, \699 );
and \U$5020 ( \5729 , \728 , RIaaa5690_479);
and \U$5021 ( \5730 , RIaaa5870_483, \690 );
nor \U$5022 ( \5731 , \5729 , \5730 );
and \U$5023 ( \5732 , RIaaa55a0_477, \4572 );
and \U$5024 ( \5733 , \712 , RIaaa5528_476);
and \U$5025 ( \5734 , RIaaa5258_470, \735 );
nor \U$5026 ( \5735 , \5732 , \5733 , \5734 );
and \U$5027 ( \5736 , \733 , RIaaa5708_480);
and \U$5028 ( \5737 , RIaaa52d0_471, \730 );
nor \U$5029 ( \5738 , \5736 , \5737 );
nand \U$5030 ( \5739 , \5731 , \5735 , \5738 );
nor \U$5031 ( \5740 , \5727 , \5728 , \5739 );
and \U$5032 ( \5741 , \696 , RIaaa5960_485);
and \U$5033 ( \5742 , RIaaa53c0_473, \721 );
nor \U$5034 ( \5743 , \5741 , \5742 );
and \U$5035 ( \5744 , \738 , RIaaa5348_472);
and \U$5036 ( \5745 , RIaaa57f8_482, \702 );
nor \U$5037 ( \5746 , \5744 , \5745 );
and \U$5038 ( \5747 , \723 , RIaaa5618_478);
and \U$5039 ( \5748 , RIaaa5780_481, \682 );
nor \U$5040 ( \5749 , \5747 , \5748 );
nand \U$5041 ( \5750 , \5740 , \5743 , \5746 , \5749 );
_DC gabb ( \5751_nGabb , \5750 , \4592 );
nand \U$5042 ( \5752 , \5751_nGabb , \4565 );
not \U$5043 ( \5753 , \5752 );
and \U$5044 ( \5754 , \5726 , \5753 );
nor \U$5045 ( \5755 , \5717 , \5724 );
nor \U$5046 ( \5756 , \5754 , \5755 );
and \U$5047 ( \5757 , \5710 , \5756 );
and \U$5048 ( \5758 , \5693 , \5709 );
or \U$5049 ( \5759 , \5757 , \5758 );
xor \U$5050 ( \5760 , \5595 , \5600 );
xor \U$5051 ( \5761 , \5760 , \5602 );
and \U$5052 ( \5762 , \5759 , \5761 );
and \U$5053 ( \5763 , \5665 , \5759 );
or \U$5054 ( \5764 , \5668 , \5762 , \5763 );
not \U$5055 ( \5765 , \5605 );
not \U$5056 ( \5766 , \5592 );
and \U$5057 ( \5767 , \5765 , \5766 );
and \U$5058 ( \5768 , \5605 , \5592 );
nor \U$5059 ( \5769 , \5767 , \5768 );
xor \U$5060 ( \5770 , \5764 , \5769 );
not \U$5061 ( \5771 , \5545 );
not \U$5062 ( \5772 , \5537 );
and \U$5063 ( \5773 , \5771 , \5772 );
and \U$5064 ( \5774 , \5545 , \5537 );
nor \U$5065 ( \5775 , \5773 , \5774 );
and \U$5066 ( \5776 , \5770 , \5775 );
and \U$5067 ( \5777 , \5764 , \5769 );
or \U$5068 ( \5778 , \5776 , \5777 );
and \U$5069 ( \5779 , \5630 , \5778 );
nor \U$5070 ( \5780 , \5629 , \5627 );
nor \U$5071 ( \5781 , \5779 , \5780 );
xor \U$5072 ( \5782 , \5626 , \5781 );
not \U$5073 ( \5783 , \5778 );
not \U$5074 ( \5784 , \5780 );
nand \U$5075 ( \5785 , \5784 , \5630 );
not \U$5076 ( \5786 , \5785 );
or \U$5077 ( \5787 , \5783 , \5786 );
or \U$5078 ( \5788 , \5785 , \5778 );
nand \U$5079 ( \5789 , \5787 , \5788 );
nand \U$5080 ( \5790 , \5119_nG10fb , \4857 );
or \U$5081 ( \5791 , \4771 , \5351_nGffe );
nand \U$5082 ( \5792 , \5791 , \4863 );
and \U$5083 ( \5793 , \5790 , \5792 );
and \U$5084 ( \5794 , \4859 , \5351_nGffe );
and \U$5085 ( \5795 , \5119_nG10fb , \4918 );
nor \U$5086 ( \5796 , \5793 , \5794 , \5795 );
and \U$5087 ( \5797 , \4960_nG12e2 , \5125 );
or \U$5088 ( \5798 , \4934 , \4960_nG12e2 );
nand \U$5089 ( \5799 , \5798 , \5128 );
nand \U$5090 ( \5800 , \5055_nG11dc , \4997 );
and \U$5091 ( \5801 , \5799 , \5800 );
and \U$5092 ( \5802 , \5055_nG11dc , \5000 );
nor \U$5093 ( \5803 , \5797 , \5801 , \5802 );
xor \U$5094 ( \5804 , \5796 , \5803 );
nand \U$5095 ( \5805 , \5526_nGe53 , \4698 );
or \U$5096 ( \5806 , \4659 , \5471_nGf21 );
nand \U$5097 ( \5807 , \5806 , \4725 );
and \U$5098 ( \5808 , \5805 , \5807 );
and \U$5099 ( \5809 , \4728 , \5471_nGf21 );
and \U$5100 ( \5810 , \5526_nGe53 , \4701 );
nor \U$5101 ( \5811 , \5808 , \5809 , \5810 );
and \U$5102 ( \5812 , \5804 , \5811 );
and \U$5103 ( \5813 , \5796 , \5803 );
or \U$5104 ( \5814 , \5812 , \5813 );
nand \U$5105 ( \5815 , \4757_nG15ca , \5392 );
or \U$5106 ( \5816 , \5288 , \4686_nG16f0 );
nand \U$5107 ( \5817 , \5816 , \5574 );
and \U$5108 ( \5818 , \5815 , \5817 );
and \U$5109 ( \5819 , \5577 , \4686_nG16f0 );
and \U$5110 ( \5820 , \4757_nG15ca , \5395 );
nor \U$5111 ( \5821 , \5818 , \5819 , \5820 );
not \U$5112 ( \5822 , \5707 );
and \U$5113 ( \5823 , \4634 , \5822 );
and \U$5114 ( \5824 , \5705 , \4594 );
and \U$5115 ( \5825 , \5282 , \5704 );
and \U$5116 ( \5826 , \4632_nG1905 , \5825 );
nor \U$5117 ( \5827 , \5823 , \5824 , \5826 );
xor \U$5118 ( \5828 , \5821 , \5827 );
nand \U$5119 ( \5829 , \4891_nG13e1 , \5200 );
or \U$5120 ( \5830 , \5149 , \4836_nG14e1 );
nand \U$5121 ( \5831 , \5830 , \5292 );
and \U$5122 ( \5832 , \5829 , \5831 );
and \U$5123 ( \5833 , \5295 , \4836_nG14e1 );
and \U$5124 ( \5834 , \4891_nG13e1 , \5203 );
nor \U$5125 ( \5835 , \5832 , \5833 , \5834 );
and \U$5126 ( \5836 , \5828 , \5835 );
and \U$5127 ( \5837 , \5821 , \5827 );
or \U$5128 ( \5838 , \5836 , \5837 );
nor \U$5129 ( \5839 , \5814 , \5838 );
xor \U$5130 ( \5840 , \5553 , \5560 );
xor \U$5131 ( \5841 , \5840 , \5568 );
not \U$5132 ( \5842 , \5841 );
and \U$5133 ( \5843 , \5839 , \5842 );
not \U$5134 ( \5844 , \5839 );
nand \U$5135 ( \5845 , \5844 , \5841 );
not \U$5136 ( \5846 , \5752 );
nor \U$5137 ( \5847 , \5725 , \5755 );
not \U$5138 ( \5848 , \5847 );
or \U$5139 ( \5849 , \5846 , \5848 );
or \U$5140 ( \5850 , \5847 , \5752 );
nand \U$5141 ( \5851 , \5849 , \5850 );
not \U$5142 ( \5852 , \5851 );
xor \U$5143 ( \5853 , \5675 , \5682 );
xor \U$5144 ( \5854 , \5853 , \5690 );
nor \U$5145 ( \5855 , \5852 , \5854 );
and \U$5146 ( \5856 , \5845 , \5855 );
nor \U$5147 ( \5857 , \5843 , \5856 );
not \U$5148 ( \5858 , \5665 );
xor \U$5149 ( \5859 , \5580 , \5283 );
xor \U$5150 ( \5860 , \5859 , \5588 );
xor \U$5151 ( \5861 , \5858 , \5860 );
xor \U$5152 ( \5862 , \5693 , \5709 );
xor \U$5153 ( \5863 , \5862 , \5756 );
and \U$5154 ( \5864 , \5861 , \5863 );
and \U$5155 ( \5865 , \5858 , \5860 );
or \U$5156 ( \5866 , \5864 , \5865 );
and \U$5157 ( \5867 , \5857 , \5866 );
xor \U$5158 ( \5868 , \5595 , \5600 );
xor \U$5159 ( \5869 , \5868 , \5602 );
xor \U$5160 ( \5870 , \5665 , \5759 );
xor \U$5161 ( \5871 , \5869 , \5870 );
not \U$5162 ( \5872 , \5871 );
or \U$5163 ( \5873 , \5664 , \5657 );
not \U$5164 ( \5874 , \5591 );
or \U$5165 ( \5875 , \5874 , \5571 );
not \U$5166 ( \5876 , \5571 );
or \U$5167 ( \5877 , \5591 , \5876 );
nand \U$5168 ( \5878 , \5873 , \5875 , \5877 );
nand \U$5169 ( \5879 , \5872 , \5878 );
xor \U$5170 ( \5880 , \5867 , \5879 );
xor \U$5171 ( \5881 , \5764 , \5769 );
xor \U$5172 ( \5882 , \5881 , \5775 );
and \U$5173 ( \5883 , \5880 , \5882 );
and \U$5174 ( \5884 , \5867 , \5879 );
or \U$5175 ( \5885 , \5883 , \5884 );
xor \U$5176 ( \5886 , \5789 , \5885 );
xor \U$5177 ( \5887 , \5857 , \5866 );
not \U$5178 ( \5888 , \5700 );
not \U$5179 ( \5889 , \5708 );
and \U$5180 ( \5890 , \5888 , \5889 );
and \U$5181 ( \5891 , \5700 , \5708 );
nor \U$5182 ( \5892 , \5890 , \5891 );
and \U$5183 ( \5893 , \5055_nG11dc , \5125 );
or \U$5184 ( \5894 , \4934 , \5055_nG11dc );
nand \U$5185 ( \5895 , \5894 , \5128 );
nand \U$5186 ( \5896 , \5119_nG10fb , \4997 );
and \U$5187 ( \5897 , \5895 , \5896 );
and \U$5188 ( \5898 , \5119_nG10fb , \5000 );
nor \U$5189 ( \5899 , \5893 , \5897 , \5898 );
nand \U$5190 ( \5900 , \4960_nG12e2 , \5200 );
or \U$5191 ( \5901 , \5149 , \4891_nG13e1 );
nand \U$5192 ( \5902 , \5901 , \5292 );
and \U$5193 ( \5903 , \5900 , \5902 );
and \U$5194 ( \5904 , \5295 , \4891_nG13e1 );
and \U$5195 ( \5905 , \4960_nG12e2 , \5203 );
nor \U$5196 ( \5906 , \5903 , \5904 , \5905 );
xor \U$5197 ( \5907 , \5899 , \5906 );
nand \U$5198 ( \5908 , \5351_nGffe , \4857 );
or \U$5199 ( \5909 , \4771 , \5471_nGf21 );
nand \U$5200 ( \5910 , \5909 , \4863 );
and \U$5201 ( \5911 , \5908 , \5910 );
and \U$5202 ( \5912 , \4859 , \5471_nGf21 );
and \U$5203 ( \5913 , \5351_nGffe , \4918 );
nor \U$5204 ( \5914 , \5911 , \5912 , \5913 );
and \U$5205 ( \5915 , \5907 , \5914 );
and \U$5206 ( \5916 , \5899 , \5906 );
or \U$5207 ( \5917 , \5915 , \5916 );
nand \U$5208 ( \5918 , \5656_nGaf0 , \4698 );
or \U$5209 ( \5919 , \4659 , \5526_nGe53 );
nand \U$5210 ( \5920 , \5919 , \4725 );
and \U$5211 ( \5921 , \5918 , \5920 );
and \U$5212 ( \5922 , \4728 , \5526_nGe53 );
and \U$5213 ( \5923 , \5656_nGaf0 , \4701 );
nor \U$5214 ( \5924 , \5921 , \5922 , \5923 );
and \U$5215 ( \5925 , \712 , RIaaa5f00_497);
and \U$5216 ( \5926 , \723 , RIaaa59d8_486);
and \U$5217 ( \5927 , RIaaa5a50_487, \728 );
nor \U$5218 ( \5928 , \5926 , \5927 );
and \U$5219 ( \5929 , \733 , RIaaa60e0_501);
and \U$5220 ( \5930 , RIaaa5bb8_490, \735 );
nor \U$5221 ( \5931 , \5929 , \5930 );
and \U$5222 ( \5932 , \738 , RIaaa5c30_491);
and \U$5223 ( \5933 , RIaaa5ff0_499, \696 );
nor \U$5224 ( \5934 , \5932 , \5933 );
and \U$5225 ( \5935 , \721 , RIaaa6068_500);
and \U$5226 ( \5936 , RIaaa6158_502, \682 );
nor \U$5227 ( \5937 , \5935 , \5936 );
nand \U$5228 ( \5938 , \5928 , \5931 , \5934 , \5937 );
nor \U$5229 ( \5939 , \5925 , \5938 );
and \U$5230 ( \5940 , \686 , RIaaa5f78_498);
and \U$5231 ( \5941 , RIaaa5d20_493, \690 );
nor \U$5232 ( \5942 , \5940 , \5941 );
and \U$5233 ( \5943 , \702 , RIaaa5ca8_492);
and \U$5234 ( \5944 , RIaaa5b40_489, \730 );
nor \U$5235 ( \5945 , \5943 , \5944 );
and \U$5236 ( \5946 , \4572 , RIaaa5e88_496);
and \U$5237 ( \5947 , RIaaa5ac8_488, \699 );
nor \U$5238 ( \5948 , \5946 , \5947 );
nand \U$5239 ( \5949 , \5939 , \5942 , \5945 , \5948 );
_DC ga4b ( \5950_nGa4b , \5949 , \4592 );
nand \U$5240 ( \5951 , \5950_nGa4b , \4565 );
xor \U$5241 ( \5952 , \5924 , \5951 );
and \U$5242 ( \5953 , \5751_nGabb , \4645 );
and \U$5243 ( \5954 , RIaaa5168_468, \682 );
and \U$5244 ( \5955 , RIaaa5078_466, \738 );
and \U$5245 ( \5956 , \686 , RIaaa4cb8_458);
and \U$5246 ( \5957 , RIaaa4a60_453, \690 );
nor \U$5247 ( \5958 , \5956 , \5957 );
and \U$5248 ( \5959 , RIaaa4bc8_456, \4572 );
and \U$5249 ( \5960 , \735 , RIaaa5000_465);
and \U$5250 ( \5961 , RIaaa4d30_459, \696 );
nor \U$5251 ( \5962 , \5959 , \5960 , \5961 );
and \U$5252 ( \5963 , \699 , RIaaa4f10_463);
and \U$5253 ( \5964 , RIaaa4c40_457, \712 );
nor \U$5254 ( \5965 , \5963 , \5964 );
nand \U$5255 ( \5966 , \5958 , \5962 , \5965 );
nor \U$5256 ( \5967 , \5954 , \5955 , \5966 );
and \U$5257 ( \5968 , \702 , RIaaa49e8_452);
and \U$5258 ( \5969 , RIaaa4e20_461, \728 );
nor \U$5259 ( \5970 , \5968 , \5969 );
and \U$5260 ( \5971 , \733 , RIaaa50f0_467);
and \U$5261 ( \5972 , RIaaa4f88_464, \730 );
nor \U$5262 ( \5973 , \5971 , \5972 );
and \U$5263 ( \5974 , \721 , RIaaa4da8_460);
and \U$5264 ( \5975 , RIaaa4e98_462, \723 );
nor \U$5265 ( \5976 , \5974 , \5975 );
nand \U$5266 ( \5977 , \5967 , \5970 , \5973 , \5976 );
_DC ga7f ( \5978_nGa7f , \5977 , \4592 );
or \U$5267 ( \5979 , \4606 , \5978_nGa7f );
nand \U$5268 ( \5980 , \5979 , \4642 );
nand \U$5269 ( \5981 , \5751_nGabb , \4638 );
and \U$5270 ( \5982 , \5980 , \5981 );
and \U$5271 ( \5983 , \5978_nGa7f , \4762 );
nor \U$5272 ( \5984 , \5953 , \5982 , \5983 );
and \U$5273 ( \5985 , \5952 , \5984 );
and \U$5274 ( \5986 , \5924 , \5951 );
or \U$5275 ( \5987 , \5985 , \5986 );
nand \U$5276 ( \5988 , \5917 , \5987 );
not \U$5277 ( \5989 , \5825 );
or \U$5278 ( \5990 , \5989 , \4594 );
or \U$5279 ( \5991 , \4593_nG17f6 , \5707 );
or \U$5280 ( \5992 , \4686_nG16f0 , \5706 );
nand \U$5281 ( \5993 , \5990 , \5991 , \5992 );
not \U$5282 ( \5994 , \5993 );
nand \U$5283 ( \5995 , \4836_nG14e1 , \5392 );
or \U$5284 ( \5996 , \5288 , \4757_nG15ca );
nand \U$5285 ( \5997 , \5996 , \5574 );
and \U$5286 ( \5998 , \5995 , \5997 );
and \U$5287 ( \5999 , \5577 , \4757_nG15ca );
and \U$5288 ( \6000 , \4836_nG14e1 , \5395 );
nor \U$5289 ( \6001 , \5998 , \5999 , \6000 );
nor \U$5290 ( \6002 , \5994 , \6001 );
and \U$5291 ( \6003 , \5988 , \6002 );
nor \U$5292 ( \6004 , \5987 , \5917 );
nor \U$5293 ( \6005 , \6003 , \6004 );
nand \U$5294 ( \6006 , \5892 , \6005 );
nand \U$5295 ( \6007 , \5978_nGa7f , \4565 );
and \U$5296 ( \6008 , \5656_nGaf0 , \4645 );
or \U$5297 ( \6009 , \4606 , \5751_nGabb );
nand \U$5298 ( \6010 , \6009 , \4642 );
nand \U$5299 ( \6011 , \5656_nGaf0 , \4638 );
and \U$5300 ( \6012 , \6010 , \6011 );
and \U$5301 ( \6013 , \5751_nGabb , \4762 );
nor \U$5302 ( \6014 , \6008 , \6012 , \6013 );
xor \U$5303 ( \6015 , \6007 , \6014 );
not \U$5304 ( \6016 , \6015 );
xor \U$5305 ( \6017 , \5796 , \5803 );
xor \U$5306 ( \6018 , \6017 , \5811 );
nor \U$5307 ( \6019 , \6016 , \6018 );
and \U$5308 ( \6020 , \6006 , \6019 );
nor \U$5309 ( \6021 , \6005 , \5892 );
nor \U$5310 ( \6022 , \6020 , \6021 );
not \U$5311 ( \6023 , \5851 );
not \U$5312 ( \6024 , \5854 );
and \U$5313 ( \6025 , \6023 , \6024 );
and \U$5314 ( \6026 , \5851 , \5854 );
nor \U$5315 ( \6027 , \6025 , \6026 );
not \U$5316 ( \6028 , \6027 );
or \U$5317 ( \6029 , \6014 , \6007 );
not \U$5318 ( \6030 , \5838 );
or \U$5319 ( \6031 , \6030 , \5814 );
not \U$5320 ( \6032 , \5814 );
or \U$5321 ( \6033 , \5838 , \6032 );
nand \U$5322 ( \6034 , \6029 , \6031 , \6033 );
nand \U$5323 ( \6035 , \6028 , \6034 );
xor \U$5324 ( \6036 , \6022 , \6035 );
xor \U$5325 ( \6037 , \5858 , \5860 );
xor \U$5326 ( \6038 , \6037 , \5863 );
and \U$5327 ( \6039 , \6036 , \6038 );
and \U$5328 ( \6040 , \6022 , \6035 );
or \U$5329 ( \6041 , \6039 , \6040 );
nand \U$5330 ( \6042 , \5887 , \6041 );
not \U$5331 ( \6043 , \6042 );
nor \U$5332 ( \6044 , \6041 , \5887 );
nor \U$5333 ( \6045 , \6043 , \6044 );
not \U$5334 ( \6046 , \6045 );
not \U$5335 ( \6047 , \5878 );
not \U$5336 ( \6048 , \5871 );
or \U$5337 ( \6049 , \6047 , \6048 );
or \U$5338 ( \6050 , \5871 , \5878 );
nand \U$5339 ( \6051 , \6049 , \6050 );
not \U$5340 ( \6052 , \6051 );
and \U$5341 ( \6053 , \6046 , \6052 );
and \U$5342 ( \6054 , \6045 , \6051 );
nor \U$5343 ( \6055 , \6053 , \6054 );
xor \U$5344 ( \6056 , \6022 , \6035 );
xor \U$5345 ( \6057 , \6056 , \6038 );
not \U$5346 ( \6058 , \5841 );
xor \U$5347 ( \6059 , \5839 , \5855 );
not \U$5348 ( \6060 , \6059 );
or \U$5349 ( \6061 , \6058 , \6060 );
or \U$5350 ( \6062 , \6059 , \5841 );
nand \U$5351 ( \6063 , \6061 , \6062 );
not \U$5352 ( \6064 , \6034 );
not \U$5353 ( \6065 , \6027 );
or \U$5354 ( \6066 , \6064 , \6065 );
or \U$5355 ( \6067 , \6027 , \6034 );
nand \U$5356 ( \6068 , \6066 , \6067 );
not \U$5357 ( \6069 , \6068 );
xor \U$5358 ( \6070 , \5821 , \5827 );
xor \U$5359 ( \6071 , \6070 , \5835 );
not \U$5360 ( \6072 , \6071 );
nand \U$5361 ( \6073 , \5471_nGf21 , \4857 );
or \U$5362 ( \6074 , \4771 , \5526_nGe53 );
nand \U$5363 ( \6075 , \6074 , \4863 );
and \U$5364 ( \6076 , \6073 , \6075 );
and \U$5365 ( \6077 , \4859 , \5526_nGe53 );
and \U$5366 ( \6078 , \5471_nGf21 , \4918 );
nor \U$5367 ( \6079 , \6076 , \6077 , \6078 );
and \U$5368 ( \6080 , \5119_nG10fb , \5125 );
or \U$5369 ( \6081 , \4934 , \5119_nG10fb );
nand \U$5370 ( \6082 , \6081 , \5128 );
nand \U$5371 ( \6083 , \5351_nGffe , \4997 );
and \U$5372 ( \6084 , \6082 , \6083 );
and \U$5373 ( \6085 , \5351_nGffe , \5000 );
nor \U$5374 ( \6086 , \6080 , \6084 , \6085 );
xor \U$5375 ( \6087 , \6079 , \6086 );
nand \U$5376 ( \6088 , \5751_nGabb , \4698 );
or \U$5377 ( \6089 , \4659 , \5656_nGaf0 );
nand \U$5378 ( \6090 , \6089 , \4725 );
and \U$5379 ( \6091 , \6088 , \6090 );
and \U$5380 ( \6092 , \4728 , \5656_nGaf0 );
and \U$5381 ( \6093 , \5751_nGabb , \4701 );
nor \U$5382 ( \6094 , \6091 , \6092 , \6093 );
and \U$5383 ( \6095 , \6087 , \6094 );
and \U$5384 ( \6096 , \6079 , \6086 );
or \U$5385 ( \6097 , \6095 , \6096 );
nand \U$5386 ( \6098 , \4891_nG13e1 , \5392 );
or \U$5387 ( \6099 , \5288 , \4836_nG14e1 );
nand \U$5388 ( \6100 , \6099 , \5574 );
and \U$5389 ( \6101 , \6098 , \6100 );
and \U$5390 ( \6102 , \5577 , \4836_nG14e1 );
and \U$5391 ( \6103 , \4891_nG13e1 , \5395 );
nor \U$5392 ( \6104 , \6101 , \6102 , \6103 );
and \U$5393 ( \6105 , \4687 , \5822 );
not \U$5394 ( \6106 , \4757_nG15ca );
and \U$5395 ( \6107 , \5705 , \6106 );
and \U$5396 ( \6108 , \4686_nG16f0 , \5825 );
nor \U$5397 ( \6109 , \6105 , \6107 , \6108 );
xor \U$5398 ( \6110 , \6104 , \6109 );
nand \U$5399 ( \6111 , \5055_nG11dc , \5200 );
or \U$5400 ( \6112 , \5149 , \4960_nG12e2 );
nand \U$5401 ( \6113 , \6112 , \5292 );
and \U$5402 ( \6114 , \6111 , \6113 );
and \U$5403 ( \6115 , \5295 , \4960_nG12e2 );
and \U$5404 ( \6116 , \5055_nG11dc , \5203 );
nor \U$5405 ( \6117 , \6114 , \6115 , \6116 );
and \U$5406 ( \6118 , \6110 , \6117 );
and \U$5407 ( \6119 , \6104 , \6109 );
or \U$5408 ( \6120 , \6118 , \6119 );
nor \U$5409 ( \6121 , \6097 , \6120 );
nand \U$5410 ( \6122 , \6072 , \6121 );
or \U$5411 ( \6123 , \6069 , \6122 );
not \U$5412 ( \6124 , \6122 );
not \U$5413 ( \6125 , \6069 );
or \U$5414 ( \6126 , \6124 , \6125 );
not \U$5415 ( \6127 , \6019 );
not \U$5416 ( \6128 , \6021 );
nand \U$5417 ( \6129 , \6128 , \6006 );
not \U$5418 ( \6130 , \6129 );
or \U$5419 ( \6131 , \6127 , \6130 );
or \U$5420 ( \6132 , \6129 , \6019 );
nand \U$5421 ( \6133 , \6131 , \6132 );
nand \U$5422 ( \6134 , \6126 , \6133 );
nand \U$5423 ( \6135 , \6123 , \6134 );
nand \U$5424 ( \6136 , \6063 , \6135 );
and \U$5425 ( \6137 , \6057 , \6136 );
nor \U$5426 ( \6138 , \6135 , \6063 );
nor \U$5427 ( \6139 , \6137 , \6138 );
xor \U$5428 ( \6140 , \6055 , \6139 );
not \U$5429 ( \6141 , \6138 );
nand \U$5430 ( \6142 , \6141 , \6136 );
not \U$5431 ( \6143 , \6142 );
not \U$5432 ( \6144 , \6057 );
or \U$5433 ( \6145 , \6143 , \6144 );
or \U$5434 ( \6146 , \6142 , \6057 );
nand \U$5435 ( \6147 , \6145 , \6146 );
not \U$5436 ( \6148 , \6097 );
and \U$5437 ( \6149 , \6148 , \6120 );
and \U$5438 ( \6150 , \5978_nGa7f , \4645 );
or \U$5439 ( \6151 , \4606 , \5950_nGa4b );
nand \U$5440 ( \6152 , \6151 , \4642 );
nand \U$5441 ( \6153 , \5978_nGa7f , \4638 );
and \U$5442 ( \6154 , \6152 , \6153 );
and \U$5443 ( \6155 , \5950_nGa4b , \4762 );
nor \U$5444 ( \6156 , \6150 , \6154 , \6155 );
and \U$5445 ( \6157 , RIaaa6e00_529, \682 );
and \U$5446 ( \6158 , RIaaa6ba8_524, \738 );
and \U$5447 ( \6159 , \686 , RIaaa6d10_527);
and \U$5448 ( \6160 , RIaaa6f68_532, \690 );
nor \U$5449 ( \6161 , \6159 , \6160 );
and \U$5450 ( \6162 , RIaaa7058_534, \4572 );
and \U$5451 ( \6163 , \735 , RIaaa6c20_525);
and \U$5452 ( \6164 , RIaaa6c98_526, \696 );
nor \U$5453 ( \6165 , \6162 , \6163 , \6164 );
and \U$5454 ( \6166 , \699 , RIaaa6a40_521);
and \U$5455 ( \6167 , RIaaa70d0_535, \712 );
nor \U$5456 ( \6168 , \6166 , \6167 );
nand \U$5457 ( \6169 , \6161 , \6165 , \6168 );
nor \U$5458 ( \6170 , \6157 , \6158 , \6169 );
and \U$5459 ( \6171 , \721 , RIaaa6e78_530);
and \U$5460 ( \6172 , RIaaa6d88_528, \733 );
nor \U$5461 ( \6173 , \6171 , \6172 );
and \U$5462 ( \6174 , \702 , RIaaa6ef0_531);
and \U$5463 ( \6175 , RIaaa69c8_520, \730 );
nor \U$5464 ( \6176 , \6174 , \6175 );
and \U$5465 ( \6177 , \723 , RIaaa6b30_523);
and \U$5466 ( \6178 , RIaaa6ab8_522, \728 );
nor \U$5467 ( \6179 , \6177 , \6178 );
nand \U$5468 ( \6180 , \6170 , \6173 , \6176 , \6179 );
_DC ga0e ( \6181_nGa0e , \6180 , \4592 );
nand \U$5469 ( \6182 , \6181_nGa0e , \4565 );
or \U$5470 ( \6183 , \6156 , \6182 );
or \U$5471 ( \6184 , \6120 , \6148 );
nand \U$5472 ( \6185 , \6183 , \6184 );
nor \U$5473 ( \6186 , \6149 , \6185 );
not \U$5474 ( \6187 , \6001 );
not \U$5475 ( \6188 , \5993 );
and \U$5476 ( \6189 , \6187 , \6188 );
and \U$5477 ( \6190 , \6001 , \5993 );
nor \U$5478 ( \6191 , \6189 , \6190 );
xor \U$5479 ( \6192 , \6186 , \6191 );
xor \U$5480 ( \6193 , \5924 , \5951 );
xor \U$5481 ( \6194 , \6193 , \5984 );
and \U$5482 ( \6195 , \6192 , \6194 );
and \U$5483 ( \6196 , \6186 , \6191 );
or \U$5484 ( \6197 , \6195 , \6196 );
not \U$5485 ( \6198 , \6015 );
not \U$5486 ( \6199 , \6018 );
and \U$5487 ( \6200 , \6198 , \6199 );
and \U$5488 ( \6201 , \6015 , \6018 );
nor \U$5489 ( \6202 , \6200 , \6201 );
xor \U$5490 ( \6203 , \6197 , \6202 );
xor \U$5491 ( \6204 , \6079 , \6086 );
xor \U$5492 ( \6205 , \6204 , \6094 );
xor \U$5493 ( \6206 , \6104 , \6109 );
xor \U$5494 ( \6207 , \6206 , \6117 );
xor \U$5495 ( \6208 , \6205 , \6207 );
xnor \U$5496 ( \6209 , \6182 , \6156 );
and \U$5497 ( \6210 , \6208 , \6209 );
and \U$5498 ( \6211 , \6205 , \6207 );
or \U$5499 ( \6212 , \6210 , \6211 );
xor \U$5500 ( \6213 , \5899 , \5906 );
xor \U$5501 ( \6214 , \6213 , \5914 );
xor \U$5502 ( \6215 , \6212 , \6214 );
and \U$5503 ( \6216 , \5351_nGffe , \5125 );
or \U$5504 ( \6217 , \4934 , \5351_nGffe );
nand \U$5505 ( \6218 , \6217 , \5128 );
nand \U$5506 ( \6219 , \5471_nGf21 , \4997 );
and \U$5507 ( \6220 , \6218 , \6219 );
and \U$5508 ( \6221 , \5471_nGf21 , \5000 );
nor \U$5509 ( \6222 , \6216 , \6220 , \6221 );
nand \U$5510 ( \6223 , \5119_nG10fb , \5200 );
or \U$5511 ( \6224 , \5149 , \5055_nG11dc );
nand \U$5512 ( \6225 , \6224 , \5292 );
and \U$5513 ( \6226 , \6223 , \6225 );
and \U$5514 ( \6227 , \5295 , \5055_nG11dc );
and \U$5515 ( \6228 , \5119_nG10fb , \5203 );
nor \U$5516 ( \6229 , \6226 , \6227 , \6228 );
xor \U$5517 ( \6230 , \6222 , \6229 );
nand \U$5518 ( \6231 , \5526_nGe53 , \4857 );
or \U$5519 ( \6232 , \4771 , \5656_nGaf0 );
nand \U$5520 ( \6233 , \6232 , \4863 );
and \U$5521 ( \6234 , \6231 , \6233 );
and \U$5522 ( \6235 , \4859 , \5656_nGaf0 );
and \U$5523 ( \6236 , \5526_nGe53 , \4918 );
nor \U$5524 ( \6237 , \6234 , \6235 , \6236 );
and \U$5525 ( \6238 , \6230 , \6237 );
and \U$5526 ( \6239 , \6222 , \6229 );
or \U$5527 ( \6240 , \6238 , \6239 );
nand \U$5528 ( \6241 , \4960_nG12e2 , \5392 );
or \U$5529 ( \6242 , \5288 , \4891_nG13e1 );
nand \U$5530 ( \6243 , \6242 , \5574 );
and \U$5531 ( \6244 , \6241 , \6243 );
and \U$5532 ( \6245 , \5577 , \4891_nG13e1 );
and \U$5533 ( \6246 , \4960_nG12e2 , \5395 );
nor \U$5534 ( \6247 , \6244 , \6245 , \6246 );
not \U$5535 ( \6248 , \6247 );
or \U$5536 ( \6249 , \5989 , \6106 );
or \U$5537 ( \6250 , \4757_nG15ca , \5707 );
or \U$5538 ( \6251 , \4836_nG14e1 , \5706 );
nand \U$5539 ( \6252 , \6249 , \6250 , \6251 );
nand \U$5540 ( \6253 , \6248 , \6252 );
xor \U$5541 ( \6254 , \6240 , \6253 );
and \U$5542 ( \6255 , \5950_nGa4b , \4645 );
or \U$5543 ( \6256 , \4606 , \6181_nGa0e );
nand \U$5544 ( \6257 , \6256 , \4642 );
nand \U$5545 ( \6258 , \5950_nGa4b , \4638 );
and \U$5546 ( \6259 , \6257 , \6258 );
and \U$5547 ( \6260 , \6181_nGa0e , \4762 );
nor \U$5548 ( \6261 , \6255 , \6259 , \6260 );
nand \U$5549 ( \6262 , \5978_nGa7f , \4698 );
or \U$5550 ( \6263 , \4659 , \5751_nGabb );
nand \U$5551 ( \6264 , \6263 , \4725 );
and \U$5552 ( \6265 , \6262 , \6264 );
and \U$5553 ( \6266 , \4728 , \5751_nGabb );
and \U$5554 ( \6267 , \5978_nGa7f , \4701 );
nor \U$5555 ( \6268 , \6265 , \6266 , \6267 );
and \U$5556 ( \6269 , \6261 , \6268 );
not \U$5557 ( \6270 , \6269 );
and \U$5558 ( \6271 , RIaaa77d8_550, \733 );
and \U$5559 ( \6272 , RIaaa7490_543, \730 );
and \U$5560 ( \6273 , \686 , RIaaa7760_549);
and \U$5561 ( \6274 , RIaaa7940_553, \690 );
nor \U$5562 ( \6275 , \6273 , \6274 );
and \U$5563 ( \6276 , RIaaa72b0_539, \4572 );
and \U$5564 ( \6277 , \735 , RIaaa73a0_541);
and \U$5565 ( \6278 , RIaaa76e8_548, \696 );
nor \U$5566 ( \6279 , \6276 , \6277 , \6278 );
and \U$5567 ( \6280 , \699 , RIaaa7580_545);
and \U$5568 ( \6281 , RIaaa7328_540, \712 );
nor \U$5569 ( \6282 , \6280 , \6281 );
nand \U$5570 ( \6283 , \6275 , \6279 , \6282 );
nor \U$5571 ( \6284 , \6271 , \6272 , \6283 );
and \U$5572 ( \6285 , \738 , RIaaa7418_542);
and \U$5573 ( \6286 , RIaaa7850_551, \682 );
nor \U$5574 ( \6287 , \6285 , \6286 );
and \U$5575 ( \6288 , \702 , RIaaa78c8_552);
and \U$5576 ( \6289 , RIaaa7508_544, \721 );
nor \U$5577 ( \6290 , \6288 , \6289 );
and \U$5578 ( \6291 , \723 , RIaaa75f8_546);
and \U$5579 ( \6292 , RIaaa7670_547, \728 );
nor \U$5580 ( \6293 , \6291 , \6292 );
nand \U$5581 ( \6294 , \6284 , \6287 , \6290 , \6293 );
_DC g9d6 ( \6295_nG9d6 , \6294 , \4592 );
nand \U$5582 ( \6296 , \6295_nG9d6 , \4565 );
not \U$5583 ( \6297 , \6296 );
and \U$5584 ( \6298 , \6270 , \6297 );
nor \U$5585 ( \6299 , \6261 , \6268 );
nor \U$5586 ( \6300 , \6298 , \6299 );
and \U$5587 ( \6301 , \6254 , \6300 );
and \U$5588 ( \6302 , \6240 , \6253 );
or \U$5589 ( \6303 , \6301 , \6302 );
and \U$5590 ( \6304 , \6215 , \6303 );
and \U$5591 ( \6305 , \6212 , \6214 );
or \U$5592 ( \6306 , \6304 , \6305 );
and \U$5593 ( \6307 , \6203 , \6306 );
and \U$5594 ( \6308 , \6197 , \6202 );
or \U$5595 ( \6309 , \6307 , \6308 );
not \U$5596 ( \6310 , \6121 );
not \U$5597 ( \6311 , \6071 );
and \U$5598 ( \6312 , \6310 , \6311 );
and \U$5599 ( \6313 , \6121 , \6071 );
nor \U$5600 ( \6314 , \6312 , \6313 );
not \U$5601 ( \6315 , \6314 );
not \U$5602 ( \6316 , \6002 );
not \U$5603 ( \6317 , \6004 );
nand \U$5604 ( \6318 , \6317 , \5988 );
not \U$5605 ( \6319 , \6318 );
or \U$5606 ( \6320 , \6316 , \6319 );
or \U$5607 ( \6321 , \6318 , \6002 );
nand \U$5608 ( \6322 , \6320 , \6321 );
nand \U$5609 ( \6323 , \6315 , \6322 );
xor \U$5610 ( \6324 , \6309 , \6323 );
not \U$5611 ( \6325 , \6133 );
not \U$5612 ( \6326 , \6122 );
and \U$5613 ( \6327 , \6325 , \6326 );
and \U$5614 ( \6328 , \6133 , \6122 );
nor \U$5615 ( \6329 , \6327 , \6328 );
not \U$5616 ( \6330 , \6329 );
not \U$5617 ( \6331 , \6068 );
and \U$5618 ( \6332 , \6330 , \6331 );
and \U$5619 ( \6333 , \6329 , \6068 );
nor \U$5620 ( \6334 , \6332 , \6333 );
and \U$5621 ( \6335 , \6324 , \6334 );
and \U$5622 ( \6336 , \6309 , \6323 );
or \U$5623 ( \6337 , \6335 , \6336 );
xor \U$5624 ( \6338 , \6147 , \6337 );
xor \U$5625 ( \6339 , \6186 , \6191 );
xor \U$5626 ( \6340 , \6339 , \6194 );
xor \U$5627 ( \6341 , \6212 , \6214 );
xor \U$5628 ( \6342 , \6341 , \6303 );
and \U$5629 ( \6343 , \6340 , \6342 );
xor \U$5630 ( \6344 , \6222 , \6229 );
xor \U$5631 ( \6345 , \6344 , \6237 );
not \U$5632 ( \6346 , \6345 );
not \U$5633 ( \6347 , \6296 );
nor \U$5634 ( \6348 , \6269 , \6299 );
not \U$5635 ( \6349 , \6348 );
or \U$5636 ( \6350 , \6347 , \6349 );
or \U$5637 ( \6351 , \6348 , \6296 );
nand \U$5638 ( \6352 , \6350 , \6351 );
nand \U$5639 ( \6353 , \6346 , \6352 );
nand \U$5640 ( \6354 , \5055_nG11dc , \5392 );
or \U$5641 ( \6355 , \5288 , \4960_nG12e2 );
nand \U$5642 ( \6356 , \6355 , \5574 );
and \U$5643 ( \6357 , \6354 , \6356 );
and \U$5644 ( \6358 , \5577 , \4960_nG12e2 );
and \U$5645 ( \6359 , \5055_nG11dc , \5395 );
nor \U$5646 ( \6360 , \6357 , \6358 , \6359 );
and \U$5647 ( \6361 , \4837 , \5822 );
and \U$5648 ( \6362 , \5705 , \4964 );
and \U$5649 ( \6363 , \4836_nG14e1 , \5825 );
nor \U$5650 ( \6364 , \6361 , \6362 , \6363 );
xor \U$5651 ( \6365 , \6360 , \6364 );
nand \U$5652 ( \6366 , \5351_nGffe , \5200 );
or \U$5653 ( \6367 , \5149 , \5119_nG10fb );
nand \U$5654 ( \6368 , \6367 , \5292 );
and \U$5655 ( \6369 , \6366 , \6368 );
and \U$5656 ( \6370 , \5295 , \5119_nG10fb );
and \U$5657 ( \6371 , \5351_nGffe , \5203 );
nor \U$5658 ( \6372 , \6369 , \6370 , \6371 );
and \U$5659 ( \6373 , \6365 , \6372 );
and \U$5660 ( \6374 , \6360 , \6364 );
or \U$5661 ( \6375 , \6373 , \6374 );
not \U$5662 ( \6376 , \6375 );
nand \U$5663 ( \6377 , \5656_nGaf0 , \4857 );
or \U$5664 ( \6378 , \4771 , \5751_nGabb );
nand \U$5665 ( \6379 , \6378 , \4863 );
and \U$5666 ( \6380 , \6377 , \6379 );
and \U$5667 ( \6381 , \4859 , \5751_nGabb );
and \U$5668 ( \6382 , \5656_nGaf0 , \4918 );
nor \U$5669 ( \6383 , \6380 , \6381 , \6382 );
and \U$5670 ( \6384 , \5471_nGf21 , \5125 );
or \U$5671 ( \6385 , \4934 , \5471_nGf21 );
nand \U$5672 ( \6386 , \6385 , \5128 );
nand \U$5673 ( \6387 , \5526_nGe53 , \4997 );
and \U$5674 ( \6388 , \6386 , \6387 );
and \U$5675 ( \6389 , \5526_nGe53 , \5000 );
nor \U$5676 ( \6390 , \6384 , \6388 , \6389 );
xor \U$5677 ( \6391 , \6383 , \6390 );
nand \U$5678 ( \6392 , \5950_nGa4b , \4698 );
or \U$5679 ( \6393 , \4659 , \5978_nGa7f );
nand \U$5680 ( \6394 , \6393 , \4725 );
and \U$5681 ( \6395 , \6392 , \6394 );
and \U$5682 ( \6396 , \4728 , \5978_nGa7f );
and \U$5683 ( \6397 , \5950_nGa4b , \4701 );
nor \U$5684 ( \6398 , \6395 , \6396 , \6397 );
and \U$5685 ( \6399 , \6391 , \6398 );
and \U$5686 ( \6400 , \6383 , \6390 );
or \U$5687 ( \6401 , \6399 , \6400 );
not \U$5688 ( \6402 , \6401 );
nand \U$5689 ( \6403 , \6376 , \6402 );
xor \U$5690 ( \6404 , \6353 , \6403 );
xor \U$5691 ( \6405 , \6205 , \6207 );
xor \U$5692 ( \6406 , \6405 , \6209 );
and \U$5693 ( \6407 , \6404 , \6406 );
and \U$5694 ( \6408 , \6353 , \6403 );
or \U$5695 ( \6409 , \6407 , \6408 );
xor \U$5696 ( \6410 , \6212 , \6214 );
xor \U$5697 ( \6411 , \6410 , \6303 );
and \U$5698 ( \6412 , \6409 , \6411 );
and \U$5699 ( \6413 , \6340 , \6409 );
or \U$5700 ( \6414 , \6343 , \6412 , \6413 );
not \U$5701 ( \6415 , \6322 );
not \U$5702 ( \6416 , \6314 );
and \U$5703 ( \6417 , \6415 , \6416 );
and \U$5704 ( \6418 , \6322 , \6314 );
nor \U$5705 ( \6419 , \6417 , \6418 );
xor \U$5706 ( \6420 , \6414 , \6419 );
xor \U$5707 ( \6421 , \6197 , \6202 );
xor \U$5708 ( \6422 , \6421 , \6306 );
xor \U$5709 ( \6423 , \6420 , \6422 );
not \U$5710 ( \6424 , \6423 );
xor \U$5711 ( \6425 , \6212 , \6214 );
xor \U$5712 ( \6426 , \6425 , \6303 );
xor \U$5713 ( \6427 , \6340 , \6409 );
xor \U$5714 ( \6428 , \6426 , \6427 );
not \U$5715 ( \6429 , \6352 );
not \U$5716 ( \6430 , \6345 );
and \U$5717 ( \6431 , \6429 , \6430 );
and \U$5718 ( \6432 , \6352 , \6345 );
nor \U$5719 ( \6433 , \6431 , \6432 );
not \U$5720 ( \6434 , \6433 );
and \U$5721 ( \6435 , \6181_nGa0e , \4645 );
or \U$5722 ( \6436 , \4606 , \6295_nG9d6 );
nand \U$5723 ( \6437 , \6436 , \4642 );
nand \U$5724 ( \6438 , \6181_nGa0e , \4638 );
and \U$5725 ( \6439 , \6437 , \6438 );
and \U$5726 ( \6440 , \6295_nG9d6 , \4762 );
nor \U$5727 ( \6441 , \6435 , \6439 , \6440 );
and \U$5728 ( \6442 , \712 , RIaaa8318_574);
and \U$5729 ( \6443 , \682 , RIaaa8840_585);
and \U$5730 ( \6444 , RIaaa8660_581, \728 );
nor \U$5731 ( \6445 , \6443 , \6444 );
and \U$5732 ( \6446 , \702 , RIaaa88b8_586);
and \U$5733 ( \6447 , RIaaa84f8_578, \721 );
nor \U$5734 ( \6448 , \6446 , \6447 );
and \U$5735 ( \6449 , \738 , RIaaa8480_577);
and \U$5736 ( \6450 , RIaaa87c8_584, \733 );
nor \U$5737 ( \6451 , \6449 , \6450 );
and \U$5738 ( \6452 , \723 , RIaaa85e8_580);
and \U$5739 ( \6453 , RIaaa8408_576, \730 );
nor \U$5740 ( \6454 , \6452 , \6453 );
nand \U$5741 ( \6455 , \6445 , \6448 , \6451 , \6454 );
nor \U$5742 ( \6456 , \6442 , \6455 );
and \U$5743 ( \6457 , \686 , RIaaa8750_583);
and \U$5744 ( \6458 , RIaaa8930_587, \690 );
nor \U$5745 ( \6459 , \6457 , \6458 );
and \U$5746 ( \6460 , \699 , RIaaa8570_579);
and \U$5747 ( \6461 , RIaaa8390_575, \735 );
nor \U$5748 ( \6462 , \6460 , \6461 );
and \U$5749 ( \6463 , \4572 , RIaaa82a0_573);
and \U$5750 ( \6464 , RIaaa86d8_582, \696 );
nor \U$5751 ( \6465 , \6463 , \6464 );
nand \U$5752 ( \6466 , \6456 , \6459 , \6462 , \6465 );
_DC g99e ( \6467_nG99e , \6466 , \4592 );
nand \U$5753 ( \6468 , \6467_nG99e , \4565 );
or \U$5754 ( \6469 , \6441 , \6468 );
or \U$5755 ( \6470 , \6376 , \6401 );
or \U$5756 ( \6471 , \6375 , \6402 );
nand \U$5757 ( \6472 , \6469 , \6470 , \6471 );
nand \U$5758 ( \6473 , \6434 , \6472 );
xor \U$5759 ( \6474 , \6240 , \6253 );
xor \U$5760 ( \6475 , \6474 , \6300 );
xor \U$5761 ( \6476 , \6473 , \6475 );
xor \U$5762 ( \6477 , \6383 , \6390 );
xor \U$5763 ( \6478 , \6477 , \6398 );
xor \U$5764 ( \6479 , \6360 , \6364 );
xor \U$5765 ( \6480 , \6479 , \6372 );
xor \U$5766 ( \6481 , \6478 , \6480 );
xnor \U$5767 ( \6482 , \6468 , \6441 );
and \U$5768 ( \6483 , \6481 , \6482 );
and \U$5769 ( \6484 , \6478 , \6480 );
or \U$5770 ( \6485 , \6483 , \6484 );
not \U$5771 ( \6486 , \6247 );
not \U$5772 ( \6487 , \6252 );
and \U$5773 ( \6488 , \6486 , \6487 );
and \U$5774 ( \6489 , \6247 , \6252 );
nor \U$5775 ( \6490 , \6488 , \6489 );
xor \U$5776 ( \6491 , \6485 , \6490 );
and \U$5777 ( \6492 , \5526_nGe53 , \5125 );
or \U$5778 ( \6493 , \4934 , \5526_nGe53 );
nand \U$5779 ( \6494 , \6493 , \5128 );
nand \U$5780 ( \6495 , \5656_nGaf0 , \4997 );
and \U$5781 ( \6496 , \6494 , \6495 );
and \U$5782 ( \6497 , \5656_nGaf0 , \5000 );
nor \U$5783 ( \6498 , \6492 , \6496 , \6497 );
nand \U$5784 ( \6499 , \5471_nGf21 , \5200 );
or \U$5785 ( \6500 , \5149 , \5351_nGffe );
nand \U$5786 ( \6501 , \6500 , \5292 );
and \U$5787 ( \6502 , \6499 , \6501 );
and \U$5788 ( \6503 , \5295 , \5351_nGffe );
and \U$5789 ( \6504 , \5471_nGf21 , \5203 );
nor \U$5790 ( \6505 , \6502 , \6503 , \6504 );
xor \U$5791 ( \6506 , \6498 , \6505 );
nand \U$5792 ( \6507 , \5751_nGabb , \4857 );
or \U$5793 ( \6508 , \4771 , \5978_nGa7f );
nand \U$5794 ( \6509 , \6508 , \4863 );
and \U$5795 ( \6510 , \6507 , \6509 );
and \U$5796 ( \6511 , \4859 , \5978_nGa7f );
and \U$5797 ( \6512 , \5751_nGabb , \4918 );
nor \U$5798 ( \6513 , \6510 , \6511 , \6512 );
and \U$5799 ( \6514 , \6506 , \6513 );
and \U$5800 ( \6515 , \6498 , \6505 );
or \U$5801 ( \6516 , \6514 , \6515 );
nand \U$5802 ( \6517 , \5119_nG10fb , \5392 );
or \U$5803 ( \6518 , \5288 , \5055_nG11dc );
nand \U$5804 ( \6519 , \6518 , \5574 );
and \U$5805 ( \6520 , \6517 , \6519 );
and \U$5806 ( \6521 , \5577 , \5055_nG11dc );
and \U$5807 ( \6522 , \5119_nG10fb , \5395 );
nor \U$5808 ( \6523 , \6520 , \6521 , \6522 );
not \U$5809 ( \6524 , \6523 );
or \U$5810 ( \6525 , \5989 , \4964 );
or \U$5811 ( \6526 , \4891_nG13e1 , \5707 );
or \U$5812 ( \6527 , \4960_nG12e2 , \5706 );
nand \U$5813 ( \6528 , \6525 , \6526 , \6527 );
nand \U$5814 ( \6529 , \6524 , \6528 );
xor \U$5815 ( \6530 , \6516 , \6529 );
nand \U$5816 ( \6531 , \6181_nGa0e , \4698 );
or \U$5817 ( \6532 , \4659 , \5950_nGa4b );
nand \U$5818 ( \6533 , \6532 , \4725 );
and \U$5819 ( \6534 , \6531 , \6533 );
and \U$5820 ( \6535 , \4728 , \5950_nGa4b );
and \U$5821 ( \6536 , \6181_nGa0e , \4701 );
nor \U$5822 ( \6537 , \6534 , \6535 , \6536 );
and \U$5823 ( \6538 , RIaaa79b8_554, \723 );
and \U$5824 ( \6539 , RIaaa7c10_559, \738 );
and \U$5825 ( \6540 , \686 , RIaaa7fd0_567);
and \U$5826 ( \6541 , RIaaa7c88_560, \690 );
nor \U$5827 ( \6542 , \6540 , \6541 );
and \U$5828 ( \6543 , RIaaa7e68_564, \4572 );
and \U$5829 ( \6544 , \735 , RIaaa7b98_558);
and \U$5830 ( \6545 , RIaaa8048_568, \721 );
nor \U$5831 ( \6546 , \6543 , \6544 , \6545 );
and \U$5832 ( \6547 , \696 , RIaaa7f58_566);
and \U$5833 ( \6548 , RIaaa7df0_563, \712 );
nor \U$5834 ( \6549 , \6547 , \6548 );
nand \U$5835 ( \6550 , \6542 , \6546 , \6549 );
nor \U$5836 ( \6551 , \6538 , \6539 , \6550 );
and \U$5837 ( \6552 , \702 , RIaaa7d00_561);
and \U$5838 ( \6553 , RIaaa8138_570, \682 );
nor \U$5839 ( \6554 , \6552 , \6553 );
and \U$5840 ( \6555 , \733 , RIaaa80c0_569);
and \U$5841 ( \6556 , RIaaa7a30_555, \728 );
nor \U$5842 ( \6557 , \6555 , \6556 );
and \U$5843 ( \6558 , \699 , RIaaa7b20_557);
and \U$5844 ( \6559 , RIaaa7aa8_556, \730 );
nor \U$5845 ( \6560 , \6558 , \6559 );
nand \U$5846 ( \6561 , \6551 , \6554 , \6557 , \6560 );
_DC g964 ( \6562_nG964 , \6561 , \4592 );
nand \U$5847 ( \6563 , \6562_nG964 , \4565 );
xor \U$5848 ( \6564 , \6537 , \6563 );
and \U$5849 ( \6565 , \6295_nG9d6 , \4645 );
or \U$5850 ( \6566 , \4606 , \6467_nG99e );
nand \U$5851 ( \6567 , \6566 , \4642 );
nand \U$5852 ( \6568 , \6295_nG9d6 , \4638 );
and \U$5853 ( \6569 , \6567 , \6568 );
and \U$5854 ( \6570 , \6467_nG99e , \4762 );
nor \U$5855 ( \6571 , \6565 , \6569 , \6570 );
and \U$5856 ( \6572 , \6564 , \6571 );
and \U$5857 ( \6573 , \6537 , \6563 );
or \U$5858 ( \6574 , \6572 , \6573 );
and \U$5859 ( \6575 , \6530 , \6574 );
and \U$5860 ( \6576 , \6516 , \6529 );
or \U$5861 ( \6577 , \6575 , \6576 );
and \U$5862 ( \6578 , \6491 , \6577 );
and \U$5863 ( \6579 , \6485 , \6490 );
or \U$5864 ( \6580 , \6578 , \6579 );
and \U$5865 ( \6581 , \6476 , \6580 );
and \U$5866 ( \6582 , \6473 , \6475 );
or \U$5867 ( \6583 , \6581 , \6582 );
nor \U$5868 ( \6584 , \6428 , \6583 );
xor \U$5869 ( \6585 , \6424 , \6584 );
and \U$5870 ( \6586 , \6428 , \6583 );
nor \U$5871 ( \6587 , \6586 , \6584 );
xor \U$5872 ( \6588 , \6473 , \6475 );
xor \U$5873 ( \6589 , \6588 , \6580 );
xor \U$5874 ( \6590 , \6353 , \6403 );
xor \U$5875 ( \6591 , \6590 , \6406 );
nor \U$5876 ( \6592 , \6589 , \6591 );
xor \U$5877 ( \6593 , \6587 , \6592 );
and \U$5878 ( \6594 , \6589 , \6591 );
nor \U$5879 ( \6595 , \6594 , \6592 );
nand \U$5880 ( \6596 , \5978_nGa7f , \4857 );
or \U$5881 ( \6597 , \4771 , \5950_nGa4b );
nand \U$5882 ( \6598 , \6597 , \4863 );
and \U$5883 ( \6599 , \6596 , \6598 );
and \U$5884 ( \6600 , \4859 , \5950_nGa4b );
and \U$5885 ( \6601 , \5978_nGa7f , \4918 );
nor \U$5886 ( \6602 , \6599 , \6600 , \6601 );
and \U$5887 ( \6603 , \5656_nGaf0 , \5125 );
or \U$5888 ( \6604 , \4934 , \5656_nGaf0 );
nand \U$5889 ( \6605 , \6604 , \5128 );
nand \U$5890 ( \6606 , \5751_nGabb , \4997 );
and \U$5891 ( \6607 , \6605 , \6606 );
and \U$5892 ( \6608 , \5751_nGabb , \5000 );
nor \U$5893 ( \6609 , \6603 , \6607 , \6608 );
xor \U$5894 ( \6610 , \6602 , \6609 );
nand \U$5895 ( \6611 , \6295_nG9d6 , \4698 );
or \U$5896 ( \6612 , \4659 , \6181_nGa0e );
nand \U$5897 ( \6613 , \6612 , \4725 );
and \U$5898 ( \6614 , \6611 , \6613 );
and \U$5899 ( \6615 , \4728 , \6181_nGa0e );
and \U$5900 ( \6616 , \6295_nG9d6 , \4701 );
nor \U$5901 ( \6617 , \6614 , \6615 , \6616 );
and \U$5902 ( \6618 , \6610 , \6617 );
and \U$5903 ( \6619 , \6602 , \6609 );
or \U$5904 ( \6620 , \6618 , \6619 );
not \U$5905 ( \6621 , \5526_nGe53 );
or \U$5906 ( \6622 , \5204 , \6621 );
or \U$5907 ( \6623 , \5149 , \5471_nGf21 );
nand \U$5908 ( \6624 , \6623 , \5292 );
nand \U$5909 ( \6625 , \5526_nGe53 , \5200 );
and \U$5910 ( \6626 , \6624 , \6625 );
and \U$5911 ( \6627 , \5471_nGf21 , \5295 );
nor \U$5912 ( \6628 , \6626 , \6627 );
nand \U$5913 ( \6629 , \6622 , \6628 );
and \U$5914 ( \6630 , \4961 , \5822 );
not \U$5915 ( \6631 , \5055_nG11dc );
and \U$5916 ( \6632 , \5705 , \6631 );
and \U$5917 ( \6633 , \4960_nG12e2 , \5825 );
nor \U$5918 ( \6634 , \6630 , \6632 , \6633 );
nand \U$5919 ( \6635 , \5351_nGffe , \5392 );
or \U$5920 ( \6636 , \5288 , \5119_nG10fb );
nand \U$5921 ( \6637 , \6636 , \5574 );
and \U$5922 ( \6638 , \6635 , \6637 );
and \U$5923 ( \6639 , \5577 , \5119_nG10fb );
and \U$5924 ( \6640 , \5351_nGffe , \5395 );
nor \U$5925 ( \6641 , \6638 , \6639 , \6640 );
nand \U$5926 ( \6642 , \6634 , \6641 );
and \U$5927 ( \6643 , \6629 , \6642 );
nor \U$5928 ( \6644 , \6641 , \6634 );
nor \U$5929 ( \6645 , \6643 , \6644 );
xor \U$5930 ( \6646 , \6620 , \6645 );
xor \U$5931 ( \6647 , \6537 , \6563 );
xor \U$5932 ( \6648 , \6647 , \6571 );
and \U$5933 ( \6649 , \6646 , \6648 );
and \U$5934 ( \6650 , \6620 , \6645 );
or \U$5935 ( \6651 , \6649 , \6650 );
xor \U$5936 ( \6652 , \6498 , \6505 );
xor \U$5937 ( \6653 , \6652 , \6513 );
not \U$5938 ( \6654 , \6653 );
not \U$5939 ( \6655 , \6528 );
not \U$5940 ( \6656 , \6523 );
or \U$5941 ( \6657 , \6655 , \6656 );
or \U$5942 ( \6658 , \6523 , \6528 );
nand \U$5943 ( \6659 , \6657 , \6658 );
nand \U$5944 ( \6660 , \6654 , \6659 );
xor \U$5945 ( \6661 , \6651 , \6660 );
xor \U$5946 ( \6662 , \6478 , \6480 );
xor \U$5947 ( \6663 , \6662 , \6482 );
and \U$5948 ( \6664 , \6661 , \6663 );
and \U$5949 ( \6665 , \6651 , \6660 );
or \U$5950 ( \6666 , \6664 , \6665 );
not \U$5951 ( \6667 , \6433 );
not \U$5952 ( \6668 , \6472 );
and \U$5953 ( \6669 , \6667 , \6668 );
and \U$5954 ( \6670 , \6433 , \6472 );
nor \U$5955 ( \6671 , \6669 , \6670 );
xor \U$5956 ( \6672 , \6666 , \6671 );
xor \U$5957 ( \6673 , \6485 , \6490 );
xor \U$5958 ( \6674 , \6673 , \6577 );
and \U$5959 ( \6675 , \6672 , \6674 );
and \U$5960 ( \6676 , \6666 , \6671 );
or \U$5961 ( \6677 , \6675 , \6676 );
not \U$5962 ( \6678 , \6677 );
xor \U$5963 ( \6679 , \6595 , \6678 );
nand \U$5964 ( \6680 , \5471_nGf21 , \5392 );
or \U$5965 ( \6681 , \5288 , \5351_nGffe );
nand \U$5966 ( \6682 , \6681 , \5574 );
and \U$5967 ( \6683 , \6680 , \6682 );
and \U$5968 ( \6684 , \5577 , \5351_nGffe );
and \U$5969 ( \6685 , \5471_nGf21 , \5395 );
nor \U$5970 ( \6686 , \6683 , \6684 , \6685 );
and \U$5971 ( \6687 , \6631 , \5822 );
not \U$5972 ( \6688 , \5119_nG10fb );
and \U$5973 ( \6689 , \5705 , \6688 );
and \U$5974 ( \6690 , \5055_nG11dc , \5825 );
nor \U$5975 ( \6691 , \6687 , \6689 , \6690 );
xor \U$5976 ( \6692 , \6686 , \6691 );
and \U$5977 ( \6693 , \6692 , \4606 );
and \U$5978 ( \6694 , \6686 , \6691 );
or \U$5979 ( \6695 , \6693 , \6694 );
and \U$5980 ( \6696 , \5751_nGabb , \5125 );
or \U$5981 ( \6697 , \4934 , \5751_nGabb );
nand \U$5982 ( \6698 , \6697 , \5128 );
nand \U$5983 ( \6699 , \5978_nGa7f , \4997 );
and \U$5984 ( \6700 , \6698 , \6699 );
and \U$5985 ( \6701 , \5978_nGa7f , \5000 );
nor \U$5986 ( \6702 , \6696 , \6700 , \6701 );
nand \U$5987 ( \6703 , \5656_nGaf0 , \5200 );
or \U$5988 ( \6704 , \5149 , \5526_nGe53 );
nand \U$5989 ( \6705 , \6704 , \5292 );
and \U$5990 ( \6706 , \6703 , \6705 );
and \U$5991 ( \6707 , \5295 , \5526_nGe53 );
and \U$5992 ( \6708 , \5656_nGaf0 , \5203 );
nor \U$5993 ( \6709 , \6706 , \6707 , \6708 );
xor \U$5994 ( \6710 , \6702 , \6709 );
nand \U$5995 ( \6711 , \5950_nGa4b , \4857 );
or \U$5996 ( \6712 , \4771 , \6181_nGa0e );
nand \U$5997 ( \6713 , \6712 , \4863 );
and \U$5998 ( \6714 , \6711 , \6713 );
and \U$5999 ( \6715 , \4859 , \6181_nGa0e );
and \U$6000 ( \6716 , \5950_nGa4b , \4918 );
nor \U$6001 ( \6717 , \6714 , \6715 , \6716 );
and \U$6002 ( \6718 , \6710 , \6717 );
and \U$6003 ( \6719 , \6702 , \6709 );
or \U$6004 ( \6720 , \6718 , \6719 );
xor \U$6005 ( \6721 , \6695 , \6720 );
and \U$6006 ( \6722 , \6467_nG99e , \4645 );
or \U$6007 ( \6723 , \4606 , \6562_nG964 );
nand \U$6008 ( \6724 , \6723 , \4642 );
nand \U$6009 ( \6725 , \6467_nG99e , \4638 );
and \U$6010 ( \6726 , \6724 , \6725 );
and \U$6011 ( \6727 , \6562_nG964 , \4762 );
nor \U$6012 ( \6728 , \6722 , \6726 , \6727 );
and \U$6013 ( \6729 , \6721 , \6728 );
and \U$6014 ( \6730 , \6695 , \6720 );
or \U$6015 ( \6731 , \6729 , \6730 );
not \U$6016 ( \6732 , \6653 );
not \U$6017 ( \6733 , \6659 );
and \U$6018 ( \6734 , \6732 , \6733 );
and \U$6019 ( \6735 , \6653 , \6659 );
nor \U$6020 ( \6736 , \6734 , \6735 );
xor \U$6021 ( \6737 , \6731 , \6736 );
xor \U$6022 ( \6738 , \6620 , \6645 );
xor \U$6023 ( \6739 , \6738 , \6648 );
and \U$6024 ( \6740 , \6737 , \6739 );
and \U$6025 ( \6741 , \6731 , \6736 );
or \U$6026 ( \6742 , \6740 , \6741 );
xor \U$6027 ( \6743 , \6516 , \6529 );
xor \U$6028 ( \6744 , \6743 , \6574 );
xor \U$6029 ( \6745 , \6742 , \6744 );
xor \U$6030 ( \6746 , \6651 , \6660 );
xor \U$6031 ( \6747 , \6746 , \6663 );
and \U$6032 ( \6748 , \6745 , \6747 );
and \U$6033 ( \6749 , \6742 , \6744 );
or \U$6034 ( \6750 , \6748 , \6749 );
xor \U$6035 ( \6751 , \6666 , \6671 );
xor \U$6036 ( \6752 , \6751 , \6674 );
and \U$6037 ( \6753 , \6750 , \6752 );
xor \U$6038 ( \6754 , \6695 , \6720 );
xor \U$6039 ( \6755 , \6754 , \6728 );
not \U$6040 ( \6756 , \6755 );
not \U$6041 ( \6757 , \6644 );
nand \U$6042 ( \6758 , \6757 , \6642 );
not \U$6043 ( \6759 , \6758 );
not \U$6044 ( \6760 , \6629 );
or \U$6045 ( \6761 , \6759 , \6760 );
or \U$6046 ( \6762 , \6629 , \6758 );
nand \U$6047 ( \6763 , \6761 , \6762 );
nand \U$6048 ( \6764 , \6756 , \6763 );
nand \U$6049 ( \6765 , \6467_nG99e , \4698 );
or \U$6050 ( \6766 , \4659 , \6295_nG9d6 );
nand \U$6051 ( \6767 , \6766 , \4725 );
and \U$6052 ( \6768 , \6765 , \6767 );
and \U$6053 ( \6769 , \4728 , \6295_nG9d6 );
and \U$6054 ( \6770 , \6467_nG99e , \4701 );
nor \U$6055 ( \6771 , \6768 , \6769 , \6770 );
nand \U$6056 ( \6772 , \5526_nGe53 , \5392 );
or \U$6057 ( \6773 , \5288 , \5471_nGf21 );
nand \U$6058 ( \6774 , \6773 , \5574 );
and \U$6059 ( \6775 , \6772 , \6774 );
and \U$6060 ( \6776 , \5577 , \5471_nGf21 );
and \U$6061 ( \6777 , \5526_nGe53 , \5395 );
nor \U$6062 ( \6778 , \6775 , \6776 , \6777 );
and \U$6063 ( \6779 , \6688 , \5822 );
not \U$6064 ( \6780 , \5351_nGffe );
and \U$6065 ( \6781 , \5705 , \6780 );
and \U$6066 ( \6782 , \5119_nG10fb , \5825 );
nor \U$6067 ( \6783 , \6779 , \6781 , \6782 );
xor \U$6068 ( \6784 , \6778 , \6783 );
nand \U$6069 ( \6785 , \5751_nGabb , \5200 );
or \U$6070 ( \6786 , \5149 , \5656_nGaf0 );
nand \U$6071 ( \6787 , \6786 , \5292 );
and \U$6072 ( \6788 , \6785 , \6787 );
and \U$6073 ( \6789 , \5295 , \5656_nGaf0 );
and \U$6074 ( \6790 , \5751_nGabb , \5203 );
nor \U$6075 ( \6791 , \6788 , \6789 , \6790 );
and \U$6076 ( \6792 , \6784 , \6791 );
and \U$6077 ( \6793 , \6778 , \6783 );
or \U$6078 ( \6794 , \6792 , \6793 );
xor \U$6079 ( \6795 , \6771 , \6794 );
nand \U$6080 ( \6796 , \6181_nGa0e , \4857 );
or \U$6081 ( \6797 , \4771 , \6295_nG9d6 );
nand \U$6082 ( \6798 , \6797 , \4863 );
and \U$6083 ( \6799 , \6796 , \6798 );
and \U$6084 ( \6800 , \4859 , \6295_nG9d6 );
and \U$6085 ( \6801 , \6181_nGa0e , \4918 );
nor \U$6086 ( \6802 , \6799 , \6800 , \6801 );
and \U$6087 ( \6803 , \5978_nGa7f , \5125 );
or \U$6088 ( \6804 , \4934 , \5978_nGa7f );
nand \U$6089 ( \6805 , \6804 , \5128 );
nand \U$6090 ( \6806 , \5950_nGa4b , \4997 );
and \U$6091 ( \6807 , \6805 , \6806 );
and \U$6092 ( \6808 , \5950_nGa4b , \5000 );
nor \U$6093 ( \6809 , \6803 , \6807 , \6808 );
xor \U$6094 ( \6810 , \6802 , \6809 );
nand \U$6095 ( \6811 , \6562_nG964 , \4698 );
or \U$6096 ( \6812 , \4659 , \6467_nG99e );
nand \U$6097 ( \6813 , \6812 , \4725 );
and \U$6098 ( \6814 , \6811 , \6813 );
and \U$6099 ( \6815 , \4728 , \6467_nG99e );
and \U$6100 ( \6816 , \6562_nG964 , \4701 );
nor \U$6101 ( \6817 , \6814 , \6815 , \6816 );
and \U$6102 ( \6818 , \6810 , \6817 );
and \U$6103 ( \6819 , \6802 , \6809 );
or \U$6104 ( \6820 , \6818 , \6819 );
and \U$6105 ( \6821 , \6795 , \6820 );
and \U$6106 ( \6822 , \6771 , \6794 );
or \U$6107 ( \6823 , \6821 , \6822 );
xor \U$6108 ( \6824 , \6602 , \6609 );
xor \U$6109 ( \6825 , \6824 , \6617 );
xor \U$6110 ( \6826 , \6823 , \6825 );
xor \U$6111 ( \6827 , \6702 , \6709 );
xor \U$6112 ( \6828 , \6827 , \6717 );
xor \U$6113 ( \6829 , \6686 , \6691 );
xor \U$6114 ( \6830 , \6829 , \4606 );
and \U$6115 ( \6831 , \6828 , \6830 );
and \U$6116 ( \6832 , \4645 , \6562_nG964 );
nand \U$6117 ( \6833 , \6562_nG964 , \4638 );
and \U$6118 ( \6834 , \6833 , \4605 );
nor \U$6119 ( \6835 , \6832 , \6834 );
xor \U$6120 ( \6836 , \6686 , \6691 );
xor \U$6121 ( \6837 , \6836 , \4606 );
and \U$6122 ( \6838 , \6835 , \6837 );
and \U$6123 ( \6839 , \6828 , \6835 );
or \U$6124 ( \6840 , \6831 , \6838 , \6839 );
and \U$6125 ( \6841 , \6826 , \6840 );
and \U$6126 ( \6842 , \6823 , \6825 );
or \U$6127 ( \6843 , \6841 , \6842 );
xor \U$6128 ( \6844 , \6764 , \6843 );
xor \U$6129 ( \6845 , \6731 , \6736 );
xor \U$6130 ( \6846 , \6845 , \6739 );
and \U$6131 ( \6847 , \6844 , \6846 );
and \U$6132 ( \6848 , \6764 , \6843 );
or \U$6133 ( \6849 , \6847 , \6848 );
xor \U$6134 ( \6850 , \6742 , \6744 );
xor \U$6135 ( \6851 , \6850 , \6747 );
and \U$6136 ( \6852 , \6849 , \6851 );
and \U$6137 ( \6853 , \5950_nGa4b , \5125 );
or \U$6138 ( \6854 , \4934 , \5950_nGa4b );
nand \U$6139 ( \6855 , \6854 , \5128 );
nand \U$6140 ( \6856 , \6181_nGa0e , \4997 );
and \U$6141 ( \6857 , \6855 , \6856 );
and \U$6142 ( \6858 , \6181_nGa0e , \5000 );
nor \U$6143 ( \6859 , \6853 , \6857 , \6858 );
nand \U$6144 ( \6860 , \5978_nGa7f , \5200 );
or \U$6145 ( \6861 , \5149 , \5751_nGabb );
nand \U$6146 ( \6862 , \6861 , \5292 );
and \U$6147 ( \6863 , \6860 , \6862 );
and \U$6148 ( \6864 , \5295 , \5751_nGabb );
and \U$6149 ( \6865 , \5978_nGa7f , \5203 );
nor \U$6150 ( \6866 , \6863 , \6864 , \6865 );
xor \U$6151 ( \6867 , \6859 , \6866 );
nand \U$6152 ( \6868 , \6295_nG9d6 , \4857 );
or \U$6153 ( \6869 , \4771 , \6467_nG99e );
nand \U$6154 ( \6870 , \6869 , \4863 );
and \U$6155 ( \6871 , \6868 , \6870 );
and \U$6156 ( \6872 , \4859 , \6467_nG99e );
and \U$6157 ( \6873 , \6295_nG9d6 , \4918 );
nor \U$6158 ( \6874 , \6871 , \6872 , \6873 );
and \U$6159 ( \6875 , \6867 , \6874 );
and \U$6160 ( \6876 , \6859 , \6866 );
or \U$6161 ( \6877 , \6875 , \6876 );
nand \U$6162 ( \6878 , \5656_nGaf0 , \5392 );
or \U$6163 ( \6879 , \5288 , \5526_nGe53 );
nand \U$6164 ( \6880 , \6879 , \5574 );
and \U$6165 ( \6881 , \6878 , \6880 );
and \U$6166 ( \6882 , \5577 , \5526_nGe53 );
and \U$6167 ( \6883 , \5656_nGaf0 , \5395 );
nor \U$6168 ( \6884 , \6881 , \6882 , \6883 );
and \U$6169 ( \6885 , \6780 , \5822 );
not \U$6170 ( \6886 , \5471_nGf21 );
and \U$6171 ( \6887 , \5705 , \6886 );
and \U$6172 ( \6888 , \5351_nGffe , \5825 );
nor \U$6173 ( \6889 , \6885 , \6887 , \6888 );
xor \U$6174 ( \6890 , \6884 , \6889 );
and \U$6175 ( \6891 , \6890 , \4659 );
and \U$6176 ( \6892 , \6884 , \6889 );
or \U$6177 ( \6893 , \6891 , \6892 );
xor \U$6178 ( \6894 , \6877 , \6893 );
xor \U$6179 ( \6895 , \6802 , \6809 );
xor \U$6180 ( \6896 , \6895 , \6817 );
and \U$6181 ( \6897 , \6894 , \6896 );
and \U$6182 ( \6898 , \6877 , \6893 );
or \U$6183 ( \6899 , \6897 , \6898 );
xor \U$6184 ( \6900 , \6771 , \6794 );
xor \U$6185 ( \6901 , \6900 , \6820 );
xor \U$6186 ( \6902 , \6899 , \6901 );
xor \U$6187 ( \6903 , \6686 , \6691 );
xor \U$6188 ( \6904 , \6903 , \4606 );
xor \U$6189 ( \6905 , \6828 , \6835 );
xor \U$6190 ( \6906 , \6904 , \6905 );
and \U$6191 ( \6907 , \6902 , \6906 );
and \U$6192 ( \6908 , \6899 , \6901 );
or \U$6193 ( \6909 , \6907 , \6908 );
xor \U$6194 ( \6910 , \6823 , \6825 );
xor \U$6195 ( \6911 , \6910 , \6840 );
xor \U$6196 ( \6912 , \6909 , \6911 );
not \U$6197 ( \6913 , \6755 );
not \U$6198 ( \6914 , \6763 );
and \U$6199 ( \6915 , \6913 , \6914 );
and \U$6200 ( \6916 , \6755 , \6763 );
nor \U$6201 ( \6917 , \6915 , \6916 );
xor \U$6202 ( \6918 , \6912 , \6917 );
not \U$6203 ( \6919 , \6918 );
xor \U$6204 ( \6920 , \6899 , \6901 );
xor \U$6205 ( \6921 , \6920 , \6906 );
nand \U$6206 ( \6922 , \5751_nGabb , \5392 );
or \U$6207 ( \6923 , \5288 , \5656_nGaf0 );
nand \U$6208 ( \6924 , \6923 , \5574 );
and \U$6209 ( \6925 , \6922 , \6924 );
and \U$6210 ( \6926 , \5577 , \5656_nGaf0 );
and \U$6211 ( \6927 , \5751_nGabb , \5395 );
nor \U$6212 ( \6928 , \6925 , \6926 , \6927 );
and \U$6213 ( \6929 , \6886 , \5822 );
and \U$6214 ( \6930 , \5705 , \6621 );
and \U$6215 ( \6931 , \5471_nGf21 , \5825 );
nor \U$6216 ( \6932 , \6929 , \6930 , \6931 );
xor \U$6217 ( \6933 , \6928 , \6932 );
nand \U$6218 ( \6934 , \5950_nGa4b , \5200 );
or \U$6219 ( \6935 , \5149 , \5978_nGa7f );
nand \U$6220 ( \6936 , \6935 , \5292 );
and \U$6221 ( \6937 , \6934 , \6936 );
and \U$6222 ( \6938 , \5295 , \5978_nGa7f );
and \U$6223 ( \6939 , \5950_nGa4b , \5203 );
nor \U$6224 ( \6940 , \6937 , \6938 , \6939 );
and \U$6225 ( \6941 , \6933 , \6940 );
and \U$6226 ( \6942 , \6928 , \6932 );
or \U$6227 ( \6943 , \6941 , \6942 );
xor \U$6228 ( \6944 , \6859 , \6866 );
xor \U$6229 ( \6945 , \6944 , \6874 );
and \U$6230 ( \6946 , \6943 , \6945 );
and \U$6231 ( \6947 , \6562_nG964 , \4728 );
not \U$6232 ( \6948 , \6562_nG964 );
and \U$6233 ( \6949 , \6948 , \4700 );
not \U$6234 ( \6950 , \4725 );
nor \U$6235 ( \6951 , \6947 , \6949 , \6950 );
xor \U$6236 ( \6952 , \6859 , \6866 );
xor \U$6237 ( \6953 , \6952 , \6874 );
and \U$6238 ( \6954 , \6951 , \6953 );
and \U$6239 ( \6955 , \6943 , \6951 );
or \U$6240 ( \6956 , \6946 , \6954 , \6955 );
xor \U$6241 ( \6957 , \6778 , \6783 );
xor \U$6242 ( \6958 , \6957 , \6791 );
xor \U$6243 ( \6959 , \6956 , \6958 );
xor \U$6244 ( \6960 , \6877 , \6893 );
xor \U$6245 ( \6961 , \6960 , \6896 );
and \U$6246 ( \6962 , \6959 , \6961 );
and \U$6247 ( \6963 , \6956 , \6958 );
or \U$6248 ( \6964 , \6962 , \6963 );
nor \U$6249 ( \6965 , \6921 , \6964 );
xor \U$6250 ( \6966 , \6919 , \6965 );
and \U$6251 ( \6967 , \6921 , \6964 );
nor \U$6252 ( \6968 , \6967 , \6965 );
xor \U$6253 ( \6969 , \6956 , \6958 );
xor \U$6254 ( \6970 , \6969 , \6961 );
nand \U$6255 ( \6971 , \5978_nGa7f , \5392 );
or \U$6256 ( \6972 , \5288 , \5751_nGabb );
nand \U$6257 ( \6973 , \6972 , \5574 );
and \U$6258 ( \6974 , \6971 , \6973 );
and \U$6259 ( \6975 , \5577 , \5751_nGabb );
and \U$6260 ( \6976 , \5978_nGa7f , \5395 );
nor \U$6261 ( \6977 , \6974 , \6975 , \6976 );
and \U$6262 ( \6978 , \6621 , \5822 );
not \U$6263 ( \6979 , \5656_nGaf0 );
and \U$6264 ( \6980 , \5705 , \6979 );
and \U$6265 ( \6981 , \5526_nGe53 , \5825 );
nor \U$6266 ( \6982 , \6978 , \6980 , \6981 );
xor \U$6267 ( \6983 , \6977 , \6982 );
and \U$6268 ( \6984 , \6983 , \4771 );
and \U$6269 ( \6985 , \6977 , \6982 );
or \U$6270 ( \6986 , \6984 , \6985 );
and \U$6271 ( \6987 , \6181_nGa0e , \5125 );
or \U$6272 ( \6988 , \4934 , \6181_nGa0e );
nand \U$6273 ( \6989 , \6988 , \5128 );
nand \U$6274 ( \6990 , \6295_nG9d6 , \4997 );
and \U$6275 ( \6991 , \6989 , \6990 );
and \U$6276 ( \6992 , \6295_nG9d6 , \5000 );
nor \U$6277 ( \6993 , \6987 , \6991 , \6992 );
xor \U$6278 ( \6994 , \6986 , \6993 );
and \U$6279 ( \6995 , \6295_nG9d6 , \5125 );
or \U$6280 ( \6996 , \4934 , \6295_nG9d6 );
nand \U$6281 ( \6997 , \6996 , \5128 );
nand \U$6282 ( \6998 , \6467_nG99e , \4997 );
and \U$6283 ( \6999 , \6997 , \6998 );
and \U$6284 ( \7000 , \6467_nG99e , \5000 );
nor \U$6285 ( \7001 , \6995 , \6999 , \7000 );
nand \U$6286 ( \7002 , \6181_nGa0e , \5200 );
or \U$6287 ( \7003 , \5149 , \5950_nGa4b );
nand \U$6288 ( \7004 , \7003 , \5292 );
and \U$6289 ( \7005 , \7002 , \7004 );
and \U$6290 ( \7006 , \5295 , \5950_nGa4b );
and \U$6291 ( \7007 , \6181_nGa0e , \5203 );
nor \U$6292 ( \7008 , \7005 , \7006 , \7007 );
xor \U$6293 ( \7009 , \7001 , \7008 );
and \U$6294 ( \7010 , \4918 , \6562_nG964 );
nand \U$6295 ( \7011 , \6562_nG964 , \4857 );
and \U$6296 ( \7012 , \7011 , \4861 );
nor \U$6297 ( \7013 , \7010 , \7012 );
and \U$6298 ( \7014 , \7009 , \7013 );
and \U$6299 ( \7015 , \7001 , \7008 );
or \U$6300 ( \7016 , \7014 , \7015 );
and \U$6301 ( \7017 , \6994 , \7016 );
and \U$6302 ( \7018 , \6986 , \6993 );
or \U$6303 ( \7019 , \7017 , \7018 );
xor \U$6304 ( \7020 , \6884 , \6889 );
xor \U$6305 ( \7021 , \7020 , \4659 );
nand \U$6306 ( \7022 , \7019 , \7021 );
not \U$6307 ( \7023 , \6467_nG99e );
or \U$6308 ( \7024 , \5006 , \7023 );
or \U$6309 ( \7025 , \6948 , \5008 );
or \U$6310 ( \7026 , \4917 , \7023 );
or \U$6311 ( \7027 , \4771 , \6562_nG964 );
nand \U$6312 ( \7028 , \7027 , \4863 );
nand \U$6313 ( \7029 , \7026 , \7028 );
nand \U$6314 ( \7030 , \7024 , \7025 , \7029 );
not \U$6315 ( \7031 , \7030 );
xor \U$6316 ( \7032 , \6928 , \6932 );
xor \U$6317 ( \7033 , \7032 , \6940 );
nor \U$6318 ( \7034 , \7031 , \7033 );
and \U$6319 ( \7035 , \7022 , \7034 );
nor \U$6320 ( \7036 , \7019 , \7021 );
nor \U$6321 ( \7037 , \7035 , \7036 );
nor \U$6322 ( \7038 , \6970 , \7037 );
xor \U$6323 ( \7039 , \6968 , \7038 );
not \U$6324 ( \7040 , \7034 );
not \U$6325 ( \7041 , \7036 );
nand \U$6326 ( \7042 , \7041 , \7022 );
not \U$6327 ( \7043 , \7042 );
or \U$6328 ( \7044 , \7040 , \7043 );
or \U$6329 ( \7045 , \7042 , \7034 );
nand \U$6330 ( \7046 , \7044 , \7045 );
xor \U$6331 ( \7047 , \6859 , \6866 );
xor \U$6332 ( \7048 , \7047 , \6874 );
xor \U$6333 ( \7049 , \6943 , \6951 );
xor \U$6334 ( \7050 , \7048 , \7049 );
not \U$6335 ( \7051 , \7050 );
xor \U$6336 ( \7052 , \7046 , \7051 );
not \U$6337 ( \7053 , \6295_nG9d6 );
or \U$6338 ( \7054 , \5204 , \7053 );
or \U$6339 ( \7055 , \5149 , \6181_nGa0e );
nand \U$6340 ( \7056 , \7055 , \5292 );
nand \U$6341 ( \7057 , \6295_nG9d6 , \5200 );
and \U$6342 ( \7058 , \7056 , \7057 );
and \U$6343 ( \7059 , \6181_nGa0e , \5295 );
nor \U$6344 ( \7060 , \7058 , \7059 );
nand \U$6345 ( \7061 , \7054 , \7060 );
and \U$6346 ( \7062 , \6979 , \5822 );
not \U$6347 ( \7063 , \5751_nGabb );
and \U$6348 ( \7064 , \5705 , \7063 );
and \U$6349 ( \7065 , \5656_nGaf0 , \5825 );
nor \U$6350 ( \7066 , \7062 , \7064 , \7065 );
nand \U$6351 ( \7067 , \5950_nGa4b , \5392 );
or \U$6352 ( \7068 , \5288 , \5978_nGa7f );
nand \U$6353 ( \7069 , \7068 , \5574 );
and \U$6354 ( \7070 , \7067 , \7069 );
and \U$6355 ( \7071 , \5577 , \5978_nGa7f );
and \U$6356 ( \7072 , \5950_nGa4b , \5395 );
nor \U$6357 ( \7073 , \7070 , \7071 , \7072 );
nand \U$6358 ( \7074 , \7066 , \7073 );
and \U$6359 ( \7075 , \7061 , \7074 );
nor \U$6360 ( \7076 , \7073 , \7066 );
nor \U$6361 ( \7077 , \7075 , \7076 );
xor \U$6362 ( \7078 , \6977 , \6982 );
xor \U$6363 ( \7079 , \7078 , \4771 );
and \U$6364 ( \7080 , \7077 , \7079 );
xor \U$6365 ( \7081 , \7001 , \7008 );
xor \U$6366 ( \7082 , \7081 , \7013 );
xor \U$6367 ( \7083 , \6977 , \6982 );
xor \U$6368 ( \7084 , \7083 , \4771 );
and \U$6369 ( \7085 , \7082 , \7084 );
and \U$6370 ( \7086 , \7077 , \7082 );
or \U$6371 ( \7087 , \7080 , \7085 , \7086 );
xor \U$6372 ( \7088 , \6986 , \6993 );
xor \U$6373 ( \7089 , \7088 , \7016 );
and \U$6374 ( \7090 , \7087 , \7089 );
not \U$6375 ( \7091 , \7090 );
not \U$6376 ( \7092 , \7030 );
not \U$6377 ( \7093 , \7033 );
and \U$6378 ( \7094 , \7092 , \7093 );
and \U$6379 ( \7095 , \7030 , \7033 );
nor \U$6380 ( \7096 , \7094 , \7095 );
not \U$6381 ( \7097 , \7096 );
and \U$6382 ( \7098 , \7091 , \7097 );
nor \U$6383 ( \7099 , \7087 , \7089 );
nor \U$6384 ( \7100 , \7098 , \7099 );
not \U$6385 ( \7101 , \7100 );
xor \U$6386 ( \7102 , \7052 , \7101 );
or \U$6387 ( \7103 , \7099 , \7090 );
not \U$6388 ( \7104 , \7103 );
not \U$6389 ( \7105 , \7096 );
and \U$6390 ( \7106 , \7104 , \7105 );
and \U$6391 ( \7107 , \7103 , \7096 );
nor \U$6392 ( \7108 , \7106 , \7107 );
xor \U$6393 ( \7109 , \6977 , \6982 );
xor \U$6394 ( \7110 , \7109 , \4771 );
xor \U$6395 ( \7111 , \7077 , \7082 );
xor \U$6396 ( \7112 , \7110 , \7111 );
nand \U$6397 ( \7113 , \6181_nGa0e , \5392 );
or \U$6398 ( \7114 , \5288 , \5950_nGa4b );
nand \U$6399 ( \7115 , \7114 , \5574 );
and \U$6400 ( \7116 , \7113 , \7115 );
and \U$6401 ( \7117 , \5577 , \5950_nGa4b );
and \U$6402 ( \7118 , \6181_nGa0e , \5395 );
nor \U$6403 ( \7119 , \7116 , \7117 , \7118 );
and \U$6404 ( \7120 , \7063 , \5822 );
not \U$6405 ( \7121 , \5978_nGa7f );
and \U$6406 ( \7122 , \5705 , \7121 );
and \U$6407 ( \7123 , \5751_nGabb , \5825 );
nor \U$6408 ( \7124 , \7120 , \7122 , \7123 );
xor \U$6409 ( \7125 , \7119 , \7124 );
and \U$6410 ( \7126 , \7125 , \4934 );
and \U$6411 ( \7127 , \7119 , \7124 );
or \U$6412 ( \7128 , \7126 , \7127 );
and \U$6413 ( \7129 , \6467_nG99e , \5125 );
or \U$6414 ( \7130 , \4934 , \6467_nG99e );
nand \U$6415 ( \7131 , \7130 , \5128 );
nand \U$6416 ( \7132 , \6562_nG964 , \4997 );
and \U$6417 ( \7133 , \7131 , \7132 );
and \U$6418 ( \7134 , \6562_nG964 , \5000 );
nor \U$6419 ( \7135 , \7129 , \7133 , \7134 );
nand \U$6420 ( \7136 , \7128 , \7135 );
or \U$6421 ( \7137 , \5209 , \6948 );
or \U$6422 ( \7138 , \6562_nG964 , \4934 );
nand \U$6423 ( \7139 , \7137 , \7138 , \5128 );
not \U$6424 ( \7140 , \7139 );
nand \U$6425 ( \7141 , \6467_nG99e , \5200 );
or \U$6426 ( \7142 , \5149 , \6295_nG9d6 );
nand \U$6427 ( \7143 , \7142 , \5292 );
and \U$6428 ( \7144 , \7141 , \7143 );
and \U$6429 ( \7145 , \5295 , \6295_nG9d6 );
and \U$6430 ( \7146 , \6467_nG99e , \5203 );
nor \U$6431 ( \7147 , \7144 , \7145 , \7146 );
nor \U$6432 ( \7148 , \7140 , \7147 );
and \U$6433 ( \7149 , \7136 , \7148 );
nor \U$6434 ( \7150 , \7135 , \7128 );
nor \U$6435 ( \7151 , \7149 , \7150 );
nor \U$6436 ( \7152 , \7112 , \7151 );
xor \U$6437 ( \7153 , \7108 , \7152 );
nand \U$6438 ( \7154 , \6295_nG9d6 , \5392 );
or \U$6439 ( \7155 , \5288 , \6181_nGa0e );
nand \U$6440 ( \7156 , \7155 , \5574 );
and \U$6441 ( \7157 , \7154 , \7156 );
and \U$6442 ( \7158 , \5577 , \6181_nGa0e );
and \U$6443 ( \7159 , \6295_nG9d6 , \5395 );
nor \U$6444 ( \7160 , \7157 , \7158 , \7159 );
and \U$6445 ( \7161 , \7121 , \5822 );
not \U$6446 ( \7162 , \5950_nGa4b );
and \U$6447 ( \7163 , \5705 , \7162 );
and \U$6448 ( \7164 , \5978_nGa7f , \5825 );
nor \U$6449 ( \7165 , \7161 , \7163 , \7164 );
xor \U$6450 ( \7166 , \7160 , \7165 );
nand \U$6451 ( \7167 , \6562_nG964 , \5200 );
or \U$6452 ( \7168 , \5149 , \6467_nG99e );
nand \U$6453 ( \7169 , \7168 , \5292 );
and \U$6454 ( \7170 , \7167 , \7169 );
and \U$6455 ( \7171 , \5295 , \6467_nG99e );
and \U$6456 ( \7172 , \6562_nG964 , \5203 );
nor \U$6457 ( \7173 , \7170 , \7171 , \7172 );
xor \U$6458 ( \7174 , \7166 , \7173 );
and \U$6459 ( \7175 , \7162 , \5822 );
not \U$6460 ( \7176 , \6181_nGa0e );
and \U$6461 ( \7177 , \5705 , \7176 );
and \U$6462 ( \7178 , \5950_nGa4b , \5825 );
nor \U$6463 ( \7179 , \7175 , \7177 , \7178 );
xor \U$6464 ( \7180 , \5149 , \7179 );
nand \U$6465 ( \7181 , \6467_nG99e , \5392 );
or \U$6466 ( \7182 , \5288 , \6295_nG9d6 );
nand \U$6467 ( \7183 , \7182 , \5574 );
and \U$6468 ( \7184 , \7181 , \7183 );
and \U$6469 ( \7185 , \5577 , \6295_nG9d6 );
and \U$6470 ( \7186 , \6467_nG99e , \5395 );
nor \U$6471 ( \7187 , \7184 , \7185 , \7186 );
and \U$6472 ( \7188 , \7180 , \7187 );
and \U$6473 ( \7189 , \5149 , \7179 );
or \U$6474 ( \7190 , \7188 , \7189 );
nor \U$6475 ( \7191 , \7174 , \7190 );
not \U$6476 ( \7192 , \7191 );
xor \U$6477 ( \7193 , \5149 , \7179 );
xor \U$6478 ( \7194 , \7193 , \7187 );
not \U$6479 ( \7195 , \7194 );
not \U$6480 ( \7196 , \5295 );
or \U$6481 ( \7197 , \7196 , \6948 );
or \U$6482 ( \7198 , \6562_nG964 , \5149 );
nand \U$6483 ( \7199 , \7197 , \7198 , \5292 );
not \U$6484 ( \7200 , \7199 );
or \U$6485 ( \7201 , \7195 , \7200 );
or \U$6486 ( \7202 , \7199 , \7194 );
nand \U$6487 ( \7203 , \7201 , \7202 );
nand \U$6488 ( \7204 , \6562_nG964 , \5392 );
or \U$6489 ( \7205 , \5288 , \6467_nG99e );
nand \U$6490 ( \7206 , \7205 , \5574 );
and \U$6491 ( \7207 , \7204 , \7206 );
and \U$6492 ( \7208 , \5577 , \6467_nG99e );
and \U$6493 ( \7209 , \6562_nG964 , \5395 );
nor \U$6494 ( \7210 , \7207 , \7208 , \7209 );
and \U$6495 ( \7211 , \7176 , \5822 );
and \U$6496 ( \7212 , \5705 , \7053 );
and \U$6497 ( \7213 , \6181_nGa0e , \5825 );
nor \U$6498 ( \7214 , \7211 , \7212 , \7213 );
nor \U$6499 ( \7215 , \7210 , \7214 );
not \U$6500 ( \7216 , \7215 );
and \U$6501 ( \7217 , \5704 , \6467_nG99e );
nor \U$6502 ( \7218 , \7217 , \5282 , \6562_nG964 );
not \U$6503 ( \7219 , \7218 );
not \U$6504 ( \7220 , \5577 );
or \U$6505 ( \7221 , \7220 , \6948 );
or \U$6506 ( \7222 , \6562_nG964 , \5288 );
nand \U$6507 ( \7223 , \7221 , \7222 , \5574 );
not \U$6508 ( \7224 , \7223 );
or \U$6509 ( \7225 , \7219 , \7224 );
or \U$6510 ( \7226 , \7223 , \7218 );
or \U$6511 ( \7227 , \5989 , \7053 );
or \U$6512 ( \7228 , \6295_nG9d6 , \5707 );
or \U$6513 ( \7229 , \6467_nG99e , \5706 );
nand \U$6514 ( \7230 , \7227 , \7228 , \7229 );
xor \U$6515 ( \7231 , \7230 , \5394 );
nand \U$6516 ( \7232 , \7226 , \7231 );
nand \U$6517 ( \7233 , \7225 , \7232 );
and \U$6518 ( \7234 , \7233 , \7230 , \5394 );
and \U$6519 ( \7235 , \7210 , \7214 );
and \U$6520 ( \7236 , \7230 , \5394 );
nor \U$6521 ( \7237 , \7233 , \7236 );
nor \U$6522 ( \7238 , \7235 , \7237 );
nor \U$6523 ( \7239 , \7234 , \7238 );
nand \U$6524 ( \7240 , \7216 , \7239 );
and \U$6525 ( \7241 , \7203 , \7240 );
and \U$6526 ( \7242 , \7233 , \7236 );
and \U$6527 ( \7243 , \7215 , \7242 );
nor \U$6528 ( \7244 , \7241 , \7243 );
not \U$6529 ( \7245 , \7194 );
nand \U$6530 ( \7246 , \7245 , \7199 );
or \U$6531 ( \7247 , \7192 , \7244 , \7246 );
and \U$6532 ( \7248 , \7174 , \7190 , \7246 );
nor \U$6533 ( \7249 , \7248 , \7244 );
and \U$6534 ( \7250 , \7174 , \7190 );
nor \U$6535 ( \7251 , \7250 , \7246 );
nor \U$6536 ( \7252 , \7249 , \7251 , \7191 );
xor \U$6537 ( \7253 , \7160 , \7165 );
and \U$6538 ( \7254 , \7253 , \7173 );
and \U$6539 ( \7255 , \7160 , \7165 );
or \U$6540 ( \7256 , \7254 , \7255 );
xor \U$6541 ( \7257 , \7119 , \7124 );
xor \U$6542 ( \7258 , \7257 , \4934 );
xor \U$6543 ( \7259 , \7256 , \7258 );
not \U$6544 ( \7260 , \7139 );
not \U$6545 ( \7261 , \7147 );
and \U$6546 ( \7262 , \7260 , \7261 );
and \U$6547 ( \7263 , \7139 , \7147 );
nor \U$6548 ( \7264 , \7262 , \7263 );
xor \U$6549 ( \7265 , \7259 , \7264 );
or \U$6550 ( \7266 , \7252 , \7265 );
nand \U$6551 ( \7267 , \7247 , \7266 );
xor \U$6552 ( \7268 , \7256 , \7258 );
and \U$6553 ( \7269 , \7268 , \7264 );
and \U$6554 ( \7270 , \7256 , \7258 );
or \U$6555 ( \7271 , \7269 , \7270 );
not \U$6556 ( \7272 , \7271 );
xor \U$6557 ( \7273 , \7267 , \7272 );
not \U$6558 ( \7274 , \7076 );
nand \U$6559 ( \7275 , \7274 , \7074 );
not \U$6560 ( \7276 , \7275 );
not \U$6561 ( \7277 , \7061 );
or \U$6562 ( \7278 , \7276 , \7277 );
or \U$6563 ( \7279 , \7061 , \7275 );
nand \U$6564 ( \7280 , \7278 , \7279 );
not \U$6565 ( \7281 , \7148 );
not \U$6566 ( \7282 , \7150 );
nand \U$6567 ( \7283 , \7282 , \7136 );
not \U$6568 ( \7284 , \7283 );
or \U$6569 ( \7285 , \7281 , \7284 );
or \U$6570 ( \7286 , \7283 , \7148 );
nand \U$6571 ( \7287 , \7285 , \7286 );
xor \U$6572 ( \7288 , \7280 , \7287 );
and \U$6573 ( \7289 , \7273 , \7288 );
and \U$6574 ( \7290 , \7267 , \7272 );
or \U$6575 ( \7291 , \7289 , \7290 );
and \U$6576 ( \7292 , \7280 , \7287 );
xor \U$6577 ( \7293 , \7291 , \7292 );
and \U$6578 ( \7294 , \7112 , \7151 );
nor \U$6579 ( \7295 , \7294 , \7152 );
and \U$6580 ( \7296 , \7293 , \7295 );
and \U$6581 ( \7297 , \7291 , \7292 );
or \U$6582 ( \7298 , \7296 , \7297 );
and \U$6583 ( \7299 , \7153 , \7298 );
and \U$6584 ( \7300 , \7108 , \7152 );
or \U$6585 ( \7301 , \7299 , \7300 );
and \U$6586 ( \7302 , \7102 , \7301 );
and \U$6587 ( \7303 , \7052 , \7101 );
or \U$6588 ( \7304 , \7302 , \7303 );
and \U$6589 ( \7305 , \7046 , \7051 );
xor \U$6590 ( \7306 , \7304 , \7305 );
and \U$6591 ( \7307 , \6970 , \7037 );
nor \U$6592 ( \7308 , \7307 , \7038 );
and \U$6593 ( \7309 , \7306 , \7308 );
and \U$6594 ( \7310 , \7304 , \7305 );
or \U$6595 ( \7311 , \7309 , \7310 );
and \U$6596 ( \7312 , \7039 , \7311 );
and \U$6597 ( \7313 , \6968 , \7038 );
or \U$6598 ( \7314 , \7312 , \7313 );
and \U$6599 ( \7315 , \6966 , \7314 );
and \U$6600 ( \7316 , \6919 , \6965 );
or \U$6601 ( \7317 , \7315 , \7316 );
xor \U$6602 ( \7318 , \6909 , \6911 );
and \U$6603 ( \7319 , \7318 , \6917 );
and \U$6604 ( \7320 , \6909 , \6911 );
or \U$6605 ( \7321 , \7319 , \7320 );
xor \U$6606 ( \7322 , \6764 , \6843 );
xor \U$6607 ( \7323 , \7322 , \6846 );
nand \U$6608 ( \7324 , \7321 , \7323 );
and \U$6609 ( \7325 , \7317 , \7324 );
nor \U$6610 ( \7326 , \7323 , \7321 );
nor \U$6611 ( \7327 , \7325 , \7326 );
xor \U$6612 ( \7328 , \6742 , \6744 );
xor \U$6613 ( \7329 , \7328 , \6747 );
and \U$6614 ( \7330 , \7327 , \7329 );
and \U$6615 ( \7331 , \6849 , \7327 );
or \U$6616 ( \7332 , \6852 , \7330 , \7331 );
xor \U$6617 ( \7333 , \6666 , \6671 );
xor \U$6618 ( \7334 , \7333 , \6674 );
and \U$6619 ( \7335 , \7332 , \7334 );
and \U$6620 ( \7336 , \6750 , \7332 );
or \U$6621 ( \7337 , \6753 , \7335 , \7336 );
not \U$6622 ( \7338 , \7337 );
and \U$6623 ( \7339 , \6679 , \7338 );
and \U$6624 ( \7340 , \6595 , \6678 );
or \U$6625 ( \7341 , \7339 , \7340 );
and \U$6626 ( \7342 , \6593 , \7341 );
and \U$6627 ( \7343 , \6587 , \6592 );
or \U$6628 ( \7344 , \7342 , \7343 );
and \U$6629 ( \7345 , \6585 , \7344 );
and \U$6630 ( \7346 , \6424 , \6584 );
or \U$6631 ( \7347 , \7345 , \7346 );
xor \U$6632 ( \7348 , \6414 , \6419 );
and \U$6633 ( \7349 , \7348 , \6422 );
and \U$6634 ( \7350 , \6414 , \6419 );
or \U$6635 ( \7351 , \7349 , \7350 );
xor \U$6636 ( \7352 , \6309 , \6323 );
xor \U$6637 ( \7353 , \7352 , \6334 );
nand \U$6638 ( \7354 , \7351 , \7353 );
and \U$6639 ( \7355 , \7347 , \7354 );
nor \U$6640 ( \7356 , \7353 , \7351 );
nor \U$6641 ( \7357 , \7355 , \7356 );
and \U$6642 ( \7358 , \6338 , \7357 );
and \U$6643 ( \7359 , \6147 , \6337 );
or \U$6644 ( \7360 , \7358 , \7359 );
not \U$6645 ( \7361 , \7360 );
and \U$6646 ( \7362 , \6140 , \7361 );
and \U$6647 ( \7363 , \6055 , \6139 );
or \U$6648 ( \7364 , \7362 , \7363 );
xor \U$6649 ( \7365 , \5867 , \5879 );
xor \U$6650 ( \7366 , \7365 , \5882 );
or \U$6651 ( \7367 , \6044 , \6051 );
nand \U$6652 ( \7368 , \7367 , \6042 );
nand \U$6653 ( \7369 , \7366 , \7368 );
and \U$6654 ( \7370 , \7364 , \7369 );
nor \U$6655 ( \7371 , \7368 , \7366 );
nor \U$6656 ( \7372 , \7370 , \7371 );
and \U$6657 ( \7373 , \5886 , \7372 );
and \U$6658 ( \7374 , \5789 , \5885 );
or \U$6659 ( \7375 , \7373 , \7374 );
not \U$6660 ( \7376 , \7375 );
and \U$6661 ( \7377 , \5782 , \7376 );
and \U$6662 ( \7378 , \5626 , \5781 );
or \U$6663 ( \7379 , \7377 , \7378 );
and \U$6664 ( \7380 , \5622 , \7379 );
and \U$6665 ( \7381 , \5489 , \5621 );
or \U$6666 ( \7382 , \7380 , \7381 );
and \U$6667 ( \7383 , \5487 , \7382 );
and \U$6668 ( \7384 , \5381 , \5486 );
or \U$6669 ( \7385 , \7383 , \7384 );
and \U$6670 ( \7386 , \5379 , \7385 );
and \U$6671 ( \7387 , \5376 , \5378 );
or \U$6672 ( \7388 , \7386 , \7387 );
and \U$6673 ( \7389 , \5272 , \7388 );
and \U$6674 ( \7390 , \5186 , \5271 );
or \U$6675 ( \7391 , \7389 , \7390 );
and \U$6676 ( \7392 , \5184 , \7391 );
and \U$6677 ( \7393 , \5181 , \5183 );
or \U$6678 ( \7394 , \7392 , \7393 );
and \U$6679 ( \7395 , \5078 , \7394 );
and \U$6680 ( \7396 , \4910 , \5077 );
or \U$6681 ( \7397 , \7395 , \7396 );
and \U$6682 ( \7398 , \4908 , \7397 );
and \U$6683 ( \7399 , \4906 , \4907 );
or \U$6684 ( \7400 , \7398 , \7399 );
not \U$6685 ( \7401 , \7400 );
or \U$6686 ( \7402 , \4804 , \7401 );
or \U$6687 ( \7403 , \7400 , \4803 );
nand \U$6688 ( \7404 , \7402 , \7403 );
buf \U$6689 ( \7405 , \4293 );
buf \U$6690 ( \7406 , \749 );
_DC g4e5 ( \7407_nG4e5 , \7405 , \7406 );
not \U$6691 ( \7408 , \7407_nG4e5 );
buf \U$6692 ( \7409 , \4322 );
_DC g506 ( \7410_nG506 , \7409 , \7406 );
not \U$6693 ( \7411 , \7410_nG506 );
buf \U$6694 ( \7412 , \1146 );
buf \U$6695 ( \7413 , \749 );
_DC g5c2 ( \7414_nG5c2 , \7412 , \7413 );
not \U$6696 ( \7415 , \7414_nG5c2 );
not \U$6697 ( \7416 , \7415 );
buf \U$6698 ( \7417 , \4496 );
_DC g5c4 ( \7418_nG5c4 , \7417 , \7406 );
not \U$6699 ( \7419 , \7418_nG5c4 );
and \U$6700 ( \7420 , \7416 , \7419 );
buf \U$6701 ( \7421 , \1179 );
_DC g5e3 ( \7422_nG5e3 , \7421 , \7413 );
nor \U$6702 ( \7423 , \7420 , \7422_nG5e3 );
buf \U$6703 ( \7424 , \4524 );
_DC g5e5 ( \7425_nG5e5 , \7424 , \7406 );
and \U$6704 ( \7426 , \7423 , \7425_nG5e5 );
and \U$6705 ( \7427 , \7418_nG5c4 , \7415 );
nor \U$6706 ( \7428 , \7426 , \7427 );
buf \U$6707 ( \7429 , \4467 );
_DC g5a5 ( \7430_nG5a5 , \7429 , \7406 );
not \U$6708 ( \7431 , \7430_nG5a5 );
and \U$6709 ( \7432 , \7428 , \7431 );
buf \U$6710 ( \7433 , \1115 );
_DC g5a3 ( \7434_nG5a3 , \7433 , \7413 );
or \U$6711 ( \7435 , \7432 , \7434_nG5a3 );
or \U$6712 ( \7436 , \7431 , \7428 );
nand \U$6713 ( \7437 , \7435 , \7436 );
buf \U$6714 ( \7438 , \4438 );
_DC g586 ( \7439_nG586 , \7438 , \7406 );
and \U$6715 ( \7440 , \7437 , \7439_nG586 );
not \U$6716 ( \7441 , \7437 );
not \U$6717 ( \7442 , \7439_nG586 );
and \U$6718 ( \7443 , \7441 , \7442 );
buf \U$6719 ( \7444 , \1079 );
_DC g584 ( \7445_nG584 , \7444 , \7413 );
nor \U$6720 ( \7446 , \7443 , \7445_nG584 );
nor \U$6721 ( \7447 , \7440 , \7446 );
buf \U$6722 ( \7448 , \4409 );
_DC g567 ( \7449_nG567 , \7448 , \7406 );
not \U$6723 ( \7450 , \7449_nG567 );
buf \U$6724 ( \7451 , \1047 );
_DC g565 ( \7452_nG565 , \7451 , \7413 );
and \U$6725 ( \7453 , \7450 , \7452_nG565 );
or \U$6726 ( \7454 , \7447 , \7453 );
or \U$6727 ( \7455 , \7452_nG565 , \7450 );
nand \U$6728 ( \7456 , \7454 , \7455 );
buf \U$6729 ( \7457 , \4380 );
_DC g546 ( \7458_nG546 , \7457 , \7406 );
and \U$6730 ( \7459 , \7456 , \7458_nG546 );
not \U$6731 ( \7460 , \7456 );
not \U$6732 ( \7461 , \7458_nG546 );
and \U$6733 ( \7462 , \7460 , \7461 );
buf \U$6734 ( \7463 , \1009 );
_DC g544 ( \7464_nG544 , \7463 , \7413 );
nor \U$6735 ( \7465 , \7462 , \7464_nG544 );
nor \U$6736 ( \7466 , \7459 , \7465 );
buf \U$6737 ( \7467 , \4351 );
_DC g527 ( \7468_nG527 , \7467 , \7406 );
not \U$6738 ( \7469 , \7468_nG527 );
buf \U$6739 ( \7470 , \973 );
_DC g525 ( \7471_nG525 , \7470 , \7413 );
and \U$6740 ( \7472 , \7469 , \7471_nG525 );
or \U$6741 ( \7473 , \7466 , \7472 );
or \U$6742 ( \7474 , \7471_nG525 , \7469 );
nand \U$6743 ( \7475 , \7473 , \7474 );
not \U$6744 ( \7476 , \7475 );
or \U$6745 ( \7477 , \7411 , \7476 );
nor \U$6746 ( \7478 , \7475 , \7410_nG506 );
buf \U$6747 ( \7479 , \935 );
_DC g504 ( \7480_nG504 , \7479 , \7413 );
or \U$6748 ( \7481 , \7478 , \7480_nG504 );
nand \U$6749 ( \7482 , \7477 , \7481 );
not \U$6750 ( \7483 , \7482 );
or \U$6751 ( \7484 , \7408 , \7483 );
nor \U$6752 ( \7485 , \7482 , \7407_nG4e5 );
buf \U$6753 ( \7486 , \897 );
_DC g4e3 ( \7487_nG4e3 , \7486 , \7413 );
or \U$6754 ( \7488 , \7485 , \7487_nG4e3 );
nand \U$6755 ( \7489 , \7484 , \7488 );
buf \U$6756 ( \7490 , \4264 );
_DC g4c4 ( \7491_nG4c4 , \7490 , \7406 );
and \U$6757 ( \7492 , \7489 , \7491_nG4c4 );
not \U$6758 ( \7493 , \7489 );
not \U$6759 ( \7494 , \7491_nG4c4 );
and \U$6760 ( \7495 , \7493 , \7494 );
buf \U$6761 ( \7496 , \859 );
_DC g4c2 ( \7497_nG4c2 , \7496 , \7413 );
nor \U$6762 ( \7498 , \7495 , \7497_nG4c2 );
nor \U$6763 ( \7499 , \7492 , \7498 );
buf \U$6764 ( \7500 , \4236 );
_DC g4a3 ( \7501_nG4a3 , \7500 , \7406 );
not \U$6765 ( \7502 , \7501_nG4a3 );
buf \U$6766 ( \7503 , \821 );
_DC g4a1 ( \7504_nG4a1 , \7503 , \7413 );
and \U$6767 ( \7505 , \7502 , \7504_nG4a1 );
or \U$6768 ( \7506 , \7499 , \7505 );
or \U$6769 ( \7507 , \7504_nG4a1 , \7502 );
nand \U$6770 ( \7508 , \7506 , \7507 );
buf \U$6771 ( \7509 , \4207 );
_DC g484 ( \7510_nG484 , \7509 , \7406 );
and \U$6772 ( \7511 , \7508 , \7510_nG484 );
not \U$6773 ( \7512 , \7508 );
not \U$6774 ( \7513 , \7510_nG484 );
and \U$6775 ( \7514 , \7512 , \7513 );
buf \U$6776 ( \7515 , \785 );
_DC g482 ( \7516_nG482 , \7515 , \7413 );
nor \U$6777 ( \7517 , \7514 , \7516_nG482 );
nor \U$6778 ( \7518 , \7511 , \7517 );
buf \U$6779 ( \7519 , \4177 );
_DC g465 ( \7520_nG465 , \7519 , \7406 );
not \U$6780 ( \7521 , \7520_nG465 );
buf \U$6781 ( \7522 , \745 );
_DC g462 ( \7523_nG462 , \7522 , \7413 );
and \U$6782 ( \7524 , \7521 , \7523_nG462 );
or \U$6783 ( \7525 , \7518 , \7524 );
or \U$6784 ( \7526 , \7523_nG462 , \7521 );
nand \U$6785 ( \7527 , \7525 , \7526 );
nor \U$6786 ( \7528 , \652 , RIaaa89a8_588);
and \U$6787 ( \7529 , RIaa97860_5, \7528 );
nand \U$6788 ( \7530 , RIaa978d8_6, \7529 );
not \U$6789 ( \7531 , \7530 );
nand \U$6790 ( \7532 , RIaa97950_7, \7531 );
not \U$6791 ( \7533 , \7532 );
nand \U$6792 ( \7534 , RIaa979c8_8, \7533 );
not \U$6793 ( \7535 , \7534 );
nand \U$6794 ( \7536 , RIaa97ba8_12, \7535 );
nor \U$6795 ( \7537 , \7536 , \827 );
nand \U$6796 ( \7538 , RIaa97ab8_10, \7537 );
not \U$6797 ( \7539 , \7538 );
or \U$6798 ( \7540 , \7539 , RIaa97a40_9);
nand \U$6799 ( \7541 , RIaa97a40_9, \7539 );
nand \U$6800 ( \7542 , \7540 , \7541 );
not \U$6801 ( \7543 , \7542 );
buf \U$6802 ( \7544 , \4207 );
buf \U$6803 ( \7545 , \749 );
_DC g301 ( \7546_nG301 , \7544 , \7545 );
not \U$6804 ( \7547 , \7546_nG301 );
and \U$6805 ( \7548 , \7543 , \7547 );
and \U$6806 ( \7549 , \7546_nG301 , \7542 );
buf \U$6807 ( \7550 , \4264 );
_DC g33a ( \7551_nG33a , \7550 , \7545 );
not \U$6808 ( \7552 , \7551_nG33a );
not \U$6809 ( \7553 , \7536 );
not \U$6810 ( \7554 , RIaa97b30_11);
and \U$6811 ( \7555 , \7553 , \7554 );
and \U$6812 ( \7556 , \7536 , RIaa97b30_11);
nor \U$6813 ( \7557 , \7555 , \7556 );
not \U$6814 ( \7558 , \7557 );
or \U$6815 ( \7559 , \7552 , \7558 );
or \U$6816 ( \7560 , \7557 , \7551_nG33a );
buf \U$6817 ( \7561 , \4293 );
_DC g357 ( \7562_nG357 , \7561 , \7545 );
or \U$6818 ( \7563 , \7535 , RIaa97ba8_12);
nand \U$6819 ( \7564 , \7563 , \7536 );
or \U$6820 ( \7565 , \7562_nG357 , \7564 );
not \U$6821 ( \7566 , \7562_nG357 );
not \U$6822 ( \7567 , \7564 );
or \U$6823 ( \7568 , \7566 , \7567 );
buf \U$6824 ( \7569 , \4351 );
_DC g391 ( \7570_nG391 , \7569 , \7545 );
not \U$6825 ( \7571 , \7570_nG391 );
buf \U$6826 ( \7572 , \4380 );
_DC g3ae ( \7573_nG3ae , \7572 , \7545 );
not \U$6827 ( \7574 , \7573_nG3ae );
xor \U$6828 ( \7575 , RIaa97860_5, \7528 );
buf \U$6829 ( \7576 , \4409 );
_DC g3cb ( \7577_nG3cb , \7576 , \7545 );
not \U$6830 ( \7578 , \7577_nG3cb );
or \U$6831 ( \7579 , \7575 , \7578 );
not \U$6832 ( \7580 , \7578 );
not \U$6833 ( \7581 , \7575 );
or \U$6834 ( \7582 , \7580 , \7581 );
buf \U$6835 ( \7583 , \4438 );
_DC g3e8 ( \7584_nG3e8 , \7583 , \7545 );
not \U$6836 ( \7585 , \7584_nG3e8 );
buf \U$6837 ( \7586 , \4467 );
_DC g405 ( \7587_nG405 , \7586 , \7545 );
not \U$6838 ( \7588 , \7587_nG405 );
nor \U$6839 ( \7589 , \1083 , RIaaa89a8_588);
xnor \U$6840 ( \7590 , RIaa97770_3, \7589 );
not \U$6841 ( \7591 , \7590 );
or \U$6842 ( \7592 , \7588 , \7591 );
buf \U$6843 ( \7593 , \4496 );
_DC g422 ( \7594_nG422 , \7593 , \7545 );
buf \U$6844 ( \7595 , \4524 );
_DC g43e ( \7596_nG43e , \7595 , \7545 );
and \U$6845 ( \7597 , \1182 , \7596_nG43e );
and \U$6846 ( \7598 , \7594_nG422 , \7597 );
and \U$6847 ( \7599 , RIaaa89a8_588, \1083 );
nor \U$6848 ( \7600 , \7598 , \7599 , \7589 );
or \U$6849 ( \7601 , \7590 , \7587_nG405 );
or \U$6850 ( \7602 , \7594_nG422 , \7597 );
nand \U$6851 ( \7603 , \7601 , \7602 );
or \U$6852 ( \7604 , \7600 , \7603 );
nand \U$6853 ( \7605 , \7592 , \7604 );
not \U$6854 ( \7606 , \7605 );
or \U$6855 ( \7607 , \7585 , \7606 );
or \U$6856 ( \7608 , \7605 , \7584_nG3e8 );
not \U$6857 ( \7609 , RIaaa89a8_588);
and \U$6858 ( \7610 , \651 , \7609 );
nor \U$6859 ( \7611 , \7610 , RIaa976f8_2);
or \U$6860 ( \7612 , \7611 , \7528 );
nand \U$6861 ( \7613 , \7608 , \7612 );
nand \U$6862 ( \7614 , \7607 , \7613 );
nand \U$6863 ( \7615 , \7582 , \7614 );
nand \U$6864 ( \7616 , \7579 , \7615 );
not \U$6865 ( \7617 , \7616 );
or \U$6866 ( \7618 , \7574 , \7617 );
or \U$6867 ( \7619 , \7616 , \7573_nG3ae );
or \U$6868 ( \7620 , \7529 , RIaa978d8_6);
nand \U$6869 ( \7621 , \7620 , \7530 );
nand \U$6870 ( \7622 , \7619 , \7621 );
nand \U$6871 ( \7623 , \7618 , \7622 );
not \U$6872 ( \7624 , \7623 );
or \U$6873 ( \7625 , \7571 , \7624 );
or \U$6874 ( \7626 , \7623 , \7570_nG391 );
or \U$6875 ( \7627 , \7531 , RIaa97950_7);
nand \U$6876 ( \7628 , \7627 , \7532 );
nand \U$6877 ( \7629 , \7626 , \7628 );
nand \U$6878 ( \7630 , \7625 , \7629 );
buf \U$6879 ( \7631 , \4322 );
_DC g374 ( \7632_nG374 , \7631 , \7545 );
or \U$6880 ( \7633 , \7630 , \7632_nG374 );
or \U$6881 ( \7634 , \7533 , RIaa979c8_8);
nand \U$6882 ( \7635 , \7634 , \7534 );
and \U$6883 ( \7636 , \7633 , \7635 );
and \U$6884 ( \7637 , \7632_nG374 , \7630 );
nor \U$6885 ( \7638 , \7636 , \7637 );
nand \U$6886 ( \7639 , \7568 , \7638 );
nand \U$6887 ( \7640 , \7560 , \7565 , \7639 );
nand \U$6888 ( \7641 , \7559 , \7640 );
or \U$6889 ( \7642 , \7537 , RIaa97ab8_10);
nand \U$6890 ( \7643 , \7642 , \7538 );
or \U$6891 ( \7644 , \7641 , \7643 );
buf \U$6892 ( \7645 , \4236 );
_DC g31e ( \7646_nG31e , \7645 , \7545 );
and \U$6893 ( \7647 , \7644 , \7646_nG31e );
and \U$6894 ( \7648 , \7643 , \7641 );
nor \U$6895 ( \7649 , \7549 , \7647 , \7648 );
nor \U$6896 ( \7650 , \7548 , \7649 );
buf \U$6897 ( \7651 , \4177 );
_DC g2e4 ( \7652_nG2e4 , \7651 , \7545 );
or \U$6898 ( \7653 , \7650 , \7652_nG2e4 );
not \U$6899 ( \7654 , \7652_nG2e4 );
not \U$6900 ( \7655 , \7650 );
or \U$6901 ( \7656 , \7654 , \7655 );
not \U$6902 ( \7657 , RIaa97680_1);
not \U$6903 ( \7658 , \7541 );
or \U$6904 ( \7659 , \7657 , \7658 );
or \U$6905 ( \7660 , \7541 , RIaa97680_1);
nand \U$6906 ( \7661 , \7659 , \7660 );
nand \U$6907 ( \7662 , \7656 , \7661 );
nand \U$6908 ( \7663 , \7653 , \7662 );
and \U$6909 ( \7664 , \7527 , \7663 , \677 , \716 );
_HMUX g21fd_GF_PartitionCandidate ( \7665_nG21fd , \4152 , \7404 , \7664 );
buf \U$6910 ( \7666 , \7665_nG21fd );
xor \U$6911 ( \7667 , \4145 , \4144 );
xor \U$6912 ( \7668 , \4906 , \4907 );
xor \U$6913 ( \7669 , \7668 , \7397 );
_HMUX g21c3_GF_PartitionCandidate ( \7670_nG21c3 , \7667 , \7669 , \7664 );
buf \U$6914 ( \7671 , \7670_nG21c3 );
xor \U$6915 ( \7672 , \1572 , \1743 );
xor \U$6916 ( \7673 , \7672 , \4136 );
xor \U$6917 ( \7674 , \4910 , \5077 );
xor \U$6918 ( \7675 , \7674 , \7394 );
_HMUX g2194_GF_PartitionCandidate ( \7676_nG2194 , \7673 , \7675 , \7664 );
buf \U$6919 ( \7677 , \7676_nG2194 );
xor \U$6920 ( \7678 , \1852 , \1854 );
xor \U$6921 ( \7679 , \7678 , \4133 );
xor \U$6922 ( \7680 , \5181 , \5183 );
xor \U$6923 ( \7681 , \7680 , \7391 );
_HMUX g215b_GF_PartitionCandidate ( \7682_nG215b , \7679 , \7681 , \7664 );
buf \U$6924 ( \7683 , \7682_nG215b );
xor \U$6925 ( \7684 , \1857 , \1943 );
xor \U$6926 ( \7685 , \7684 , \4130 );
xor \U$6927 ( \7686 , \5186 , \5271 );
xor \U$6928 ( \7687 , \7686 , \7388 );
_HMUX g20f7_GF_PartitionCandidate ( \7688_nG20f7 , \7685 , \7687 , \7664 );
buf \U$6929 ( \7689 , \7688_nG20f7 );
xor \U$6930 ( \7690 , \2057 , \2059 );
xor \U$6931 ( \7691 , \7690 , \4127 );
xor \U$6932 ( \7692 , \5376 , \5378 );
xor \U$6933 ( \7693 , \7692 , \7385 );
_HMUX g208a_GF_PartitionCandidate ( \7694_nG208a , \7691 , \7693 , \7664 );
buf \U$6934 ( \7695 , \7694_nG208a );
xor \U$6935 ( \7696 , \2171 , \2175 );
xor \U$6936 ( \7697 , \7696 , \4124 );
xor \U$6937 ( \7698 , \5381 , \5486 );
xor \U$6938 ( \7699 , \7698 , \7382 );
_HMUX g2017_GF_PartitionCandidate ( \7700_nG2017 , \7697 , \7699 , \7664 );
buf \U$6939 ( \7701 , \7700_nG2017 );
xor \U$6940 ( \7702 , \2183 , \2322 );
xor \U$6941 ( \7703 , \7702 , \4120 );
not \U$6942 ( \7704 , \7703 );
xor \U$6943 ( \7705 , \5489 , \5621 );
xor \U$6944 ( \7706 , \7705 , \7379 );
_HMUX g1f99_GF_PartitionCandidate ( \7707_nG1f99 , \7704 , \7706 , \7664 );
buf \U$6945 ( \7708 , \7707_nG1f99 );
xor \U$6946 ( \7709 , \2185 , \2192 );
xor \U$6947 ( \7710 , \7709 , \2319 );
xor \U$6948 ( \7711 , \2485 , \4115 );
xor \U$6949 ( \7712 , \7710 , \7711 );
not \U$6950 ( \7713 , \7712 );
xor \U$6951 ( \7714 , \5626 , \5781 );
xor \U$6952 ( \7715 , \7714 , \7376 );
_HMUX g1eee_GF_PartitionCandidate ( \7716_nG1eee , \7713 , \7715 , \7664 );
buf \U$6953 ( \7717 , \7716_nG1eee );
xor \U$6954 ( \7718 , \2474 , \2479 );
xor \U$6955 ( \7719 , \7718 , \2482 );
xor \U$6956 ( \7720 , \2587 , \4110 );
xor \U$6957 ( \7721 , \7719 , \7720 );
not \U$6958 ( \7722 , \7721 );
xor \U$6959 ( \7723 , \5789 , \5885 );
xor \U$6960 ( \7724 , \7723 , \7372 );
not \U$6961 ( \7725 , \7724 );
_HMUX g1e36_GF_PartitionCandidate ( \7726_nG1e36 , \7722 , \7725 , \7664 );
buf \U$6962 ( \7727 , \7726_nG1e36 );
not \U$6963 ( \7728 , \4109 );
nand \U$6964 ( \7729 , \7728 , \4107 );
not \U$6965 ( \7730 , \7729 );
not \U$6966 ( \7731 , \4102 );
or \U$6967 ( \7732 , \7730 , \7731 );
or \U$6968 ( \7733 , \4102 , \7729 );
nand \U$6969 ( \7734 , \7732 , \7733 );
not \U$6970 ( \7735 , \7371 );
nand \U$6971 ( \7736 , \7735 , \7369 );
not \U$6972 ( \7737 , \7736 );
not \U$6973 ( \7738 , \7364 );
or \U$6974 ( \7739 , \7737 , \7738 );
or \U$6975 ( \7740 , \7364 , \7736 );
nand \U$6976 ( \7741 , \7739 , \7740 );
_HMUX g1d83_GF_PartitionCandidate ( \7742_nG1d83 , \7734 , \7741 , \7664 );
buf \U$6977 ( \7743 , \7742_nG1d83 );
xor \U$6978 ( \7744 , \2767 , \2847 );
xor \U$6979 ( \7745 , \7744 , \4099 );
xor \U$6980 ( \7746 , \6055 , \6139 );
xor \U$6981 ( \7747 , \7746 , \7361 );
_HMUX g1ca7_GF_PartitionCandidate ( \7748_nG1ca7 , \7745 , \7747 , \7664 );
buf \U$6982 ( \7749 , \7748_nG1ca7 );
xor \U$6983 ( \7750 , \2855 , \3049 );
xor \U$6984 ( \7751 , \7750 , \4095 );
not \U$6985 ( \7752 , \7751 );
xor \U$6986 ( \7753 , \6147 , \6337 );
xor \U$6987 ( \7754 , \7753 , \7357 );
not \U$6988 ( \7755 , \7754 );
_HMUX g1bcd_GF_PartitionCandidate ( \7756_nG1bcd , \7752 , \7755 , \7664 );
buf \U$6989 ( \7757 , \7756_nG1bcd );
not \U$6990 ( \7758 , \4094 );
nand \U$6991 ( \7759 , \7758 , \4091 );
not \U$6992 ( \7760 , \7759 );
not \U$6993 ( \7761 , \4083 );
or \U$6994 ( \7762 , \7760 , \7761 );
or \U$6995 ( \7763 , \4083 , \7759 );
nand \U$6996 ( \7764 , \7762 , \7763 );
not \U$6997 ( \7765 , \7356 );
nand \U$6998 ( \7766 , \7765 , \7354 );
not \U$6999 ( \7767 , \7766 );
not \U$7000 ( \7768 , \7347 );
or \U$7001 ( \7769 , \7767 , \7768 );
or \U$7002 ( \7770 , \7347 , \7766 );
nand \U$7003 ( \7771 , \7769 , \7770 );
_HMUX g1af9_GF_PartitionCandidate ( \7772_nG1af9 , \7764 , \7771 , \7664 );
buf \U$7004 ( \7773 , \7772_nG1af9 );
xor \U$7005 ( \7774 , \3143 , \3313 );
xor \U$7006 ( \7775 , \7774 , \4080 );
xor \U$7007 ( \7776 , \6424 , \6584 );
xor \U$7008 ( \7777 , \7776 , \7344 );
_HMUX g19e9_GF_PartitionCandidate ( \7778_nG19e9 , \7775 , \7777 , \7664 );
buf \U$7009 ( \7779 , \7778_nG19e9 );
xor \U$7010 ( \7780 , \3316 , \3326 );
xor \U$7011 ( \7781 , \7780 , \4077 );
xor \U$7012 ( \7782 , \6587 , \6592 );
xor \U$7013 ( \7783 , \7782 , \7341 );
_HMUX g18d0_GF_PartitionCandidate ( \7784_nG18d0 , \7781 , \7783 , \7664 );
buf \U$7014 ( \7785 , \7784_nG18d0 );
xor \U$7015 ( \7786 , \3329 , \3411 );
xor \U$7016 ( \7787 , \7786 , \4073 );
not \U$7017 ( \7788 , \7787 );
xor \U$7018 ( \7789 , \6595 , \6678 );
xor \U$7019 ( \7790 , \7789 , \7338 );
_HMUX g17c2_GF_PartitionCandidate ( \7791_nG17c2 , \7788 , \7790 , \7664 );
buf \U$7020 ( \7792 , \7791_nG17c2 );
xor \U$7021 ( \7793 , \3331 , \3336 );
xor \U$7022 ( \7794 , \7793 , \3408 );
xor \U$7023 ( \7795 , \3485 , \4068 );
xor \U$7024 ( \7796 , \7794 , \7795 );
not \U$7025 ( \7797 , \7796 );
xor \U$7026 ( \7798 , \6666 , \6671 );
xor \U$7027 ( \7799 , \7798 , \6674 );
xor \U$7028 ( \7800 , \6750 , \7332 );
xor \U$7029 ( \7801 , \7799 , \7800 );
not \U$7030 ( \7802 , \7801 );
_HMUX g16bb_GF_PartitionCandidate ( \7803_nG16bb , \7797 , \7802 , \7664 );
buf \U$7031 ( \7804 , \7803_nG16bb );
xor \U$7032 ( \7805 , \3475 , \3477 );
xor \U$7033 ( \7806 , \7805 , \3482 );
xor \U$7034 ( \7807 , \3577 , \4063 );
xor \U$7035 ( \7808 , \7806 , \7807 );
not \U$7036 ( \7809 , \7808 );
xor \U$7037 ( \7810 , \6742 , \6744 );
xor \U$7038 ( \7811 , \7810 , \6747 );
xor \U$7039 ( \7812 , \6849 , \7327 );
xor \U$7040 ( \7813 , \7811 , \7812 );
not \U$7041 ( \7814 , \7813 );
_HMUX g1596_GF_PartitionCandidate ( \7815_nG1596 , \7809 , \7814 , \7664 );
buf \U$7042 ( \7816 , \7815_nG1596 );
not \U$7043 ( \7817 , \4062 );
nand \U$7044 ( \7818 , \7817 , \4060 );
not \U$7045 ( \7819 , \7818 );
not \U$7046 ( \7820 , \4053 );
or \U$7047 ( \7821 , \7819 , \7820 );
or \U$7048 ( \7822 , \4053 , \7818 );
nand \U$7049 ( \7823 , \7821 , \7822 );
not \U$7050 ( \7824 , \7326 );
nand \U$7051 ( \7825 , \7824 , \7324 );
not \U$7052 ( \7826 , \7825 );
not \U$7053 ( \7827 , \7317 );
or \U$7054 ( \7828 , \7826 , \7827 );
or \U$7055 ( \7829 , \7317 , \7825 );
nand \U$7056 ( \7830 , \7828 , \7829 );
_HMUX g14ad_GF_PartitionCandidate ( \7831_nG14ad , \7823 , \7830 , \7664 );
buf \U$7057 ( \7832 , \7831_nG14ad );
xor \U$7058 ( \7833 , \3643 , \3690 );
xor \U$7059 ( \7834 , \7833 , \4050 );
xor \U$7060 ( \7835 , \6919 , \6965 );
xor \U$7061 ( \7836 , \7835 , \7314 );
_HMUX g13ad_GF_PartitionCandidate ( \7837_nG13ad , \7834 , \7836 , \7664 );
buf \U$7062 ( \7838 , \7837_nG13ad );
xor \U$7063 ( \7839 , \3693 , \3763 );
xor \U$7064 ( \7840 , \7839 , \4047 );
xor \U$7065 ( \7841 , \6968 , \7038 );
xor \U$7066 ( \7842 , \7841 , \7311 );
_HMUX g12ae_GF_PartitionCandidate ( \7843_nG12ae , \7840 , \7842 , \7664 );
buf \U$7067 ( \7844 , \7843_nG12ae );
xor \U$7068 ( \7845 , \4040 , \4041 );
xor \U$7069 ( \7846 , \7845 , \4044 );
xor \U$7070 ( \7847 , \7304 , \7305 );
xor \U$7071 ( \7848 , \7847 , \7308 );
_HMUX g11a4_GF_PartitionCandidate ( \7849_nG11a4 , \7846 , \7848 , \7664 );
buf \U$7072 ( \7850 , \7849_nG11a4 );
xor \U$7073 ( \7851 , \3777 , \3826 );
xor \U$7074 ( \7852 , \7851 , \4037 );
xor \U$7075 ( \7853 , \7052 , \7101 );
xor \U$7076 ( \7854 , \7853 , \7301 );
_HMUX g10c7_GF_PartitionCandidate ( \7855_nG10c7 , \7852 , \7854 , \7664 );
buf \U$7077 ( \7856 , \7855_nG10c7 );
xor \U$7078 ( \7857 , \3833 , \3877 );
xor \U$7079 ( \7858 , \7857 , \4034 );
xor \U$7080 ( \7859 , \7108 , \7152 );
xor \U$7081 ( \7860 , \7859 , \7298 );
_HMUX gfc2_GF_PartitionCandidate ( \7861_nGfc2 , \7858 , \7860 , \7664 );
buf \U$7082 ( \7862 , \7861_nGfc2 );
xor \U$7083 ( \7863 , \4027 , \4028 );
xor \U$7084 ( \7864 , \7863 , \4031 );
xor \U$7085 ( \7865 , \7291 , \7292 );
xor \U$7086 ( \7866 , \7865 , \7295 );
_HMUX geed_GF_PartitionCandidate ( \7867_nGeed , \7864 , \7866 , \7664 );
buf \U$7087 ( \7868 , \7867_nGeed );
xor \U$7088 ( \7869 , \3892 , \3928 );
xor \U$7089 ( \7870 , \7869 , \4024 );
xor \U$7090 ( \7871 , \7267 , \7272 );
xor \U$7091 ( \7872 , \7871 , \7288 );
_HMUX ge16_GF_PartitionCandidate ( \7873_nGe16 , \7870 , \7872 , \7664 );
buf \U$7092 ( \7874 , \7873_nGe16 );
and \U$7093 ( \7875 , RIaaa9128_604, RIaaa91a0_605);
nand \U$7094 ( \7876 , RIaaa90b0_603, \7875 );
not \U$7095 ( \7877 , \7876 );
nand \U$7096 ( \7878 , \7877 , RIaaa9218_606);
not \U$7097 ( \7879 , \7878 );
nand \U$7098 ( \7880 , \7879 , RIaaa9290_607);
not \U$7099 ( \7881 , \7880 );
nand \U$7100 ( \7882 , \7881 , RIaaa9308_608);
not \U$7101 ( \7883 , \7882 );
nand \U$7102 ( \7884 , \7883 , RIaaa9380_609);
not \U$7103 ( \7885 , \7884 );
nand \U$7104 ( \7886 , \7885 , RIaaa93f8_610);
not \U$7105 ( \7887 , \7886 );
nand \U$7106 ( \7888 , \7887 , RIaaa9038_602);
not \U$7107 ( \7889 , \7888 );
nand \U$7108 ( \7890 , \7889 , RIaaa9470_611);
not \U$7109 ( \7891 , \7890 );
nand \U$7110 ( \7892 , \7891 , RIaaa94e8_612);
not \U$7111 ( \7893 , \7892 );
not \U$7112 ( \7894 , RIaaa95d8_614);
and \U$7113 ( \7895 , \7893 , \7894 );
and \U$7114 ( \7896 , \7892 , RIaaa95d8_614);
nor \U$7115 ( \7897 , \7895 , \7896 );
nor \U$7116 ( \7898 , RIaaa8de0_597, RIaaa8b88_592);
not \U$7117 ( \7899 , \7898 );
or \U$7118 ( \7900 , RIaaa8cf0_595, RIaaa8c78_594, RIaaa8b10_591, RIaaa8c00_593);
nor \U$7119 ( \7901 , \7899 , \7900 , RIaaa8d68_596, RIaaa8a98_590);
not \U$7120 ( \7902 , \7901 );
nor \U$7121 ( \7903 , \7902 , RIaaa8a20_589);
nand \U$7122 ( \7904 , RIaaa8f48_600, \7903 );
not \U$7123 ( \7905 , RIaaa8fc0_601);
nor \U$7124 ( \7906 , \7904 , \7905 );
not \U$7125 ( \7907 , RIaaa8e58_598);
nor \U$7126 ( \7908 , \7907 , RIaaa8ed0_599);
and \U$7127 ( \7909 , \7906 , \7908 );
and \U$7128 ( \7910 , RIaa98418_30, \7909 );
nor \U$7129 ( \7911 , RIaaa8ed0_599, RIaaa8e58_598);
not \U$7130 ( \7912 , \7911 );
nor \U$7131 ( \7913 , \7912 , RIaaa8fc0_601, RIaaa8f48_600);
and \U$7132 ( \7914 , \7903 , \7913 );
and \U$7133 ( \7915 , RIaa97e78_18, \7914 );
not \U$7134 ( \7916 , RIaaa8f48_600);
nand \U$7135 ( \7917 , \7916 , \7903 );
nor \U$7136 ( \7918 , \7917 , \7905 );
and \U$7137 ( \7919 , \7918 , \7908 );
and \U$7138 ( \7920 , \7919 , RIaa98238_26);
and \U$7139 ( \7921 , RIaaa8ed0_599, RIaaa8e58_598);
not \U$7140 ( \7922 , \7921 );
nor \U$7141 ( \7923 , \7922 , \7904 );
and \U$7142 ( \7924 , \7923 , \7905 );
and \U$7143 ( \7925 , RIaa980d0_23, \7924 );
nor \U$7144 ( \7926 , \7920 , \7925 );
nor \U$7145 ( \7927 , \7917 , RIaaa8fc0_601);
and \U$7146 ( \7928 , \7927 , \7921 );
and \U$7147 ( \7929 , \7928 , RIaa982b0_27);
and \U$7148 ( \7930 , \7918 , \7921 );
and \U$7149 ( \7931 , RIaa98328_28, \7930 );
nor \U$7150 ( \7932 , \7929 , \7931 );
not \U$7151 ( \7933 , RIaaa8ed0_599);
nor \U$7152 ( \7934 , \7933 , RIaaa8e58_598);
and \U$7153 ( \7935 , \7918 , \7934 );
and \U$7154 ( \7936 , \7935 , RIaa98508_32);
not \U$7155 ( \7937 , \7903 );
nand \U$7156 ( \7938 , RIaaa8fc0_601, \7921 , RIaaa8f48_600);
nor \U$7157 ( \7939 , \7937 , \7938 );
and \U$7158 ( \7940 , RIaa98148_24, \7939 );
nor \U$7159 ( \7941 , \7936 , \7940 );
and \U$7160 ( \7942 , \7927 , \7908 );
and \U$7161 ( \7943 , \7942 , RIaa981c0_25);
and \U$7162 ( \7944 , \7906 , \7934 );
and \U$7163 ( \7945 , RIaa985f8_34, \7944 );
nor \U$7164 ( \7946 , \7943 , \7945 );
nand \U$7165 ( \7947 , \7926 , \7932 , \7941 , \7946 );
nor \U$7166 ( \7948 , \7910 , \7915 , \7947 );
and \U$7167 ( \7949 , \7918 , \7911 );
and \U$7168 ( \7950 , \7949 , RIaa97ef0_19);
nor \U$7169 ( \7951 , \7904 , RIaaa8fc0_601);
and \U$7170 ( \7952 , \7951 , \7911 );
and \U$7171 ( \7953 , RIaa97fe0_21, \7952 );
nor \U$7172 ( \7954 , \7950 , \7953 );
and \U$7173 ( \7955 , \7913 , \7901 , RIaaa8a20_589);
nand \U$7174 ( \7956 , RIaa97f68_20, \7955 );
and \U$7175 ( \7957 , \7951 , \7934 );
and \U$7176 ( \7958 , RIaa98490_31, \7957 );
and \U$7177 ( \7959 , \7951 , \7908 );
and \U$7178 ( \7960 , RIaa983a0_29, \7959 );
and \U$7179 ( \7961 , \7927 , \7934 );
and \U$7180 ( \7962 , \7961 , RIaa98580_33);
and \U$7181 ( \7963 , \7906 , \7911 );
and \U$7182 ( \7964 , RIaa98058_22, \7963 );
nor \U$7183 ( \7965 , \7962 , \7964 );
not \U$7184 ( \7966 , \7965 );
nor \U$7185 ( \7967 , \7958 , \7960 , \7966 );
nand \U$7186 ( \7968 , \7948 , \7954 , \7956 , \7967 );
buf \U$7187 ( \7969 , \7968 );
not \U$7188 ( \7970 , \7913 );
nand \U$7189 ( \7971 , \7970 , RIaaa8a20_589);
nand \U$7190 ( \7972 , \7971 , \7901 );
buf \U$7191 ( \7973 , \7972 );
_DC g2a78 ( \7974_nG2a78 , \7969 , \7973 );
xor \U$7192 ( \7975 , \7897 , \7974_nG2a78 );
not \U$7193 ( \7976 , \7890 );
not \U$7194 ( \7977 , RIaaa94e8_612);
and \U$7195 ( \7978 , \7976 , \7977 );
and \U$7196 ( \7979 , \7890 , RIaaa94e8_612);
nor \U$7197 ( \7980 , \7978 , \7979 );
and \U$7198 ( \7981 , \7959 , RIaa98b98_46);
and \U$7199 ( \7982 , \7928 , RIaa98c88_48);
and \U$7200 ( \7983 , RIaa98c10_47, \7909 );
nor \U$7201 ( \7984 , \7982 , \7983 );
and \U$7202 ( \7985 , \7935 , RIaa98df0_51);
nand \U$7203 ( \7986 , RIaa98760_37, \7955 );
not \U$7204 ( \7987 , \7986 );
nor \U$7205 ( \7988 , \7985 , \7987 );
and \U$7206 ( \7989 , \7930 , RIaa98aa8_44);
and \U$7207 ( \7990 , RIaa98850_39, \7939 );
nor \U$7208 ( \7991 , \7989 , \7990 );
and \U$7209 ( \7992 , \7942 , RIaa989b8_42);
and \U$7210 ( \7993 , RIaa98d00_49, \7944 );
nor \U$7211 ( \7994 , \7992 , \7993 );
nand \U$7212 ( \7995 , \7984 , \7988 , \7991 , \7994 );
and \U$7213 ( \7996 , \7952 , RIaa988c8_40);
and \U$7214 ( \7997 , RIaa98d78_50, \7957 );
nor \U$7215 ( \7998 , \7996 , \7997 );
not \U$7216 ( \7999 , \7998 );
nor \U$7217 ( \8000 , \7981 , \7995 , \7999 );
and \U$7218 ( \8001 , \7949 , RIaa98670_35);
and \U$7219 ( \8002 , RIaa98940_41, \7963 );
nor \U$7220 ( \8003 , \8001 , \8002 );
and \U$7221 ( \8004 , \7961 , RIaa98b20_45);
and \U$7222 ( \8005 , RIaa98a30_43, \7919 );
nor \U$7223 ( \8006 , \8004 , \8005 );
and \U$7224 ( \8007 , \7914 , RIaa986e8_36);
and \U$7225 ( \8008 , RIaa987d8_38, \7924 );
nor \U$7226 ( \8009 , \8007 , \8008 );
nand \U$7227 ( \8010 , \8000 , \8003 , \8006 , \8009 );
buf \U$7228 ( \8011 , \8010 );
_DC g2898 ( \8012_nG2898 , \8011 , \7973 );
xor \U$7229 ( \8013 , \7980 , \8012_nG2898 );
not \U$7230 ( \8014 , \7888 );
not \U$7231 ( \8015 , RIaaa9470_611);
and \U$7232 ( \8016 , \8014 , \8015 );
and \U$7233 ( \8017 , \7888 , RIaaa9470_611);
nor \U$7234 ( \8018 , \8016 , \8017 );
and \U$7235 ( \8019 , \7959 , RIaa9e3b8_234);
and \U$7236 ( \8020 , \7928 , RIaa9e2c8_232);
and \U$7237 ( \8021 , RIaa9e430_235, \7909 );
nor \U$7238 ( \8022 , \8020 , \8021 );
and \U$7239 ( \8023 , \7949 , RIaa9de90_223);
nand \U$7240 ( \8024 , RIaa9df80_225, \7955 );
not \U$7241 ( \8025 , \8024 );
nor \U$7242 ( \8026 , \8023 , \8025 );
and \U$7243 ( \8027 , \7930 , RIaa9e340_233);
and \U$7244 ( \8028 , RIaa9e160_229, \7939 );
nor \U$7245 ( \8029 , \8027 , \8028 );
and \U$7246 ( \8030 , \7961 , RIaa9e598_238);
and \U$7247 ( \8031 , RIaa9e070_227, \7963 );
nor \U$7248 ( \8032 , \8030 , \8031 );
nand \U$7249 ( \8033 , \8022 , \8026 , \8029 , \8032 );
and \U$7250 ( \8034 , \7952 , RIaa9dff8_226);
and \U$7251 ( \8035 , RIaa9e4a8_236, \7957 );
nor \U$7252 ( \8036 , \8034 , \8035 );
not \U$7253 ( \8037 , \8036 );
nor \U$7254 ( \8038 , \8019 , \8033 , \8037 );
and \U$7255 ( \8039 , \7935 , RIaa9e520_237);
and \U$7256 ( \8040 , RIaa9e610_239, \7944 );
nor \U$7257 ( \8041 , \8039 , \8040 );
and \U$7258 ( \8042 , \7942 , RIaa9e1d8_230);
and \U$7259 ( \8043 , RIaa9e250_231, \7919 );
nor \U$7260 ( \8044 , \8042 , \8043 );
and \U$7261 ( \8045 , \7914 , RIaa9df08_224);
and \U$7262 ( \8046 , RIaa9e0e8_228, \7924 );
nor \U$7263 ( \8047 , \8045 , \8046 );
nand \U$7264 ( \8048 , \8038 , \8041 , \8044 , \8047 );
buf \U$7265 ( \8049 , \8048 );
_DC g2896 ( \8050_nG2896 , \8049 , \7973 );
xor \U$7266 ( \8051 , \8018 , \8050_nG2896 );
and \U$7267 ( \8052 , \7886 , RIaaa9038_602);
not \U$7268 ( \8053 , \7886 );
not \U$7269 ( \8054 , RIaaa9038_602);
and \U$7270 ( \8055 , \8053 , \8054 );
nor \U$7271 ( \8056 , \8052 , \8055 );
and \U$7272 ( \8057 , \7959 , RIaa9d878_210);
and \U$7273 ( \8058 , \7928 , RIaa9d698_206);
and \U$7274 ( \8059 , RIaa9d8f0_211, \7909 );
nor \U$7275 ( \8060 , \8058 , \8059 );
and \U$7276 ( \8061 , \7949 , RIaa9da58_214);
nand \U$7277 ( \8062 , RIaa9db48_216, \7955 );
not \U$7278 ( \8063 , \8062 );
nor \U$7279 ( \8064 , \8061 , \8063 );
and \U$7280 ( \8065 , \7930 , RIaa9d710_207);
and \U$7281 ( \8066 , RIaa9de18_222, \7939 );
nor \U$7282 ( \8067 , \8065 , \8066 );
and \U$7283 ( \8068 , \7961 , RIaa9d788_208);
and \U$7284 ( \8069 , RIaa9dc38_218, \7963 );
nor \U$7285 ( \8070 , \8068 , \8069 );
nand \U$7286 ( \8071 , \8060 , \8064 , \8067 , \8070 );
and \U$7287 ( \8072 , \7952 , RIaa9dbc0_217);
and \U$7288 ( \8073 , RIaa9d968_212, \7957 );
nor \U$7289 ( \8074 , \8072 , \8073 );
not \U$7290 ( \8075 , \8074 );
nor \U$7291 ( \8076 , \8057 , \8071 , \8075 );
and \U$7292 ( \8077 , \7935 , RIaa9d9e0_213);
and \U$7293 ( \8078 , RIaa9d800_209, \7944 );
nor \U$7294 ( \8079 , \8077 , \8078 );
and \U$7295 ( \8080 , \7942 , RIaa9dcb0_219);
and \U$7296 ( \8081 , RIaa9dd28_220, \7919 );
nor \U$7297 ( \8082 , \8080 , \8081 );
and \U$7298 ( \8083 , \7914 , RIaa9dad0_215);
and \U$7299 ( \8084 , RIaa9dda0_221, \7924 );
nor \U$7300 ( \8085 , \8083 , \8084 );
nand \U$7301 ( \8086 , \8076 , \8079 , \8082 , \8085 );
buf \U$7302 ( \8087 , \8086 );
_DC g26eb ( \8088_nG26eb , \8087 , \7973 );
xor \U$7303 ( \8089 , \8056 , \8088_nG26eb );
not \U$7304 ( \8090 , \7884 );
not \U$7305 ( \8091 , RIaaa93f8_610);
and \U$7306 ( \8092 , \8090 , \8091 );
and \U$7307 ( \8093 , \7884 , RIaaa93f8_610);
nor \U$7308 ( \8094 , \8092 , \8093 );
and \U$7309 ( \8095 , \7939 , RIaa99048_56);
and \U$7310 ( \8096 , RIaa995e8_68, \7957 );
and \U$7311 ( \8097 , \7959 , RIaa991b0_59);
and \U$7312 ( \8098 , RIaa99570_67, \7935 );
nor \U$7313 ( \8099 , \8096 , \8097 , \8098 );
and \U$7314 ( \8100 , \7914 , RIaa98ee0_53);
and \U$7315 ( \8101 , RIaa99318_62, \7952 );
nor \U$7316 ( \8102 , \8100 , \8101 );
and \U$7317 ( \8103 , \7942 , RIaa99390_63);
and \U$7318 ( \8104 , RIaa994f8_66, \7944 );
nor \U$7319 ( \8105 , \8103 , \8104 );
and \U$7320 ( \8106 , \7919 , RIaa99408_64);
and \U$7321 ( \8107 , RIaa98fd0_55, \7924 );
nor \U$7322 ( \8108 , \8106 , \8107 );
nand \U$7323 ( \8109 , \8099 , \8102 , \8105 , \8108 );
and \U$7324 ( \8110 , \7928 , RIaa99480_65);
and \U$7325 ( \8111 , RIaa990c0_57, \7930 );
nor \U$7326 ( \8112 , \8110 , \8111 );
not \U$7327 ( \8113 , \8112 );
nor \U$7328 ( \8114 , \8095 , \8109 , \8113 );
and \U$7329 ( \8115 , \7961 , RIaa99138_58);
and \U$7330 ( \8116 , RIaa99228_60, \7909 );
nor \U$7331 ( \8117 , \8115 , \8116 );
nand \U$7332 ( \8118 , RIaa98f58_54, \7955 );
and \U$7333 ( \8119 , \7949 , RIaa98e68_52);
and \U$7334 ( \8120 , RIaa992a0_61, \7963 );
nor \U$7335 ( \8121 , \8119 , \8120 );
nand \U$7336 ( \8122 , \8114 , \8117 , \8118 , \8121 );
buf \U$7337 ( \8123 , \8122 );
_DC g26e9 ( \8124_nG26e9 , \8123 , \7973 );
xor \U$7338 ( \8125 , \8094 , \8124_nG26e9 );
and \U$7339 ( \8126 , \7882 , RIaaa9380_609);
not \U$7340 ( \8127 , \7882 );
not \U$7341 ( \8128 , RIaaa9380_609);
and \U$7342 ( \8129 , \8127 , \8128 );
nor \U$7343 ( \8130 , \8126 , \8129 );
and \U$7344 ( \8131 , \7959 , RIaa99750_71);
and \U$7345 ( \8132 , \7928 , RIaa99cf0_83);
and \U$7346 ( \8133 , RIaa997c8_72, \7909 );
nor \U$7347 ( \8134 , \8132 , \8133 );
and \U$7348 ( \8135 , \7949 , RIaa99840_73);
nand \U$7349 ( \8136 , RIaa99930_75, \7955 );
not \U$7350 ( \8137 , \8136 );
nor \U$7351 ( \8138 , \8135 , \8137 );
and \U$7352 ( \8139 , \7930 , RIaa99c78_82);
and \U$7353 ( \8140 , RIaa99a20_77, \7939 );
nor \U$7354 ( \8141 , \8139 , \8140 );
and \U$7355 ( \8142 , \7961 , RIaa99d68_84);
and \U$7356 ( \8143 , RIaa99a98_78, \7963 );
nor \U$7357 ( \8144 , \8142 , \8143 );
nand \U$7358 ( \8145 , \8134 , \8138 , \8141 , \8144 );
and \U$7359 ( \8146 , \7952 , RIaa99b10_79);
and \U$7360 ( \8147 , RIaa996d8_70, \7957 );
nor \U$7361 ( \8148 , \8146 , \8147 );
not \U$7362 ( \8149 , \8148 );
nor \U$7363 ( \8150 , \8131 , \8145 , \8149 );
and \U$7364 ( \8151 , \7935 , RIaa99660_69);
and \U$7365 ( \8152 , RIaa99de0_85, \7944 );
nor \U$7366 ( \8153 , \8151 , \8152 );
and \U$7367 ( \8154 , \7942 , RIaa99b88_80);
and \U$7368 ( \8155 , RIaa99c00_81, \7919 );
nor \U$7369 ( \8156 , \8154 , \8155 );
and \U$7370 ( \8157 , \7914 , RIaa998b8_74);
and \U$7371 ( \8158 , RIaa999a8_76, \7924 );
nor \U$7372 ( \8159 , \8157 , \8158 );
nand \U$7373 ( \8160 , \8150 , \8153 , \8156 , \8159 );
buf \U$7374 ( \8161 , \8160 );
_DC g2358 ( \8162_nG2358 , \8161 , \7973 );
xor \U$7375 ( \8163 , \8130 , \8162_nG2358 );
not \U$7376 ( \8164 , \7880 );
not \U$7377 ( \8165 , RIaaa9308_608);
and \U$7378 ( \8166 , \8164 , \8165 );
and \U$7379 ( \8167 , \7880 , RIaaa9308_608);
nor \U$7380 ( \8168 , \8166 , \8167 );
and \U$7381 ( \8169 , \7939 , RIaa9a038_90);
and \U$7382 ( \8170 , RIaa9a3f8_98, \7957 );
and \U$7383 ( \8171 , \7959 , RIaa9a4e8_100);
and \U$7384 ( \8172 , RIaa9a380_97, \7935 );
nor \U$7385 ( \8173 , \8170 , \8171 , \8172 );
and \U$7386 ( \8174 , \7914 , RIaa99fc0_89);
and \U$7387 ( \8175 , RIaa9a1a0_93, \7952 );
nor \U$7388 ( \8176 , \8174 , \8175 );
and \U$7389 ( \8177 , \7942 , RIaa9a0b0_91);
and \U$7390 ( \8178 , RIaa9a5d8_102, \7944 );
nor \U$7391 ( \8179 , \8177 , \8178 );
and \U$7392 ( \8180 , \7919 , RIaa9a218_94);
and \U$7393 ( \8181 , RIaa99f48_88, \7924 );
nor \U$7394 ( \8182 , \8180 , \8181 );
nand \U$7395 ( \8183 , \8173 , \8176 , \8179 , \8182 );
and \U$7396 ( \8184 , \7928 , RIaa9a470_99);
and \U$7397 ( \8185 , RIaa9a308_96, \7930 );
nor \U$7398 ( \8186 , \8184 , \8185 );
not \U$7399 ( \8187 , \8186 );
nor \U$7400 ( \8188 , \8169 , \8183 , \8187 );
and \U$7401 ( \8189 , \7961 , RIaa9a290_95);
and \U$7402 ( \8190 , RIaa9a560_101, \7909 );
nor \U$7403 ( \8191 , \8189 , \8190 );
nand \U$7404 ( \8192 , RIaa99ed0_87, \7955 );
and \U$7405 ( \8193 , \7949 , RIaa99e58_86);
and \U$7406 ( \8194 , RIaa9a128_92, \7963 );
nor \U$7407 ( \8195 , \8193 , \8194 );
nand \U$7408 ( \8196 , \8188 , \8191 , \8192 , \8195 );
buf \U$7409 ( \8197 , \8196 );
_DC g2356 ( \8198_nG2356 , \8197 , \7973 );
xor \U$7410 ( \8199 , \8168 , \8198_nG2356 );
not \U$7411 ( \8200 , \7878 );
not \U$7412 ( \8201 , RIaaa9290_607);
and \U$7413 ( \8202 , \8200 , \8201 );
and \U$7414 ( \8203 , \7878 , RIaaa9290_607);
nor \U$7415 ( \8204 , \8202 , \8203 );
and \U$7416 ( \8205 , \7939 , RIaa9a830_107);
and \U$7417 ( \8206 , RIaa9aa10_111, \7957 );
and \U$7418 ( \8207 , \7959 , RIaa9ab78_114);
and \U$7419 ( \8208 , RIaa9a998_110, \7935 );
nor \U$7420 ( \8209 , \8206 , \8207 , \8208 );
and \U$7421 ( \8210 , \7914 , RIaa9a6c8_104);
and \U$7422 ( \8211 , RIaa9ac68_116, \7952 );
nor \U$7423 ( \8212 , \8210 , \8211 );
and \U$7424 ( \8213 , \7942 , RIaa9ad58_118);
and \U$7425 ( \8214 , RIaa9abf0_115, \7944 );
nor \U$7426 ( \8215 , \8213 , \8214 );
and \U$7427 ( \8216 , \7919 , RIaa9add0_119);
and \U$7428 ( \8217 , RIaa9a7b8_106, \7924 );
nor \U$7429 ( \8218 , \8216 , \8217 );
nand \U$7430 ( \8219 , \8209 , \8212 , \8215 , \8218 );
nand \U$7431 ( \8220 , RIaa9a740_105, \7955 );
not \U$7432 ( \8221 , \8220 );
nor \U$7433 ( \8222 , \8205 , \8219 , \8221 );
and \U$7434 ( \8223 , \7961 , RIaa9a8a8_108);
and \U$7435 ( \8224 , RIaa9ab00_113, \7909 );
nor \U$7436 ( \8225 , \8223 , \8224 );
and \U$7437 ( \8226 , \7928 , RIaa9aa88_112);
and \U$7438 ( \8227 , RIaa9a920_109, \7930 );
nor \U$7439 ( \8228 , \8226 , \8227 );
and \U$7440 ( \8229 , \7949 , RIaa9a650_103);
and \U$7441 ( \8230 , RIaa9ace0_117, \7963 );
nor \U$7442 ( \8231 , \8229 , \8230 );
nand \U$7443 ( \8232 , \8222 , \8225 , \8228 , \8231 );
buf \U$7444 ( \8233 , \8232 );
_DC g22e8 ( \8234_nG22e8 , \8233 , \7973 );
xor \U$7445 ( \8235 , \8204 , \8234_nG22e8 );
not \U$7446 ( \8236 , \7876 );
not \U$7447 ( \8237 , RIaaa9218_606);
and \U$7448 ( \8238 , \8236 , \8237 );
and \U$7449 ( \8239 , \7876 , RIaaa9218_606);
nor \U$7450 ( \8240 , \8238 , \8239 );
and \U$7451 ( \8241 , \7939 , RIaa9cf90_191);
and \U$7452 ( \8242 , RIaa9d260_197, \7957 );
and \U$7453 ( \8243 , \7959 , RIaa9d3c8_200);
and \U$7454 ( \8244 , RIaa9d1e8_196, \7935 );
nor \U$7455 ( \8245 , \8242 , \8243 , \8244 );
and \U$7456 ( \8246 , \7914 , RIaa9d080_193);
and \U$7457 ( \8247 , RIaa9d530_203, \7952 );
nor \U$7458 ( \8248 , \8246 , \8247 );
and \U$7459 ( \8249 , \7942 , RIaa9d5a8_204);
and \U$7460 ( \8250 , RIaa9d440_201, \7944 );
nor \U$7461 ( \8251 , \8249 , \8250 );
and \U$7462 ( \8252 , \7919 , RIaa9d620_205);
and \U$7463 ( \8253 , RIaa9cf18_190, \7924 );
nor \U$7464 ( \8254 , \8252 , \8253 );
nand \U$7465 ( \8255 , \8245 , \8248 , \8251 , \8254 );
and \U$7466 ( \8256 , \7928 , RIaa9d2d8_198);
and \U$7467 ( \8257 , RIaa9d0f8_194, \7930 );
nor \U$7468 ( \8258 , \8256 , \8257 );
not \U$7469 ( \8259 , \8258 );
nor \U$7470 ( \8260 , \8241 , \8255 , \8259 );
and \U$7471 ( \8261 , \7961 , RIaa9d170_195);
and \U$7472 ( \8262 , RIaa9d350_199, \7909 );
nor \U$7473 ( \8263 , \8261 , \8262 );
nand \U$7474 ( \8264 , RIaa9cea0_189, \7955 );
and \U$7475 ( \8265 , \7949 , RIaa9d008_192);
and \U$7476 ( \8266 , RIaa9d4b8_202, \7963 );
nor \U$7477 ( \8267 , \8265 , \8266 );
nand \U$7478 ( \8268 , \8260 , \8263 , \8264 , \8267 );
buf \U$7479 ( \8269 , \8268 );
_DC g22e6 ( \8270_nG22e6 , \8269 , \7973 );
xor \U$7480 ( \8271 , \8240 , \8270_nG22e6 );
xnor \U$7481 ( \8272 , RIaaa90b0_603, \7875 );
and \U$7482 ( \8273 , \7939 , RIaa9b028_124);
and \U$7483 ( \8274 , RIaa9b4d8_134, \7919 );
and \U$7484 ( \8275 , \7959 , RIaa9b370_131);
and \U$7485 ( \8276 , RIaa9aec0_121, \7914 );
nor \U$7486 ( \8277 , \8274 , \8275 , \8276 );
and \U$7487 ( \8278 , \7952 , RIaa9b5c8_136);
and \U$7488 ( \8279 , RIaa9b208_128, \7957 );
nor \U$7489 ( \8280 , \8278 , \8279 );
and \U$7490 ( \8281 , \7935 , RIaa9b190_127);
and \U$7491 ( \8282 , RIaa9b3e8_132, \7944 );
nor \U$7492 ( \8283 , \8281 , \8282 );
and \U$7493 ( \8284 , \7942 , RIaa9b460_133);
and \U$7494 ( \8285 , RIaa9afb0_123, \7924 );
nor \U$7495 ( \8286 , \8284 , \8285 );
nand \U$7496 ( \8287 , \8277 , \8280 , \8283 , \8286 );
nand \U$7497 ( \8288 , RIaa9af38_122, \7955 );
not \U$7498 ( \8289 , \8288 );
nor \U$7499 ( \8290 , \8273 , \8287 , \8289 );
and \U$7500 ( \8291 , \7961 , RIaa9b0a0_125);
and \U$7501 ( \8292 , RIaa9b2f8_130, \7909 );
nor \U$7502 ( \8293 , \8291 , \8292 );
and \U$7503 ( \8294 , \7928 , RIaa9b280_129);
and \U$7504 ( \8295 , RIaa9b118_126, \7930 );
nor \U$7505 ( \8296 , \8294 , \8295 );
and \U$7506 ( \8297 , \7949 , RIaa9ae48_120);
and \U$7507 ( \8298 , RIaa9b550_135, \7963 );
nor \U$7508 ( \8299 , \8297 , \8298 );
nand \U$7509 ( \8300 , \8290 , \8293 , \8296 , \8299 );
buf \U$7510 ( \8301 , \8300 );
_DC g2290 ( \8302_nG2290 , \8301 , \7973 );
xor \U$7511 ( \8303 , \8272 , \8302_nG2290 );
not \U$7512 ( \8304 , RIaaa91a0_605);
and \U$7513 ( \8305 , RIaaa9128_604, \8304 );
not \U$7514 ( \8306 , RIaaa9128_604);
and \U$7515 ( \8307 , \8306 , RIaaa91a0_605);
nor \U$7516 ( \8308 , \8305 , \8307 );
and \U$7517 ( \8309 , \7939 , RIaa9ba00_145);
and \U$7518 ( \8310 , RIaa9b7a8_140, \7957 );
and \U$7519 ( \8311 , \7959 , RIaa9bb68_148);
and \U$7520 ( \8312 , RIaa9b820_141, \7949 );
nor \U$7521 ( \8313 , \8310 , \8311 , \8312 );
and \U$7522 ( \8314 , \7914 , RIaa9b898_142);
and \U$7523 ( \8315 , RIaa9bcd0_151, \7952 );
nor \U$7524 ( \8316 , \8314 , \8315 );
and \U$7525 ( \8317 , \7942 , RIaa9bd48_152);
and \U$7526 ( \8318 , RIaa9bbe0_149, \7944 );
nor \U$7527 ( \8319 , \8317 , \8318 );
and \U$7528 ( \8320 , \7919 , RIaa9bdc0_153);
and \U$7529 ( \8321 , RIaa9b988_144, \7924 );
nor \U$7530 ( \8322 , \8320 , \8321 );
nand \U$7531 ( \8323 , \8313 , \8316 , \8319 , \8322 );
and \U$7532 ( \8324 , \7928 , RIaa9ba78_146);
and \U$7533 ( \8325 , RIaa9b640_137, \7930 );
nor \U$7534 ( \8326 , \8324 , \8325 );
not \U$7535 ( \8327 , \8326 );
nor \U$7536 ( \8328 , \8309 , \8323 , \8327 );
and \U$7537 ( \8329 , \7961 , RIaa9b6b8_138);
and \U$7538 ( \8330 , RIaa9bc58_150, \7963 );
nor \U$7539 ( \8331 , \8329 , \8330 );
nand \U$7540 ( \8332 , RIaa9b910_143, \7955 );
and \U$7541 ( \8333 , \7935 , RIaa9b730_139);
and \U$7542 ( \8334 , RIaa9baf0_147, \7909 );
nor \U$7543 ( \8335 , \8333 , \8334 );
nand \U$7544 ( \8336 , \8328 , \8331 , \8332 , \8335 );
buf \U$7545 ( \8337 , \8336 );
_DC g2292 ( \8338_nG2292 , \8337 , \7973 );
xor \U$7546 ( \8339 , \8308 , \8338_nG2292 );
and \U$7547 ( \8340 , \7959 , RIaa9c360_165);
and \U$7548 ( \8341 , \7928 , RIaa9be38_154);
and \U$7549 ( \8342 , RIaa9c3d8_166, \7909 );
nor \U$7550 ( \8343 , \8341 , \8342 );
and \U$7551 ( \8344 , \7949 , RIaa9c018_158);
nand \U$7552 ( \8345 , RIaa9c108_160, \7955 );
not \U$7553 ( \8346 , \8345 );
nor \U$7554 ( \8347 , \8344 , \8346 );
and \U$7555 ( \8348 , \7930 , RIaa9c5b8_170);
and \U$7556 ( \8349 , RIaa9c180_161, \7939 );
nor \U$7557 ( \8350 , \8348 , \8349 );
and \U$7558 ( \8351 , \7961 , RIaa9c2e8_164);
and \U$7559 ( \8352 , RIaa9bfa0_157, \7963 );
nor \U$7560 ( \8353 , \8351 , \8352 );
nand \U$7561 ( \8354 , \8343 , \8347 , \8350 , \8353 );
and \U$7562 ( \8355 , \7952 , RIaa9bf28_156);
and \U$7563 ( \8356 , RIaa9c540_169, \7957 );
nor \U$7564 ( \8357 , \8355 , \8356 );
not \U$7565 ( \8358 , \8357 );
nor \U$7566 ( \8359 , \8340 , \8354 , \8358 );
and \U$7567 ( \8360 , \7935 , RIaa9c270_163);
and \U$7568 ( \8361 , RIaa9beb0_155, \7944 );
nor \U$7569 ( \8362 , \8360 , \8361 );
and \U$7570 ( \8363 , \7942 , RIaa9c450_167);
and \U$7571 ( \8364 , RIaa9c4c8_168, \7919 );
nor \U$7572 ( \8365 , \8363 , \8364 );
and \U$7573 ( \8366 , \7914 , RIaa9c090_159);
and \U$7574 ( \8367 , RIaa9c1f8_162, \7924 );
nor \U$7575 ( \8368 , \8366 , \8367 );
nand \U$7576 ( \8369 , \8359 , \8362 , \8365 , \8368 );
buf \U$7577 ( \8370 , \8369 );
_DC g221f ( \8371_nG221f , \8370 , \7973 );
xor \U$7578 ( \8372 , RIaaa91a0_605, \8371_nG221f );
and \U$7579 ( \8373 , \7939 , RIaa9c810_175);
and \U$7580 ( \8374 , RIaa9c900_177, \7957 );
and \U$7581 ( \8375 , \7959 , RIaa9c9f0_179);
and \U$7582 ( \8376 , RIaa9cc48_184, \7935 );
nor \U$7583 ( \8377 , \8374 , \8375 , \8376 );
and \U$7584 ( \8378 , \7914 , RIaa9c798_174);
and \U$7585 ( \8379 , RIaa9cae0_181, \7952 );
nor \U$7586 ( \8380 , \8378 , \8379 );
and \U$7587 ( \8381 , \7942 , RIaa9ca68_180);
and \U$7588 ( \8382 , RIaa9cdb0_187, \7944 );
nor \U$7589 ( \8383 , \8381 , \8382 );
and \U$7590 ( \8384 , \7919 , RIaa9cb58_182);
and \U$7591 ( \8385 , RIaa9c630_171, \7924 );
nor \U$7592 ( \8386 , \8384 , \8385 );
nand \U$7593 ( \8387 , \8377 , \8380 , \8383 , \8386 );
and \U$7594 ( \8388 , \7928 , RIaa9cd38_186);
and \U$7595 ( \8389 , RIaa9c888_176, \7930 );
nor \U$7596 ( \8390 , \8388 , \8389 );
not \U$7597 ( \8391 , \8390 );
nor \U$7598 ( \8392 , \8373 , \8387 , \8391 );
and \U$7599 ( \8393 , \7961 , RIaa9ccc0_185);
and \U$7600 ( \8394 , RIaa9cbd0_183, \7909 );
nor \U$7601 ( \8395 , \8393 , \8394 );
nand \U$7602 ( \8396 , RIaa9c720_173, \7955 );
and \U$7603 ( \8397 , \7949 , RIaa9c6a8_172);
and \U$7604 ( \8398 , RIaa9c978_178, \7963 );
nor \U$7605 ( \8399 , \8397 , \8398 );
nand \U$7606 ( \8400 , \8392 , \8395 , \8396 , \8399 );
buf \U$7607 ( \8401 , \8400 );
_DC g221d ( \8402_nG221d , \8401 , \7973 );
not \U$7608 ( \8403 , RIaaa9560_613);
nand \U$7609 ( \8404 , \8402_nG221d , \8403 );
not \U$7610 ( \8405 , \8404 );
and \U$7611 ( \8406 , \8372 , \8405 );
and \U$7612 ( \8407 , RIaaa91a0_605, \8371_nG221f );
or \U$7613 ( \8408 , \8406 , \8407 );
and \U$7614 ( \8409 , \8339 , \8408 );
and \U$7615 ( \8410 , \8308 , \8338_nG2292 );
or \U$7616 ( \8411 , \8409 , \8410 );
and \U$7617 ( \8412 , \8303 , \8411 );
and \U$7618 ( \8413 , \8272 , \8302_nG2290 );
or \U$7619 ( \8414 , \8412 , \8413 );
and \U$7620 ( \8415 , \8271 , \8414 );
and \U$7621 ( \8416 , \8240 , \8270_nG22e6 );
or \U$7622 ( \8417 , \8415 , \8416 );
and \U$7623 ( \8418 , \8235 , \8417 );
and \U$7624 ( \8419 , \8204 , \8234_nG22e8 );
or \U$7625 ( \8420 , \8418 , \8419 );
and \U$7626 ( \8421 , \8199 , \8420 );
and \U$7627 ( \8422 , \8168 , \8198_nG2356 );
or \U$7628 ( \8423 , \8421 , \8422 );
and \U$7629 ( \8424 , \8163 , \8423 );
and \U$7630 ( \8425 , \8130 , \8162_nG2358 );
or \U$7631 ( \8426 , \8424 , \8425 );
and \U$7632 ( \8427 , \8125 , \8426 );
and \U$7633 ( \8428 , \8094 , \8124_nG26e9 );
or \U$7634 ( \8429 , \8427 , \8428 );
and \U$7635 ( \8430 , \8089 , \8429 );
and \U$7636 ( \8431 , \8056 , \8088_nG26eb );
or \U$7637 ( \8432 , \8430 , \8431 );
and \U$7638 ( \8433 , \8051 , \8432 );
and \U$7639 ( \8434 , \8018 , \8050_nG2896 );
or \U$7640 ( \8435 , \8433 , \8434 );
and \U$7641 ( \8436 , \8013 , \8435 );
and \U$7642 ( \8437 , \7980 , \8012_nG2898 );
or \U$7643 ( \8438 , \8436 , \8437 );
and \U$7644 ( \8439 , \7975 , \8438 );
and \U$7645 ( \8440 , \7897 , \7974_nG2a78 );
or \U$7646 ( \8441 , \8439 , \8440 );
not \U$7647 ( \8442 , \7892 );
nand \U$7648 ( \8443 , \8442 , RIaaa95d8_614);
nor \U$7649 ( \8444 , \8441 , \8443 );
not \U$7650 ( \8445 , \8444 );
and \U$7651 ( \8446 , RIaa9f2b8_266, \7957 );
and \U$7652 ( \8447 , RIaa9f768_276, \7944 );
and \U$7653 ( \8448 , \7924 , RIaa9f600_273);
and \U$7654 ( \8449 , RIaa9f9c0_281, \7930 );
nor \U$7655 ( \8450 , \8448 , \8449 );
and \U$7656 ( \8451 , \7961 , RIaa9f498_270);
and \U$7657 ( \8452 , RIaa9f858_278, \7963 );
nor \U$7658 ( \8453 , \8451 , \8452 );
or \U$7659 ( \8454 , \7955 , \7939 );
and \U$7660 ( \8455 , \8454 , RIaa9f588_272);
and \U$7661 ( \8456 , RIaa9f948_280, \7935 );
nor \U$7662 ( \8457 , \8455 , \8456 );
and \U$7663 ( \8458 , \7928 , RIaa9f8d0_279);
and \U$7664 ( \8459 , RIaa9f7e0_277, \7909 );
nor \U$7665 ( \8460 , \8458 , \8459 );
nand \U$7666 ( \8461 , \8450 , \8453 , \8457 , \8460 );
nor \U$7667 ( \8462 , \8446 , \8447 , \8461 );
and \U$7668 ( \8463 , \7942 , RIaa9f3a8_268);
and \U$7669 ( \8464 , RIaa9f6f0_275, \7959 );
nor \U$7670 ( \8465 , \8463 , \8464 );
and \U$7671 ( \8466 , \7914 , RIaa9f510_271);
and \U$7672 ( \8467 , RIaa9f678_274, \7919 );
nor \U$7673 ( \8468 , \8466 , \8467 );
and \U$7674 ( \8469 , \7949 , RIaa9f330_267);
and \U$7675 ( \8470 , RIaa9f420_269, \7952 );
nor \U$7676 ( \8471 , \8469 , \8470 );
nand \U$7677 ( \8472 , \8462 , \8465 , \8468 , \8471 );
buf \U$7678 ( \8473 , \7972 );
_DC g30a2 ( \8474_nG30a2 , \8472 , \8473 );
not \U$7679 ( \8475 , \8474_nG30a2 );
nor \U$7680 ( \8476 , \8445 , \8475 );
xor \U$7681 ( \8477 , \7897 , \7974_nG2a78 );
xor \U$7682 ( \8478 , \8477 , \8438 );
not \U$7683 ( \8479 , \8478 );
xor \U$7684 ( \8480 , \7980 , \8012_nG2898 );
xor \U$7685 ( \8481 , \8480 , \8435 );
not \U$7686 ( \8482 , \8481 );
and \U$7687 ( \8483 , \8479 , \8482 );
and \U$7688 ( \8484 , \8441 , \8443 );
nor \U$7689 ( \8485 , \8484 , \8444 );
nor \U$7690 ( \8486 , \8483 , \8485 );
not \U$7691 ( \8487 , \8486 );
and \U$7692 ( \8488 , RIaa9eb38_250, \7924 );
and \U$7693 ( \8489 , RIaa9f060_261, \7909 );
and \U$7694 ( \8490 , \7959 , RIaa9eef8_258);
and \U$7695 ( \8491 , RIaa9f0d8_262, \7944 );
nor \U$7696 ( \8492 , \8490 , \8491 );
and \U$7697 ( \8493 , \7914 , RIaa9eac0_249);
and \U$7698 ( \8494 , RIaa9ec28_252, \7957 );
nor \U$7699 ( \8495 , \8493 , \8494 );
and \U$7700 ( \8496 , \7942 , RIaa9ed18_254);
and \U$7701 ( \8497 , RIaa9ee80_257, \7919 );
nor \U$7702 ( \8498 , \8496 , \8497 );
and \U$7703 ( \8499 , \7949 , RIaa9eca0_253);
and \U$7704 ( \8500 , RIaa9ee08_256, \7952 );
nor \U$7705 ( \8501 , \8499 , \8500 );
nand \U$7706 ( \8502 , \8492 , \8495 , \8498 , \8501 );
nor \U$7707 ( \8503 , \8488 , \8489 , \8502 );
and \U$7708 ( \8504 , \7928 , RIaa9f1c8_264);
and \U$7709 ( \8505 , RIaa9ef70_259, \7935 );
nor \U$7710 ( \8506 , \8504 , \8505 );
and \U$7711 ( \8507 , \7961 , RIaa9ed90_255);
and \U$7712 ( \8508 , RIaa9efe8_260, \7930 );
nor \U$7713 ( \8509 , \8507 , \8508 );
and \U$7714 ( \8510 , \8454 , RIaa9ebb0_251);
and \U$7715 ( \8511 , RIaa9f150_263, \7963 );
nor \U$7716 ( \8512 , \8510 , \8511 );
nand \U$7717 ( \8513 , \8503 , \8506 , \8509 , \8512 );
_DC g31b0 ( \8514_nG31b0 , \8513 , \8473 );
or \U$7718 ( \8515 , \8487 , \8514_nG31b0 );
not \U$7719 ( \8516 , \8514_nG31b0 );
and \U$7720 ( \8517 , \8485 , \8478 );
nor \U$7721 ( \8518 , \8485 , \8478 );
xnor \U$7722 ( \8519 , \8481 , \8478 );
not \U$7723 ( \8520 , \8519 );
nor \U$7724 ( \8521 , \8517 , \8518 , \8520 );
nand \U$7725 ( \8522 , \8487 , \8521 );
or \U$7726 ( \8523 , \8516 , \8522 );
or \U$7727 ( \8524 , \8521 , \8487 );
nand \U$7728 ( \8525 , \8515 , \8523 , \8524 );
xnor \U$7729 ( \8526 , \8476 , \8525 );
nand \U$7730 ( \8527 , \8520 , \8487 );
or \U$7731 ( \8528 , \8527 , \8516 );
or \U$7732 ( \8529 , \8475 , \8522 );
or \U$7733 ( \8530 , \8519 , \8516 );
or \U$7734 ( \8531 , \8487 , \8474_nG30a2 );
nand \U$7735 ( \8532 , \8531 , \8524 );
nand \U$7736 ( \8533 , \8530 , \8532 );
nand \U$7737 ( \8534 , \8528 , \8529 , \8533 );
xor \U$7738 ( \8535 , \8018 , \8050_nG2896 );
xor \U$7739 ( \8536 , \8535 , \8432 );
xor \U$7740 ( \8537 , \8056 , \8088_nG26eb );
xor \U$7741 ( \8538 , \8537 , \8429 );
nor \U$7742 ( \8539 , \8536 , \8538 );
or \U$7743 ( \8540 , \8481 , \8539 );
and \U$7744 ( \8541 , \8534 , \8540 );
and \U$7745 ( \8542 , RIaa9fc18_286, \8454 );
and \U$7746 ( \8543 , RIaa9fd80_289, \7930 );
and \U$7747 ( \8544 , \7959 , RIaa9ffd8_294);
and \U$7748 ( \8545 , RIaa9fe70_291, \7944 );
nor \U$7749 ( \8546 , \8544 , \8545 );
and \U$7750 ( \8547 , \7914 , RIaa9fba0_285);
and \U$7751 ( \8548 , RIaaa01b8_298, \7957 );
nor \U$7752 ( \8549 , \8547 , \8548 );
and \U$7753 ( \8550 , \7942 , RIaaa0050_295);
and \U$7754 ( \8551 , RIaa9ff60_293, \7919 );
nor \U$7755 ( \8552 , \8550 , \8551 );
and \U$7756 ( \8553 , \7949 , RIaaa0140_297);
and \U$7757 ( \8554 , RIaa9fdf8_290, \7952 );
nor \U$7758 ( \8555 , \8553 , \8554 );
nand \U$7759 ( \8556 , \8546 , \8549 , \8552 , \8555 );
nor \U$7760 ( \8557 , \8542 , \8543 , \8556 );
and \U$7761 ( \8558 , \7928 , RIaa9fab0_283);
and \U$7762 ( \8559 , RIaa9fee8_292, \7909 );
nor \U$7763 ( \8560 , \8558 , \8559 );
and \U$7764 ( \8561 , \7961 , RIaaa00c8_296);
and \U$7765 ( \8562 , RIaa9fd08_288, \7935 );
nor \U$7766 ( \8563 , \8561 , \8562 );
and \U$7767 ( \8564 , \7963 , RIaa9fa38_282);
and \U$7768 ( \8565 , RIaa9fc90_287, \7924 );
nor \U$7769 ( \8566 , \8564 , \8565 );
nand \U$7770 ( \8567 , \8557 , \8560 , \8563 , \8566 );
_DC g2f9c ( \8568_nG2f9c , \8567 , \8473 );
nand \U$7771 ( \8569 , \8568_nG2f9c , \8444 );
not \U$7772 ( \8570 , \8569 );
nor \U$7773 ( \8571 , \8541 , \8570 );
xor \U$7774 ( \8572 , \8526 , \8571 );
not \U$7775 ( \8573 , \8572 );
not \U$7776 ( \8574 , \8536 );
not \U$7777 ( \8575 , \8481 );
or \U$7778 ( \8576 , \8574 , \8575 );
or \U$7779 ( \8577 , \8481 , \8536 );
nand \U$7780 ( \8578 , \8576 , \8577 );
xor \U$7781 ( \8579 , \8538 , \8536 );
nor \U$7782 ( \8580 , \8578 , \8579 );
not \U$7783 ( \8581 , \8580 );
not \U$7784 ( \8582 , \8540 );
nor \U$7785 ( \8583 , \8581 , \8582 );
not \U$7786 ( \8584 , \8583 );
or \U$7787 ( \8585 , \8584 , \8516 );
or \U$7788 ( \8586 , \8581 , \8516 );
nand \U$7789 ( \8587 , \8586 , \8582 );
nand \U$7790 ( \8588 , \8585 , \8587 );
or \U$7791 ( \8589 , \8527 , \8475 );
not \U$7792 ( \8590 , \8568_nG2f9c );
or \U$7793 ( \8591 , \8590 , \8522 );
or \U$7794 ( \8592 , \8519 , \8475 );
or \U$7795 ( \8593 , \8487 , \8568_nG2f9c );
nand \U$7796 ( \8594 , \8593 , \8524 );
nand \U$7797 ( \8595 , \8592 , \8594 );
nand \U$7798 ( \8596 , \8589 , \8591 , \8595 );
and \U$7799 ( \8597 , \8588 , \8596 );
not \U$7800 ( \8598 , \8569 );
and \U$7801 ( \8599 , \8534 , \8540 );
not \U$7802 ( \8600 , \8534 );
and \U$7803 ( \8601 , \8600 , \8582 );
nor \U$7804 ( \8602 , \8599 , \8601 );
not \U$7805 ( \8603 , \8602 );
or \U$7806 ( \8604 , \8598 , \8603 );
or \U$7807 ( \8605 , \8602 , \8569 );
nand \U$7808 ( \8606 , \8604 , \8605 );
and \U$7809 ( \8607 , \8597 , \8606 );
xor \U$7810 ( \8608 , \8573 , \8607 );
or \U$7811 ( \8609 , \8584 , \8475 );
and \U$7812 ( \8610 , \8540 , \8579 );
not \U$7813 ( \8611 , \8610 );
or \U$7814 ( \8612 , \8516 , \8611 );
or \U$7815 ( \8613 , \8581 , \8475 );
or \U$7816 ( \8614 , \8540 , \8514_nG31b0 );
or \U$7817 ( \8615 , \8540 , \8579 );
nand \U$7818 ( \8616 , \8614 , \8615 );
nand \U$7819 ( \8617 , \8613 , \8616 );
nand \U$7820 ( \8618 , \8609 , \8612 , \8617 );
xor \U$7821 ( \8619 , \8094 , \8124_nG26e9 );
xor \U$7822 ( \8620 , \8619 , \8426 );
xor \U$7823 ( \8621 , \8130 , \8162_nG2358 );
xor \U$7824 ( \8622 , \8621 , \8423 );
nor \U$7825 ( \8623 , \8620 , \8622 );
or \U$7826 ( \8624 , \8538 , \8623 );
and \U$7827 ( \8625 , \8618 , \8624 );
not \U$7828 ( \8626 , \8618 );
not \U$7829 ( \8627 , \8624 );
and \U$7830 ( \8628 , \8626 , \8627 );
not \U$7831 ( \8629 , \8527 );
and \U$7832 ( \8630 , \8568_nG2f9c , \8629 );
and \U$7833 ( \8631 , RIaaa06e0_309, \7957 );
and \U$7834 ( \8632 , RIaaa0230_299, \7944 );
and \U$7835 ( \8633 , \7924 , RIaaa0848_312);
and \U$7836 ( \8634 , RIaaa0398_302, \7930 );
nor \U$7837 ( \8635 , \8633 , \8634 );
and \U$7838 ( \8636 , \7961 , RIaaa0500_305);
and \U$7839 ( \8637 , RIaaa0938_314, \7963 );
nor \U$7840 ( \8638 , \8636 , \8637 );
and \U$7841 ( \8639 , \8454 , RIaaa07d0_311);
and \U$7842 ( \8640 , RIaaa0320_301, \7935 );
nor \U$7843 ( \8641 , \8639 , \8640 );
and \U$7844 ( \8642 , \7928 , RIaaa08c0_313);
and \U$7845 ( \8643 , RIaaa02a8_300, \7909 );
nor \U$7846 ( \8644 , \8642 , \8643 );
nand \U$7847 ( \8645 , \8635 , \8638 , \8641 , \8644 );
nor \U$7848 ( \8646 , \8631 , \8632 , \8645 );
and \U$7849 ( \8647 , \7942 , RIaaa0488_304);
and \U$7850 ( \8648 , RIaaa05f0_307, \7959 );
nor \U$7851 ( \8649 , \8647 , \8648 );
and \U$7852 ( \8650 , \7914 , RIaaa0758_310);
and \U$7853 ( \8651 , RIaaa0578_306, \7919 );
nor \U$7854 ( \8652 , \8650 , \8651 );
and \U$7855 ( \8653 , \7949 , RIaaa0668_308);
and \U$7856 ( \8654 , RIaaa0410_303, \7952 );
nor \U$7857 ( \8655 , \8653 , \8654 );
nand \U$7858 ( \8656 , \8646 , \8649 , \8652 , \8655 );
_DC g2e7a ( \8657_nG2e7a , \8656 , \8473 );
or \U$7859 ( \8658 , \8487 , \8657_nG2e7a );
nand \U$7860 ( \8659 , \8658 , \8524 );
nand \U$7861 ( \8660 , \8568_nG2f9c , \8520 );
and \U$7862 ( \8661 , \8659 , \8660 );
not \U$7863 ( \8662 , \8522 );
and \U$7864 ( \8663 , \8657_nG2e7a , \8662 );
nor \U$7865 ( \8664 , \8630 , \8661 , \8663 );
nor \U$7866 ( \8665 , \8628 , \8664 );
nor \U$7867 ( \8666 , \8625 , \8665 );
xor \U$7868 ( \8667 , \8588 , \8596 );
not \U$7869 ( \8668 , \8667 );
nand \U$7870 ( \8669 , \8657_nG2e7a , \8444 );
not \U$7871 ( \8670 , \8669 );
and \U$7872 ( \8671 , \8668 , \8670 );
and \U$7873 ( \8672 , \8667 , \8669 );
nor \U$7874 ( \8673 , \8671 , \8672 );
nand \U$7875 ( \8674 , \8666 , \8673 );
xor \U$7876 ( \8675 , \8597 , \8606 );
and \U$7877 ( \8676 , \8674 , \8675 );
and \U$7878 ( \8677 , \8608 , \8676 );
not \U$7879 ( \8678 , \8677 );
and \U$7880 ( \8679 , \8573 , \8607 );
or \U$7881 ( \8680 , \8679 , \8486 );
and \U$7882 ( \8681 , \8679 , \8486 );
and \U$7883 ( \8682 , \8476 , \8525 );
nor \U$7884 ( \8683 , \8681 , \8682 );
nand \U$7885 ( \8684 , \8680 , \8683 );
not \U$7886 ( \8685 , \8684 );
and \U$7887 ( \8686 , \8444 , \8514_nG31b0 );
and \U$7888 ( \8687 , \8526 , \8571 );
nor \U$7889 ( \8688 , \8686 , \8687 );
not \U$7890 ( \8689 , \8688 );
and \U$7891 ( \8690 , \8685 , \8689 );
and \U$7892 ( \8691 , \8684 , \8688 );
nor \U$7893 ( \8692 , \8690 , \8691 );
not \U$7894 ( \8693 , \8692 );
or \U$7895 ( \8694 , \8678 , \8693 );
or \U$7896 ( \8695 , \8692 , \8677 );
nand \U$7897 ( \8696 , \8694 , \8695 );
not \U$7898 ( \8697 , \8696 );
xor \U$7899 ( \8698 , \8674 , \8675 );
not \U$7900 ( \8699 , \8667 );
nor \U$7901 ( \8700 , \8699 , \8669 );
xor \U$7902 ( \8701 , \8698 , \8700 );
and \U$7903 ( \8702 , \8657_nG2e7a , \8629 );
and \U$7904 ( \8703 , RIaaa10b8_330, \7928 );
and \U$7905 ( \8704 , RIaaa0e60_325, \7930 );
and \U$7906 ( \8705 , \7959 , RIaaa0b90_319);
and \U$7907 ( \8706 , RIaaa0cf8_322, \7944 );
nor \U$7908 ( \8707 , \8705 , \8706 );
and \U$7909 ( \8708 , \7914 , RIaaa0f50_327);
and \U$7910 ( \8709 , RIaaa0c80_321, \7957 );
nor \U$7911 ( \8710 , \8708 , \8709 );
and \U$7912 ( \8711 , \7942 , RIaaa0a28_316);
and \U$7913 ( \8712 , RIaaa0b18_318, \7919 );
nor \U$7914 ( \8713 , \8711 , \8712 );
and \U$7915 ( \8714 , \7949 , RIaaa0c08_320);
and \U$7916 ( \8715 , RIaaa0ed8_326, \7952 );
nor \U$7917 ( \8716 , \8714 , \8715 );
nand \U$7918 ( \8717 , \8707 , \8710 , \8713 , \8716 );
nor \U$7919 ( \8718 , \8703 , \8704 , \8717 );
and \U$7920 ( \8719 , \7961 , RIaaa0aa0_317);
and \U$7921 ( \8720 , RIaaa0d70_323, \7909 );
nor \U$7922 ( \8721 , \8719 , \8720 );
and \U$7923 ( \8722 , \8454 , RIaaa0fc8_328);
and \U$7924 ( \8723 , RIaaa1130_331, \7963 );
nor \U$7925 ( \8724 , \8722 , \8723 );
and \U$7926 ( \8725 , \7935 , RIaaa0de8_324);
and \U$7927 ( \8726 , RIaaa1040_329, \7924 );
nor \U$7928 ( \8727 , \8725 , \8726 );
nand \U$7929 ( \8728 , \8718 , \8721 , \8724 , \8727 );
_DC g2d90 ( \8729_nG2d90 , \8728 , \8473 );
or \U$7930 ( \8730 , \8487 , \8729_nG2d90 );
nand \U$7931 ( \8731 , \8730 , \8524 );
nand \U$7932 ( \8732 , \8657_nG2e7a , \8520 );
and \U$7933 ( \8733 , \8731 , \8732 );
and \U$7934 ( \8734 , \8729_nG2d90 , \8662 );
nor \U$7935 ( \8735 , \8702 , \8733 , \8734 );
and \U$7936 ( \8736 , RIaaa2198_366, \7928 );
and \U$7937 ( \8737 , RIaaa1fb8_362, \7930 );
and \U$7938 ( \8738 , \7952 , RIaaa1d60_357);
and \U$7939 ( \8739 , RIaaa1bf8_354, \7957 );
nor \U$7940 ( \8740 , \8738 , \8739 );
and \U$7941 ( \8741 , \7942 , RIaaa1ce8_356);
and \U$7942 ( \8742 , RIaaa1e50_359, \7919 );
nor \U$7943 ( \8743 , \8741 , \8742 );
and \U$7944 ( \8744 , \7914 , RIaaa1a90_351);
and \U$7945 ( \8745 , RIaaa1c70_355, \7949 );
nor \U$7946 ( \8746 , \8744 , \8745 );
and \U$7947 ( \8747 , \7959 , RIaaa1ec8_360);
and \U$7948 ( \8748 , RIaaa2030_363, \7944 );
nor \U$7949 ( \8749 , \8747 , \8748 );
nand \U$7950 ( \8750 , \8740 , \8743 , \8746 , \8749 );
nor \U$7951 ( \8751 , \8736 , \8737 , \8750 );
and \U$7952 ( \8752 , \7961 , RIaaa1dd8_358);
and \U$7953 ( \8753 , RIaaa20a8_364, \7909 );
nor \U$7954 ( \8754 , \8752 , \8753 );
and \U$7955 ( \8755 , \8454 , RIaaa1b08_352);
and \U$7956 ( \8756 , RIaaa2120_365, \7963 );
nor \U$7957 ( \8757 , \8755 , \8756 );
and \U$7958 ( \8758 , \7935 , RIaaa1f40_361);
and \U$7959 ( \8759 , RIaaa1b80_353, \7924 );
nor \U$7960 ( \8760 , \8758 , \8759 );
nand \U$7961 ( \8761 , \8751 , \8754 , \8757 , \8760 );
_DC g2c8f ( \8762_nG2c8f , \8761 , \8473 );
nand \U$7962 ( \8763 , \8762_nG2c8f , \8444 );
or \U$7963 ( \8764 , \8735 , \8763 );
and \U$7964 ( \8765 , \8538 , \8620 );
nor \U$7965 ( \8766 , \8538 , \8620 );
xor \U$7966 ( \8767 , \8620 , \8622 );
nor \U$7967 ( \8768 , \8765 , \8766 , \8767 );
and \U$7968 ( \8769 , \8768 , \8624 );
and \U$7969 ( \8770 , \8514_nG31b0 , \8769 );
not \U$7970 ( \8771 , \8624 );
and \U$7971 ( \8772 , \8516 , \8771 );
or \U$7972 ( \8773 , \8768 , \8624 );
not \U$7973 ( \8774 , \8773 );
nor \U$7974 ( \8775 , \8770 , \8772 , \8774 );
nand \U$7975 ( \8776 , \8568_nG2f9c , \8580 );
or \U$7976 ( \8777 , \8540 , \8474_nG30a2 );
nand \U$7977 ( \8778 , \8777 , \8615 );
and \U$7978 ( \8779 , \8776 , \8778 );
and \U$7979 ( \8780 , \8610 , \8474_nG30a2 );
and \U$7980 ( \8781 , \8568_nG2f9c , \8583 );
nor \U$7981 ( \8782 , \8779 , \8780 , \8781 );
or \U$7982 ( \8783 , \8775 , \8782 );
nand \U$7983 ( \8784 , \8764 , \8783 );
not \U$7984 ( \8785 , \8729_nG2d90 );
nor \U$7985 ( \8786 , \8445 , \8785 );
and \U$7986 ( \8787 , \8618 , \8624 );
not \U$7987 ( \8788 , \8618 );
and \U$7988 ( \8789 , \8788 , \8771 );
nor \U$7989 ( \8790 , \8787 , \8789 );
not \U$7990 ( \8791 , \8790 );
not \U$7991 ( \8792 , \8664 );
or \U$7992 ( \8793 , \8791 , \8792 );
or \U$7993 ( \8794 , \8664 , \8790 );
nand \U$7994 ( \8795 , \8793 , \8794 );
xor \U$7995 ( \8796 , \8786 , \8795 );
and \U$7996 ( \8797 , \8784 , \8796 );
or \U$7997 ( \8798 , \8673 , \8666 );
nand \U$7998 ( \8799 , \8798 , \8674 );
and \U$7999 ( \8800 , \8797 , \8799 );
and \U$8000 ( \8801 , \8701 , \8800 );
and \U$8001 ( \8802 , \8698 , \8700 );
or \U$8002 ( \8803 , \8801 , \8802 );
xor \U$8003 ( \8804 , \8608 , \8676 );
xor \U$8004 ( \8805 , \8803 , \8804 );
xor \U$8005 ( \8806 , \8698 , \8700 );
xor \U$8006 ( \8807 , \8806 , \8800 );
xor \U$8007 ( \8808 , \8797 , \8799 );
and \U$8008 ( \8809 , \8786 , \8795 );
xor \U$8009 ( \8810 , \8808 , \8809 );
xor \U$8010 ( \8811 , \8168 , \8198_nG2356 );
xor \U$8011 ( \8812 , \8811 , \8420 );
xor \U$8012 ( \8813 , \8204 , \8234_nG22e8 );
xor \U$8013 ( \8814 , \8813 , \8417 );
nor \U$8014 ( \8815 , \8812 , \8814 );
or \U$8015 ( \8816 , \8622 , \8815 );
not \U$8016 ( \8817 , \8816 );
nand \U$8017 ( \8818 , \8657_nG2e7a , \8580 );
or \U$8018 ( \8819 , \8540 , \8568_nG2f9c );
nand \U$8019 ( \8820 , \8819 , \8615 );
and \U$8020 ( \8821 , \8818 , \8820 );
and \U$8021 ( \8822 , \8610 , \8568_nG2f9c );
and \U$8022 ( \8823 , \8657_nG2e7a , \8583 );
nor \U$8023 ( \8824 , \8821 , \8822 , \8823 );
nand \U$8024 ( \8825 , \8514_nG31b0 , \8767 );
or \U$8025 ( \8826 , \8624 , \8474_nG30a2 );
nand \U$8026 ( \8827 , \8826 , \8773 );
and \U$8027 ( \8828 , \8825 , \8827 );
and \U$8028 ( \8829 , \8769 , \8474_nG30a2 );
not \U$8029 ( \8830 , \8767 );
nor \U$8030 ( \8831 , \8771 , \8830 );
and \U$8031 ( \8832 , \8514_nG31b0 , \8831 );
nor \U$8032 ( \8833 , \8828 , \8829 , \8832 );
nor \U$8033 ( \8834 , \8824 , \8833 );
not \U$8034 ( \8835 , \8834 );
nand \U$8035 ( \8836 , \8833 , \8824 );
nand \U$8036 ( \8837 , \8835 , \8836 );
not \U$8037 ( \8838 , \8837 );
or \U$8038 ( \8839 , \8817 , \8838 );
or \U$8039 ( \8840 , \8837 , \8816 );
nand \U$8040 ( \8841 , \8839 , \8840 );
and \U$8041 ( \8842 , RIaaa1310_335, \8454 );
and \U$8042 ( \8843 , RIaaa17c0_345, \7930 );
and \U$8043 ( \8844 , \7959 , RIaaa16d0_343);
and \U$8044 ( \8845 , RIaaa1838_346, \7944 );
nor \U$8045 ( \8846 , \8844 , \8845 );
and \U$8046 ( \8847 , \7914 , RIaaa1298_334);
and \U$8047 ( \8848 , RIaaa1400_337, \7957 );
nor \U$8048 ( \8849 , \8847 , \8848 );
and \U$8049 ( \8850 , \7942 , RIaaa14f0_339);
and \U$8050 ( \8851 , RIaaa1658_342, \7919 );
nor \U$8051 ( \8852 , \8850 , \8851 );
and \U$8052 ( \8853 , \7949 , RIaaa1478_338);
and \U$8053 ( \8854 , RIaaa1568_340, \7952 );
nor \U$8054 ( \8855 , \8853 , \8854 );
nand \U$8055 ( \8856 , \8846 , \8849 , \8852 , \8855 );
nor \U$8056 ( \8857 , \8842 , \8843 , \8856 );
and \U$8057 ( \8858 , \7928 , RIaaa19a0_349);
and \U$8058 ( \8859 , RIaaa1928_348, \7963 );
nor \U$8059 ( \8860 , \8858 , \8859 );
and \U$8060 ( \8861 , \7961 , RIaaa15e0_341);
and \U$8061 ( \8862 , RIaaa1748_344, \7935 );
nor \U$8062 ( \8863 , \8861 , \8862 );
and \U$8063 ( \8864 , \7924 , RIaaa1388_336);
and \U$8064 ( \8865 , RIaaa18b0_347, \7909 );
nor \U$8065 ( \8866 , \8864 , \8865 );
nand \U$8066 ( \8867 , \8857 , \8860 , \8863 , \8866 );
_DC g2b9c ( \8868_nG2b9c , \8867 , \8473 );
not \U$8067 ( \8869 , \8868_nG2b9c );
nor \U$8068 ( \8870 , \8445 , \8869 );
or \U$8069 ( \8871 , \8527 , \8785 );
not \U$8070 ( \8872 , \8762_nG2c8f );
or \U$8071 ( \8873 , \8872 , \8522 );
or \U$8072 ( \8874 , \8519 , \8785 );
or \U$8073 ( \8875 , \8487 , \8762_nG2c8f );
nand \U$8074 ( \8876 , \8875 , \8524 );
nand \U$8075 ( \8877 , \8874 , \8876 );
nand \U$8076 ( \8878 , \8871 , \8873 , \8877 );
xor \U$8077 ( \8879 , \8870 , \8878 );
and \U$8078 ( \8880 , \8841 , \8879 );
not \U$8079 ( \8881 , \8812 );
not \U$8080 ( \8882 , \8622 );
or \U$8081 ( \8883 , \8881 , \8882 );
or \U$8082 ( \8884 , \8622 , \8812 );
nand \U$8083 ( \8885 , \8883 , \8884 );
xor \U$8084 ( \8886 , \8814 , \8812 );
nor \U$8085 ( \8887 , \8885 , \8886 );
not \U$8086 ( \8888 , \8887 );
not \U$8087 ( \8889 , \8816 );
nor \U$8088 ( \8890 , \8888 , \8889 );
not \U$8089 ( \8891 , \8890 );
or \U$8090 ( \8892 , \8891 , \8516 );
or \U$8091 ( \8893 , \8888 , \8516 );
nand \U$8092 ( \8894 , \8893 , \8889 );
nand \U$8093 ( \8895 , \8892 , \8894 );
not \U$8094 ( \8896 , \8831 );
or \U$8095 ( \8897 , \8896 , \8475 );
not \U$8096 ( \8898 , \8769 );
or \U$8097 ( \8899 , \8590 , \8898 );
or \U$8098 ( \8900 , \8830 , \8475 );
or \U$8099 ( \8901 , \8624 , \8568_nG2f9c );
nand \U$8100 ( \8902 , \8901 , \8773 );
nand \U$8101 ( \8903 , \8900 , \8902 );
nand \U$8102 ( \8904 , \8897 , \8899 , \8903 );
and \U$8103 ( \8905 , \8895 , \8904 );
and \U$8104 ( \8906 , \8762_nG2c8f , \8629 );
or \U$8105 ( \8907 , \8487 , \8868_nG2b9c );
nand \U$8106 ( \8908 , \8907 , \8524 );
nand \U$8107 ( \8909 , \8762_nG2c8f , \8520 );
and \U$8108 ( \8910 , \8908 , \8909 );
and \U$8109 ( \8911 , \8868_nG2b9c , \8662 );
nor \U$8110 ( \8912 , \8906 , \8910 , \8911 );
nand \U$8111 ( \8913 , \8729_nG2d90 , \8580 );
or \U$8112 ( \8914 , \8540 , \8657_nG2e7a );
nand \U$8113 ( \8915 , \8914 , \8615 );
and \U$8114 ( \8916 , \8913 , \8915 );
and \U$8115 ( \8917 , \8610 , \8657_nG2e7a );
and \U$8116 ( \8918 , \8729_nG2d90 , \8583 );
nor \U$8117 ( \8919 , \8916 , \8917 , \8918 );
and \U$8118 ( \8920 , \8912 , \8919 );
and \U$8119 ( \8921 , RIaaa2be8_388, \7957 );
and \U$8120 ( \8922 , RIaaa2a80_385, \7919 );
and \U$8121 ( \8923 , \7924 , RIaaa3098_398);
and \U$8122 ( \8924 , RIaaa2dc8_392, \7930 );
nor \U$8123 ( \8925 , \8923 , \8924 );
and \U$8124 ( \8926 , \7961 , RIaaa2af8_386);
and \U$8125 ( \8927 , RIaaa2fa8_396, \7963 );
nor \U$8126 ( \8928 , \8926 , \8927 );
and \U$8127 ( \8929 , \8454 , RIaaa3110_399);
and \U$8128 ( \8930 , RIaaa2e40_393, \7935 );
nor \U$8129 ( \8931 , \8929 , \8930 );
and \U$8130 ( \8932 , \7928 , RIaaa2f30_395);
and \U$8131 ( \8933 , RIaaa2cd8_390, \7909 );
nor \U$8132 ( \8934 , \8932 , \8933 );
nand \U$8133 ( \8935 , \8925 , \8928 , \8931 , \8934 );
nor \U$8134 ( \8936 , \8921 , \8922 , \8935 );
and \U$8135 ( \8937 , \7949 , RIaaa2c60_389);
and \U$8136 ( \8938 , RIaaa2eb8_394, \7952 );
nor \U$8137 ( \8939 , \8937 , \8938 );
and \U$8138 ( \8940 , \7914 , RIaaa3020_397);
and \U$8139 ( \8941 , RIaaa2b70_387, \7942 );
nor \U$8140 ( \8942 , \8940 , \8941 );
and \U$8141 ( \8943 , \7959 , RIaaa2a08_384);
and \U$8142 ( \8944 , RIaaa2d50_391, \7944 );
nor \U$8143 ( \8945 , \8943 , \8944 );
nand \U$8144 ( \8946 , \8936 , \8939 , \8942 , \8945 );
_DC g2a93 ( \8947_nG2a93 , \8946 , \8473 );
nand \U$8145 ( \8948 , \8947_nG2a93 , \8444 );
or \U$8146 ( \8949 , \8920 , \8948 );
or \U$8147 ( \8950 , \8912 , \8919 );
nand \U$8148 ( \8951 , \8949 , \8950 );
and \U$8149 ( \8952 , \8905 , \8951 );
and \U$8150 ( \8953 , \8880 , \8952 );
and \U$8151 ( \8954 , \8836 , \8816 );
and \U$8152 ( \8955 , \8870 , \8878 );
nor \U$8153 ( \8956 , \8954 , \8955 , \8834 );
xnor \U$8154 ( \8957 , \8763 , \8735 );
not \U$8155 ( \8958 , \8957 );
xor \U$8156 ( \8959 , \8775 , \8782 );
not \U$8157 ( \8960 , \8959 );
and \U$8158 ( \8961 , \8958 , \8960 );
and \U$8159 ( \8962 , \8957 , \8959 );
nor \U$8160 ( \8963 , \8961 , \8962 );
nand \U$8161 ( \8964 , \8956 , \8963 );
xor \U$8162 ( \8965 , \8953 , \8964 );
xor \U$8163 ( \8966 , \8784 , \8796 );
and \U$8164 ( \8967 , \8965 , \8966 );
and \U$8165 ( \8968 , \8953 , \8964 );
or \U$8166 ( \8969 , \8967 , \8968 );
and \U$8167 ( \8970 , \8810 , \8969 );
and \U$8168 ( \8971 , \8808 , \8809 );
or \U$8169 ( \8972 , \8970 , \8971 );
xor \U$8170 ( \8973 , \8807 , \8972 );
xor \U$8171 ( \8974 , \8808 , \8809 );
xor \U$8172 ( \8975 , \8974 , \8969 );
and \U$8173 ( \8976 , \8868_nG2b9c , \8629 );
or \U$8174 ( \8977 , \8487 , \8947_nG2a93 );
nand \U$8175 ( \8978 , \8977 , \8524 );
nand \U$8176 ( \8979 , \8868_nG2b9c , \8520 );
and \U$8177 ( \8980 , \8978 , \8979 );
and \U$8178 ( \8981 , \8947_nG2a93 , \8662 );
nor \U$8179 ( \8982 , \8976 , \8980 , \8981 );
nand \U$8180 ( \8983 , \8762_nG2c8f , \8580 );
or \U$8181 ( \8984 , \8540 , \8729_nG2d90 );
nand \U$8182 ( \8985 , \8984 , \8615 );
and \U$8183 ( \8986 , \8983 , \8985 );
and \U$8184 ( \8987 , \8610 , \8729_nG2d90 );
and \U$8185 ( \8988 , \8762_nG2c8f , \8583 );
nor \U$8186 ( \8989 , \8986 , \8987 , \8988 );
and \U$8187 ( \8990 , \8982 , \8989 );
not \U$8188 ( \8991 , \8990 );
and \U$8189 ( \8992 , RIaaa26c0_377, \7957 );
and \U$8190 ( \8993 , RIaaa2300_369, \7944 );
and \U$8191 ( \8994 , \7924 , RIaaa2918_382);
and \U$8192 ( \8995 , RIaaa2210_367, \7930 );
nor \U$8193 ( \8996 , \8994 , \8995 );
and \U$8194 ( \8997 , \7961 , RIaaa25d0_375);
and \U$8195 ( \8998 , RIaaa2738_378, \7963 );
nor \U$8196 ( \8999 , \8997 , \8998 );
and \U$8197 ( \9000 , \8454 , RIaaa28a0_381);
and \U$8198 ( \9001 , RIaaa2288_368, \7935 );
nor \U$8199 ( \9002 , \9000 , \9001 );
and \U$8200 ( \9003 , \7928 , RIaaa27b0_379);
and \U$8201 ( \9004 , RIaaa2378_370, \7909 );
nor \U$8202 ( \9005 , \9003 , \9004 );
nand \U$8203 ( \9006 , \8996 , \8999 , \9002 , \9005 );
nor \U$8204 ( \9007 , \8992 , \8993 , \9006 );
and \U$8205 ( \9008 , \7942 , RIaaa2558_374);
and \U$8206 ( \9009 , RIaaa24e0_373, \7959 );
nor \U$8207 ( \9010 , \9008 , \9009 );
and \U$8208 ( \9011 , \7914 , RIaaa2828_380);
and \U$8209 ( \9012 , RIaaa2468_372, \7919 );
nor \U$8210 ( \9013 , \9011 , \9012 );
and \U$8211 ( \9014 , \7949 , RIaaa2648_376);
and \U$8212 ( \9015 , RIaaa23f0_371, \7952 );
nor \U$8213 ( \9016 , \9014 , \9015 );
nand \U$8214 ( \9017 , \9007 , \9010 , \9013 , \9016 );
_DC g29b3 ( \9018_nG29b3 , \9017 , \8473 );
nand \U$8215 ( \9019 , \9018_nG29b3 , \8444 );
not \U$8216 ( \9020 , \9019 );
and \U$8217 ( \9021 , \8991 , \9020 );
nor \U$8218 ( \9022 , \8982 , \8989 );
nor \U$8219 ( \9023 , \9021 , \9022 );
and \U$8220 ( \9024 , \8474_nG30a2 , \8890 );
or \U$8221 ( \9025 , \8816 , \8514_nG31b0 );
or \U$8222 ( \9026 , \8816 , \8886 );
nand \U$8223 ( \9027 , \9025 , \9026 );
nand \U$8224 ( \9028 , \8474_nG30a2 , \8887 );
and \U$8225 ( \9029 , \9027 , \9028 );
and \U$8226 ( \9030 , \8816 , \8886 );
and \U$8227 ( \9031 , \8514_nG31b0 , \9030 );
nor \U$8228 ( \9032 , \9024 , \9029 , \9031 );
nand \U$8229 ( \9033 , \8568_nG2f9c , \8767 );
or \U$8230 ( \9034 , \8624 , \8657_nG2e7a );
nand \U$8231 ( \9035 , \9034 , \8773 );
and \U$8232 ( \9036 , \9033 , \9035 );
and \U$8233 ( \9037 , \8769 , \8657_nG2e7a );
and \U$8234 ( \9038 , \8568_nG2f9c , \8831 );
nor \U$8235 ( \9039 , \9036 , \9037 , \9038 );
nand \U$8236 ( \9040 , \9032 , \9039 );
xor \U$8237 ( \9041 , \8272 , \8302_nG2290 );
xor \U$8238 ( \9042 , \9041 , \8411 );
not \U$8239 ( \9043 , \9042 );
xor \U$8240 ( \9044 , \8240 , \8270_nG22e6 );
xor \U$8241 ( \9045 , \9044 , \8414 );
not \U$8242 ( \9046 , \9045 );
and \U$8243 ( \9047 , \9043 , \9046 );
or \U$8244 ( \9048 , \8814 , \9047 );
and \U$8245 ( \9049 , \9040 , \9048 );
nor \U$8246 ( \9050 , \9039 , \9032 );
nor \U$8247 ( \9051 , \9049 , \9050 );
nor \U$8248 ( \9052 , \9023 , \9051 );
xor \U$8249 ( \9053 , \8895 , \8904 );
not \U$8250 ( \9054 , \9053 );
not \U$8251 ( \9055 , \8950 );
nor \U$8252 ( \9056 , \9055 , \8920 );
not \U$8253 ( \9057 , \9056 );
not \U$8254 ( \9058 , \8948 );
and \U$8255 ( \9059 , \9057 , \9058 );
and \U$8256 ( \9060 , \9056 , \8948 );
nor \U$8257 ( \9061 , \9059 , \9060 );
nor \U$8258 ( \9062 , \9054 , \9061 );
and \U$8259 ( \9063 , \9052 , \9062 );
xor \U$8260 ( \9064 , \8841 , \8879 );
xor \U$8261 ( \9065 , \8905 , \8951 );
and \U$8262 ( \9066 , \9064 , \9065 );
xor \U$8263 ( \9067 , \9063 , \9066 );
or \U$8264 ( \9068 , \8963 , \8956 );
nand \U$8265 ( \9069 , \9068 , \8964 );
and \U$8266 ( \9070 , \9067 , \9069 );
and \U$8267 ( \9071 , \9063 , \9066 );
or \U$8268 ( \9072 , \9070 , \9071 );
not \U$8269 ( \9073 , \8959 );
nor \U$8270 ( \9074 , \9073 , \8957 );
xor \U$8271 ( \9075 , \9072 , \9074 );
xor \U$8272 ( \9076 , \8953 , \8964 );
xor \U$8273 ( \9077 , \9076 , \8966 );
and \U$8274 ( \9078 , \9075 , \9077 );
and \U$8275 ( \9079 , \9072 , \9074 );
or \U$8276 ( \9080 , \9078 , \9079 );
xor \U$8277 ( \9081 , \8975 , \9080 );
xor \U$8278 ( \9082 , \9072 , \9074 );
xor \U$8279 ( \9083 , \9082 , \9077 );
xor \U$8280 ( \9084 , \9064 , \9065 );
not \U$8281 ( \9085 , \9045 );
not \U$8282 ( \9086 , \8814 );
or \U$8283 ( \9087 , \9085 , \9086 );
or \U$8284 ( \9088 , \8814 , \9045 );
nand \U$8285 ( \9089 , \9087 , \9088 );
xor \U$8286 ( \9090 , \9043 , \9046 );
nor \U$8287 ( \9091 , \9089 , \9090 );
not \U$8288 ( \9092 , \9091 );
not \U$8289 ( \9093 , \9048 );
nor \U$8290 ( \9094 , \9092 , \9093 );
not \U$8291 ( \9095 , \9094 );
or \U$8292 ( \9096 , \9095 , \8516 );
or \U$8293 ( \9097 , \9092 , \8516 );
nand \U$8294 ( \9098 , \9097 , \9093 );
nand \U$8295 ( \9099 , \9096 , \9098 );
or \U$8296 ( \9100 , \8891 , \8590 );
not \U$8297 ( \9101 , \9030 );
or \U$8298 ( \9102 , \8475 , \9101 );
or \U$8299 ( \9103 , \8888 , \8590 );
or \U$8300 ( \9104 , \8816 , \8474_nG30a2 );
nand \U$8301 ( \9105 , \9104 , \9026 );
nand \U$8302 ( \9106 , \9103 , \9105 );
nand \U$8303 ( \9107 , \9100 , \9102 , \9106 );
and \U$8304 ( \9108 , \9099 , \9107 );
not \U$8305 ( \9109 , \8947_nG2a93 );
or \U$8306 ( \9110 , \8527 , \9109 );
not \U$8307 ( \9111 , \9018_nG29b3 );
or \U$8308 ( \9112 , \9111 , \8522 );
or \U$8309 ( \9113 , \8519 , \9109 );
or \U$8310 ( \9114 , \8487 , \9018_nG29b3 );
nand \U$8311 ( \9115 , \9114 , \8524 );
nand \U$8312 ( \9116 , \9113 , \9115 );
nand \U$8313 ( \9117 , \9110 , \9112 , \9116 );
nand \U$8314 ( \9118 , \8657_nG2e7a , \8767 );
or \U$8315 ( \9119 , \8624 , \8729_nG2d90 );
nand \U$8316 ( \9120 , \9119 , \8773 );
and \U$8317 ( \9121 , \9118 , \9120 );
and \U$8318 ( \9122 , \8769 , \8729_nG2d90 );
and \U$8319 ( \9123 , \8657_nG2e7a , \8831 );
nor \U$8320 ( \9124 , \9121 , \9122 , \9123 );
nand \U$8321 ( \9125 , \8868_nG2b9c , \8580 );
or \U$8322 ( \9126 , \8540 , \8762_nG2c8f );
nand \U$8323 ( \9127 , \9126 , \8615 );
and \U$8324 ( \9128 , \9125 , \9127 );
and \U$8325 ( \9129 , \8610 , \8762_nG2c8f );
and \U$8326 ( \9130 , \8868_nG2b9c , \8583 );
nor \U$8327 ( \9131 , \9128 , \9129 , \9130 );
nand \U$8328 ( \9132 , \9124 , \9131 );
and \U$8329 ( \9133 , \9117 , \9132 );
nor \U$8330 ( \9134 , \9131 , \9124 );
nor \U$8331 ( \9135 , \9133 , \9134 );
not \U$8332 ( \9136 , \9135 );
and \U$8333 ( \9137 , \9108 , \9136 );
not \U$8334 ( \9138 , \9048 );
not \U$8335 ( \9139 , \9050 );
nand \U$8336 ( \9140 , \9139 , \9040 );
not \U$8337 ( \9141 , \9140 );
or \U$8338 ( \9142 , \9138 , \9141 );
or \U$8339 ( \9143 , \9140 , \9048 );
nand \U$8340 ( \9144 , \9142 , \9143 );
not \U$8341 ( \9145 , \9019 );
nor \U$8342 ( \9146 , \8990 , \9022 );
not \U$8343 ( \9147 , \9146 );
or \U$8344 ( \9148 , \9145 , \9147 );
or \U$8345 ( \9149 , \9146 , \9019 );
nand \U$8346 ( \9150 , \9148 , \9149 );
and \U$8347 ( \9151 , \9144 , \9150 );
and \U$8348 ( \9152 , \9137 , \9151 );
xor \U$8349 ( \9153 , \9084 , \9152 );
xnor \U$8350 ( \9154 , \9051 , \9023 );
not \U$8351 ( \9155 , \9061 );
not \U$8352 ( \9156 , \9053 );
and \U$8353 ( \9157 , \9155 , \9156 );
and \U$8354 ( \9158 , \9061 , \9053 );
nor \U$8355 ( \9159 , \9157 , \9158 );
nand \U$8356 ( \9160 , \9154 , \9159 );
and \U$8357 ( \9161 , \9153 , \9160 );
and \U$8358 ( \9162 , \9084 , \9152 );
or \U$8359 ( \9163 , \9161 , \9162 );
xor \U$8360 ( \9164 , \8880 , \8952 );
xor \U$8361 ( \9165 , \9163 , \9164 );
xor \U$8362 ( \9166 , \9063 , \9066 );
xor \U$8363 ( \9167 , \9166 , \9069 );
and \U$8364 ( \9168 , \9165 , \9167 );
and \U$8365 ( \9169 , \9163 , \9164 );
or \U$8366 ( \9170 , \9168 , \9169 );
xor \U$8367 ( \9171 , \9083 , \9170 );
xor \U$8368 ( \9172 , \9052 , \9062 );
xor \U$8369 ( \9173 , \9084 , \9152 );
xor \U$8370 ( \9174 , \9173 , \9160 );
and \U$8371 ( \9175 , \9172 , \9174 );
xor \U$8372 ( \9176 , \9108 , \9136 );
xor \U$8373 ( \9177 , \9144 , \9150 );
and \U$8374 ( \9178 , \9176 , \9177 );
xor \U$8375 ( \9179 , \9099 , \9107 );
not \U$8376 ( \9180 , \9134 );
nand \U$8377 ( \9181 , \9180 , \9132 );
not \U$8378 ( \9182 , \9181 );
not \U$8379 ( \9183 , \9117 );
or \U$8380 ( \9184 , \9182 , \9183 );
or \U$8381 ( \9185 , \9117 , \9181 );
nand \U$8382 ( \9186 , \9184 , \9185 );
and \U$8383 ( \9187 , \9179 , \9186 );
and \U$8384 ( \9188 , \9048 , \9090 );
and \U$8385 ( \9189 , \8514_nG31b0 , \9188 );
or \U$8386 ( \9190 , \9048 , \8514_nG31b0 );
or \U$8387 ( \9191 , \9048 , \9090 );
nand \U$8388 ( \9192 , \9190 , \9191 );
nand \U$8389 ( \9193 , \8474_nG30a2 , \9091 );
and \U$8390 ( \9194 , \9192 , \9193 );
and \U$8391 ( \9195 , \8474_nG30a2 , \9094 );
nor \U$8392 ( \9196 , \9189 , \9194 , \9195 );
xor \U$8393 ( \9197 , RIaaa91a0_605, \8371_nG221f );
xor \U$8394 ( \9198 , \9197 , \8405 );
not \U$8395 ( \9199 , \9198 );
xor \U$8396 ( \9200 , \8308 , \8338_nG2292 );
xor \U$8397 ( \9201 , \9200 , \8408 );
not \U$8398 ( \9202 , \9201 );
and \U$8399 ( \9203 , \9199 , \9202 );
or \U$8400 ( \9204 , \9042 , \9203 );
not \U$8401 ( \9205 , \9204 );
xor \U$8402 ( \9206 , \9196 , \9205 );
and \U$8403 ( \9207 , \8657_nG2e7a , \8890 );
or \U$8404 ( \9208 , \8816 , \8568_nG2f9c );
nand \U$8405 ( \9209 , \9208 , \9026 );
nand \U$8406 ( \9210 , \8657_nG2e7a , \8887 );
and \U$8407 ( \9211 , \9209 , \9210 );
and \U$8408 ( \9212 , \8568_nG2f9c , \9030 );
nor \U$8409 ( \9213 , \9207 , \9211 , \9212 );
and \U$8410 ( \9214 , \9206 , \9213 );
and \U$8411 ( \9215 , \9196 , \9205 );
or \U$8412 ( \9216 , \9214 , \9215 );
not \U$8413 ( \9217 , \9216 );
nand \U$8414 ( \9218 , \8947_nG2a93 , \8580 );
or \U$8415 ( \9219 , \8540 , \8868_nG2b9c );
nand \U$8416 ( \9220 , \9219 , \8615 );
and \U$8417 ( \9221 , \9218 , \9220 );
and \U$8418 ( \9222 , \8610 , \8868_nG2b9c );
and \U$8419 ( \9223 , \8947_nG2a93 , \8583 );
nor \U$8420 ( \9224 , \9221 , \9222 , \9223 );
nand \U$8421 ( \9225 , \8729_nG2d90 , \8767 );
or \U$8422 ( \9226 , \8624 , \8762_nG2c8f );
nand \U$8423 ( \9227 , \9226 , \8773 );
and \U$8424 ( \9228 , \9225 , \9227 );
and \U$8425 ( \9229 , \8769 , \8762_nG2c8f );
and \U$8426 ( \9230 , \8729_nG2d90 , \8831 );
nor \U$8427 ( \9231 , \9228 , \9229 , \9230 );
xor \U$8428 ( \9232 , \9224 , \9231 );
and \U$8429 ( \9233 , \9018_nG29b3 , \8629 );
and \U$8430 ( \9234 , RIaaa3c50_423, \7928 );
and \U$8431 ( \9235 , RIaaa3d40_425, \7930 );
and \U$8432 ( \9236 , \7952 , RIaaa3f98_430);
and \U$8433 ( \9237 , RIaaa3e30_427, \7957 );
nor \U$8434 ( \9238 , \9236 , \9237 );
and \U$8435 ( \9239 , \7942 , RIaaa3ea8_428);
and \U$8436 ( \9240 , RIaaa3b60_421, \7909 );
nor \U$8437 ( \9241 , \9239 , \9240 );
and \U$8438 ( \9242 , \7914 , RIaaa4088_432);
and \U$8439 ( \9243 , RIaaa3f20_429, \7949 );
nor \U$8440 ( \9244 , \9242 , \9243 );
and \U$8441 ( \9245 , \7959 , RIaaa3a70_419);
and \U$8442 ( \9246 , RIaaa3ae8_420, \7944 );
nor \U$8443 ( \9247 , \9245 , \9246 );
nand \U$8444 ( \9248 , \9238 , \9241 , \9244 , \9247 );
nor \U$8445 ( \9249 , \9234 , \9235 , \9248 );
and \U$8446 ( \9250 , \8454 , RIaaa4100_433);
and \U$8447 ( \9251 , RIaaa3bd8_422, \7963 );
nor \U$8448 ( \9252 , \9250 , \9251 );
and \U$8449 ( \9253 , \7961 , RIaaa4010_431);
and \U$8450 ( \9254 , RIaaa39f8_418, \7919 );
nor \U$8451 ( \9255 , \9253 , \9254 );
and \U$8452 ( \9256 , \7935 , RIaaa3cc8_424);
and \U$8453 ( \9257 , RIaaa4178_434, \7924 );
nor \U$8454 ( \9258 , \9256 , \9257 );
nand \U$8455 ( \9259 , \9249 , \9252 , \9255 , \9258 );
_DC g28b3 ( \9260_nG28b3 , \9259 , \8473 );
or \U$8456 ( \9261 , \8487 , \9260_nG28b3 );
nand \U$8457 ( \9262 , \9261 , \8524 );
nand \U$8458 ( \9263 , \9018_nG29b3 , \8520 );
and \U$8459 ( \9264 , \9262 , \9263 );
and \U$8460 ( \9265 , \9260_nG28b3 , \8662 );
nor \U$8461 ( \9266 , \9233 , \9264 , \9265 );
and \U$8462 ( \9267 , \9232 , \9266 );
and \U$8463 ( \9268 , \9224 , \9231 );
or \U$8464 ( \9269 , \9267 , \9268 );
not \U$8465 ( \9270 , \9269 );
and \U$8466 ( \9271 , \9217 , \9270 );
and \U$8467 ( \9272 , \9187 , \9271 );
xor \U$8468 ( \9273 , \9178 , \9272 );
or \U$8469 ( \9274 , \9159 , \9154 );
nand \U$8470 ( \9275 , \9274 , \9160 );
and \U$8471 ( \9276 , \9273 , \9275 );
and \U$8472 ( \9277 , \9178 , \9272 );
or \U$8473 ( \9278 , \9276 , \9277 );
xor \U$8474 ( \9279 , \9084 , \9152 );
xor \U$8475 ( \9280 , \9279 , \9160 );
and \U$8476 ( \9281 , \9278 , \9280 );
and \U$8477 ( \9282 , \9172 , \9278 );
or \U$8478 ( \9283 , \9175 , \9281 , \9282 );
xor \U$8479 ( \9284 , \9163 , \9164 );
xor \U$8480 ( \9285 , \9284 , \9167 );
xor \U$8481 ( \9286 , \9283 , \9285 );
xor \U$8482 ( \9287 , \9084 , \9152 );
xor \U$8483 ( \9288 , \9287 , \9160 );
xor \U$8484 ( \9289 , \9172 , \9278 );
xor \U$8485 ( \9290 , \9288 , \9289 );
and \U$8486 ( \9291 , RIaaa3278_402, \7957 );
and \U$8487 ( \9292 , RIaaa32f0_403, \7942 );
and \U$8488 ( \9293 , \7924 , RIaaa35c0_409);
and \U$8489 ( \9294 , RIaaa3980_417, \7930 );
nor \U$8490 ( \9295 , \9293 , \9294 );
and \U$8491 ( \9296 , \7961 , RIaaa3458_406);
and \U$8492 ( \9297 , RIaaa3638_410, \7963 );
nor \U$8493 ( \9298 , \9296 , \9297 );
and \U$8494 ( \9299 , \8454 , RIaaa3548_408);
and \U$8495 ( \9300 , RIaaa3908_416, \7935 );
nor \U$8496 ( \9301 , \9299 , \9300 );
and \U$8497 ( \9302 , \7928 , RIaaa36b0_411);
and \U$8498 ( \9303 , RIaaa37a0_413, \7909 );
nor \U$8499 ( \9304 , \9302 , \9303 );
nand \U$8500 ( \9305 , \9295 , \9298 , \9301 , \9304 );
nor \U$8501 ( \9306 , \9291 , \9292 , \9305 );
and \U$8502 ( \9307 , \7949 , RIaaa3368_404);
and \U$8503 ( \9308 , RIaaa33e0_405, \7952 );
nor \U$8504 ( \9309 , \9307 , \9308 );
and \U$8505 ( \9310 , \7914 , RIaaa34d0_407);
and \U$8506 ( \9311 , RIaaa3890_415, \7959 );
nor \U$8507 ( \9312 , \9310 , \9311 );
and \U$8508 ( \9313 , \7919 , RIaaa3818_414);
and \U$8509 ( \9314 , RIaaa3728_412, \7944 );
nor \U$8510 ( \9315 , \9313 , \9314 );
nand \U$8511 ( \9316 , \9306 , \9309 , \9312 , \9315 );
_DC g27da ( \9317_nG27da , \9316 , \8473 );
nand \U$8512 ( \9318 , \9317_nG27da , \8444 );
not \U$8513 ( \9319 , \9318 );
xor \U$8514 ( \9320 , \9224 , \9231 );
xor \U$8515 ( \9321 , \9320 , \9266 );
xor \U$8516 ( \9322 , \9196 , \9205 );
xor \U$8517 ( \9323 , \9322 , \9213 );
nor \U$8518 ( \9324 , \9321 , \9323 );
nor \U$8519 ( \9325 , \9319 , \9324 );
not \U$8520 ( \9326 , \9325 );
or \U$8521 ( \9327 , \9042 , \9201 );
nand \U$8522 ( \9328 , \9201 , \9042 );
nand \U$8523 ( \9329 , \9327 , \9328 );
xor \U$8524 ( \9330 , \9199 , \9202 );
nor \U$8525 ( \9331 , \9329 , \9330 );
not \U$8526 ( \9332 , \9331 );
nor \U$8527 ( \9333 , \9332 , \9205 );
not \U$8528 ( \9334 , \9333 );
or \U$8529 ( \9335 , \9334 , \8516 );
or \U$8530 ( \9336 , \9332 , \8516 );
nand \U$8531 ( \9337 , \9336 , \9205 );
nand \U$8532 ( \9338 , \9335 , \9337 );
not \U$8533 ( \9339 , \9338 );
and \U$8534 ( \9340 , \8474_nG30a2 , \9188 );
or \U$8535 ( \9341 , \9048 , \8474_nG30a2 );
nand \U$8536 ( \9342 , \9341 , \9191 );
nand \U$8537 ( \9343 , \8568_nG2f9c , \9091 );
and \U$8538 ( \9344 , \9342 , \9343 );
and \U$8539 ( \9345 , \8568_nG2f9c , \9094 );
nor \U$8540 ( \9346 , \9340 , \9344 , \9345 );
nor \U$8541 ( \9347 , \9339 , \9346 );
not \U$8542 ( \9348 , \9347 );
nand \U$8543 ( \9349 , \8762_nG2c8f , \8767 );
or \U$8544 ( \9350 , \8624 , \8868_nG2b9c );
nand \U$8545 ( \9351 , \9350 , \8773 );
and \U$8546 ( \9352 , \9349 , \9351 );
and \U$8547 ( \9353 , \8769 , \8868_nG2b9c );
and \U$8548 ( \9354 , \8762_nG2c8f , \8831 );
nor \U$8549 ( \9355 , \9352 , \9353 , \9354 );
and \U$8550 ( \9356 , \8729_nG2d90 , \8890 );
or \U$8551 ( \9357 , \8816 , \8657_nG2e7a );
nand \U$8552 ( \9358 , \9357 , \9026 );
nand \U$8553 ( \9359 , \8729_nG2d90 , \8887 );
and \U$8554 ( \9360 , \9358 , \9359 );
and \U$8555 ( \9361 , \8657_nG2e7a , \9030 );
nor \U$8556 ( \9362 , \9356 , \9360 , \9361 );
xor \U$8557 ( \9363 , \9355 , \9362 );
nand \U$8558 ( \9364 , \9018_nG29b3 , \8580 );
or \U$8559 ( \9365 , \8540 , \8947_nG2a93 );
nand \U$8560 ( \9366 , \9365 , \8615 );
and \U$8561 ( \9367 , \9364 , \9366 );
and \U$8562 ( \9368 , \8610 , \8947_nG2a93 );
and \U$8563 ( \9369 , \9018_nG29b3 , \8583 );
nor \U$8564 ( \9370 , \9367 , \9368 , \9369 );
and \U$8565 ( \9371 , \9363 , \9370 );
and \U$8566 ( \9372 , \9355 , \9362 );
or \U$8567 ( \9373 , \9371 , \9372 );
nor \U$8568 ( \9374 , \9348 , \9373 );
nand \U$8569 ( \9375 , \9326 , \9374 );
xor \U$8570 ( \9376 , \9179 , \9186 );
nand \U$8571 ( \9377 , \9260_nG28b3 , \8444 );
and \U$8572 ( \9378 , \9376 , \9377 );
xor \U$8573 ( \9379 , \9217 , \9270 );
nor \U$8574 ( \9380 , \9378 , \9379 );
or \U$8575 ( \9381 , \9375 , \9380 );
not \U$8576 ( \9382 , \9380 );
not \U$8577 ( \9383 , \9375 );
or \U$8578 ( \9384 , \9382 , \9383 );
xor \U$8579 ( \9385 , \9176 , \9177 );
nand \U$8580 ( \9386 , \9384 , \9385 );
nand \U$8581 ( \9387 , \9381 , \9386 );
xor \U$8582 ( \9388 , \9137 , \9151 );
xor \U$8583 ( \9389 , \9387 , \9388 );
xor \U$8584 ( \9390 , \9178 , \9272 );
xor \U$8585 ( \9391 , \9390 , \9275 );
and \U$8586 ( \9392 , \9389 , \9391 );
and \U$8587 ( \9393 , \9387 , \9388 );
or \U$8588 ( \9394 , \9392 , \9393 );
xor \U$8589 ( \9395 , \9290 , \9394 );
xor \U$8590 ( \9396 , \9387 , \9388 );
xor \U$8591 ( \9397 , \9396 , \9391 );
xor \U$8592 ( \9398 , \9377 , \9376 );
xor \U$8593 ( \9399 , \9379 , \9398 );
nand \U$8594 ( \9400 , \8868_nG2b9c , \8767 );
or \U$8595 ( \9401 , \8624 , \8947_nG2a93 );
nand \U$8596 ( \9402 , \9401 , \8773 );
and \U$8597 ( \9403 , \9400 , \9402 );
and \U$8598 ( \9404 , \8769 , \8947_nG2a93 );
and \U$8599 ( \9405 , \8868_nG2b9c , \8831 );
nor \U$8600 ( \9406 , \9403 , \9404 , \9405 );
and \U$8601 ( \9407 , \8762_nG2c8f , \8890 );
or \U$8602 ( \9408 , \8816 , \8729_nG2d90 );
nand \U$8603 ( \9409 , \9408 , \9026 );
nand \U$8604 ( \9410 , \8762_nG2c8f , \8887 );
and \U$8605 ( \9411 , \9409 , \9410 );
and \U$8606 ( \9412 , \8729_nG2d90 , \9030 );
nor \U$8607 ( \9413 , \9407 , \9411 , \9412 );
xor \U$8608 ( \9414 , \9406 , \9413 );
nand \U$8609 ( \9415 , \9260_nG28b3 , \8580 );
or \U$8610 ( \9416 , \8540 , \9018_nG29b3 );
nand \U$8611 ( \9417 , \9416 , \8615 );
and \U$8612 ( \9418 , \9415 , \9417 );
and \U$8613 ( \9419 , \8610 , \9018_nG29b3 );
and \U$8614 ( \9420 , \9260_nG28b3 , \8583 );
nor \U$8615 ( \9421 , \9418 , \9419 , \9420 );
and \U$8616 ( \9422 , \9414 , \9421 );
and \U$8617 ( \9423 , \9406 , \9413 );
or \U$8618 ( \9424 , \9422 , \9423 );
nand \U$8619 ( \9425 , \8474_nG30a2 , \9331 );
or \U$8620 ( \9426 , \9204 , \8514_nG31b0 );
or \U$8621 ( \9427 , \9204 , \9330 );
nand \U$8622 ( \9428 , \9426 , \9427 );
and \U$8623 ( \9429 , \9425 , \9428 );
and \U$8624 ( \9430 , \9204 , \9330 );
and \U$8625 ( \9431 , \9430 , \8514_nG31b0 );
and \U$8626 ( \9432 , \8474_nG30a2 , \9333 );
nor \U$8627 ( \9433 , \9429 , \9431 , \9432 );
xor \U$8628 ( \9434 , \9433 , \9199 );
and \U$8629 ( \9435 , \8568_nG2f9c , \9188 );
or \U$8630 ( \9436 , \9048 , \8568_nG2f9c );
nand \U$8631 ( \9437 , \9436 , \9191 );
nand \U$8632 ( \9438 , \8657_nG2e7a , \9091 );
and \U$8633 ( \9439 , \9437 , \9438 );
and \U$8634 ( \9440 , \8657_nG2e7a , \9094 );
nor \U$8635 ( \9441 , \9435 , \9439 , \9440 );
and \U$8636 ( \9442 , \9434 , \9441 );
and \U$8637 ( \9443 , \9433 , \9199 );
or \U$8638 ( \9444 , \9442 , \9443 );
nor \U$8639 ( \9445 , \9424 , \9444 );
not \U$8640 ( \9446 , \9445 );
xor \U$8641 ( \9447 , \9355 , \9362 );
xor \U$8642 ( \9448 , \9447 , \9370 );
not \U$8643 ( \9449 , \9346 );
not \U$8644 ( \9450 , \9338 );
and \U$8645 ( \9451 , \9449 , \9450 );
and \U$8646 ( \9452 , \9346 , \9338 );
nor \U$8647 ( \9453 , \9451 , \9452 );
xor \U$8648 ( \9454 , \9448 , \9453 );
and \U$8649 ( \9455 , RIaaa42e0_437, \8454 );
and \U$8650 ( \9456 , RIaaa4790_447, \7930 );
and \U$8651 ( \9457 , \7963 , RIaaa48f8_450);
and \U$8652 ( \9458 , RIaaa4808_448, \7944 );
nor \U$8653 ( \9459 , \9457 , \9458 );
and \U$8654 ( \9460 , \7949 , RIaaa4448_440);
and \U$8655 ( \9461 , RIaaa4538_442, \7952 );
nor \U$8656 ( \9462 , \9460 , \9461 );
and \U$8657 ( \9463 , \7914 , RIaaa4268_436);
and \U$8658 ( \9464 , RIaaa44c0_441, \7942 );
nor \U$8659 ( \9465 , \9463 , \9464 );
and \U$8660 ( \9466 , \7919 , RIaaa4628_444);
and \U$8661 ( \9467 , RIaaa46a0_445, \7959 );
nor \U$8662 ( \9468 , \9466 , \9467 );
nand \U$8663 ( \9469 , \9459 , \9462 , \9465 , \9468 );
nor \U$8664 ( \9470 , \9455 , \9456 , \9469 );
and \U$8665 ( \9471 , \7935 , RIaaa4718_446);
and \U$8666 ( \9472 , RIaaa43d0_439, \7957 );
nor \U$8667 ( \9473 , \9471 , \9472 );
and \U$8668 ( \9474 , \7961 , RIaaa45b0_443);
and \U$8669 ( \9475 , RIaaa4970_451, \7928 );
nor \U$8670 ( \9476 , \9474 , \9475 );
and \U$8671 ( \9477 , \7924 , RIaaa4358_438);
and \U$8672 ( \9478 , RIaaa4880_449, \7909 );
nor \U$8673 ( \9479 , \9477 , \9478 );
nand \U$8674 ( \9480 , \9470 , \9473 , \9476 , \9479 );
_DC g2706 ( \9481_nG2706 , \9480 , \8473 );
nand \U$8675 ( \9482 , \9481_nG2706 , \8444 );
and \U$8676 ( \9483 , \9260_nG28b3 , \8629 );
or \U$8677 ( \9484 , \8487 , \9317_nG27da );
nand \U$8678 ( \9485 , \9484 , \8524 );
nand \U$8679 ( \9486 , \9260_nG28b3 , \8520 );
and \U$8680 ( \9487 , \9485 , \9486 );
and \U$8681 ( \9488 , \9317_nG27da , \8662 );
nor \U$8682 ( \9489 , \9483 , \9487 , \9488 );
xnor \U$8683 ( \9490 , \9482 , \9489 );
and \U$8684 ( \9491 , \9454 , \9490 );
and \U$8685 ( \9492 , \9448 , \9453 );
or \U$8686 ( \9493 , \9491 , \9492 );
nor \U$8687 ( \9494 , \9446 , \9493 );
nor \U$8688 ( \9495 , \9399 , \9494 );
and \U$8689 ( \9496 , \9321 , \9323 );
nor \U$8690 ( \9497 , \9496 , \9324 );
not \U$8691 ( \9498 , \9497 );
not \U$8692 ( \9499 , \9318 );
and \U$8693 ( \9500 , \9498 , \9499 );
and \U$8694 ( \9501 , \9497 , \9318 );
nor \U$8695 ( \9502 , \9500 , \9501 );
not \U$8696 ( \9503 , \9502 );
or \U$8697 ( \9504 , \9373 , \9347 );
or \U$8698 ( \9505 , \9482 , \9489 );
nand \U$8699 ( \9506 , \9347 , \9373 );
nand \U$8700 ( \9507 , \9504 , \9505 , \9506 );
nand \U$8701 ( \9508 , \9503 , \9507 );
or \U$8702 ( \9509 , \9495 , \9508 );
nand \U$8703 ( \9510 , \9494 , \9399 );
nand \U$8704 ( \9511 , \9509 , \9510 );
not \U$8705 ( \9512 , \9187 );
not \U$8706 ( \9513 , \9377 );
nor \U$8707 ( \9514 , \9513 , \9271 );
not \U$8708 ( \9515 , \9514 );
or \U$8709 ( \9516 , \9512 , \9515 );
or \U$8710 ( \9517 , \9514 , \9187 );
nand \U$8711 ( \9518 , \9516 , \9517 );
nor \U$8712 ( \9519 , \9511 , \9518 );
xnor \U$8713 ( \9520 , \9380 , \9375 );
not \U$8714 ( \9521 , \9520 );
not \U$8715 ( \9522 , \9385 );
and \U$8716 ( \9523 , \9521 , \9522 );
and \U$8717 ( \9524 , \9520 , \9385 );
nor \U$8718 ( \9525 , \9523 , \9524 );
or \U$8719 ( \9526 , \9519 , \9525 );
nand \U$8720 ( \9527 , \9518 , \9511 );
nand \U$8721 ( \9528 , \9526 , \9527 );
xor \U$8722 ( \9529 , \9397 , \9528 );
not \U$8723 ( \9530 , \9525 );
not \U$8724 ( \9531 , \9519 );
nand \U$8725 ( \9532 , \9531 , \9527 );
not \U$8726 ( \9533 , \9532 );
or \U$8727 ( \9534 , \9530 , \9533 );
or \U$8728 ( \9535 , \9532 , \9525 );
nand \U$8729 ( \9536 , \9534 , \9535 );
and \U$8730 ( \9537 , RIaaa6860_517, \7919 );
and \U$8731 ( \9538 , RIaaa6680_513, \7944 );
and \U$8732 ( \9539 , \7924 , RIaaa6338_506);
and \U$8733 ( \9540 , RIaaa6950_519, \7930 );
nor \U$8734 ( \9541 , \9539 , \9540 );
and \U$8735 ( \9542 , \7961 , RIaaa6518_510);
and \U$8736 ( \9543 , RIaaa66f8_514, \7963 );
nor \U$8737 ( \9544 , \9542 , \9543 );
and \U$8738 ( \9545 , \8454 , RIaaa62c0_505);
and \U$8739 ( \9546 , RIaaa68d8_518, \7935 );
nor \U$8740 ( \9547 , \9545 , \9546 );
and \U$8741 ( \9548 , \7928 , RIaaa6770_515);
and \U$8742 ( \9549 , RIaaa6608_512, \7909 );
nor \U$8743 ( \9550 , \9548 , \9549 );
nand \U$8744 ( \9551 , \9541 , \9544 , \9547 , \9550 );
nor \U$8745 ( \9552 , \9537 , \9538 , \9551 );
and \U$8746 ( \9553 , \7942 , RIaaa64a0_509);
and \U$8747 ( \9554 , RIaaa63b0_507, \7957 );
nor \U$8748 ( \9555 , \9553 , \9554 );
and \U$8749 ( \9556 , \7914 , RIaaa6248_504);
and \U$8750 ( \9557 , RIaaa6590_511, \7952 );
nor \U$8751 ( \9558 , \9556 , \9557 );
and \U$8752 ( \9559 , \7949 , RIaaa6428_508);
and \U$8753 ( \9560 , RIaaa67e8_516, \7959 );
nor \U$8754 ( \9561 , \9559 , \9560 );
nand \U$8755 ( \9562 , \9552 , \9555 , \9558 , \9561 );
_DC g23ac ( \9563_nG23ac , \9562 , \8473 );
nand \U$8756 ( \9564 , \9563_nG23ac , \8444 );
and \U$8757 ( \9565 , \9317_nG27da , \8629 );
or \U$8758 ( \9566 , \8487 , \9481_nG2706 );
nand \U$8759 ( \9567 , \9566 , \8524 );
nand \U$8760 ( \9568 , \9317_nG27da , \8520 );
and \U$8761 ( \9569 , \9567 , \9568 );
and \U$8762 ( \9570 , \9481_nG2706 , \8662 );
nor \U$8763 ( \9571 , \9565 , \9569 , \9570 );
xnor \U$8764 ( \9572 , \9564 , \9571 );
xor \U$8765 ( \9573 , \9448 , \9453 );
xor \U$8766 ( \9574 , \9573 , \9490 );
and \U$8767 ( \9575 , \9572 , \9574 );
and \U$8768 ( \9576 , \8868_nG2b9c , \8890 );
or \U$8769 ( \9577 , \8816 , \8762_nG2c8f );
nand \U$8770 ( \9578 , \9577 , \9026 );
nand \U$8771 ( \9579 , \8868_nG2b9c , \8887 );
and \U$8772 ( \9580 , \9578 , \9579 );
and \U$8773 ( \9581 , \8762_nG2c8f , \9030 );
nor \U$8774 ( \9582 , \9576 , \9580 , \9581 );
and \U$8775 ( \9583 , \8657_nG2e7a , \9188 );
or \U$8776 ( \9584 , \9048 , \8657_nG2e7a );
nand \U$8777 ( \9585 , \9584 , \9191 );
nand \U$8778 ( \9586 , \8729_nG2d90 , \9091 );
and \U$8779 ( \9587 , \9585 , \9586 );
and \U$8780 ( \9588 , \8729_nG2d90 , \9094 );
nor \U$8781 ( \9589 , \9583 , \9587 , \9588 );
xor \U$8782 ( \9590 , \9582 , \9589 );
nand \U$8783 ( \9591 , \8947_nG2a93 , \8767 );
or \U$8784 ( \9592 , \8624 , \9018_nG29b3 );
nand \U$8785 ( \9593 , \9592 , \8773 );
and \U$8786 ( \9594 , \9591 , \9593 );
and \U$8787 ( \9595 , \8769 , \9018_nG29b3 );
and \U$8788 ( \9596 , \8947_nG2a93 , \8831 );
nor \U$8789 ( \9597 , \9594 , \9595 , \9596 );
and \U$8790 ( \9598 , \9590 , \9597 );
and \U$8791 ( \9599 , \9582 , \9589 );
or \U$8792 ( \9600 , \9598 , \9599 );
nand \U$8793 ( \9601 , \8568_nG2f9c , \9331 );
or \U$8794 ( \9602 , \9204 , \8474_nG30a2 );
nand \U$8795 ( \9603 , \9602 , \9427 );
and \U$8796 ( \9604 , \9601 , \9603 );
and \U$8797 ( \9605 , \9430 , \8474_nG30a2 );
and \U$8798 ( \9606 , \8568_nG2f9c , \9333 );
nor \U$8799 ( \9607 , \9604 , \9605 , \9606 );
not \U$8800 ( \9608 , \9607 );
or \U$8801 ( \9609 , \9198 , \8514_nG31b0 );
or \U$8802 ( \9610 , \8403 , \8402_nG221d );
nand \U$8803 ( \9611 , \9610 , \8404 );
nor \U$8804 ( \9612 , \9198 , \9611 );
not \U$8805 ( \9613 , \9612 );
nand \U$8806 ( \9614 , \9199 , \9613 );
nand \U$8807 ( \9615 , \9609 , \9614 );
nand \U$8808 ( \9616 , \9608 , \9615 );
xor \U$8809 ( \9617 , \9600 , \9616 );
and \U$8810 ( \9618 , \9481_nG2706 , \8629 );
or \U$8811 ( \9619 , \8487 , \9563_nG23ac );
nand \U$8812 ( \9620 , \9619 , \8524 );
nand \U$8813 ( \9621 , \9481_nG2706 , \8520 );
and \U$8814 ( \9622 , \9620 , \9621 );
and \U$8815 ( \9623 , \9563_nG23ac , \8662 );
nor \U$8816 ( \9624 , \9618 , \9622 , \9623 );
nand \U$8817 ( \9625 , \9317_nG27da , \8580 );
or \U$8818 ( \9626 , \8540 , \9260_nG28b3 );
nand \U$8819 ( \9627 , \9626 , \8615 );
and \U$8820 ( \9628 , \9625 , \9627 );
and \U$8821 ( \9629 , \8610 , \9260_nG28b3 );
and \U$8822 ( \9630 , \9317_nG27da , \8583 );
nor \U$8823 ( \9631 , \9628 , \9629 , \9630 );
and \U$8824 ( \9632 , \9624 , \9631 );
not \U$8825 ( \9633 , \9632 );
and \U$8826 ( \9634 , RIaaa5870_483, \7928 );
and \U$8827 ( \9635 , RIaaa58e8_484, \7930 );
and \U$8828 ( \9636 , \7952 , RIaaa53c0_473);
and \U$8829 ( \9637 , RIaaa5258_470, \7957 );
nor \U$8830 ( \9638 , \9636 , \9637 );
and \U$8831 ( \9639 , \7942 , RIaaa52d0_471);
and \U$8832 ( \9640 , RIaaa5618_478, \7919 );
nor \U$8833 ( \9641 , \9639 , \9640 );
and \U$8834 ( \9642 , \7914 , RIaaa54b0_475);
and \U$8835 ( \9643 , RIaaa5348_472, \7949 );
nor \U$8836 ( \9644 , \9642 , \9643 );
and \U$8837 ( \9645 , \7959 , RIaaa5690_479);
and \U$8838 ( \9646 , RIaaa5708_480, \7944 );
nor \U$8839 ( \9647 , \9645 , \9646 );
nand \U$8840 ( \9648 , \9638 , \9641 , \9644 , \9647 );
nor \U$8841 ( \9649 , \9634 , \9635 , \9648 );
and \U$8842 ( \9650 , \7961 , RIaaa5438_474);
and \U$8843 ( \9651 , RIaaa5780_481, \7909 );
nor \U$8844 ( \9652 , \9650 , \9651 );
and \U$8845 ( \9653 , \8454 , RIaaa55a0_477);
and \U$8846 ( \9654 , RIaaa57f8_482, \7963 );
nor \U$8847 ( \9655 , \9653 , \9654 );
and \U$8848 ( \9656 , \7935 , RIaaa5960_485);
and \U$8849 ( \9657 , RIaaa5528_476, \7924 );
nor \U$8850 ( \9658 , \9656 , \9657 );
nand \U$8851 ( \9659 , \9649 , \9652 , \9655 , \9658 );
_DC g2373 ( \9660_nG2373 , \9659 , \8473 );
nand \U$8852 ( \9661 , \9660_nG2373 , \8444 );
not \U$8853 ( \9662 , \9661 );
and \U$8854 ( \9663 , \9633 , \9662 );
nor \U$8855 ( \9664 , \9624 , \9631 );
nor \U$8856 ( \9665 , \9663 , \9664 );
and \U$8857 ( \9666 , \9617 , \9665 );
and \U$8858 ( \9667 , \9600 , \9616 );
or \U$8859 ( \9668 , \9666 , \9667 );
xor \U$8860 ( \9669 , \9448 , \9453 );
xor \U$8861 ( \9670 , \9669 , \9490 );
and \U$8862 ( \9671 , \9668 , \9670 );
and \U$8863 ( \9672 , \9572 , \9668 );
or \U$8864 ( \9673 , \9575 , \9671 , \9672 );
not \U$8865 ( \9674 , \9493 );
not \U$8866 ( \9675 , \9445 );
and \U$8867 ( \9676 , \9674 , \9675 );
and \U$8868 ( \9677 , \9493 , \9445 );
nor \U$8869 ( \9678 , \9676 , \9677 );
xor \U$8870 ( \9679 , \9673 , \9678 );
not \U$8871 ( \9680 , \9502 );
not \U$8872 ( \9681 , \9507 );
and \U$8873 ( \9682 , \9680 , \9681 );
and \U$8874 ( \9683 , \9502 , \9507 );
nor \U$8875 ( \9684 , \9682 , \9683 );
and \U$8876 ( \9685 , \9679 , \9684 );
and \U$8877 ( \9686 , \9673 , \9678 );
or \U$8878 ( \9687 , \9685 , \9686 );
not \U$8879 ( \9688 , \9325 );
not \U$8880 ( \9689 , \9374 );
and \U$8881 ( \9690 , \9688 , \9689 );
and \U$8882 ( \9691 , \9325 , \9374 );
nor \U$8883 ( \9692 , \9690 , \9691 );
xor \U$8884 ( \9693 , \9687 , \9692 );
not \U$8885 ( \9694 , \9510 );
nor \U$8886 ( \9695 , \9694 , \9495 );
not \U$8887 ( \9696 , \9695 );
not \U$8888 ( \9697 , \9508 );
and \U$8889 ( \9698 , \9696 , \9697 );
and \U$8890 ( \9699 , \9695 , \9508 );
nor \U$8891 ( \9700 , \9698 , \9699 );
and \U$8892 ( \9701 , \9693 , \9700 );
and \U$8893 ( \9702 , \9687 , \9692 );
or \U$8894 ( \9703 , \9701 , \9702 );
xor \U$8895 ( \9704 , \9536 , \9703 );
nand \U$8896 ( \9705 , \9018_nG29b3 , \8767 );
or \U$8897 ( \9706 , \8624 , \9260_nG28b3 );
nand \U$8898 ( \9707 , \9706 , \8773 );
and \U$8899 ( \9708 , \9705 , \9707 );
and \U$8900 ( \9709 , \8769 , \9260_nG28b3 );
and \U$8901 ( \9710 , \9018_nG29b3 , \8831 );
nor \U$8902 ( \9711 , \9708 , \9709 , \9710 );
and \U$8903 ( \9712 , \8947_nG2a93 , \8890 );
or \U$8904 ( \9713 , \8816 , \8868_nG2b9c );
nand \U$8905 ( \9714 , \9713 , \9026 );
nand \U$8906 ( \9715 , \8947_nG2a93 , \8887 );
and \U$8907 ( \9716 , \9714 , \9715 );
and \U$8908 ( \9717 , \8868_nG2b9c , \9030 );
nor \U$8909 ( \9718 , \9712 , \9716 , \9717 );
xor \U$8910 ( \9719 , \9711 , \9718 );
nand \U$8911 ( \9720 , \9481_nG2706 , \8580 );
or \U$8912 ( \9721 , \8540 , \9317_nG27da );
nand \U$8913 ( \9722 , \9721 , \8615 );
and \U$8914 ( \9723 , \9720 , \9722 );
and \U$8915 ( \9724 , \8610 , \9317_nG27da );
and \U$8916 ( \9725 , \9481_nG2706 , \8583 );
nor \U$8917 ( \9726 , \9723 , \9724 , \9725 );
and \U$8918 ( \9727 , \9719 , \9726 );
and \U$8919 ( \9728 , \9711 , \9718 );
or \U$8920 ( \9729 , \9727 , \9728 );
nand \U$8921 ( \9730 , \8657_nG2e7a , \9331 );
or \U$8922 ( \9731 , \9204 , \8568_nG2f9c );
nand \U$8923 ( \9732 , \9731 , \9427 );
and \U$8924 ( \9733 , \9730 , \9732 );
and \U$8925 ( \9734 , \9430 , \8568_nG2f9c );
and \U$8926 ( \9735 , \8657_nG2e7a , \9333 );
nor \U$8927 ( \9736 , \9733 , \9734 , \9735 );
not \U$8928 ( \9737 , \9614 );
and \U$8929 ( \9738 , \8516 , \9737 );
and \U$8930 ( \9739 , \9612 , \8475 );
nand \U$8931 ( \9740 , \9611 , \9198 );
not \U$8932 ( \9741 , \9740 );
and \U$8933 ( \9742 , \8514_nG31b0 , \9741 );
nor \U$8934 ( \9743 , \9738 , \9739 , \9742 );
xor \U$8935 ( \9744 , \9736 , \9743 );
and \U$8936 ( \9745 , \8729_nG2d90 , \9188 );
or \U$8937 ( \9746 , \9048 , \8729_nG2d90 );
nand \U$8938 ( \9747 , \9746 , \9191 );
nand \U$8939 ( \9748 , \8762_nG2c8f , \9091 );
and \U$8940 ( \9749 , \9747 , \9748 );
and \U$8941 ( \9750 , \8762_nG2c8f , \9094 );
nor \U$8942 ( \9751 , \9745 , \9749 , \9750 );
and \U$8943 ( \9752 , \9744 , \9751 );
and \U$8944 ( \9753 , \9736 , \9743 );
or \U$8945 ( \9754 , \9752 , \9753 );
nor \U$8946 ( \9755 , \9729 , \9754 );
xor \U$8947 ( \9756 , \9406 , \9413 );
xor \U$8948 ( \9757 , \9756 , \9421 );
not \U$8949 ( \9758 , \9757 );
and \U$8950 ( \9759 , \9755 , \9758 );
not \U$8951 ( \9760 , \9755 );
not \U$8952 ( \9761 , \9758 );
and \U$8953 ( \9762 , \9760 , \9761 );
xor \U$8954 ( \9763 , \9582 , \9589 );
xor \U$8955 ( \9764 , \9763 , \9597 );
not \U$8956 ( \9765 , \9764 );
not \U$8957 ( \9766 , \9661 );
nor \U$8958 ( \9767 , \9632 , \9664 );
not \U$8959 ( \9768 , \9767 );
or \U$8960 ( \9769 , \9766 , \9768 );
or \U$8961 ( \9770 , \9767 , \9661 );
nand \U$8962 ( \9771 , \9769 , \9770 );
nand \U$8963 ( \9772 , \9765 , \9771 );
nor \U$8964 ( \9773 , \9762 , \9772 );
nor \U$8965 ( \9774 , \9759 , \9773 );
xor \U$8966 ( \9775 , \9433 , \9199 );
xor \U$8967 ( \9776 , \9775 , \9441 );
xor \U$8968 ( \9777 , \9600 , \9616 );
xor \U$8969 ( \9778 , \9777 , \9665 );
nand \U$8970 ( \9779 , \9776 , \9778 );
and \U$8971 ( \9780 , \9779 , \9572 );
nor \U$8972 ( \9781 , \9778 , \9776 );
nor \U$8973 ( \9782 , \9780 , \9781 );
and \U$8974 ( \9783 , \9774 , \9782 );
xor \U$8975 ( \9784 , \9448 , \9453 );
xor \U$8976 ( \9785 , \9784 , \9490 );
xor \U$8977 ( \9786 , \9572 , \9668 );
xor \U$8978 ( \9787 , \9785 , \9786 );
not \U$8979 ( \9788 , \9787 );
or \U$8980 ( \9789 , \9571 , \9564 );
not \U$8981 ( \9790 , \9444 );
or \U$8982 ( \9791 , \9790 , \9424 );
not \U$8983 ( \9792 , \9424 );
or \U$8984 ( \9793 , \9444 , \9792 );
nand \U$8985 ( \9794 , \9789 , \9791 , \9793 );
nand \U$8986 ( \9795 , \9788 , \9794 );
xor \U$8987 ( \9796 , \9783 , \9795 );
xor \U$8988 ( \9797 , \9673 , \9678 );
xor \U$8989 ( \9798 , \9797 , \9684 );
and \U$8990 ( \9799 , \9796 , \9798 );
and \U$8991 ( \9800 , \9783 , \9795 );
or \U$8992 ( \9801 , \9799 , \9800 );
xor \U$8993 ( \9802 , \9687 , \9692 );
xor \U$8994 ( \9803 , \9802 , \9700 );
and \U$8995 ( \9804 , \9801 , \9803 );
not \U$8996 ( \9805 , \9607 );
not \U$8997 ( \9806 , \9615 );
and \U$8998 ( \9807 , \9805 , \9806 );
and \U$8999 ( \9808 , \9607 , \9615 );
nor \U$9000 ( \9809 , \9807 , \9808 );
and \U$9001 ( \9810 , \9018_nG29b3 , \8890 );
or \U$9002 ( \9811 , \8816 , \8947_nG2a93 );
nand \U$9003 ( \9812 , \9811 , \9026 );
nand \U$9004 ( \9813 , \9018_nG29b3 , \8887 );
and \U$9005 ( \9814 , \9812 , \9813 );
and \U$9006 ( \9815 , \8947_nG2a93 , \9030 );
nor \U$9007 ( \9816 , \9810 , \9814 , \9815 );
and \U$9008 ( \9817 , \8762_nG2c8f , \9188 );
or \U$9009 ( \9818 , \9048 , \8762_nG2c8f );
nand \U$9010 ( \9819 , \9818 , \9191 );
nand \U$9011 ( \9820 , \8868_nG2b9c , \9091 );
and \U$9012 ( \9821 , \9819 , \9820 );
and \U$9013 ( \9822 , \8868_nG2b9c , \9094 );
nor \U$9014 ( \9823 , \9817 , \9821 , \9822 );
xor \U$9015 ( \9824 , \9816 , \9823 );
nand \U$9016 ( \9825 , \9260_nG28b3 , \8767 );
or \U$9017 ( \9826 , \8624 , \9317_nG27da );
nand \U$9018 ( \9827 , \9826 , \8773 );
and \U$9019 ( \9828 , \9825 , \9827 );
and \U$9020 ( \9829 , \8769 , \9317_nG27da );
and \U$9021 ( \9830 , \9260_nG28b3 , \8831 );
nor \U$9022 ( \9831 , \9828 , \9829 , \9830 );
and \U$9023 ( \9832 , \9824 , \9831 );
and \U$9024 ( \9833 , \9816 , \9823 );
or \U$9025 ( \9834 , \9832 , \9833 );
nand \U$9026 ( \9835 , \9563_nG23ac , \8580 );
or \U$9027 ( \9836 , \8540 , \9481_nG2706 );
nand \U$9028 ( \9837 , \9836 , \8615 );
and \U$9029 ( \9838 , \9835 , \9837 );
and \U$9030 ( \9839 , \8610 , \9481_nG2706 );
and \U$9031 ( \9840 , \9563_nG23ac , \8583 );
nor \U$9032 ( \9841 , \9838 , \9839 , \9840 );
and \U$9033 ( \9842 , RIaaa59d8_486, \7919 );
and \U$9034 ( \9843 , RIaaa60e0_501, \7944 );
and \U$9035 ( \9844 , \7924 , RIaaa5f00_497);
and \U$9036 ( \9845 , RIaaa5f78_498, \7930 );
nor \U$9037 ( \9846 , \9844 , \9845 );
and \U$9038 ( \9847 , \7961 , RIaaa5ac8_488);
and \U$9039 ( \9848 , RIaaa5ca8_492, \7963 );
nor \U$9040 ( \9849 , \9847 , \9848 );
and \U$9041 ( \9850 , \8454 , RIaaa5e88_496);
and \U$9042 ( \9851 , RIaaa5ff0_499, \7935 );
nor \U$9043 ( \9852 , \9850 , \9851 );
and \U$9044 ( \9853 , \7928 , RIaaa5d20_493);
and \U$9045 ( \9854 , RIaaa6158_502, \7909 );
nor \U$9046 ( \9855 , \9853 , \9854 );
nand \U$9047 ( \9856 , \9846 , \9849 , \9852 , \9855 );
nor \U$9048 ( \9857 , \9842 , \9843 , \9856 );
and \U$9049 ( \9858 , \7942 , RIaaa5b40_489);
and \U$9050 ( \9859 , RIaaa5bb8_490, \7957 );
nor \U$9051 ( \9860 , \9858 , \9859 );
and \U$9052 ( \9861 , \7914 , RIaaa5e10_495);
and \U$9053 ( \9862 , RIaaa6068_500, \7952 );
nor \U$9054 ( \9863 , \9861 , \9862 );
and \U$9055 ( \9864 , \7949 , RIaaa5c30_491);
and \U$9056 ( \9865 , RIaaa5a50_487, \7959 );
nor \U$9057 ( \9866 , \9864 , \9865 );
nand \U$9058 ( \9867 , \9857 , \9860 , \9863 , \9866 );
_DC g2303 ( \9868_nG2303 , \9867 , \8473 );
nand \U$9059 ( \9869 , \9868_nG2303 , \8444 );
xor \U$9060 ( \9870 , \9841 , \9869 );
and \U$9061 ( \9871 , \9660_nG2373 , \8629 );
and \U$9062 ( \9872 , RIaaa4e20_461, \7959 );
and \U$9063 ( \9873 , RIaaa4e98_462, \7919 );
and \U$9064 ( \9874 , \7924 , RIaaa4c40_457);
and \U$9065 ( \9875 , RIaaa4cb8_458, \7930 );
nor \U$9066 ( \9876 , \9874 , \9875 );
and \U$9067 ( \9877 , \8454 , RIaaa4bc8_456);
and \U$9068 ( \9878 , RIaaa5000_465, \7957 );
nor \U$9069 ( \9879 , \9877 , \9878 );
and \U$9070 ( \9880 , \7928 , RIaaa4a60_453);
and \U$9071 ( \9881 , RIaaa4d30_459, \7935 );
nor \U$9072 ( \9882 , \9880 , \9881 );
and \U$9073 ( \9883 , \7961 , RIaaa4f10_463);
and \U$9074 ( \9884 , RIaaa49e8_452, \7963 );
nor \U$9075 ( \9885 , \9883 , \9884 );
nand \U$9076 ( \9886 , \9876 , \9879 , \9882 , \9885 );
nor \U$9077 ( \9887 , \9872 , \9873 , \9886 );
and \U$9078 ( \9888 , \7949 , RIaaa5078_466);
and \U$9079 ( \9889 , RIaaa4da8_460, \7952 );
nor \U$9080 ( \9890 , \9888 , \9889 );
and \U$9081 ( \9891 , \7914 , RIaaa4b50_455);
and \U$9082 ( \9892 , RIaaa4f88_464, \7942 );
nor \U$9083 ( \9893 , \9891 , \9892 );
and \U$9084 ( \9894 , \7944 , RIaaa50f0_467);
and \U$9085 ( \9895 , RIaaa5168_468, \7909 );
nor \U$9086 ( \9896 , \9894 , \9895 );
nand \U$9087 ( \9897 , \9887 , \9890 , \9893 , \9896 );
_DC g233b ( \9898_nG233b , \9897 , \8473 );
or \U$9088 ( \9899 , \8487 , \9898_nG233b );
nand \U$9089 ( \9900 , \9899 , \8524 );
nand \U$9090 ( \9901 , \9660_nG2373 , \8520 );
and \U$9091 ( \9902 , \9900 , \9901 );
and \U$9092 ( \9903 , \9898_nG233b , \8662 );
nor \U$9093 ( \9904 , \9871 , \9902 , \9903 );
and \U$9094 ( \9905 , \9870 , \9904 );
and \U$9095 ( \9906 , \9841 , \9869 );
or \U$9096 ( \9907 , \9905 , \9906 );
nand \U$9097 ( \9908 , \9834 , \9907 );
or \U$9098 ( \9909 , \9740 , \8475 );
or \U$9099 ( \9910 , \8474_nG30a2 , \9614 );
or \U$9100 ( \9911 , \8568_nG2f9c , \9613 );
nand \U$9101 ( \9912 , \9909 , \9910 , \9911 );
not \U$9102 ( \9913 , \9912 );
nand \U$9103 ( \9914 , \8729_nG2d90 , \9331 );
or \U$9104 ( \9915 , \9204 , \8657_nG2e7a );
nand \U$9105 ( \9916 , \9915 , \9427 );
and \U$9106 ( \9917 , \9914 , \9916 );
and \U$9107 ( \9918 , \9430 , \8657_nG2e7a );
and \U$9108 ( \9919 , \8729_nG2d90 , \9333 );
nor \U$9109 ( \9920 , \9917 , \9918 , \9919 );
nor \U$9110 ( \9921 , \9913 , \9920 );
and \U$9111 ( \9922 , \9908 , \9921 );
nor \U$9112 ( \9923 , \9907 , \9834 );
nor \U$9113 ( \9924 , \9922 , \9923 );
nand \U$9114 ( \9925 , \9809 , \9924 );
nand \U$9115 ( \9926 , \9898_nG233b , \8444 );
and \U$9116 ( \9927 , \9563_nG23ac , \8629 );
or \U$9117 ( \9928 , \8487 , \9660_nG2373 );
nand \U$9118 ( \9929 , \9928 , \8524 );
nand \U$9119 ( \9930 , \9563_nG23ac , \8520 );
and \U$9120 ( \9931 , \9929 , \9930 );
and \U$9121 ( \9932 , \9660_nG2373 , \8662 );
nor \U$9122 ( \9933 , \9927 , \9931 , \9932 );
xor \U$9123 ( \9934 , \9926 , \9933 );
not \U$9124 ( \9935 , \9934 );
xor \U$9125 ( \9936 , \9711 , \9718 );
xor \U$9126 ( \9937 , \9936 , \9726 );
nor \U$9127 ( \9938 , \9935 , \9937 );
and \U$9128 ( \9939 , \9925 , \9938 );
nor \U$9129 ( \9940 , \9924 , \9809 );
nor \U$9130 ( \9941 , \9939 , \9940 );
not \U$9131 ( \9942 , \9941 );
not \U$9132 ( \9943 , \9572 );
not \U$9133 ( \9944 , \9781 );
nand \U$9134 ( \9945 , \9944 , \9779 );
not \U$9135 ( \9946 , \9945 );
or \U$9136 ( \9947 , \9943 , \9946 );
or \U$9137 ( \9948 , \9945 , \9572 );
nand \U$9138 ( \9949 , \9947 , \9948 );
nand \U$9139 ( \9950 , \9942 , \9949 );
not \U$9140 ( \9951 , \9950 );
not \U$9141 ( \9952 , \9941 );
nor \U$9142 ( \9953 , \9952 , \9949 );
nor \U$9143 ( \9954 , \9951 , \9953 );
not \U$9144 ( \9955 , \9954 );
not \U$9145 ( \9956 , \9771 );
not \U$9146 ( \9957 , \9764 );
and \U$9147 ( \9958 , \9956 , \9957 );
and \U$9148 ( \9959 , \9771 , \9764 );
nor \U$9149 ( \9960 , \9958 , \9959 );
not \U$9150 ( \9961 , \9960 );
or \U$9151 ( \9962 , \9933 , \9926 );
not \U$9152 ( \9963 , \9754 );
or \U$9153 ( \9964 , \9963 , \9729 );
not \U$9154 ( \9965 , \9729 );
or \U$9155 ( \9966 , \9754 , \9965 );
nand \U$9156 ( \9967 , \9962 , \9964 , \9966 );
nand \U$9157 ( \9968 , \9961 , \9967 );
not \U$9158 ( \9969 , \9968 );
and \U$9159 ( \9970 , \9955 , \9969 );
and \U$9160 ( \9971 , \9954 , \9968 );
nor \U$9161 ( \9972 , \9970 , \9971 );
not \U$9162 ( \9973 , \9757 );
not \U$9163 ( \9974 , \9755 );
not \U$9164 ( \9975 , \9772 );
or \U$9165 ( \9976 , \9974 , \9975 );
or \U$9166 ( \9977 , \9772 , \9755 );
nand \U$9167 ( \9978 , \9976 , \9977 );
not \U$9168 ( \9979 , \9978 );
or \U$9169 ( \9980 , \9973 , \9979 );
or \U$9170 ( \9981 , \9978 , \9757 );
nand \U$9171 ( \9982 , \9980 , \9981 );
not \U$9172 ( \9983 , \9967 );
not \U$9173 ( \9984 , \9960 );
or \U$9174 ( \9985 , \9983 , \9984 );
or \U$9175 ( \9986 , \9960 , \9967 );
nand \U$9176 ( \9987 , \9985 , \9986 );
not \U$9177 ( \9988 , \9987 );
xor \U$9178 ( \9989 , \9736 , \9743 );
xor \U$9179 ( \9990 , \9989 , \9751 );
not \U$9180 ( \9991 , \9990 );
nand \U$9181 ( \9992 , \9317_nG27da , \8767 );
or \U$9182 ( \9993 , \8624 , \9481_nG2706 );
nand \U$9183 ( \9994 , \9993 , \8773 );
and \U$9184 ( \9995 , \9992 , \9994 );
and \U$9185 ( \9996 , \8769 , \9481_nG2706 );
and \U$9186 ( \9997 , \9317_nG27da , \8831 );
nor \U$9187 ( \9998 , \9995 , \9996 , \9997 );
and \U$9188 ( \9999 , \9260_nG28b3 , \8890 );
or \U$9189 ( \10000 , \8816 , \9018_nG29b3 );
nand \U$9190 ( \10001 , \10000 , \9026 );
nand \U$9191 ( \10002 , \9260_nG28b3 , \8887 );
and \U$9192 ( \10003 , \10001 , \10002 );
and \U$9193 ( \10004 , \9018_nG29b3 , \9030 );
nor \U$9194 ( \10005 , \9999 , \10003 , \10004 );
xor \U$9195 ( \10006 , \9998 , \10005 );
nand \U$9196 ( \10007 , \9660_nG2373 , \8580 );
or \U$9197 ( \10008 , \8540 , \9563_nG23ac );
nand \U$9198 ( \10009 , \10008 , \8615 );
and \U$9199 ( \10010 , \10007 , \10009 );
and \U$9200 ( \10011 , \8610 , \9563_nG23ac );
and \U$9201 ( \10012 , \9660_nG2373 , \8583 );
nor \U$9202 ( \10013 , \10010 , \10011 , \10012 );
and \U$9203 ( \10014 , \10006 , \10013 );
and \U$9204 ( \10015 , \9998 , \10005 );
or \U$9205 ( \10016 , \10014 , \10015 );
nand \U$9206 ( \10017 , \8762_nG2c8f , \9331 );
or \U$9207 ( \10018 , \9204 , \8729_nG2d90 );
nand \U$9208 ( \10019 , \10018 , \9427 );
and \U$9209 ( \10020 , \10017 , \10019 );
and \U$9210 ( \10021 , \9430 , \8729_nG2d90 );
and \U$9211 ( \10022 , \8762_nG2c8f , \9333 );
nor \U$9212 ( \10023 , \10020 , \10021 , \10022 );
and \U$9213 ( \10024 , \8590 , \9737 );
not \U$9214 ( \10025 , \8657_nG2e7a );
and \U$9215 ( \10026 , \9612 , \10025 );
and \U$9216 ( \10027 , \8568_nG2f9c , \9741 );
nor \U$9217 ( \10028 , \10024 , \10026 , \10027 );
xor \U$9218 ( \10029 , \10023 , \10028 );
and \U$9219 ( \10030 , \8868_nG2b9c , \9188 );
or \U$9220 ( \10031 , \9048 , \8868_nG2b9c );
nand \U$9221 ( \10032 , \10031 , \9191 );
nand \U$9222 ( \10033 , \8947_nG2a93 , \9091 );
and \U$9223 ( \10034 , \10032 , \10033 );
and \U$9224 ( \10035 , \8947_nG2a93 , \9094 );
nor \U$9225 ( \10036 , \10030 , \10034 , \10035 );
and \U$9226 ( \10037 , \10029 , \10036 );
and \U$9227 ( \10038 , \10023 , \10028 );
or \U$9228 ( \10039 , \10037 , \10038 );
nor \U$9229 ( \10040 , \10016 , \10039 );
nand \U$9230 ( \10041 , \9991 , \10040 );
or \U$9231 ( \10042 , \9988 , \10041 );
not \U$9232 ( \10043 , \10041 );
not \U$9233 ( \10044 , \9988 );
or \U$9234 ( \10045 , \10043 , \10044 );
not \U$9235 ( \10046 , \9938 );
not \U$9236 ( \10047 , \9940 );
nand \U$9237 ( \10048 , \10047 , \9925 );
not \U$9238 ( \10049 , \10048 );
or \U$9239 ( \10050 , \10046 , \10049 );
or \U$9240 ( \10051 , \10048 , \9938 );
nand \U$9241 ( \10052 , \10050 , \10051 );
nand \U$9242 ( \10053 , \10045 , \10052 );
nand \U$9243 ( \10054 , \10042 , \10053 );
nand \U$9244 ( \10055 , \9982 , \10054 );
and \U$9245 ( \10056 , \9972 , \10055 );
nor \U$9246 ( \10057 , \10054 , \9982 );
nor \U$9247 ( \10058 , \10056 , \10057 );
not \U$9248 ( \10059 , \9787 );
not \U$9249 ( \10060 , \9794 );
and \U$9250 ( \10061 , \10059 , \10060 );
and \U$9251 ( \10062 , \9787 , \9794 );
nor \U$9252 ( \10063 , \10061 , \10062 );
xor \U$9253 ( \10064 , \9774 , \9782 );
nand \U$9254 ( \10065 , \10063 , \10064 );
not \U$9255 ( \10066 , \10065 );
nor \U$9256 ( \10067 , \10064 , \10063 );
nor \U$9257 ( \10068 , \10066 , \10067 );
not \U$9258 ( \10069 , \10068 );
or \U$9259 ( \10070 , \9953 , \9968 );
nand \U$9260 ( \10071 , \10070 , \9950 );
not \U$9261 ( \10072 , \10071 );
and \U$9262 ( \10073 , \10069 , \10072 );
and \U$9263 ( \10074 , \10068 , \10071 );
nor \U$9264 ( \10075 , \10073 , \10074 );
xor \U$9265 ( \10076 , \10058 , \10075 );
not \U$9266 ( \10077 , \9972 );
not \U$9267 ( \10078 , \10057 );
nand \U$9268 ( \10079 , \10078 , \10055 );
not \U$9269 ( \10080 , \10079 );
or \U$9270 ( \10081 , \10077 , \10080 );
or \U$9271 ( \10082 , \10079 , \9972 );
nand \U$9272 ( \10083 , \10081 , \10082 );
not \U$9273 ( \10084 , \10016 );
and \U$9274 ( \10085 , \10084 , \10039 );
and \U$9275 ( \10086 , \9898_nG233b , \8629 );
or \U$9276 ( \10087 , \8487 , \9868_nG2303 );
nand \U$9277 ( \10088 , \10087 , \8524 );
nand \U$9278 ( \10089 , \9898_nG233b , \8520 );
and \U$9279 ( \10090 , \10088 , \10089 );
and \U$9280 ( \10091 , \9868_nG2303 , \8662 );
nor \U$9281 ( \10092 , \10086 , \10090 , \10091 );
and \U$9282 ( \10093 , RIaaa6c20_525, \7957 );
and \U$9283 ( \10094 , RIaaa69c8_520, \7942 );
and \U$9284 ( \10095 , \7924 , RIaaa70d0_535);
and \U$9285 ( \10096 , RIaaa6d10_527, \7930 );
nor \U$9286 ( \10097 , \10095 , \10096 );
and \U$9287 ( \10098 , \7961 , RIaaa6a40_521);
and \U$9288 ( \10099 , RIaaa6ef0_531, \7963 );
nor \U$9289 ( \10100 , \10098 , \10099 );
and \U$9290 ( \10101 , \8454 , RIaaa7058_534);
and \U$9291 ( \10102 , RIaaa6c98_526, \7935 );
nor \U$9292 ( \10103 , \10101 , \10102 );
and \U$9293 ( \10104 , \7928 , RIaaa6f68_532);
and \U$9294 ( \10105 , RIaaa6e00_529, \7909 );
nor \U$9295 ( \10106 , \10104 , \10105 );
nand \U$9296 ( \10107 , \10097 , \10100 , \10103 , \10106 );
nor \U$9297 ( \10108 , \10093 , \10094 , \10107 );
and \U$9298 ( \10109 , \7949 , RIaaa6ba8_524);
and \U$9299 ( \10110 , RIaaa6e78_530, \7952 );
nor \U$9300 ( \10111 , \10109 , \10110 );
and \U$9301 ( \10112 , \7914 , RIaaa6fe0_533);
and \U$9302 ( \10113 , RIaaa6ab8_522, \7959 );
nor \U$9303 ( \10114 , \10112 , \10113 );
and \U$9304 ( \10115 , \7919 , RIaaa6b30_523);
and \U$9305 ( \10116 , RIaaa6d88_528, \7944 );
nor \U$9306 ( \10117 , \10115 , \10116 );
nand \U$9307 ( \10118 , \10108 , \10111 , \10114 , \10117 );
_DC g22ca ( \10119_nG22ca , \10118 , \8473 );
nand \U$9308 ( \10120 , \10119_nG22ca , \8444 );
or \U$9309 ( \10121 , \10092 , \10120 );
or \U$9310 ( \10122 , \10039 , \10084 );
nand \U$9311 ( \10123 , \10121 , \10122 );
nor \U$9312 ( \10124 , \10085 , \10123 );
not \U$9313 ( \10125 , \9920 );
not \U$9314 ( \10126 , \9912 );
and \U$9315 ( \10127 , \10125 , \10126 );
and \U$9316 ( \10128 , \9920 , \9912 );
nor \U$9317 ( \10129 , \10127 , \10128 );
xor \U$9318 ( \10130 , \10124 , \10129 );
xor \U$9319 ( \10131 , \9841 , \9869 );
xor \U$9320 ( \10132 , \10131 , \9904 );
and \U$9321 ( \10133 , \10130 , \10132 );
and \U$9322 ( \10134 , \10124 , \10129 );
or \U$9323 ( \10135 , \10133 , \10134 );
not \U$9324 ( \10136 , \9934 );
not \U$9325 ( \10137 , \9937 );
and \U$9326 ( \10138 , \10136 , \10137 );
and \U$9327 ( \10139 , \9934 , \9937 );
nor \U$9328 ( \10140 , \10138 , \10139 );
xor \U$9329 ( \10141 , \10135 , \10140 );
xor \U$9330 ( \10142 , \9998 , \10005 );
xor \U$9331 ( \10143 , \10142 , \10013 );
xor \U$9332 ( \10144 , \10023 , \10028 );
xor \U$9333 ( \10145 , \10144 , \10036 );
xor \U$9334 ( \10146 , \10143 , \10145 );
xnor \U$9335 ( \10147 , \10120 , \10092 );
and \U$9336 ( \10148 , \10146 , \10147 );
and \U$9337 ( \10149 , \10143 , \10145 );
or \U$9338 ( \10150 , \10148 , \10149 );
xor \U$9339 ( \10151 , \9816 , \9823 );
xor \U$9340 ( \10152 , \10151 , \9831 );
xor \U$9341 ( \10153 , \10150 , \10152 );
and \U$9342 ( \10154 , \9317_nG27da , \8890 );
or \U$9343 ( \10155 , \8816 , \9260_nG28b3 );
nand \U$9344 ( \10156 , \10155 , \9026 );
nand \U$9345 ( \10157 , \9317_nG27da , \8887 );
and \U$9346 ( \10158 , \10156 , \10157 );
and \U$9347 ( \10159 , \9260_nG28b3 , \9030 );
nor \U$9348 ( \10160 , \10154 , \10158 , \10159 );
and \U$9349 ( \10161 , \8947_nG2a93 , \9188 );
or \U$9350 ( \10162 , \9048 , \8947_nG2a93 );
nand \U$9351 ( \10163 , \10162 , \9191 );
nand \U$9352 ( \10164 , \9018_nG29b3 , \9091 );
and \U$9353 ( \10165 , \10163 , \10164 );
and \U$9354 ( \10166 , \9018_nG29b3 , \9094 );
nor \U$9355 ( \10167 , \10161 , \10165 , \10166 );
xor \U$9356 ( \10168 , \10160 , \10167 );
nand \U$9357 ( \10169 , \9481_nG2706 , \8767 );
or \U$9358 ( \10170 , \8624 , \9563_nG23ac );
nand \U$9359 ( \10171 , \10170 , \8773 );
and \U$9360 ( \10172 , \10169 , \10171 );
and \U$9361 ( \10173 , \8769 , \9563_nG23ac );
and \U$9362 ( \10174 , \9481_nG2706 , \8831 );
nor \U$9363 ( \10175 , \10172 , \10173 , \10174 );
and \U$9364 ( \10176 , \10168 , \10175 );
and \U$9365 ( \10177 , \10160 , \10167 );
or \U$9366 ( \10178 , \10176 , \10177 );
nand \U$9367 ( \10179 , \8868_nG2b9c , \9331 );
or \U$9368 ( \10180 , \9204 , \8762_nG2c8f );
nand \U$9369 ( \10181 , \10180 , \9427 );
and \U$9370 ( \10182 , \10179 , \10181 );
and \U$9371 ( \10183 , \9430 , \8762_nG2c8f );
and \U$9372 ( \10184 , \8868_nG2b9c , \9333 );
nor \U$9373 ( \10185 , \10182 , \10183 , \10184 );
not \U$9374 ( \10186 , \10185 );
or \U$9375 ( \10187 , \9740 , \10025 );
or \U$9376 ( \10188 , \8657_nG2e7a , \9614 );
or \U$9377 ( \10189 , \8729_nG2d90 , \9613 );
nand \U$9378 ( \10190 , \10187 , \10188 , \10189 );
nand \U$9379 ( \10191 , \10186 , \10190 );
xor \U$9380 ( \10192 , \10178 , \10191 );
and \U$9381 ( \10193 , \9868_nG2303 , \8629 );
or \U$9382 ( \10194 , \8487 , \10119_nG22ca );
nand \U$9383 ( \10195 , \10194 , \8524 );
nand \U$9384 ( \10196 , \9868_nG2303 , \8520 );
and \U$9385 ( \10197 , \10195 , \10196 );
and \U$9386 ( \10198 , \10119_nG22ca , \8662 );
nor \U$9387 ( \10199 , \10193 , \10197 , \10198 );
nand \U$9388 ( \10200 , \9898_nG233b , \8580 );
or \U$9389 ( \10201 , \8540 , \9660_nG2373 );
nand \U$9390 ( \10202 , \10201 , \8615 );
and \U$9391 ( \10203 , \10200 , \10202 );
and \U$9392 ( \10204 , \8610 , \9660_nG2373 );
and \U$9393 ( \10205 , \9898_nG233b , \8583 );
nor \U$9394 ( \10206 , \10203 , \10204 , \10205 );
and \U$9395 ( \10207 , \10199 , \10206 );
not \U$9396 ( \10208 , \10207 );
and \U$9397 ( \10209 , RIaaa7328_540, \7924 );
and \U$9398 ( \10210 , RIaaa76e8_548, \7935 );
and \U$9399 ( \10211 , \7952 , RIaaa7508_544);
and \U$9400 ( \10212 , RIaaa73a0_541, \7957 );
nor \U$9401 ( \10213 , \10211 , \10212 );
and \U$9402 ( \10214 , \7942 , RIaaa7490_543);
and \U$9403 ( \10215 , RIaaa75f8_546, \7919 );
nor \U$9404 ( \10216 , \10214 , \10215 );
and \U$9405 ( \10217 , \7914 , RIaaa7238_538);
and \U$9406 ( \10218 , RIaaa7418_542, \7949 );
nor \U$9407 ( \10219 , \10217 , \10218 );
and \U$9408 ( \10220 , \7959 , RIaaa7670_547);
and \U$9409 ( \10221 , RIaaa77d8_550, \7944 );
nor \U$9410 ( \10222 , \10220 , \10221 );
nand \U$9411 ( \10223 , \10213 , \10216 , \10219 , \10222 );
nor \U$9412 ( \10224 , \10209 , \10210 , \10223 );
and \U$9413 ( \10225 , \8454 , RIaaa72b0_539);
and \U$9414 ( \10226 , RIaaa78c8_552, \7963 );
nor \U$9415 ( \10227 , \10225 , \10226 );
and \U$9416 ( \10228 , \7928 , RIaaa7940_553);
and \U$9417 ( \10229 , RIaaa7760_549, \7930 );
nor \U$9418 ( \10230 , \10228 , \10229 );
and \U$9419 ( \10231 , \7961 , RIaaa7580_545);
and \U$9420 ( \10232 , RIaaa7850_551, \7909 );
nor \U$9421 ( \10233 , \10231 , \10232 );
nand \U$9422 ( \10234 , \10224 , \10227 , \10230 , \10233 );
_DC g228e ( \10235_nG228e , \10234 , \8473 );
nand \U$9423 ( \10236 , \10235_nG228e , \8444 );
not \U$9424 ( \10237 , \10236 );
and \U$9425 ( \10238 , \10208 , \10237 );
nor \U$9426 ( \10239 , \10199 , \10206 );
nor \U$9427 ( \10240 , \10238 , \10239 );
and \U$9428 ( \10241 , \10192 , \10240 );
and \U$9429 ( \10242 , \10178 , \10191 );
or \U$9430 ( \10243 , \10241 , \10242 );
and \U$9431 ( \10244 , \10153 , \10243 );
and \U$9432 ( \10245 , \10150 , \10152 );
or \U$9433 ( \10246 , \10244 , \10245 );
and \U$9434 ( \10247 , \10141 , \10246 );
and \U$9435 ( \10248 , \10135 , \10140 );
or \U$9436 ( \10249 , \10247 , \10248 );
not \U$9437 ( \10250 , \10040 );
not \U$9438 ( \10251 , \9990 );
and \U$9439 ( \10252 , \10250 , \10251 );
and \U$9440 ( \10253 , \10040 , \9990 );
nor \U$9441 ( \10254 , \10252 , \10253 );
not \U$9442 ( \10255 , \10254 );
not \U$9443 ( \10256 , \9921 );
not \U$9444 ( \10257 , \9923 );
nand \U$9445 ( \10258 , \10257 , \9908 );
not \U$9446 ( \10259 , \10258 );
or \U$9447 ( \10260 , \10256 , \10259 );
or \U$9448 ( \10261 , \10258 , \9921 );
nand \U$9449 ( \10262 , \10260 , \10261 );
nand \U$9450 ( \10263 , \10255 , \10262 );
xor \U$9451 ( \10264 , \10249 , \10263 );
not \U$9452 ( \10265 , \10052 );
not \U$9453 ( \10266 , \10041 );
and \U$9454 ( \10267 , \10265 , \10266 );
and \U$9455 ( \10268 , \10052 , \10041 );
nor \U$9456 ( \10269 , \10267 , \10268 );
not \U$9457 ( \10270 , \10269 );
not \U$9458 ( \10271 , \9987 );
and \U$9459 ( \10272 , \10270 , \10271 );
and \U$9460 ( \10273 , \10269 , \9987 );
nor \U$9461 ( \10274 , \10272 , \10273 );
and \U$9462 ( \10275 , \10264 , \10274 );
and \U$9463 ( \10276 , \10249 , \10263 );
or \U$9464 ( \10277 , \10275 , \10276 );
xor \U$9465 ( \10278 , \10083 , \10277 );
xor \U$9466 ( \10279 , \10160 , \10167 );
xor \U$9467 ( \10280 , \10279 , \10175 );
not \U$9468 ( \10281 , \10280 );
not \U$9469 ( \10282 , \10236 );
nor \U$9470 ( \10283 , \10207 , \10239 );
not \U$9471 ( \10284 , \10283 );
or \U$9472 ( \10285 , \10282 , \10284 );
or \U$9473 ( \10286 , \10283 , \10236 );
nand \U$9474 ( \10287 , \10285 , \10286 );
nand \U$9475 ( \10288 , \10281 , \10287 );
nand \U$9476 ( \10289 , \8947_nG2a93 , \9331 );
or \U$9477 ( \10290 , \9204 , \8868_nG2b9c );
nand \U$9478 ( \10291 , \10290 , \9427 );
and \U$9479 ( \10292 , \10289 , \10291 );
and \U$9480 ( \10293 , \9430 , \8868_nG2b9c );
and \U$9481 ( \10294 , \8947_nG2a93 , \9333 );
nor \U$9482 ( \10295 , \10292 , \10293 , \10294 );
and \U$9483 ( \10296 , \8785 , \9737 );
and \U$9484 ( \10297 , \9612 , \8872 );
and \U$9485 ( \10298 , \8729_nG2d90 , \9741 );
nor \U$9486 ( \10299 , \10296 , \10297 , \10298 );
xor \U$9487 ( \10300 , \10295 , \10299 );
and \U$9488 ( \10301 , \9018_nG29b3 , \9188 );
or \U$9489 ( \10302 , \9048 , \9018_nG29b3 );
nand \U$9490 ( \10303 , \10302 , \9191 );
nand \U$9491 ( \10304 , \9260_nG28b3 , \9091 );
and \U$9492 ( \10305 , \10303 , \10304 );
and \U$9493 ( \10306 , \9260_nG28b3 , \9094 );
nor \U$9494 ( \10307 , \10301 , \10305 , \10306 );
and \U$9495 ( \10308 , \10300 , \10307 );
and \U$9496 ( \10309 , \10295 , \10299 );
or \U$9497 ( \10310 , \10308 , \10309 );
not \U$9498 ( \10311 , \10310 );
nand \U$9499 ( \10312 , \9563_nG23ac , \8767 );
or \U$9500 ( \10313 , \8624 , \9660_nG2373 );
nand \U$9501 ( \10314 , \10313 , \8773 );
and \U$9502 ( \10315 , \10312 , \10314 );
and \U$9503 ( \10316 , \8769 , \9660_nG2373 );
and \U$9504 ( \10317 , \9563_nG23ac , \8831 );
nor \U$9505 ( \10318 , \10315 , \10316 , \10317 );
and \U$9506 ( \10319 , \9481_nG2706 , \8890 );
or \U$9507 ( \10320 , \8816 , \9317_nG27da );
nand \U$9508 ( \10321 , \10320 , \9026 );
nand \U$9509 ( \10322 , \9481_nG2706 , \8887 );
and \U$9510 ( \10323 , \10321 , \10322 );
and \U$9511 ( \10324 , \9317_nG27da , \9030 );
nor \U$9512 ( \10325 , \10319 , \10323 , \10324 );
xor \U$9513 ( \10326 , \10318 , \10325 );
nand \U$9514 ( \10327 , \9868_nG2303 , \8580 );
or \U$9515 ( \10328 , \8540 , \9898_nG233b );
nand \U$9516 ( \10329 , \10328 , \8615 );
and \U$9517 ( \10330 , \10327 , \10329 );
and \U$9518 ( \10331 , \8610 , \9898_nG233b );
and \U$9519 ( \10332 , \9868_nG2303 , \8583 );
nor \U$9520 ( \10333 , \10330 , \10331 , \10332 );
and \U$9521 ( \10334 , \10326 , \10333 );
and \U$9522 ( \10335 , \10318 , \10325 );
or \U$9523 ( \10336 , \10334 , \10335 );
not \U$9524 ( \10337 , \10336 );
nand \U$9525 ( \10338 , \10311 , \10337 );
xor \U$9526 ( \10339 , \10288 , \10338 );
xor \U$9527 ( \10340 , \10143 , \10145 );
xor \U$9528 ( \10341 , \10340 , \10147 );
and \U$9529 ( \10342 , \10339 , \10341 );
and \U$9530 ( \10343 , \10288 , \10338 );
or \U$9531 ( \10344 , \10342 , \10343 );
xor \U$9532 ( \10345 , \10124 , \10129 );
xor \U$9533 ( \10346 , \10345 , \10132 );
xor \U$9534 ( \10347 , \10344 , \10346 );
xor \U$9535 ( \10348 , \10150 , \10152 );
xor \U$9536 ( \10349 , \10348 , \10243 );
and \U$9537 ( \10350 , \10347 , \10349 );
and \U$9538 ( \10351 , \10344 , \10346 );
or \U$9539 ( \10352 , \10350 , \10351 );
not \U$9540 ( \10353 , \10262 );
not \U$9541 ( \10354 , \10254 );
and \U$9542 ( \10355 , \10353 , \10354 );
and \U$9543 ( \10356 , \10262 , \10254 );
nor \U$9544 ( \10357 , \10355 , \10356 );
nor \U$9545 ( \10358 , \10352 , \10357 );
and \U$9546 ( \10359 , \10352 , \10357 );
or \U$9547 ( \10360 , \10358 , \10359 );
not \U$9548 ( \10361 , \10360 );
xor \U$9549 ( \10362 , \10135 , \10140 );
xor \U$9550 ( \10363 , \10362 , \10246 );
not \U$9551 ( \10364 , \10363 );
and \U$9552 ( \10365 , \10361 , \10364 );
and \U$9553 ( \10366 , \10360 , \10363 );
nor \U$9554 ( \10367 , \10365 , \10366 );
xor \U$9555 ( \10368 , \10344 , \10346 );
xor \U$9556 ( \10369 , \10368 , \10349 );
not \U$9557 ( \10370 , \10287 );
not \U$9558 ( \10371 , \10280 );
and \U$9559 ( \10372 , \10370 , \10371 );
and \U$9560 ( \10373 , \10287 , \10280 );
nor \U$9561 ( \10374 , \10372 , \10373 );
not \U$9562 ( \10375 , \10374 );
and \U$9563 ( \10376 , \10119_nG22ca , \8629 );
or \U$9564 ( \10377 , \8487 , \10235_nG228e );
nand \U$9565 ( \10378 , \10377 , \8524 );
nand \U$9566 ( \10379 , \10119_nG22ca , \8520 );
and \U$9567 ( \10380 , \10378 , \10379 );
and \U$9568 ( \10381 , \10235_nG228e , \8662 );
nor \U$9569 ( \10382 , \10376 , \10380 , \10381 );
and \U$9570 ( \10383 , RIaaa85e8_580, \7919 );
and \U$9571 ( \10384 , RIaaa87c8_584, \7944 );
and \U$9572 ( \10385 , \7924 , RIaaa8318_574);
and \U$9573 ( \10386 , RIaaa8750_583, \7930 );
nor \U$9574 ( \10387 , \10385 , \10386 );
and \U$9575 ( \10388 , \7961 , RIaaa8570_579);
and \U$9576 ( \10389 , RIaaa88b8_586, \7963 );
nor \U$9577 ( \10390 , \10388 , \10389 );
and \U$9578 ( \10391 , \8454 , RIaaa82a0_573);
and \U$9579 ( \10392 , RIaaa86d8_582, \7935 );
nor \U$9580 ( \10393 , \10391 , \10392 );
and \U$9581 ( \10394 , \7928 , RIaaa8930_587);
and \U$9582 ( \10395 , RIaaa8840_585, \7909 );
nor \U$9583 ( \10396 , \10394 , \10395 );
nand \U$9584 ( \10397 , \10387 , \10390 , \10393 , \10396 );
nor \U$9585 ( \10398 , \10383 , \10384 , \10397 );
and \U$9586 ( \10399 , \7942 , RIaaa8408_576);
and \U$9587 ( \10400 , RIaaa8390_575, \7957 );
nor \U$9588 ( \10401 , \10399 , \10400 );
and \U$9589 ( \10402 , \7914 , RIaaa8228_572);
and \U$9590 ( \10403 , RIaaa84f8_578, \7952 );
nor \U$9591 ( \10404 , \10402 , \10403 );
and \U$9592 ( \10405 , \7949 , RIaaa8480_577);
and \U$9593 ( \10406 , RIaaa8660_581, \7959 );
nor \U$9594 ( \10407 , \10405 , \10406 );
nand \U$9595 ( \10408 , \10398 , \10401 , \10404 , \10407 );
_DC g225a ( \10409_nG225a , \10408 , \8473 );
nand \U$9596 ( \10410 , \10409_nG225a , \8444 );
or \U$9597 ( \10411 , \10382 , \10410 );
or \U$9598 ( \10412 , \10311 , \10336 );
or \U$9599 ( \10413 , \10310 , \10337 );
nand \U$9600 ( \10414 , \10411 , \10412 , \10413 );
nand \U$9601 ( \10415 , \10375 , \10414 );
xor \U$9602 ( \10416 , \10178 , \10191 );
xor \U$9603 ( \10417 , \10416 , \10240 );
xor \U$9604 ( \10418 , \10415 , \10417 );
xor \U$9605 ( \10419 , \10318 , \10325 );
xor \U$9606 ( \10420 , \10419 , \10333 );
xor \U$9607 ( \10421 , \10295 , \10299 );
xor \U$9608 ( \10422 , \10421 , \10307 );
xor \U$9609 ( \10423 , \10420 , \10422 );
xnor \U$9610 ( \10424 , \10410 , \10382 );
and \U$9611 ( \10425 , \10423 , \10424 );
and \U$9612 ( \10426 , \10420 , \10422 );
or \U$9613 ( \10427 , \10425 , \10426 );
not \U$9614 ( \10428 , \10185 );
not \U$9615 ( \10429 , \10190 );
and \U$9616 ( \10430 , \10428 , \10429 );
and \U$9617 ( \10431 , \10185 , \10190 );
nor \U$9618 ( \10432 , \10430 , \10431 );
xor \U$9619 ( \10433 , \10427 , \10432 );
and \U$9620 ( \10434 , \9563_nG23ac , \8890 );
or \U$9621 ( \10435 , \8816 , \9481_nG2706 );
nand \U$9622 ( \10436 , \10435 , \9026 );
nand \U$9623 ( \10437 , \9563_nG23ac , \8887 );
and \U$9624 ( \10438 , \10436 , \10437 );
and \U$9625 ( \10439 , \9481_nG2706 , \9030 );
nor \U$9626 ( \10440 , \10434 , \10438 , \10439 );
and \U$9627 ( \10441 , \9260_nG28b3 , \9188 );
or \U$9628 ( \10442 , \9048 , \9260_nG28b3 );
nand \U$9629 ( \10443 , \10442 , \9191 );
nand \U$9630 ( \10444 , \9317_nG27da , \9091 );
and \U$9631 ( \10445 , \10443 , \10444 );
and \U$9632 ( \10446 , \9317_nG27da , \9094 );
nor \U$9633 ( \10447 , \10441 , \10445 , \10446 );
xor \U$9634 ( \10448 , \10440 , \10447 );
nand \U$9635 ( \10449 , \9660_nG2373 , \8767 );
or \U$9636 ( \10450 , \8624 , \9898_nG233b );
nand \U$9637 ( \10451 , \10450 , \8773 );
and \U$9638 ( \10452 , \10449 , \10451 );
and \U$9639 ( \10453 , \8769 , \9898_nG233b );
and \U$9640 ( \10454 , \9660_nG2373 , \8831 );
nor \U$9641 ( \10455 , \10452 , \10453 , \10454 );
and \U$9642 ( \10456 , \10448 , \10455 );
and \U$9643 ( \10457 , \10440 , \10447 );
or \U$9644 ( \10458 , \10456 , \10457 );
nand \U$9645 ( \10459 , \9018_nG29b3 , \9331 );
or \U$9646 ( \10460 , \9204 , \8947_nG2a93 );
nand \U$9647 ( \10461 , \10460 , \9427 );
and \U$9648 ( \10462 , \10459 , \10461 );
and \U$9649 ( \10463 , \9430 , \8947_nG2a93 );
and \U$9650 ( \10464 , \9018_nG29b3 , \9333 );
nor \U$9651 ( \10465 , \10462 , \10463 , \10464 );
not \U$9652 ( \10466 , \10465 );
or \U$9653 ( \10467 , \9740 , \8872 );
or \U$9654 ( \10468 , \8762_nG2c8f , \9614 );
or \U$9655 ( \10469 , \8868_nG2b9c , \9613 );
nand \U$9656 ( \10470 , \10467 , \10468 , \10469 );
nand \U$9657 ( \10471 , \10466 , \10470 );
xor \U$9658 ( \10472 , \10458 , \10471 );
nand \U$9659 ( \10473 , \10119_nG22ca , \8580 );
or \U$9660 ( \10474 , \8540 , \9868_nG2303 );
nand \U$9661 ( \10475 , \10474 , \8615 );
and \U$9662 ( \10476 , \10473 , \10475 );
and \U$9663 ( \10477 , \8610 , \9868_nG2303 );
and \U$9664 ( \10478 , \10119_nG22ca , \8583 );
nor \U$9665 ( \10479 , \10476 , \10477 , \10478 );
and \U$9666 ( \10480 , RIaaa7df0_563, \7924 );
and \U$9667 ( \10481 , RIaaa7f58_566, \7935 );
and \U$9668 ( \10482 , \7959 , RIaaa7a30_555);
and \U$9669 ( \10483 , RIaaa80c0_569, \7944 );
nor \U$9670 ( \10484 , \10482 , \10483 );
and \U$9671 ( \10485 , \7914 , RIaaa7d78_562);
and \U$9672 ( \10486 , RIaaa7b98_558, \7957 );
nor \U$9673 ( \10487 , \10485 , \10486 );
and \U$9674 ( \10488 , \7942 , RIaaa7aa8_556);
and \U$9675 ( \10489 , RIaaa79b8_554, \7919 );
nor \U$9676 ( \10490 , \10488 , \10489 );
and \U$9677 ( \10491 , \7949 , RIaaa7c10_559);
and \U$9678 ( \10492 , RIaaa8048_568, \7952 );
nor \U$9679 ( \10493 , \10491 , \10492 );
nand \U$9680 ( \10494 , \10484 , \10487 , \10490 , \10493 );
nor \U$9681 ( \10495 , \10480 , \10481 , \10494 );
and \U$9682 ( \10496 , \8454 , RIaaa7e68_564);
and \U$9683 ( \10497 , RIaaa8138_570, \7909 );
nor \U$9684 ( \10498 , \10496 , \10497 );
and \U$9685 ( \10499 , \7961 , RIaaa7b20_557);
and \U$9686 ( \10500 , RIaaa7fd0_567, \7930 );
nor \U$9687 ( \10501 , \10499 , \10500 );
and \U$9688 ( \10502 , \7928 , RIaaa7c88_560);
and \U$9689 ( \10503 , RIaaa7d00_561, \7963 );
nor \U$9690 ( \10504 , \10502 , \10503 );
nand \U$9691 ( \10505 , \10495 , \10498 , \10501 , \10504 );
_DC g221a ( \10506_nG221a , \10505 , \8473 );
nand \U$9692 ( \10507 , \10506_nG221a , \8444 );
xor \U$9693 ( \10508 , \10479 , \10507 );
and \U$9694 ( \10509 , \10235_nG228e , \8629 );
or \U$9695 ( \10510 , \8487 , \10409_nG225a );
nand \U$9696 ( \10511 , \10510 , \8524 );
nand \U$9697 ( \10512 , \10235_nG228e , \8520 );
and \U$9698 ( \10513 , \10511 , \10512 );
and \U$9699 ( \10514 , \10409_nG225a , \8662 );
nor \U$9700 ( \10515 , \10509 , \10513 , \10514 );
and \U$9701 ( \10516 , \10508 , \10515 );
and \U$9702 ( \10517 , \10479 , \10507 );
or \U$9703 ( \10518 , \10516 , \10517 );
and \U$9704 ( \10519 , \10472 , \10518 );
and \U$9705 ( \10520 , \10458 , \10471 );
or \U$9706 ( \10521 , \10519 , \10520 );
and \U$9707 ( \10522 , \10433 , \10521 );
and \U$9708 ( \10523 , \10427 , \10432 );
or \U$9709 ( \10524 , \10522 , \10523 );
and \U$9710 ( \10525 , \10418 , \10524 );
and \U$9711 ( \10526 , \10415 , \10417 );
or \U$9712 ( \10527 , \10525 , \10526 );
nor \U$9713 ( \10528 , \10369 , \10527 );
xor \U$9714 ( \10529 , \10367 , \10528 );
and \U$9715 ( \10530 , \10369 , \10527 );
nor \U$9716 ( \10531 , \10530 , \10528 );
xor \U$9717 ( \10532 , \10415 , \10417 );
xor \U$9718 ( \10533 , \10532 , \10524 );
xor \U$9719 ( \10534 , \10288 , \10338 );
xor \U$9720 ( \10535 , \10534 , \10341 );
nor \U$9721 ( \10536 , \10533 , \10535 );
xor \U$9722 ( \10537 , \10531 , \10536 );
and \U$9723 ( \10538 , \10533 , \10535 );
nor \U$9724 ( \10539 , \10538 , \10536 );
nand \U$9725 ( \10540 , \9898_nG233b , \8767 );
or \U$9726 ( \10541 , \8624 , \9868_nG2303 );
nand \U$9727 ( \10542 , \10541 , \8773 );
and \U$9728 ( \10543 , \10540 , \10542 );
and \U$9729 ( \10544 , \8769 , \9868_nG2303 );
and \U$9730 ( \10545 , \9898_nG233b , \8831 );
nor \U$9731 ( \10546 , \10543 , \10544 , \10545 );
and \U$9732 ( \10547 , \9660_nG2373 , \8890 );
or \U$9733 ( \10548 , \8816 , \9563_nG23ac );
nand \U$9734 ( \10549 , \10548 , \9026 );
nand \U$9735 ( \10550 , \9660_nG2373 , \8887 );
and \U$9736 ( \10551 , \10549 , \10550 );
and \U$9737 ( \10552 , \9563_nG23ac , \9030 );
nor \U$9738 ( \10553 , \10547 , \10551 , \10552 );
xor \U$9739 ( \10554 , \10546 , \10553 );
nand \U$9740 ( \10555 , \10235_nG228e , \8580 );
or \U$9741 ( \10556 , \8540 , \10119_nG22ca );
nand \U$9742 ( \10557 , \10556 , \8615 );
and \U$9743 ( \10558 , \10555 , \10557 );
and \U$9744 ( \10559 , \8610 , \10119_nG22ca );
and \U$9745 ( \10560 , \10235_nG228e , \8583 );
nor \U$9746 ( \10561 , \10558 , \10559 , \10560 );
and \U$9747 ( \10562 , \10554 , \10561 );
and \U$9748 ( \10563 , \10546 , \10553 );
or \U$9749 ( \10564 , \10562 , \10563 );
nand \U$9750 ( \10565 , \9260_nG28b3 , \9331 );
or \U$9751 ( \10566 , \9204 , \9018_nG29b3 );
nand \U$9752 ( \10567 , \10566 , \9427 );
and \U$9753 ( \10568 , \10565 , \10567 );
and \U$9754 ( \10569 , \9430 , \9018_nG29b3 );
and \U$9755 ( \10570 , \9260_nG28b3 , \9333 );
nor \U$9756 ( \10571 , \10568 , \10569 , \10570 );
and \U$9757 ( \10572 , \8869 , \9737 );
and \U$9758 ( \10573 , \9612 , \9109 );
and \U$9759 ( \10574 , \8868_nG2b9c , \9741 );
nor \U$9760 ( \10575 , \10572 , \10573 , \10574 );
xor \U$9761 ( \10576 , \10571 , \10575 );
and \U$9762 ( \10577 , \9317_nG27da , \9188 );
or \U$9763 ( \10578 , \9048 , \9317_nG27da );
nand \U$9764 ( \10579 , \10578 , \9191 );
nand \U$9765 ( \10580 , \9481_nG2706 , \9091 );
and \U$9766 ( \10581 , \10579 , \10580 );
and \U$9767 ( \10582 , \9481_nG2706 , \9094 );
nor \U$9768 ( \10583 , \10577 , \10581 , \10582 );
and \U$9769 ( \10584 , \10576 , \10583 );
and \U$9770 ( \10585 , \10571 , \10575 );
or \U$9771 ( \10586 , \10584 , \10585 );
xor \U$9772 ( \10587 , \10564 , \10586 );
xor \U$9773 ( \10588 , \10479 , \10507 );
xor \U$9774 ( \10589 , \10588 , \10515 );
and \U$9775 ( \10590 , \10587 , \10589 );
and \U$9776 ( \10591 , \10564 , \10586 );
or \U$9777 ( \10592 , \10590 , \10591 );
xor \U$9778 ( \10593 , \10440 , \10447 );
xor \U$9779 ( \10594 , \10593 , \10455 );
not \U$9780 ( \10595 , \10594 );
not \U$9781 ( \10596 , \10470 );
not \U$9782 ( \10597 , \10465 );
or \U$9783 ( \10598 , \10596 , \10597 );
or \U$9784 ( \10599 , \10465 , \10470 );
nand \U$9785 ( \10600 , \10598 , \10599 );
nand \U$9786 ( \10601 , \10595 , \10600 );
xor \U$9787 ( \10602 , \10592 , \10601 );
xor \U$9788 ( \10603 , \10420 , \10422 );
xor \U$9789 ( \10604 , \10603 , \10424 );
and \U$9790 ( \10605 , \10602 , \10604 );
and \U$9791 ( \10606 , \10592 , \10601 );
or \U$9792 ( \10607 , \10605 , \10606 );
not \U$9793 ( \10608 , \10374 );
not \U$9794 ( \10609 , \10414 );
and \U$9795 ( \10610 , \10608 , \10609 );
and \U$9796 ( \10611 , \10374 , \10414 );
nor \U$9797 ( \10612 , \10610 , \10611 );
xor \U$9798 ( \10613 , \10607 , \10612 );
xor \U$9799 ( \10614 , \10427 , \10432 );
xor \U$9800 ( \10615 , \10614 , \10521 );
and \U$9801 ( \10616 , \10613 , \10615 );
and \U$9802 ( \10617 , \10607 , \10612 );
or \U$9803 ( \10618 , \10616 , \10617 );
not \U$9804 ( \10619 , \10618 );
xor \U$9805 ( \10620 , \10539 , \10619 );
nand \U$9806 ( \10621 , \9317_nG27da , \9331 );
or \U$9807 ( \10622 , \9204 , \9260_nG28b3 );
nand \U$9808 ( \10623 , \10622 , \9427 );
and \U$9809 ( \10624 , \10621 , \10623 );
and \U$9810 ( \10625 , \9430 , \9260_nG28b3 );
and \U$9811 ( \10626 , \9317_nG27da , \9333 );
nor \U$9812 ( \10627 , \10624 , \10625 , \10626 );
and \U$9813 ( \10628 , \9109 , \9737 );
and \U$9814 ( \10629 , \9612 , \9111 );
and \U$9815 ( \10630 , \8947_nG2a93 , \9741 );
nor \U$9816 ( \10631 , \10628 , \10629 , \10630 );
xor \U$9817 ( \10632 , \10627 , \10631 );
and \U$9818 ( \10633 , \10632 , \8487 );
and \U$9819 ( \10634 , \10627 , \10631 );
or \U$9820 ( \10635 , \10633 , \10634 );
and \U$9821 ( \10636 , \9898_nG233b , \8890 );
or \U$9822 ( \10637 , \8816 , \9660_nG2373 );
nand \U$9823 ( \10638 , \10637 , \9026 );
nand \U$9824 ( \10639 , \9898_nG233b , \8887 );
and \U$9825 ( \10640 , \10638 , \10639 );
and \U$9826 ( \10641 , \9660_nG2373 , \9030 );
nor \U$9827 ( \10642 , \10636 , \10640 , \10641 );
and \U$9828 ( \10643 , \9481_nG2706 , \9188 );
or \U$9829 ( \10644 , \9048 , \9481_nG2706 );
nand \U$9830 ( \10645 , \10644 , \9191 );
nand \U$9831 ( \10646 , \9563_nG23ac , \9091 );
and \U$9832 ( \10647 , \10645 , \10646 );
and \U$9833 ( \10648 , \9563_nG23ac , \9094 );
nor \U$9834 ( \10649 , \10643 , \10647 , \10648 );
xor \U$9835 ( \10650 , \10642 , \10649 );
nand \U$9836 ( \10651 , \9868_nG2303 , \8767 );
or \U$9837 ( \10652 , \8624 , \10119_nG22ca );
nand \U$9838 ( \10653 , \10652 , \8773 );
and \U$9839 ( \10654 , \10651 , \10653 );
and \U$9840 ( \10655 , \8769 , \10119_nG22ca );
and \U$9841 ( \10656 , \9868_nG2303 , \8831 );
nor \U$9842 ( \10657 , \10654 , \10655 , \10656 );
and \U$9843 ( \10658 , \10650 , \10657 );
and \U$9844 ( \10659 , \10642 , \10649 );
or \U$9845 ( \10660 , \10658 , \10659 );
xor \U$9846 ( \10661 , \10635 , \10660 );
and \U$9847 ( \10662 , \10409_nG225a , \8629 );
or \U$9848 ( \10663 , \8487 , \10506_nG221a );
nand \U$9849 ( \10664 , \10663 , \8524 );
nand \U$9850 ( \10665 , \10409_nG225a , \8520 );
and \U$9851 ( \10666 , \10664 , \10665 );
and \U$9852 ( \10667 , \10506_nG221a , \8662 );
nor \U$9853 ( \10668 , \10662 , \10666 , \10667 );
and \U$9854 ( \10669 , \10661 , \10668 );
and \U$9855 ( \10670 , \10635 , \10660 );
or \U$9856 ( \10671 , \10669 , \10670 );
not \U$9857 ( \10672 , \10594 );
not \U$9858 ( \10673 , \10600 );
and \U$9859 ( \10674 , \10672 , \10673 );
and \U$9860 ( \10675 , \10594 , \10600 );
nor \U$9861 ( \10676 , \10674 , \10675 );
xor \U$9862 ( \10677 , \10671 , \10676 );
xor \U$9863 ( \10678 , \10564 , \10586 );
xor \U$9864 ( \10679 , \10678 , \10589 );
and \U$9865 ( \10680 , \10677 , \10679 );
and \U$9866 ( \10681 , \10671 , \10676 );
or \U$9867 ( \10682 , \10680 , \10681 );
xor \U$9868 ( \10683 , \10458 , \10471 );
xor \U$9869 ( \10684 , \10683 , \10518 );
xor \U$9870 ( \10685 , \10682 , \10684 );
xor \U$9871 ( \10686 , \10592 , \10601 );
xor \U$9872 ( \10687 , \10686 , \10604 );
and \U$9873 ( \10688 , \10685 , \10687 );
and \U$9874 ( \10689 , \10682 , \10684 );
or \U$9875 ( \10690 , \10688 , \10689 );
xor \U$9876 ( \10691 , \10607 , \10612 );
xor \U$9877 ( \10692 , \10691 , \10615 );
and \U$9878 ( \10693 , \10690 , \10692 );
xor \U$9879 ( \10694 , \10635 , \10660 );
xor \U$9880 ( \10695 , \10694 , \10668 );
xor \U$9881 ( \10696 , \10571 , \10575 );
xor \U$9882 ( \10697 , \10696 , \10583 );
or \U$9883 ( \10698 , \10695 , \10697 );
nand \U$9884 ( \10699 , \10409_nG225a , \8580 );
or \U$9885 ( \10700 , \8540 , \10235_nG228e );
nand \U$9886 ( \10701 , \10700 , \8615 );
and \U$9887 ( \10702 , \10699 , \10701 );
and \U$9888 ( \10703 , \8610 , \10235_nG228e );
and \U$9889 ( \10704 , \10409_nG225a , \8583 );
nor \U$9890 ( \10705 , \10702 , \10703 , \10704 );
nand \U$9891 ( \10706 , \9481_nG2706 , \9331 );
or \U$9892 ( \10707 , \9204 , \9317_nG27da );
nand \U$9893 ( \10708 , \10707 , \9427 );
and \U$9894 ( \10709 , \10706 , \10708 );
and \U$9895 ( \10710 , \9430 , \9317_nG27da );
and \U$9896 ( \10711 , \9481_nG2706 , \9333 );
nor \U$9897 ( \10712 , \10709 , \10710 , \10711 );
and \U$9898 ( \10713 , \9111 , \9737 );
not \U$9899 ( \10714 , \9260_nG28b3 );
and \U$9900 ( \10715 , \9612 , \10714 );
and \U$9901 ( \10716 , \9018_nG29b3 , \9741 );
nor \U$9902 ( \10717 , \10713 , \10715 , \10716 );
xor \U$9903 ( \10718 , \10712 , \10717 );
and \U$9904 ( \10719 , \9563_nG23ac , \9188 );
or \U$9905 ( \10720 , \9048 , \9563_nG23ac );
nand \U$9906 ( \10721 , \10720 , \9191 );
nand \U$9907 ( \10722 , \9660_nG2373 , \9091 );
and \U$9908 ( \10723 , \10721 , \10722 );
and \U$9909 ( \10724 , \9660_nG2373 , \9094 );
nor \U$9910 ( \10725 , \10719 , \10723 , \10724 );
and \U$9911 ( \10726 , \10718 , \10725 );
and \U$9912 ( \10727 , \10712 , \10717 );
or \U$9913 ( \10728 , \10726 , \10727 );
xor \U$9914 ( \10729 , \10705 , \10728 );
nand \U$9915 ( \10730 , \10119_nG22ca , \8767 );
or \U$9916 ( \10731 , \8624 , \10235_nG228e );
nand \U$9917 ( \10732 , \10731 , \8773 );
and \U$9918 ( \10733 , \10730 , \10732 );
and \U$9919 ( \10734 , \8769 , \10235_nG228e );
and \U$9920 ( \10735 , \10119_nG22ca , \8831 );
nor \U$9921 ( \10736 , \10733 , \10734 , \10735 );
and \U$9922 ( \10737 , \9868_nG2303 , \8890 );
or \U$9923 ( \10738 , \8816 , \9898_nG233b );
nand \U$9924 ( \10739 , \10738 , \9026 );
nand \U$9925 ( \10740 , \9868_nG2303 , \8887 );
and \U$9926 ( \10741 , \10739 , \10740 );
and \U$9927 ( \10742 , \9898_nG233b , \9030 );
nor \U$9928 ( \10743 , \10737 , \10741 , \10742 );
xor \U$9929 ( \10744 , \10736 , \10743 );
nand \U$9930 ( \10745 , \10506_nG221a , \8580 );
or \U$9931 ( \10746 , \8540 , \10409_nG225a );
nand \U$9932 ( \10747 , \10746 , \8615 );
and \U$9933 ( \10748 , \10745 , \10747 );
and \U$9934 ( \10749 , \8610 , \10409_nG225a );
and \U$9935 ( \10750 , \10506_nG221a , \8583 );
nor \U$9936 ( \10751 , \10748 , \10749 , \10750 );
and \U$9937 ( \10752 , \10744 , \10751 );
and \U$9938 ( \10753 , \10736 , \10743 );
or \U$9939 ( \10754 , \10752 , \10753 );
and \U$9940 ( \10755 , \10729 , \10754 );
and \U$9941 ( \10756 , \10705 , \10728 );
or \U$9942 ( \10757 , \10755 , \10756 );
xor \U$9943 ( \10758 , \10546 , \10553 );
xor \U$9944 ( \10759 , \10758 , \10561 );
xor \U$9945 ( \10760 , \10757 , \10759 );
xor \U$9946 ( \10761 , \10642 , \10649 );
xor \U$9947 ( \10762 , \10761 , \10657 );
xor \U$9948 ( \10763 , \10627 , \10631 );
xor \U$9949 ( \10764 , \10763 , \8487 );
and \U$9950 ( \10765 , \10762 , \10764 );
nand \U$9951 ( \10766 , \10506_nG221a , \8520 );
and \U$9952 ( \10767 , \8486 , \10766 );
and \U$9953 ( \10768 , \10506_nG221a , \8629 );
nor \U$9954 ( \10769 , \10767 , \10768 );
xor \U$9955 ( \10770 , \10627 , \10631 );
xor \U$9956 ( \10771 , \10770 , \8487 );
and \U$9957 ( \10772 , \10769 , \10771 );
and \U$9958 ( \10773 , \10762 , \10769 );
or \U$9959 ( \10774 , \10765 , \10772 , \10773 );
and \U$9960 ( \10775 , \10760 , \10774 );
and \U$9961 ( \10776 , \10757 , \10759 );
or \U$9962 ( \10777 , \10775 , \10776 );
xor \U$9963 ( \10778 , \10698 , \10777 );
xor \U$9964 ( \10779 , \10671 , \10676 );
xor \U$9965 ( \10780 , \10779 , \10679 );
and \U$9966 ( \10781 , \10778 , \10780 );
and \U$9967 ( \10782 , \10698 , \10777 );
or \U$9968 ( \10783 , \10781 , \10782 );
xor \U$9969 ( \10784 , \10682 , \10684 );
xor \U$9970 ( \10785 , \10784 , \10687 );
and \U$9971 ( \10786 , \10783 , \10785 );
and \U$9972 ( \10787 , \10119_nG22ca , \8890 );
or \U$9973 ( \10788 , \8816 , \9868_nG2303 );
nand \U$9974 ( \10789 , \10788 , \9026 );
nand \U$9975 ( \10790 , \10119_nG22ca , \8887 );
and \U$9976 ( \10791 , \10789 , \10790 );
and \U$9977 ( \10792 , \9868_nG2303 , \9030 );
nor \U$9978 ( \10793 , \10787 , \10791 , \10792 );
and \U$9979 ( \10794 , \9660_nG2373 , \9188 );
or \U$9980 ( \10795 , \9048 , \9660_nG2373 );
nand \U$9981 ( \10796 , \10795 , \9191 );
nand \U$9982 ( \10797 , \9898_nG233b , \9091 );
and \U$9983 ( \10798 , \10796 , \10797 );
and \U$9984 ( \10799 , \9898_nG233b , \9094 );
nor \U$9985 ( \10800 , \10794 , \10798 , \10799 );
xor \U$9986 ( \10801 , \10793 , \10800 );
nand \U$9987 ( \10802 , \10235_nG228e , \8767 );
or \U$9988 ( \10803 , \8624 , \10409_nG225a );
nand \U$9989 ( \10804 , \10803 , \8773 );
and \U$9990 ( \10805 , \10802 , \10804 );
and \U$9991 ( \10806 , \8769 , \10409_nG225a );
and \U$9992 ( \10807 , \10235_nG228e , \8831 );
nor \U$9993 ( \10808 , \10805 , \10806 , \10807 );
and \U$9994 ( \10809 , \10801 , \10808 );
and \U$9995 ( \10810 , \10793 , \10800 );
or \U$9996 ( \10811 , \10809 , \10810 );
nand \U$9997 ( \10812 , \9563_nG23ac , \9331 );
or \U$9998 ( \10813 , \9204 , \9481_nG2706 );
nand \U$9999 ( \10814 , \10813 , \9427 );
and \U$10000 ( \10815 , \10812 , \10814 );
and \U$10001 ( \10816 , \9430 , \9481_nG2706 );
and \U$10002 ( \10817 , \9563_nG23ac , \9333 );
nor \U$10003 ( \10818 , \10815 , \10816 , \10817 );
and \U$10004 ( \10819 , \10714 , \9737 );
not \U$10005 ( \10820 , \9317_nG27da );
and \U$10006 ( \10821 , \9612 , \10820 );
and \U$10007 ( \10822 , \9260_nG28b3 , \9741 );
nor \U$10008 ( \10823 , \10819 , \10821 , \10822 );
xor \U$10009 ( \10824 , \10818 , \10823 );
and \U$10010 ( \10825 , \10824 , \8540 );
and \U$10011 ( \10826 , \10818 , \10823 );
or \U$10012 ( \10827 , \10825 , \10826 );
xor \U$10013 ( \10828 , \10811 , \10827 );
xor \U$10014 ( \10829 , \10736 , \10743 );
xor \U$10015 ( \10830 , \10829 , \10751 );
and \U$10016 ( \10831 , \10828 , \10830 );
and \U$10017 ( \10832 , \10811 , \10827 );
or \U$10018 ( \10833 , \10831 , \10832 );
xor \U$10019 ( \10834 , \10705 , \10728 );
xor \U$10020 ( \10835 , \10834 , \10754 );
xor \U$10021 ( \10836 , \10833 , \10835 );
xor \U$10022 ( \10837 , \10627 , \10631 );
xor \U$10023 ( \10838 , \10837 , \8487 );
xor \U$10024 ( \10839 , \10762 , \10769 );
xor \U$10025 ( \10840 , \10838 , \10839 );
and \U$10026 ( \10841 , \10836 , \10840 );
and \U$10027 ( \10842 , \10833 , \10835 );
or \U$10028 ( \10843 , \10841 , \10842 );
xor \U$10029 ( \10844 , \10757 , \10759 );
xor \U$10030 ( \10845 , \10844 , \10774 );
xor \U$10031 ( \10846 , \10843 , \10845 );
xnor \U$10032 ( \10847 , \10697 , \10695 );
xor \U$10033 ( \10848 , \10846 , \10847 );
not \U$10034 ( \10849 , \10848 );
xor \U$10035 ( \10850 , \10833 , \10835 );
xor \U$10036 ( \10851 , \10850 , \10840 );
nand \U$10037 ( \10852 , \9660_nG2373 , \9331 );
or \U$10038 ( \10853 , \9204 , \9563_nG23ac );
nand \U$10039 ( \10854 , \10853 , \9427 );
and \U$10040 ( \10855 , \10852 , \10854 );
and \U$10041 ( \10856 , \9430 , \9563_nG23ac );
and \U$10042 ( \10857 , \9660_nG2373 , \9333 );
nor \U$10043 ( \10858 , \10855 , \10856 , \10857 );
and \U$10044 ( \10859 , \10820 , \9737 );
not \U$10045 ( \10860 , \9481_nG2706 );
and \U$10046 ( \10861 , \9612 , \10860 );
and \U$10047 ( \10862 , \9317_nG27da , \9741 );
nor \U$10048 ( \10863 , \10859 , \10861 , \10862 );
xor \U$10049 ( \10864 , \10858 , \10863 );
and \U$10050 ( \10865 , \9898_nG233b , \9188 );
or \U$10051 ( \10866 , \9048 , \9898_nG233b );
nand \U$10052 ( \10867 , \10866 , \9191 );
nand \U$10053 ( \10868 , \9868_nG2303 , \9091 );
and \U$10054 ( \10869 , \10867 , \10868 );
and \U$10055 ( \10870 , \9868_nG2303 , \9094 );
nor \U$10056 ( \10871 , \10865 , \10869 , \10870 );
and \U$10057 ( \10872 , \10864 , \10871 );
and \U$10058 ( \10873 , \10858 , \10863 );
or \U$10059 ( \10874 , \10872 , \10873 );
xor \U$10060 ( \10875 , \10793 , \10800 );
xor \U$10061 ( \10876 , \10875 , \10808 );
and \U$10062 ( \10877 , \10874 , \10876 );
and \U$10063 ( \10878 , \10506_nG221a , \8610 );
not \U$10064 ( \10879 , \10506_nG221a );
and \U$10065 ( \10880 , \10879 , \8582 );
not \U$10066 ( \10881 , \8615 );
nor \U$10067 ( \10882 , \10878 , \10880 , \10881 );
xor \U$10068 ( \10883 , \10793 , \10800 );
xor \U$10069 ( \10884 , \10883 , \10808 );
and \U$10070 ( \10885 , \10882 , \10884 );
and \U$10071 ( \10886 , \10874 , \10882 );
or \U$10072 ( \10887 , \10877 , \10885 , \10886 );
xor \U$10073 ( \10888 , \10712 , \10717 );
xor \U$10074 ( \10889 , \10888 , \10725 );
xor \U$10075 ( \10890 , \10887 , \10889 );
xor \U$10076 ( \10891 , \10811 , \10827 );
xor \U$10077 ( \10892 , \10891 , \10830 );
and \U$10078 ( \10893 , \10890 , \10892 );
and \U$10079 ( \10894 , \10887 , \10889 );
or \U$10080 ( \10895 , \10893 , \10894 );
nor \U$10081 ( \10896 , \10851 , \10895 );
xor \U$10082 ( \10897 , \10849 , \10896 );
and \U$10083 ( \10898 , \10851 , \10895 );
nor \U$10084 ( \10899 , \10898 , \10896 );
xor \U$10085 ( \10900 , \10887 , \10889 );
xor \U$10086 ( \10901 , \10900 , \10892 );
xor \U$10087 ( \10902 , \10818 , \10823 );
xor \U$10088 ( \10903 , \10902 , \8540 );
nand \U$10089 ( \10904 , \9898_nG233b , \9331 );
or \U$10090 ( \10905 , \9204 , \9660_nG2373 );
nand \U$10091 ( \10906 , \10905 , \9427 );
and \U$10092 ( \10907 , \10904 , \10906 );
and \U$10093 ( \10908 , \9430 , \9660_nG2373 );
and \U$10094 ( \10909 , \9898_nG233b , \9333 );
nor \U$10095 ( \10910 , \10907 , \10908 , \10909 );
and \U$10096 ( \10911 , \10860 , \9737 );
not \U$10097 ( \10912 , \9563_nG23ac );
and \U$10098 ( \10913 , \9612 , \10912 );
and \U$10099 ( \10914 , \9481_nG2706 , \9741 );
nor \U$10100 ( \10915 , \10911 , \10913 , \10914 );
xor \U$10101 ( \10916 , \10910 , \10915 );
and \U$10102 ( \10917 , \10916 , \8624 );
and \U$10103 ( \10918 , \10910 , \10915 );
or \U$10104 ( \10919 , \10917 , \10918 );
and \U$10105 ( \10920 , \10235_nG228e , \8890 );
or \U$10106 ( \10921 , \8816 , \10119_nG22ca );
nand \U$10107 ( \10922 , \10921 , \9026 );
nand \U$10108 ( \10923 , \10235_nG228e , \8887 );
and \U$10109 ( \10924 , \10922 , \10923 );
and \U$10110 ( \10925 , \10119_nG22ca , \9030 );
nor \U$10111 ( \10926 , \10920 , \10924 , \10925 );
xor \U$10112 ( \10927 , \10919 , \10926 );
and \U$10113 ( \10928 , \10409_nG225a , \8890 );
or \U$10114 ( \10929 , \8816 , \10235_nG228e );
nand \U$10115 ( \10930 , \10929 , \9026 );
nand \U$10116 ( \10931 , \10409_nG225a , \8887 );
and \U$10117 ( \10932 , \10930 , \10931 );
and \U$10118 ( \10933 , \10235_nG228e , \9030 );
nor \U$10119 ( \10934 , \10928 , \10932 , \10933 );
and \U$10120 ( \10935 , \9868_nG2303 , \9188 );
or \U$10121 ( \10936 , \9048 , \9868_nG2303 );
nand \U$10122 ( \10937 , \10936 , \9191 );
nand \U$10123 ( \10938 , \10119_nG22ca , \9091 );
and \U$10124 ( \10939 , \10937 , \10938 );
and \U$10125 ( \10940 , \10119_nG22ca , \9094 );
nor \U$10126 ( \10941 , \10935 , \10939 , \10940 );
xor \U$10127 ( \10942 , \10934 , \10941 );
and \U$10128 ( \10943 , \8831 , \10506_nG221a );
nand \U$10129 ( \10944 , \10506_nG221a , \8767 );
and \U$10130 ( \10945 , \10944 , \8771 );
nor \U$10131 ( \10946 , \10943 , \10945 );
and \U$10132 ( \10947 , \10942 , \10946 );
and \U$10133 ( \10948 , \10934 , \10941 );
or \U$10134 ( \10949 , \10947 , \10948 );
and \U$10135 ( \10950 , \10927 , \10949 );
and \U$10136 ( \10951 , \10919 , \10926 );
or \U$10137 ( \10952 , \10950 , \10951 );
nand \U$10138 ( \10953 , \10903 , \10952 );
not \U$10139 ( \10954 , \10409_nG225a );
or \U$10140 ( \10955 , \8896 , \10954 );
or \U$10141 ( \10956 , \10879 , \8898 );
or \U$10142 ( \10957 , \8830 , \10954 );
or \U$10143 ( \10958 , \8624 , \10506_nG221a );
nand \U$10144 ( \10959 , \10958 , \8773 );
nand \U$10145 ( \10960 , \10957 , \10959 );
nand \U$10146 ( \10961 , \10955 , \10956 , \10960 );
not \U$10147 ( \10962 , \10961 );
xor \U$10148 ( \10963 , \10858 , \10863 );
xor \U$10149 ( \10964 , \10963 , \10871 );
nor \U$10150 ( \10965 , \10962 , \10964 );
and \U$10151 ( \10966 , \10953 , \10965 );
nor \U$10152 ( \10967 , \10952 , \10903 );
nor \U$10153 ( \10968 , \10966 , \10967 );
nor \U$10154 ( \10969 , \10901 , \10968 );
xor \U$10155 ( \10970 , \10899 , \10969 );
not \U$10156 ( \10971 , \10965 );
not \U$10157 ( \10972 , \10967 );
nand \U$10158 ( \10973 , \10972 , \10953 );
not \U$10159 ( \10974 , \10973 );
or \U$10160 ( \10975 , \10971 , \10974 );
or \U$10161 ( \10976 , \10973 , \10965 );
nand \U$10162 ( \10977 , \10975 , \10976 );
xor \U$10163 ( \10978 , \10793 , \10800 );
xor \U$10164 ( \10979 , \10978 , \10808 );
xor \U$10165 ( \10980 , \10874 , \10882 );
xor \U$10166 ( \10981 , \10979 , \10980 );
not \U$10167 ( \10982 , \10981 );
xor \U$10168 ( \10983 , \10977 , \10982 );
not \U$10169 ( \10984 , \10961 );
not \U$10170 ( \10985 , \10964 );
and \U$10171 ( \10986 , \10984 , \10985 );
and \U$10172 ( \10987 , \10961 , \10964 );
nor \U$10173 ( \10988 , \10986 , \10987 );
not \U$10174 ( \10989 , \10988 );
nand \U$10175 ( \10990 , \9868_nG2303 , \9331 );
or \U$10176 ( \10991 , \9204 , \9898_nG233b );
nand \U$10177 ( \10992 , \10991 , \9427 );
and \U$10178 ( \10993 , \10990 , \10992 );
and \U$10179 ( \10994 , \9430 , \9898_nG233b );
and \U$10180 ( \10995 , \9868_nG2303 , \9333 );
nor \U$10181 ( \10996 , \10993 , \10994 , \10995 );
not \U$10182 ( \10997 , \10996 );
and \U$10183 ( \10998 , \10912 , \9737 );
not \U$10184 ( \10999 , \9660_nG2373 );
and \U$10185 ( \11000 , \9612 , \10999 );
and \U$10186 ( \11001 , \9563_nG23ac , \9741 );
nor \U$10187 ( \11002 , \10998 , \11000 , \11001 );
not \U$10188 ( \11003 , \11002 );
and \U$10189 ( \11004 , \10997 , \11003 );
and \U$10190 ( \11005 , \10996 , \11002 );
and \U$10191 ( \11006 , \10119_nG22ca , \9188 );
or \U$10192 ( \11007 , \9048 , \10119_nG22ca );
nand \U$10193 ( \11008 , \11007 , \9191 );
nand \U$10194 ( \11009 , \10235_nG228e , \9091 );
and \U$10195 ( \11010 , \11008 , \11009 );
and \U$10196 ( \11011 , \10235_nG228e , \9094 );
nor \U$10197 ( \11012 , \11006 , \11010 , \11011 );
nor \U$10198 ( \11013 , \11005 , \11012 );
nor \U$10199 ( \11014 , \11004 , \11013 );
xor \U$10200 ( \11015 , \10910 , \10915 );
xor \U$10201 ( \11016 , \11015 , \8624 );
and \U$10202 ( \11017 , \11014 , \11016 );
xor \U$10203 ( \11018 , \10934 , \10941 );
xor \U$10204 ( \11019 , \11018 , \10946 );
xor \U$10205 ( \11020 , \10910 , \10915 );
xor \U$10206 ( \11021 , \11020 , \8624 );
and \U$10207 ( \11022 , \11019 , \11021 );
and \U$10208 ( \11023 , \11014 , \11019 );
or \U$10209 ( \11024 , \11017 , \11022 , \11023 );
xor \U$10210 ( \11025 , \10919 , \10926 );
xor \U$10211 ( \11026 , \11025 , \10949 );
or \U$10212 ( \11027 , \11024 , \11026 );
not \U$10213 ( \11028 , \11027 );
or \U$10214 ( \11029 , \10989 , \11028 );
nand \U$10215 ( \11030 , \11026 , \11024 );
nand \U$10216 ( \11031 , \11029 , \11030 );
not \U$10217 ( \11032 , \11031 );
xor \U$10218 ( \11033 , \10983 , \11032 );
nand \U$10219 ( \11034 , \11027 , \11030 );
not \U$10220 ( \11035 , \11034 );
not \U$10221 ( \11036 , \10988 );
and \U$10222 ( \11037 , \11035 , \11036 );
and \U$10223 ( \11038 , \11034 , \10988 );
nor \U$10224 ( \11039 , \11037 , \11038 );
xor \U$10225 ( \11040 , \10910 , \10915 );
xor \U$10226 ( \11041 , \11040 , \8624 );
xor \U$10227 ( \11042 , \11014 , \11019 );
xor \U$10228 ( \11043 , \11041 , \11042 );
or \U$10229 ( \11044 , \9101 , \10879 );
or \U$10230 ( \11045 , \10506_nG221a , \8816 );
nand \U$10231 ( \11046 , \11044 , \11045 , \9026 );
not \U$10232 ( \11047 , \11046 );
and \U$10233 ( \11048 , \10235_nG228e , \9188 );
or \U$10234 ( \11049 , \9048 , \10235_nG228e );
nand \U$10235 ( \11050 , \11049 , \9191 );
nand \U$10236 ( \11051 , \10409_nG225a , \9091 );
and \U$10237 ( \11052 , \11050 , \11051 );
and \U$10238 ( \11053 , \10409_nG225a , \9094 );
nor \U$10239 ( \11054 , \11048 , \11052 , \11053 );
nor \U$10240 ( \11055 , \11047 , \11054 );
nand \U$10241 ( \11056 , \10119_nG22ca , \9331 );
or \U$10242 ( \11057 , \9204 , \9868_nG2303 );
nand \U$10243 ( \11058 , \11057 , \9427 );
and \U$10244 ( \11059 , \11056 , \11058 );
and \U$10245 ( \11060 , \9430 , \9868_nG2303 );
and \U$10246 ( \11061 , \10119_nG22ca , \9333 );
nor \U$10247 ( \11062 , \11059 , \11060 , \11061 );
and \U$10248 ( \11063 , \10999 , \9737 );
not \U$10249 ( \11064 , \9898_nG233b );
and \U$10250 ( \11065 , \9612 , \11064 );
and \U$10251 ( \11066 , \9660_nG2373 , \9741 );
nor \U$10252 ( \11067 , \11063 , \11065 , \11066 );
xor \U$10253 ( \11068 , \11062 , \11067 );
and \U$10254 ( \11069 , \11068 , \8816 );
and \U$10255 ( \11070 , \11062 , \11067 );
or \U$10256 ( \11071 , \11069 , \11070 );
and \U$10257 ( \11072 , \10506_nG221a , \8890 );
or \U$10258 ( \11073 , \8816 , \10409_nG225a );
nand \U$10259 ( \11074 , \11073 , \9026 );
nand \U$10260 ( \11075 , \10506_nG221a , \8887 );
and \U$10261 ( \11076 , \11074 , \11075 );
and \U$10262 ( \11077 , \10409_nG225a , \9030 );
nor \U$10263 ( \11078 , \11072 , \11076 , \11077 );
nand \U$10264 ( \11079 , \11071 , \11078 );
and \U$10265 ( \11080 , \11055 , \11079 );
nor \U$10266 ( \11081 , \11078 , \11071 );
nor \U$10267 ( \11082 , \11080 , \11081 );
nor \U$10268 ( \11083 , \11043 , \11082 );
xor \U$10269 ( \11084 , \11039 , \11083 );
not \U$10270 ( \11085 , \10996 );
xor \U$10271 ( \11086 , \11002 , \11012 );
not \U$10272 ( \11087 , \11086 );
or \U$10273 ( \11088 , \11085 , \11087 );
or \U$10274 ( \11089 , \11086 , \10996 );
nand \U$10275 ( \11090 , \11088 , \11089 );
not \U$10276 ( \11091 , \11055 );
not \U$10277 ( \11092 , \11081 );
nand \U$10278 ( \11093 , \11092 , \11079 );
not \U$10279 ( \11094 , \11093 );
or \U$10280 ( \11095 , \11091 , \11094 );
or \U$10281 ( \11096 , \11093 , \11055 );
nand \U$10282 ( \11097 , \11095 , \11096 );
xor \U$10283 ( \11098 , \11090 , \11097 );
not \U$10284 ( \11099 , \11046 );
not \U$10285 ( \11100 , \11054 );
and \U$10286 ( \11101 , \11099 , \11100 );
and \U$10287 ( \11102 , \11046 , \11054 );
nor \U$10288 ( \11103 , \11101 , \11102 );
nand \U$10289 ( \11104 , \10235_nG228e , \9331 );
or \U$10290 ( \11105 , \9204 , \10119_nG22ca );
nand \U$10291 ( \11106 , \11105 , \9427 );
and \U$10292 ( \11107 , \11104 , \11106 );
and \U$10293 ( \11108 , \9430 , \10119_nG22ca );
and \U$10294 ( \11109 , \10235_nG228e , \9333 );
nor \U$10295 ( \11110 , \11107 , \11108 , \11109 );
and \U$10296 ( \11111 , \11064 , \9737 );
not \U$10297 ( \11112 , \9868_nG2303 );
and \U$10298 ( \11113 , \9612 , \11112 );
and \U$10299 ( \11114 , \9898_nG233b , \9741 );
nor \U$10300 ( \11115 , \11111 , \11113 , \11114 );
xor \U$10301 ( \11116 , \11110 , \11115 );
and \U$10302 ( \11117 , \10409_nG225a , \9188 );
or \U$10303 ( \11118 , \9048 , \10409_nG225a );
nand \U$10304 ( \11119 , \11118 , \9191 );
nand \U$10305 ( \11120 , \10506_nG221a , \9091 );
and \U$10306 ( \11121 , \11119 , \11120 );
and \U$10307 ( \11122 , \10506_nG221a , \9094 );
nor \U$10308 ( \11123 , \11117 , \11121 , \11122 );
and \U$10309 ( \11124 , \11116 , \11123 );
and \U$10310 ( \11125 , \11110 , \11115 );
or \U$10311 ( \11126 , \11124 , \11125 );
xor \U$10312 ( \11127 , \11062 , \11067 );
xor \U$10313 ( \11128 , \11127 , \8816 );
or \U$10314 ( \11129 , \11126 , \11128 );
and \U$10315 ( \11130 , \11103 , \11129 );
and \U$10316 ( \11131 , \11128 , \11126 );
nor \U$10317 ( \11132 , \11130 , \11131 );
xor \U$10318 ( \11133 , \11098 , \11132 );
xor \U$10319 ( \11134 , \11128 , \11103 );
and \U$10320 ( \11135 , \11134 , \11126 );
nor \U$10321 ( \11136 , \11134 , \11126 );
or \U$10322 ( \11137 , \11135 , \11136 );
or \U$10323 ( \11138 , \9740 , \11112 );
or \U$10324 ( \11139 , \9868_nG2303 , \9614 );
or \U$10325 ( \11140 , \10119_nG22ca , \9613 );
nand \U$10326 ( \11141 , \11138 , \11139 , \11140 );
xor \U$10327 ( \11142 , \9093 , \11141 );
or \U$10328 ( \11143 , \9334 , \10954 );
or \U$10329 ( \11144 , \9204 , \10235_nG228e );
nand \U$10330 ( \11145 , \11144 , \9427 );
nand \U$10331 ( \11146 , \10409_nG225a , \9331 );
and \U$10332 ( \11147 , \11145 , \11146 );
and \U$10333 ( \11148 , \10235_nG228e , \9430 );
nor \U$10334 ( \11149 , \11147 , \11148 );
nand \U$10335 ( \11150 , \11143 , \11149 );
and \U$10336 ( \11151 , \11142 , \11150 );
and \U$10337 ( \11152 , \9093 , \11141 );
or \U$10338 ( \11153 , \11151 , \11152 );
not \U$10339 ( \11154 , \11153 );
xor \U$10340 ( \11155 , \11110 , \11115 );
xor \U$10341 ( \11156 , \11155 , \11123 );
nor \U$10342 ( \11157 , \11154 , \11156 );
nand \U$10343 ( \11158 , \11137 , \11157 );
or \U$10344 ( \11159 , \11135 , \11136 , \11157 );
xor \U$10345 ( \11160 , \9093 , \11141 );
xor \U$10346 ( \11161 , \11160 , \11150 );
not \U$10347 ( \11162 , \11161 );
and \U$10348 ( \11163 , \10506_nG221a , \9188 );
and \U$10349 ( \11164 , \10879 , \9093 );
not \U$10350 ( \11165 , \9191 );
nor \U$10351 ( \11166 , \11163 , \11164 , \11165 );
not \U$10352 ( \11167 , \11166 );
or \U$10353 ( \11168 , \11162 , \11167 );
or \U$10354 ( \11169 , \11166 , \11161 );
nand \U$10355 ( \11170 , \11168 , \11169 );
nand \U$10356 ( \11171 , \10506_nG221a , \9331 );
or \U$10357 ( \11172 , \9204 , \10409_nG225a );
nand \U$10358 ( \11173 , \11172 , \9427 );
and \U$10359 ( \11174 , \11171 , \11173 );
and \U$10360 ( \11175 , \9430 , \10409_nG225a );
and \U$10361 ( \11176 , \10506_nG221a , \9333 );
nor \U$10362 ( \11177 , \11174 , \11175 , \11176 );
not \U$10363 ( \11178 , \10119_nG22ca );
and \U$10364 ( \11179 , \11178 , \9737 );
not \U$10365 ( \11180 , \10235_nG228e );
and \U$10366 ( \11181 , \9612 , \11180 );
and \U$10367 ( \11182 , \10119_nG22ca , \9741 );
nor \U$10368 ( \11183 , \11179 , \11181 , \11182 );
nor \U$10369 ( \11184 , \11177 , \11183 );
or \U$10370 ( \11185 , \11170 , \11184 );
and \U$10371 ( \11186 , \9611 , \10409_nG225a );
nor \U$10372 ( \11187 , \11186 , \9198 , \10506_nG221a );
not \U$10373 ( \11188 , \11187 );
or \U$10374 ( \11189 , \9740 , \11180 );
or \U$10375 ( \11190 , \10235_nG228e , \9614 );
or \U$10376 ( \11191 , \10409_nG225a , \9613 );
nand \U$10377 ( \11192 , \11189 , \11190 , \11191 );
xor \U$10378 ( \11193 , \11192 , \9205 );
not \U$10379 ( \11194 , \11193 );
or \U$10380 ( \11195 , \11188 , \11194 );
not \U$10381 ( \11196 , \9430 );
and \U$10382 ( \11197 , \11196 , \10506_nG221a );
and \U$10383 ( \11198 , \10879 , \9204 );
nor \U$10384 ( \11199 , \11197 , \11198 );
not \U$10385 ( \11200 , \9427 );
or \U$10386 ( \11201 , \11199 , \11200 );
or \U$10387 ( \11202 , \11187 , \11193 );
nand \U$10388 ( \11203 , \11201 , \11202 );
nand \U$10389 ( \11204 , \11195 , \11203 );
and \U$10390 ( \11205 , \11192 , \9205 );
and \U$10391 ( \11206 , \11204 , \11205 );
and \U$10392 ( \11207 , \11177 , \11183 );
nor \U$10393 ( \11208 , \11207 , \11184 );
or \U$10394 ( \11209 , \11206 , \11208 );
or \U$10395 ( \11210 , \11205 , \11204 );
nand \U$10396 ( \11211 , \11185 , \11209 , \11210 );
not \U$10397 ( \11212 , \11166 );
nand \U$10398 ( \11213 , \11212 , \11161 );
nand \U$10399 ( \11214 , \11184 , \11170 );
and \U$10400 ( \11215 , \11211 , \11213 , \11214 );
not \U$10401 ( \11216 , \11156 );
not \U$10402 ( \11217 , \11153 );
and \U$10403 ( \11218 , \11216 , \11217 );
and \U$10404 ( \11219 , \11156 , \11153 );
nor \U$10405 ( \11220 , \11218 , \11219 );
nor \U$10406 ( \11221 , \11215 , \11220 );
nor \U$10407 ( \11222 , \11211 , \11213 );
or \U$10408 ( \11223 , \11221 , \11222 );
nand \U$10409 ( \11224 , \11159 , \11223 );
nand \U$10410 ( \11225 , \11158 , \11224 );
and \U$10411 ( \11226 , \11133 , \11225 );
and \U$10412 ( \11227 , \11098 , \11132 );
or \U$10413 ( \11228 , \11226 , \11227 );
and \U$10414 ( \11229 , \11090 , \11097 );
xor \U$10415 ( \11230 , \11228 , \11229 );
and \U$10416 ( \11231 , \11043 , \11082 );
nor \U$10417 ( \11232 , \11231 , \11083 );
and \U$10418 ( \11233 , \11230 , \11232 );
and \U$10419 ( \11234 , \11228 , \11229 );
or \U$10420 ( \11235 , \11233 , \11234 );
and \U$10421 ( \11236 , \11084 , \11235 );
and \U$10422 ( \11237 , \11039 , \11083 );
or \U$10423 ( \11238 , \11236 , \11237 );
and \U$10424 ( \11239 , \11033 , \11238 );
and \U$10425 ( \11240 , \10983 , \11032 );
or \U$10426 ( \11241 , \11239 , \11240 );
and \U$10427 ( \11242 , \10977 , \10982 );
xor \U$10428 ( \11243 , \11241 , \11242 );
and \U$10429 ( \11244 , \10901 , \10968 );
nor \U$10430 ( \11245 , \11244 , \10969 );
and \U$10431 ( \11246 , \11243 , \11245 );
and \U$10432 ( \11247 , \11241 , \11242 );
or \U$10433 ( \11248 , \11246 , \11247 );
and \U$10434 ( \11249 , \10970 , \11248 );
and \U$10435 ( \11250 , \10899 , \10969 );
or \U$10436 ( \11251 , \11249 , \11250 );
and \U$10437 ( \11252 , \10897 , \11251 );
and \U$10438 ( \11253 , \10849 , \10896 );
or \U$10439 ( \11254 , \11252 , \11253 );
xor \U$10440 ( \11255 , \10843 , \10845 );
and \U$10441 ( \11256 , \11255 , \10847 );
and \U$10442 ( \11257 , \10843 , \10845 );
or \U$10443 ( \11258 , \11256 , \11257 );
xor \U$10444 ( \11259 , \10698 , \10777 );
xor \U$10445 ( \11260 , \11259 , \10780 );
nand \U$10446 ( \11261 , \11258 , \11260 );
and \U$10447 ( \11262 , \11254 , \11261 );
nor \U$10448 ( \11263 , \11260 , \11258 );
nor \U$10449 ( \11264 , \11262 , \11263 );
xor \U$10450 ( \11265 , \10682 , \10684 );
xor \U$10451 ( \11266 , \11265 , \10687 );
and \U$10452 ( \11267 , \11264 , \11266 );
and \U$10453 ( \11268 , \10783 , \11264 );
or \U$10454 ( \11269 , \10786 , \11267 , \11268 );
xor \U$10455 ( \11270 , \10607 , \10612 );
xor \U$10456 ( \11271 , \11270 , \10615 );
and \U$10457 ( \11272 , \11269 , \11271 );
and \U$10458 ( \11273 , \10690 , \11269 );
or \U$10459 ( \11274 , \10693 , \11272 , \11273 );
not \U$10460 ( \11275 , \11274 );
and \U$10461 ( \11276 , \10620 , \11275 );
and \U$10462 ( \11277 , \10539 , \10619 );
or \U$10463 ( \11278 , \11276 , \11277 );
and \U$10464 ( \11279 , \10537 , \11278 );
and \U$10465 ( \11280 , \10531 , \10536 );
or \U$10466 ( \11281 , \11279 , \11280 );
and \U$10467 ( \11282 , \10529 , \11281 );
and \U$10468 ( \11283 , \10367 , \10528 );
or \U$10469 ( \11284 , \11282 , \11283 );
xor \U$10470 ( \11285 , \10249 , \10263 );
xor \U$10471 ( \11286 , \11285 , \10274 );
not \U$10472 ( \11287 , \10359 );
not \U$10473 ( \11288 , \10363 );
and \U$10474 ( \11289 , \11287 , \11288 );
nor \U$10475 ( \11290 , \11289 , \10358 );
nand \U$10476 ( \11291 , \11286 , \11290 );
and \U$10477 ( \11292 , \11284 , \11291 );
nor \U$10478 ( \11293 , \11290 , \11286 );
nor \U$10479 ( \11294 , \11292 , \11293 );
and \U$10480 ( \11295 , \10278 , \11294 );
and \U$10481 ( \11296 , \10083 , \10277 );
or \U$10482 ( \11297 , \11295 , \11296 );
not \U$10483 ( \11298 , \11297 );
and \U$10484 ( \11299 , \10076 , \11298 );
and \U$10485 ( \11300 , \10058 , \10075 );
or \U$10486 ( \11301 , \11299 , \11300 );
xor \U$10487 ( \11302 , \9783 , \9795 );
xor \U$10488 ( \11303 , \11302 , \9798 );
or \U$10489 ( \11304 , \10071 , \10067 );
nand \U$10490 ( \11305 , \11304 , \10065 );
nand \U$10491 ( \11306 , \11303 , \11305 );
and \U$10492 ( \11307 , \11301 , \11306 );
nor \U$10493 ( \11308 , \11305 , \11303 );
nor \U$10494 ( \11309 , \11307 , \11308 );
xor \U$10495 ( \11310 , \9687 , \9692 );
xor \U$10496 ( \11311 , \11310 , \9700 );
and \U$10497 ( \11312 , \11309 , \11311 );
and \U$10498 ( \11313 , \9801 , \11309 );
or \U$10499 ( \11314 , \9804 , \11312 , \11313 );
and \U$10500 ( \11315 , \9704 , \11314 );
and \U$10501 ( \11316 , \9536 , \9703 );
or \U$10502 ( \11317 , \11315 , \11316 );
not \U$10503 ( \11318 , \11317 );
and \U$10504 ( \11319 , \9529 , \11318 );
and \U$10505 ( \11320 , \9397 , \9528 );
or \U$10506 ( \11321 , \11319 , \11320 );
and \U$10507 ( \11322 , \9395 , \11321 );
and \U$10508 ( \11323 , \9290 , \9394 );
or \U$10509 ( \11324 , \11322 , \11323 );
and \U$10510 ( \11325 , \9286 , \11324 );
and \U$10511 ( \11326 , \9283 , \9285 );
or \U$10512 ( \11327 , \11325 , \11326 );
and \U$10513 ( \11328 , \9171 , \11327 );
and \U$10514 ( \11329 , \9083 , \9170 );
or \U$10515 ( \11330 , \11328 , \11329 );
and \U$10516 ( \11331 , \9081 , \11330 );
and \U$10517 ( \11332 , \8975 , \9080 );
or \U$10518 ( \11333 , \11331 , \11332 );
and \U$10519 ( \11334 , \8973 , \11333 );
and \U$10520 ( \11335 , \8807 , \8972 );
or \U$10521 ( \11336 , \11334 , \11335 );
and \U$10522 ( \11337 , \8805 , \11336 );
and \U$10523 ( \11338 , \8803 , \8804 );
or \U$10524 ( \11339 , \11337 , \11338 );
not \U$10525 ( \11340 , \11339 );
or \U$10526 ( \11341 , \8697 , \11340 );
or \U$10527 ( \11342 , \11339 , \8696 );
nand \U$10528 ( \11343 , \11341 , \11342 );
and \U$10529 ( \11344 , \7944 , RIaa981c0_25);
and \U$10530 ( \11345 , \7959 , RIaa98418_30);
and \U$10531 ( \11346 , RIaa982b0_27, \7909 );
nor \U$10532 ( \11347 , \11345 , \11346 );
and \U$10533 ( \11348 , \7914 , RIaa97ef0_19);
and \U$10534 ( \11349 , RIaa98058_22, \7952 );
nor \U$10535 ( \11350 , \11348 , \11349 );
and \U$10536 ( \11351 , \7942 , RIaa98238_26);
and \U$10537 ( \11352 , RIaa983a0_29, \7919 );
nor \U$10538 ( \11353 , \11351 , \11352 );
and \U$10539 ( \11354 , \7961 , RIaa98508_32);
and \U$10540 ( \11355 , RIaa985f8_34, \7957 );
nor \U$10541 ( \11356 , \11354 , \11355 );
nand \U$10542 ( \11357 , \11347 , \11350 , \11353 , \11356 );
not \U$10543 ( \11358 , \7956 );
nor \U$10544 ( \11359 , \11344 , \11357 , \11358 );
and \U$10545 ( \11360 , \7928 , RIaa98328_28);
and \U$10546 ( \11361 , RIaa980d0_23, \7930 );
nor \U$10547 ( \11362 , \11360 , \11361 );
and \U$10548 ( \11363 , \7949 , RIaa97fe0_21);
and \U$10549 ( \11364 , RIaa98148_24, \7923 );
nor \U$10550 ( \11365 , \11363 , \11364 );
and \U$10551 ( \11366 , \7935 , RIaa98490_31);
and \U$10552 ( \11367 , RIaa98580_33, \7963 );
nor \U$10553 ( \11368 , \11366 , \11367 );
nand \U$10554 ( \11369 , \11359 , \11362 , \11365 , \11368 );
buf \U$10555 ( \11370 , \11369 );
buf \U$10556 ( \11371 , \7972 );
_DC g2a95 ( \11372_nG2a95 , \11370 , \11371 );
xor \U$10557 ( \11373 , \7897 , \11372_nG2a95 );
and \U$10558 ( \11374 , \7923 , RIaa98850_39);
and \U$10559 ( \11375 , \7919 , RIaa98b98_46);
and \U$10560 ( \11376 , RIaa98c10_47, \7959 );
nor \U$10561 ( \11377 , \11375 , \11376 );
and \U$10562 ( \11378 , \7942 , RIaa98a30_43);
and \U$10563 ( \11379 , RIaa98d00_49, \7957 );
nor \U$10564 ( \11380 , \11378 , \11379 );
and \U$10565 ( \11381 , \7961 , RIaa98df0_51);
and \U$10566 ( \11382 , RIaa98940_41, \7952 );
nor \U$10567 ( \11383 , \11381 , \11382 );
and \U$10568 ( \11384 , \7928 , RIaa98aa8_44);
and \U$10569 ( \11385 , RIaa98c88_48, \7909 );
nor \U$10570 ( \11386 , \11384 , \11385 );
nand \U$10571 ( \11387 , \11377 , \11380 , \11383 , \11386 );
and \U$10572 ( \11388 , \7930 , RIaa987d8_38);
and \U$10573 ( \11389 , RIaa989b8_42, \7944 );
nor \U$10574 ( \11390 , \11388 , \11389 );
not \U$10575 ( \11391 , \11390 );
nor \U$10576 ( \11392 , \11374 , \11387 , \11391 );
and \U$10577 ( \11393 , \7914 , RIaa98670_35);
and \U$10578 ( \11394 , RIaa988c8_40, \7949 );
nor \U$10579 ( \11395 , \11393 , \11394 );
and \U$10580 ( \11396 , \7935 , RIaa98d78_50);
and \U$10581 ( \11397 , RIaa98b20_45, \7963 );
nor \U$10582 ( \11398 , \11396 , \11397 );
nand \U$10583 ( \11399 , \11392 , \11395 , \7986 , \11398 );
buf \U$10584 ( \11400 , \11399 );
_DC g28b7 ( \11401_nG28b7 , \11400 , \11371 );
xor \U$10585 ( \11402 , \7980 , \11401_nG28b7 );
and \U$10586 ( \11403 , RIaa9e340_233, \7928 );
and \U$10587 ( \11404 , RIaa9e070_227, \7952 );
and \U$10588 ( \11405 , \7963 , RIaa9e598_238);
and \U$10589 ( \11406 , RIaa9e0e8_228, \7930 );
nor \U$10590 ( \11407 , \11405 , \11406 );
and \U$10591 ( \11408 , RIaa9e4a8_236, \7935 );
and \U$10592 ( \11409 , \7944 , RIaa9e1d8_230);
and \U$10593 ( \11410 , RIaa9dff8_226, \7949 );
nor \U$10594 ( \11411 , \11408 , \11409 , \11410 );
and \U$10595 ( \11412 , \7914 , RIaa9de90_223);
and \U$10596 ( \11413 , RIaa9e160_229, \7923 );
nor \U$10597 ( \11414 , \11412 , \11413 );
nand \U$10598 ( \11415 , \11407 , \11411 , \11414 );
nor \U$10599 ( \11416 , \11403 , \11404 , \11415 );
and \U$10600 ( \11417 , \7961 , RIaa9e520_237);
and \U$10601 ( \11418 , RIaa9e610_239, \7957 );
nor \U$10602 ( \11419 , \11417 , \11418 );
and \U$10603 ( \11420 , RIaa9e430_235, \7959 );
and \U$10604 ( \11421 , RIaa9e2c8_232, \7909 );
and \U$10605 ( \11422 , \7942 , RIaa9e250_231);
and \U$10606 ( \11423 , RIaa9e3b8_234, \7919 );
nor \U$10607 ( \11424 , \11422 , \11423 );
not \U$10608 ( \11425 , \11424 );
nor \U$10609 ( \11426 , \11420 , \11421 , \11425 );
nand \U$10610 ( \11427 , \11416 , \11419 , \8024 , \11426 );
buf \U$10611 ( \11428 , \11427 );
_DC g28b5 ( \11429_nG28b5 , \11428 , \11371 );
xor \U$10612 ( \11430 , \8018 , \11429_nG28b5 );
and \U$10613 ( \11431 , \7923 , RIaa9de18_222);
and \U$10614 ( \11432 , \7919 , RIaa9d878_210);
and \U$10615 ( \11433 , RIaa9d8f0_211, \7959 );
nor \U$10616 ( \11434 , \11432 , \11433 );
and \U$10617 ( \11435 , \7928 , RIaa9d710_207);
and \U$10618 ( \11436 , RIaa9d698_206, \7909 );
nor \U$10619 ( \11437 , \11435 , \11436 );
and \U$10620 ( \11438 , \7961 , RIaa9d9e0_213);
and \U$10621 ( \11439 , RIaa9dc38_218, \7952 );
nor \U$10622 ( \11440 , \11438 , \11439 );
and \U$10623 ( \11441 , \7942 , RIaa9dd28_220);
and \U$10624 ( \11442 , RIaa9d800_209, \7957 );
nor \U$10625 ( \11443 , \11441 , \11442 );
nand \U$10626 ( \11444 , \11434 , \11437 , \11440 , \11443 );
and \U$10627 ( \11445 , \7930 , RIaa9dda0_221);
and \U$10628 ( \11446 , RIaa9dcb0_219, \7944 );
nor \U$10629 ( \11447 , \11445 , \11446 );
not \U$10630 ( \11448 , \11447 );
nor \U$10631 ( \11449 , \11431 , \11444 , \11448 );
and \U$10632 ( \11450 , \7914 , RIaa9da58_214);
and \U$10633 ( \11451 , RIaa9dbc0_217, \7949 );
nor \U$10634 ( \11452 , \11450 , \11451 );
and \U$10635 ( \11453 , \7935 , RIaa9d968_212);
and \U$10636 ( \11454 , RIaa9d788_208, \7963 );
nor \U$10637 ( \11455 , \11453 , \11454 );
nand \U$10638 ( \11456 , \11449 , \11452 , \8062 , \11455 );
buf \U$10639 ( \11457 , \11456 );
_DC g270a ( \11458_nG270a , \11457 , \11371 );
xor \U$10640 ( \11459 , \8056 , \11458_nG270a );
and \U$10641 ( \11460 , RIaa99048_56, \7923 );
and \U$10642 ( \11461 , RIaa98e68_52, \7914 );
and \U$10643 ( \11462 , \7919 , RIaa991b0_59);
and \U$10644 ( \11463 , RIaa99228_60, \7959 );
nor \U$10645 ( \11464 , \11462 , \11463 );
and \U$10646 ( \11465 , \7928 , RIaa990c0_57);
and \U$10647 ( \11466 , RIaa99480_65, \7909 );
nor \U$10648 ( \11467 , \11465 , \11466 );
and \U$10649 ( \11468 , \7961 , RIaa99570_67);
and \U$10650 ( \11469 , RIaa992a0_61, \7952 );
nor \U$10651 ( \11470 , \11468 , \11469 );
and \U$10652 ( \11471 , \7942 , RIaa99408_64);
and \U$10653 ( \11472 , RIaa994f8_66, \7957 );
nor \U$10654 ( \11473 , \11471 , \11472 );
nand \U$10655 ( \11474 , \11464 , \11467 , \11470 , \11473 );
nor \U$10656 ( \11475 , \11460 , \11461 , \11474 );
and \U$10657 ( \11476 , \7963 , RIaa99138_58);
and \U$10658 ( \11477 , RIaa98fd0_55, \7930 );
nor \U$10659 ( \11478 , \11476 , \11477 );
and \U$10660 ( \11479 , \7949 , RIaa99318_62);
not \U$10661 ( \11480 , \8118 );
nor \U$10662 ( \11481 , \11479 , \11480 );
and \U$10663 ( \11482 , \7935 , RIaa995e8_68);
and \U$10664 ( \11483 , RIaa99390_63, \7944 );
nor \U$10665 ( \11484 , \11482 , \11483 );
nand \U$10666 ( \11485 , \11475 , \11478 , \11481 , \11484 );
buf \U$10667 ( \11486 , \11485 );
_DC g2708 ( \11487_nG2708 , \11486 , \11371 );
xor \U$10668 ( \11488 , \8094 , \11487_nG2708 );
and \U$10669 ( \11489 , RIaa99c00_81, \7942 );
and \U$10670 ( \11490 , RIaa99de0_85, \7957 );
and \U$10671 ( \11491 , \7961 , RIaa99660_69);
and \U$10672 ( \11492 , RIaa99a98_78, \7952 );
nor \U$10673 ( \11493 , \11491 , \11492 );
not \U$10674 ( \11494 , \11493 );
nor \U$10675 ( \11495 , \11489 , \11490 , \11494 );
and \U$10676 ( \11496 , \7944 , RIaa99b88_80);
and \U$10677 ( \11497 , RIaa99cf0_83, \7909 );
nor \U$10678 ( \11498 , \11496 , \11497 );
and \U$10679 ( \11499 , \7928 , RIaa99c78_82);
and \U$10680 ( \11500 , RIaa999a8_76, \7930 );
nor \U$10681 ( \11501 , \11499 , \11500 );
and \U$10682 ( \11502 , RIaa99750_71, \7919 );
and \U$10683 ( \11503 , \7959 , RIaa997c8_72);
and \U$10684 ( \11504 , RIaa99a20_77, \7923 );
nor \U$10685 ( \11505 , \11502 , \11503 , \11504 );
nand \U$10686 ( \11506 , \11495 , \11498 , \11501 , \11505 );
not \U$10687 ( \11507 , \11506 );
and \U$10688 ( \11508 , \7935 , RIaa996d8_70);
and \U$10689 ( \11509 , RIaa99d68_84, \7963 );
nor \U$10690 ( \11510 , \11508 , \11509 );
and \U$10691 ( \11511 , \7914 , RIaa99840_73);
and \U$10692 ( \11512 , RIaa99b10_79, \7949 );
nor \U$10693 ( \11513 , \11511 , \11512 );
nand \U$10694 ( \11514 , \11507 , \11510 , \8136 , \11513 );
buf \U$10695 ( \11515 , \11514 );
_DC g2377 ( \11516_nG2377 , \11515 , \11371 );
xor \U$10696 ( \11517 , \8130 , \11516_nG2377 );
and \U$10697 ( \11518 , RIaa9a038_90, \7923 );
and \U$10698 ( \11519 , RIaa99e58_86, \7914 );
and \U$10699 ( \11520 , \7919 , RIaa9a4e8_100);
and \U$10700 ( \11521 , RIaa9a560_101, \7959 );
nor \U$10701 ( \11522 , \11520 , \11521 );
and \U$10702 ( \11523 , \7942 , RIaa9a218_94);
and \U$10703 ( \11524 , RIaa9a5d8_102, \7957 );
nor \U$10704 ( \11525 , \11523 , \11524 );
and \U$10705 ( \11526 , \7961 , RIaa9a380_97);
and \U$10706 ( \11527 , RIaa9a128_92, \7952 );
nor \U$10707 ( \11528 , \11526 , \11527 );
and \U$10708 ( \11529 , \7928 , RIaa9a308_96);
and \U$10709 ( \11530 , RIaa9a470_99, \7909 );
nor \U$10710 ( \11531 , \11529 , \11530 );
nand \U$10711 ( \11532 , \11522 , \11525 , \11528 , \11531 );
nor \U$10712 ( \11533 , \11518 , \11519 , \11532 );
and \U$10713 ( \11534 , \7963 , RIaa9a290_95);
and \U$10714 ( \11535 , RIaa99f48_88, \7930 );
nor \U$10715 ( \11536 , \11534 , \11535 );
and \U$10716 ( \11537 , \7949 , RIaa9a1a0_93);
not \U$10717 ( \11538 , \8192 );
nor \U$10718 ( \11539 , \11537 , \11538 );
and \U$10719 ( \11540 , \7935 , RIaa9a3f8_98);
and \U$10720 ( \11541 , RIaa9a0b0_91, \7944 );
nor \U$10721 ( \11542 , \11540 , \11541 );
nand \U$10722 ( \11543 , \11533 , \11536 , \11539 , \11542 );
buf \U$10723 ( \11544 , \11543 );
_DC g2375 ( \11545_nG2375 , \11544 , \11371 );
xor \U$10724 ( \11546 , \8168 , \11545_nG2375 );
and \U$10725 ( \11547 , RIaa9a920_109, \7928 );
and \U$10726 ( \11548 , RIaa9ace0_117, \7952 );
and \U$10727 ( \11549 , \7963 , RIaa9a8a8_108);
and \U$10728 ( \11550 , RIaa9a7b8_106, \7930 );
nor \U$10729 ( \11551 , \11549 , \11550 );
and \U$10730 ( \11552 , RIaa9aa10_111, \7935 );
and \U$10731 ( \11553 , \7944 , RIaa9ad58_118);
and \U$10732 ( \11554 , RIaa9ac68_116, \7949 );
nor \U$10733 ( \11555 , \11552 , \11553 , \11554 );
and \U$10734 ( \11556 , \7914 , RIaa9a650_103);
and \U$10735 ( \11557 , RIaa9a830_107, \7923 );
nor \U$10736 ( \11558 , \11556 , \11557 );
nand \U$10737 ( \11559 , \11551 , \11555 , \11558 );
nor \U$10738 ( \11560 , \11547 , \11548 , \11559 );
and \U$10739 ( \11561 , \7961 , RIaa9a998_110);
and \U$10740 ( \11562 , RIaa9abf0_115, \7957 );
nor \U$10741 ( \11563 , \11561 , \11562 );
and \U$10742 ( \11564 , RIaa9ab00_113, \7959 );
and \U$10743 ( \11565 , RIaa9aa88_112, \7909 );
and \U$10744 ( \11566 , \7942 , RIaa9add0_119);
and \U$10745 ( \11567 , RIaa9ab78_114, \7919 );
nor \U$10746 ( \11568 , \11566 , \11567 );
not \U$10747 ( \11569 , \11568 );
nor \U$10748 ( \11570 , \11564 , \11565 , \11569 );
nand \U$10749 ( \11571 , \11560 , \11563 , \8220 , \11570 );
buf \U$10750 ( \11572 , \11571 );
_DC g2307 ( \11573_nG2307 , \11572 , \11371 );
xor \U$10751 ( \11574 , \8204 , \11573_nG2307 );
and \U$10752 ( \11575 , RIaa9cf90_191, \7923 );
and \U$10753 ( \11576 , RIaa9d008_192, \7914 );
and \U$10754 ( \11577 , \7919 , RIaa9d3c8_200);
and \U$10755 ( \11578 , RIaa9d350_199, \7959 );
nor \U$10756 ( \11579 , \11577 , \11578 );
and \U$10757 ( \11580 , \7942 , RIaa9d620_205);
and \U$10758 ( \11581 , RIaa9d440_201, \7957 );
nor \U$10759 ( \11582 , \11580 , \11581 );
and \U$10760 ( \11583 , \7961 , RIaa9d1e8_196);
and \U$10761 ( \11584 , RIaa9d4b8_202, \7952 );
nor \U$10762 ( \11585 , \11583 , \11584 );
and \U$10763 ( \11586 , \7928 , RIaa9d0f8_194);
and \U$10764 ( \11587 , RIaa9d2d8_198, \7909 );
nor \U$10765 ( \11588 , \11586 , \11587 );
nand \U$10766 ( \11589 , \11579 , \11582 , \11585 , \11588 );
nor \U$10767 ( \11590 , \11575 , \11576 , \11589 );
and \U$10768 ( \11591 , \7963 , RIaa9d170_195);
and \U$10769 ( \11592 , RIaa9cf18_190, \7930 );
nor \U$10770 ( \11593 , \11591 , \11592 );
and \U$10771 ( \11594 , \7949 , RIaa9d530_203);
not \U$10772 ( \11595 , \8264 );
nor \U$10773 ( \11596 , \11594 , \11595 );
and \U$10774 ( \11597 , \7935 , RIaa9d260_197);
and \U$10775 ( \11598 , RIaa9d5a8_204, \7944 );
nor \U$10776 ( \11599 , \11597 , \11598 );
nand \U$10777 ( \11600 , \11590 , \11593 , \11596 , \11599 );
buf \U$10778 ( \11601 , \11600 );
_DC g2305 ( \11602_nG2305 , \11601 , \11371 );
xor \U$10779 ( \11603 , \8240 , \11602_nG2305 );
and \U$10780 ( \11604 , RIaa9b118_126, \7928 );
and \U$10781 ( \11605 , RIaa9b550_135, \7952 );
and \U$10782 ( \11606 , \7963 , RIaa9b0a0_125);
and \U$10783 ( \11607 , RIaa9afb0_123, \7930 );
nor \U$10784 ( \11608 , \11606 , \11607 );
and \U$10785 ( \11609 , RIaa9b208_128, \7935 );
and \U$10786 ( \11610 , \7944 , RIaa9b460_133);
and \U$10787 ( \11611 , RIaa9b5c8_136, \7949 );
nor \U$10788 ( \11612 , \11609 , \11610 , \11611 );
and \U$10789 ( \11613 , \7914 , RIaa9ae48_120);
and \U$10790 ( \11614 , RIaa9b028_124, \7923 );
nor \U$10791 ( \11615 , \11613 , \11614 );
nand \U$10792 ( \11616 , \11608 , \11612 , \11615 );
nor \U$10793 ( \11617 , \11604 , \11605 , \11616 );
and \U$10794 ( \11618 , \7961 , RIaa9b190_127);
and \U$10795 ( \11619 , RIaa9b3e8_132, \7957 );
nor \U$10796 ( \11620 , \11618 , \11619 );
and \U$10797 ( \11621 , RIaa9b2f8_130, \7959 );
and \U$10798 ( \11622 , RIaa9b280_129, \7909 );
and \U$10799 ( \11623 , \7942 , RIaa9b4d8_134);
and \U$10800 ( \11624 , RIaa9b370_131, \7919 );
nor \U$10801 ( \11625 , \11623 , \11624 );
not \U$10802 ( \11626 , \11625 );
nor \U$10803 ( \11627 , \11621 , \11622 , \11626 );
nand \U$10804 ( \11628 , \11617 , \11620 , \8288 , \11627 );
buf \U$10805 ( \11629 , \11628 );
_DC g22ad ( \11630_nG22ad , \11629 , \11371 );
xor \U$10806 ( \11631 , \8272 , \11630_nG22ad );
and \U$10807 ( \11632 , \7919 , RIaa9bb68_148);
and \U$10808 ( \11633 , RIaa9baf0_147, \7959 );
nor \U$10809 ( \11634 , \11632 , \11633 );
and \U$10810 ( \11635 , \7961 , RIaa9b730_139);
and \U$10811 ( \11636 , RIaa9bc58_150, \7952 );
nor \U$10812 ( \11637 , \11635 , \11636 );
nand \U$10813 ( \11638 , RIaa9bcd0_151, \7949 );
and \U$10814 ( \11639 , \7963 , RIaa9b6b8_138);
and \U$10815 ( \11640 , RIaa9b988_144, \7930 );
nor \U$10816 ( \11641 , \11639 , \11640 );
nand \U$10817 ( \11642 , \11634 , \11637 , \11638 , \11641 );
not \U$10818 ( \11643 , \11642 );
and \U$10819 ( \11644 , RIaa9bdc0_153, \7942 );
and \U$10820 ( \11645 , \7957 , RIaa9bbe0_149);
and \U$10821 ( \11646 , RIaa9b640_137, \7928 );
nor \U$10822 ( \11647 , \11644 , \11645 , \11646 );
nand \U$10823 ( \11648 , RIaa9ba78_146, \7909 );
and \U$10824 ( \11649 , \11647 , \11648 , \8332 );
and \U$10825 ( \11650 , \7914 , RIaa9b820_141);
and \U$10826 ( \11651 , RIaa9ba00_145, \7923 );
nor \U$10827 ( \11652 , \11650 , \11651 );
and \U$10828 ( \11653 , \7935 , RIaa9b7a8_140);
and \U$10829 ( \11654 , RIaa9bd48_152, \7944 );
nor \U$10830 ( \11655 , \11653 , \11654 );
nand \U$10831 ( \11656 , \11643 , \11649 , \11652 , \11655 );
buf \U$10832 ( \11657 , \11656 );
_DC g22af ( \11658_nG22af , \11657 , \11371 );
xor \U$10833 ( \11659 , \8308 , \11658_nG22af );
and \U$10834 ( \11660 , \7923 , RIaa9c180_161);
and \U$10835 ( \11661 , \7919 , RIaa9c360_165);
and \U$10836 ( \11662 , RIaa9c3d8_166, \7959 );
nor \U$10837 ( \11663 , \11661 , \11662 );
and \U$10838 ( \11664 , \7942 , RIaa9c4c8_168);
and \U$10839 ( \11665 , RIaa9beb0_155, \7957 );
nor \U$10840 ( \11666 , \11664 , \11665 );
and \U$10841 ( \11667 , \7961 , RIaa9c270_163);
and \U$10842 ( \11668 , RIaa9bfa0_157, \7952 );
nor \U$10843 ( \11669 , \11667 , \11668 );
and \U$10844 ( \11670 , \7928 , RIaa9c5b8_170);
and \U$10845 ( \11671 , RIaa9be38_154, \7909 );
nor \U$10846 ( \11672 , \11670 , \11671 );
nand \U$10847 ( \11673 , \11663 , \11666 , \11669 , \11672 );
and \U$10848 ( \11674 , \7930 , RIaa9c1f8_162);
and \U$10849 ( \11675 , RIaa9c450_167, \7944 );
nor \U$10850 ( \11676 , \11674 , \11675 );
not \U$10851 ( \11677 , \11676 );
nor \U$10852 ( \11678 , \11660 , \11673 , \11677 );
and \U$10853 ( \11679 , \7914 , RIaa9c018_158);
and \U$10854 ( \11680 , RIaa9bf28_156, \7949 );
nor \U$10855 ( \11681 , \11679 , \11680 );
and \U$10856 ( \11682 , \7935 , RIaa9c540_169);
and \U$10857 ( \11683 , RIaa9c2e8_164, \7963 );
nor \U$10858 ( \11684 , \11682 , \11683 );
nand \U$10859 ( \11685 , \11678 , \11681 , \8345 , \11684 );
buf \U$10860 ( \11686 , \11685 );
_DC g223f ( \11687_nG223f , \11686 , \11371 );
xor \U$10861 ( \11688 , RIaaa91a0_605, \11687_nG223f );
and \U$10862 ( \11689 , \7963 , RIaa9ccc0_185);
and \U$10863 ( \11690 , RIaa9c630_171, \7930 );
nor \U$10864 ( \11691 , \11689 , \11690 );
and \U$10865 ( \11692 , \7961 , RIaa9cc48_184);
and \U$10866 ( \11693 , RIaa9c978_178, \7952 );
nor \U$10867 ( \11694 , \11692 , \11693 );
nand \U$10868 ( \11695 , RIaa9cae0_181, \7949 );
and \U$10869 ( \11696 , \7942 , RIaa9cb58_182);
and \U$10870 ( \11697 , RIaa9cdb0_187, \7957 );
nor \U$10871 ( \11698 , \11696 , \11697 );
nand \U$10872 ( \11699 , \11691 , \11694 , \11695 , \11698 );
not \U$10873 ( \11700 , \11699 );
and \U$10874 ( \11701 , RIaa9c9f0_179, \7919 );
and \U$10875 ( \11702 , \7959 , RIaa9cbd0_183);
and \U$10876 ( \11703 , RIaa9c888_176, \7928 );
nor \U$10877 ( \11704 , \11701 , \11702 , \11703 );
nand \U$10878 ( \11705 , RIaa9cd38_186, \7909 );
and \U$10879 ( \11706 , \11704 , \11705 , \8396 );
and \U$10880 ( \11707 , \7914 , RIaa9c6a8_172);
and \U$10881 ( \11708 , RIaa9c810_175, \7923 );
nor \U$10882 ( \11709 , \11707 , \11708 );
and \U$10883 ( \11710 , \7935 , RIaa9c900_177);
and \U$10884 ( \11711 , RIaa9ca68_180, \7944 );
nor \U$10885 ( \11712 , \11710 , \11711 );
nand \U$10886 ( \11713 , \11700 , \11706 , \11709 , \11712 );
buf \U$10887 ( \11714 , \11713 );
_DC g223d ( \11715_nG223d , \11714 , \11371 );
nand \U$10888 ( \11716 , \11715_nG223d , \8403 );
not \U$10889 ( \11717 , \11716 );
and \U$10890 ( \11718 , \11688 , \11717 );
and \U$10891 ( \11719 , RIaaa91a0_605, \11687_nG223f );
or \U$10892 ( \11720 , \11718 , \11719 );
and \U$10893 ( \11721 , \11659 , \11720 );
and \U$10894 ( \11722 , \8308 , \11658_nG22af );
or \U$10895 ( \11723 , \11721 , \11722 );
and \U$10896 ( \11724 , \11631 , \11723 );
and \U$10897 ( \11725 , \8272 , \11630_nG22ad );
or \U$10898 ( \11726 , \11724 , \11725 );
and \U$10899 ( \11727 , \11603 , \11726 );
and \U$10900 ( \11728 , \8240 , \11602_nG2305 );
or \U$10901 ( \11729 , \11727 , \11728 );
and \U$10902 ( \11730 , \11574 , \11729 );
and \U$10903 ( \11731 , \8204 , \11573_nG2307 );
or \U$10904 ( \11732 , \11730 , \11731 );
and \U$10905 ( \11733 , \11546 , \11732 );
and \U$10906 ( \11734 , \8168 , \11545_nG2375 );
or \U$10907 ( \11735 , \11733 , \11734 );
and \U$10908 ( \11736 , \11517 , \11735 );
and \U$10909 ( \11737 , \8130 , \11516_nG2377 );
or \U$10910 ( \11738 , \11736 , \11737 );
and \U$10911 ( \11739 , \11488 , \11738 );
and \U$10912 ( \11740 , \8094 , \11487_nG2708 );
or \U$10913 ( \11741 , \11739 , \11740 );
and \U$10914 ( \11742 , \11459 , \11741 );
and \U$10915 ( \11743 , \8056 , \11458_nG270a );
or \U$10916 ( \11744 , \11742 , \11743 );
and \U$10917 ( \11745 , \11430 , \11744 );
and \U$10918 ( \11746 , \8018 , \11429_nG28b5 );
or \U$10919 ( \11747 , \11745 , \11746 );
and \U$10920 ( \11748 , \11402 , \11747 );
and \U$10921 ( \11749 , \7980 , \11401_nG28b7 );
or \U$10922 ( \11750 , \11748 , \11749 );
and \U$10923 ( \11751 , \11373 , \11750 );
and \U$10924 ( \11752 , \7897 , \11372_nG2a95 );
or \U$10925 ( \11753 , \11751 , \11752 );
nor \U$10926 ( \11754 , \11753 , \8443 );
not \U$10927 ( \11755 , \11754 );
and \U$10928 ( \11756 , RIaa9f768_276, \7957 );
and \U$10929 ( \11757 , RIaa9f3a8_268, \7944 );
and \U$10930 ( \11758 , \7949 , RIaa9f420_269);
and \U$10931 ( \11759 , RIaa9f600_273, \7930 );
nor \U$10932 ( \11760 , \11758 , \11759 );
or \U$10933 ( \11761 , \7923 , \7955 );
and \U$10934 ( \11762 , RIaa9f588_272, \11761 );
and \U$10935 ( \11763 , \7935 , RIaa9f2b8_266);
and \U$10936 ( \11764 , RIaa9f948_280, \7961 );
nor \U$10937 ( \11765 , \11762 , \11763 , \11764 );
and \U$10938 ( \11766 , \7928 , RIaa9f9c0_281);
and \U$10939 ( \11767 , RIaa9f8d0_279, \7909 );
nor \U$10940 ( \11768 , \11766 , \11767 );
nand \U$10941 ( \11769 , \11760 , \11765 , \11768 );
nor \U$10942 ( \11770 , \11756 , \11757 , \11769 );
and \U$10943 ( \11771 , \7914 , RIaa9f330_267);
and \U$10944 ( \11772 , RIaa9f7e0_277, \7959 );
nor \U$10945 ( \11773 , \11771 , \11772 );
and \U$10946 ( \11774 , \7942 , RIaa9f678_274);
and \U$10947 ( \11775 , RIaa9f6f0_275, \7919 );
nor \U$10948 ( \11776 , \11774 , \11775 );
and \U$10949 ( \11777 , \7952 , RIaa9f858_278);
and \U$10950 ( \11778 , RIaa9f498_270, \7963 );
nor \U$10951 ( \11779 , \11777 , \11778 );
nand \U$10952 ( \11780 , \11770 , \11773 , \11776 , \11779 );
buf \U$10953 ( \11781 , \7972 );
_DC g30bb ( \11782_nG30bb , \11780 , \11781 );
not \U$10954 ( \11783 , \11782_nG30bb );
nor \U$10955 ( \11784 , \11755 , \11783 );
xor \U$10956 ( \11785 , \7897 , \11372_nG2a95 );
xor \U$10957 ( \11786 , \11785 , \11750 );
not \U$10958 ( \11787 , \11786 );
xor \U$10959 ( \11788 , \7980 , \11401_nG28b7 );
xor \U$10960 ( \11789 , \11788 , \11747 );
not \U$10961 ( \11790 , \11789 );
and \U$10962 ( \11791 , \11787 , \11790 );
and \U$10963 ( \11792 , \11753 , \8443 );
nor \U$10964 ( \11793 , \11792 , \11754 );
nor \U$10965 ( \11794 , \11791 , \11793 );
not \U$10966 ( \11795 , \11794 );
and \U$10967 ( \11796 , \11761 , RIaa9ebb0_251);
and \U$10968 ( \11797 , \7935 , RIaa9ec28_252);
and \U$10969 ( \11798 , RIaa9f0d8_262, \7957 );
nor \U$10970 ( \11799 , \11797 , \11798 );
and \U$10971 ( \11800 , \7942 , RIaa9ee80_257);
and \U$10972 ( \11801 , RIaa9ed18_254, \7944 );
nor \U$10973 ( \11802 , \11800 , \11801 );
and \U$10974 ( \11803 , \7914 , RIaa9eca0_253);
and \U$10975 ( \11804 , RIaa9f150_263, \7952 );
nor \U$10976 ( \11805 , \11803 , \11804 );
and \U$10977 ( \11806 , \7919 , RIaa9eef8_258);
and \U$10978 ( \11807 , RIaa9f060_261, \7959 );
nor \U$10979 ( \11808 , \11806 , \11807 );
nand \U$10980 ( \11809 , \11799 , \11802 , \11805 , \11808 );
nor \U$10981 ( \11810 , \11796 , \11809 );
and \U$10982 ( \11811 , \7928 , RIaa9efe8_260);
and \U$10983 ( \11812 , RIaa9f1c8_264, \7909 );
nor \U$10984 ( \11813 , \11811 , \11812 );
and \U$10985 ( \11814 , \7961 , RIaa9ef70_259);
and \U$10986 ( \11815 , RIaa9ed90_255, \7963 );
nor \U$10987 ( \11816 , \11814 , \11815 );
and \U$10988 ( \11817 , \7949 , RIaa9ee08_256);
and \U$10989 ( \11818 , RIaa9eb38_250, \7930 );
nor \U$10990 ( \11819 , \11817 , \11818 );
nand \U$10991 ( \11820 , \11810 , \11813 , \11816 , \11819 );
_DC g31ca ( \11821_nG31ca , \11820 , \11781 );
or \U$10992 ( \11822 , \11795 , \11821_nG31ca );
not \U$10993 ( \11823 , \11821_nG31ca );
and \U$10994 ( \11824 , \11793 , \11786 );
nor \U$10995 ( \11825 , \11793 , \11786 );
xnor \U$10996 ( \11826 , \11789 , \11786 );
not \U$10997 ( \11827 , \11826 );
nor \U$10998 ( \11828 , \11824 , \11825 , \11827 );
nand \U$10999 ( \11829 , \11795 , \11828 );
or \U$11000 ( \11830 , \11823 , \11829 );
or \U$11001 ( \11831 , \11828 , \11795 );
nand \U$11002 ( \11832 , \11822 , \11830 , \11831 );
xnor \U$11003 ( \11833 , \11784 , \11832 );
nor \U$11004 ( \11834 , \11794 , \11826 );
not \U$11005 ( \11835 , \11834 );
or \U$11006 ( \11836 , \11835 , \11823 );
or \U$11007 ( \11837 , \11783 , \11829 );
or \U$11008 ( \11838 , \11826 , \11823 );
or \U$11009 ( \11839 , \11795 , \11782_nG30bb );
nand \U$11010 ( \11840 , \11839 , \11831 );
nand \U$11011 ( \11841 , \11838 , \11840 );
nand \U$11012 ( \11842 , \11836 , \11837 , \11841 );
xor \U$11013 ( \11843 , \8018 , \11429_nG28b5 );
xor \U$11014 ( \11844 , \11843 , \11744 );
xor \U$11015 ( \11845 , \8056 , \11458_nG270a );
xor \U$11016 ( \11846 , \11845 , \11741 );
nor \U$11017 ( \11847 , \11844 , \11846 );
or \U$11018 ( \11848 , \11789 , \11847 );
and \U$11019 ( \11849 , \11842 , \11848 );
and \U$11020 ( \11850 , RIaa9ff60_293, \7942 );
and \U$11021 ( \11851 , RIaa9ffd8_294, \7919 );
and \U$11022 ( \11852 , \7963 , RIaaa00c8_296);
and \U$11023 ( \11853 , RIaa9fc90_287, \7930 );
nor \U$11024 ( \11854 , \11852 , \11853 );
and \U$11025 ( \11855 , RIaa9fc18_286, \11761 );
and \U$11026 ( \11856 , \7961 , RIaa9fd08_288);
and \U$11027 ( \11857 , RIaa9fdf8_290, \7949 );
nor \U$11028 ( \11858 , \11855 , \11856 , \11857 );
and \U$11029 ( \11859 , \7928 , RIaa9fd80_289);
and \U$11030 ( \11860 , RIaa9fab0_283, \7909 );
nor \U$11031 ( \11861 , \11859 , \11860 );
nand \U$11032 ( \11862 , \11854 , \11858 , \11861 );
nor \U$11033 ( \11863 , \11850 , \11851 , \11862 );
and \U$11034 ( \11864 , \7952 , RIaa9fa38_282);
and \U$11035 ( \11865 , RIaaa01b8_298, \7935 );
nor \U$11036 ( \11866 , \11864 , \11865 );
and \U$11037 ( \11867 , \7914 , RIaaa0140_297);
and \U$11038 ( \11868 , RIaa9fee8_292, \7959 );
nor \U$11039 ( \11869 , \11867 , \11868 );
and \U$11040 ( \11870 , \7957 , RIaa9fe70_291);
and \U$11041 ( \11871 , RIaaa0050_295, \7944 );
nor \U$11042 ( \11872 , \11870 , \11871 );
nand \U$11043 ( \11873 , \11863 , \11866 , \11869 , \11872 );
_DC g2fb5 ( \11874_nG2fb5 , \11873 , \11781 );
nand \U$11044 ( \11875 , \11874_nG2fb5 , \11754 );
not \U$11045 ( \11876 , \11875 );
nor \U$11046 ( \11877 , \11849 , \11876 );
xor \U$11047 ( \11878 , \11833 , \11877 );
not \U$11048 ( \11879 , \11878 );
not \U$11049 ( \11880 , \11844 );
not \U$11050 ( \11881 , \11789 );
or \U$11051 ( \11882 , \11880 , \11881 );
or \U$11052 ( \11883 , \11789 , \11844 );
nand \U$11053 ( \11884 , \11882 , \11883 );
xor \U$11054 ( \11885 , \11846 , \11844 );
nor \U$11055 ( \11886 , \11884 , \11885 );
not \U$11056 ( \11887 , \11886 );
not \U$11057 ( \11888 , \11848 );
nor \U$11058 ( \11889 , \11887 , \11888 );
not \U$11059 ( \11890 , \11889 );
or \U$11060 ( \11891 , \11890 , \11823 );
or \U$11061 ( \11892 , \11887 , \11823 );
nand \U$11062 ( \11893 , \11892 , \11888 );
nand \U$11063 ( \11894 , \11891 , \11893 );
or \U$11064 ( \11895 , \11835 , \11783 );
not \U$11065 ( \11896 , \11874_nG2fb5 );
or \U$11066 ( \11897 , \11896 , \11829 );
or \U$11067 ( \11898 , \11826 , \11783 );
or \U$11068 ( \11899 , \11795 , \11874_nG2fb5 );
nand \U$11069 ( \11900 , \11899 , \11831 );
nand \U$11070 ( \11901 , \11898 , \11900 );
nand \U$11071 ( \11902 , \11895 , \11897 , \11901 );
and \U$11072 ( \11903 , \11894 , \11902 );
not \U$11073 ( \11904 , \11875 );
and \U$11074 ( \11905 , \11842 , \11848 );
not \U$11075 ( \11906 , \11842 );
and \U$11076 ( \11907 , \11906 , \11888 );
nor \U$11077 ( \11908 , \11905 , \11907 );
not \U$11078 ( \11909 , \11908 );
or \U$11079 ( \11910 , \11904 , \11909 );
or \U$11080 ( \11911 , \11908 , \11875 );
nand \U$11081 ( \11912 , \11910 , \11911 );
and \U$11082 ( \11913 , \11903 , \11912 );
xor \U$11083 ( \11914 , \11879 , \11913 );
nand \U$11084 ( \11915 , \11782_nG30bb , \11886 );
or \U$11085 ( \11916 , \11848 , \11821_nG31ca );
or \U$11086 ( \11917 , \11848 , \11885 );
nand \U$11087 ( \11918 , \11916 , \11917 );
and \U$11088 ( \11919 , \11915 , \11918 );
and \U$11089 ( \11920 , \11848 , \11885 );
and \U$11090 ( \11921 , \11920 , \11821_nG31ca );
and \U$11091 ( \11922 , \11782_nG30bb , \11889 );
nor \U$11092 ( \11923 , \11919 , \11921 , \11922 );
and \U$11093 ( \11924 , \11874_nG2fb5 , \11834 );
not \U$11094 ( \11925 , \11829 );
and \U$11095 ( \11926 , \7930 , RIaaa0848_312);
and \U$11096 ( \11927 , \7952 , RIaaa0938_314);
and \U$11097 ( \11928 , RIaaa0230_299, \7957 );
nor \U$11098 ( \11929 , \11927 , \11928 );
and \U$11099 ( \11930 , \7942 , RIaaa0578_306);
and \U$11100 ( \11931 , RIaaa0488_304, \7944 );
nor \U$11101 ( \11932 , \11930 , \11931 );
and \U$11102 ( \11933 , \7914 , RIaaa0668_308);
and \U$11103 ( \11934 , RIaaa06e0_309, \7935 );
nor \U$11104 ( \11935 , \11933 , \11934 );
and \U$11105 ( \11936 , \7919 , RIaaa05f0_307);
and \U$11106 ( \11937 , RIaaa02a8_300, \7959 );
nor \U$11107 ( \11938 , \11936 , \11937 );
nand \U$11108 ( \11939 , \11929 , \11932 , \11935 , \11938 );
nor \U$11109 ( \11940 , \11926 , \11939 );
and \U$11110 ( \11941 , \7961 , RIaaa0320_301);
and \U$11111 ( \11942 , RIaaa0500_305, \7963 );
nor \U$11112 ( \11943 , \11941 , \11942 );
and \U$11113 ( \11944 , \7928 , RIaaa0398_302);
and \U$11114 ( \11945 , RIaaa08c0_313, \7909 );
nor \U$11115 ( \11946 , \11944 , \11945 );
and \U$11116 ( \11947 , \11761 , RIaaa07d0_311);
and \U$11117 ( \11948 , RIaaa0410_303, \7949 );
nor \U$11118 ( \11949 , \11947 , \11948 );
nand \U$11119 ( \11950 , \11940 , \11943 , \11946 , \11949 );
_DC g2e94 ( \11951_nG2e94 , \11950 , \11781 );
and \U$11120 ( \11952 , \11925 , \11951_nG2e94 );
nand \U$11121 ( \11953 , \11874_nG2fb5 , \11827 );
or \U$11122 ( \11954 , \11795 , \11951_nG2e94 );
nand \U$11123 ( \11955 , \11954 , \11831 );
and \U$11124 ( \11956 , \11953 , \11955 );
nor \U$11125 ( \11957 , \11924 , \11952 , \11956 );
nand \U$11126 ( \11958 , \11923 , \11957 );
xor \U$11127 ( \11959 , \8094 , \11487_nG2708 );
xor \U$11128 ( \11960 , \11959 , \11738 );
xor \U$11129 ( \11961 , \8130 , \11516_nG2377 );
xor \U$11130 ( \11962 , \11961 , \11735 );
nor \U$11131 ( \11963 , \11960 , \11962 );
or \U$11132 ( \11964 , \11846 , \11963 );
and \U$11133 ( \11965 , \11958 , \11964 );
nor \U$11134 ( \11966 , \11957 , \11923 );
nor \U$11135 ( \11967 , \11965 , \11966 );
xor \U$11136 ( \11968 , \11894 , \11902 );
not \U$11137 ( \11969 , \11968 );
nand \U$11138 ( \11970 , \11951_nG2e94 , \11754 );
not \U$11139 ( \11971 , \11970 );
and \U$11140 ( \11972 , \11969 , \11971 );
and \U$11141 ( \11973 , \11968 , \11970 );
nor \U$11142 ( \11974 , \11972 , \11973 );
nand \U$11143 ( \11975 , \11967 , \11974 );
xor \U$11144 ( \11976 , \11903 , \11912 );
and \U$11145 ( \11977 , \11975 , \11976 );
and \U$11146 ( \11978 , \11914 , \11977 );
not \U$11147 ( \11979 , \11978 );
and \U$11148 ( \11980 , \11879 , \11913 );
or \U$11149 ( \11981 , \11980 , \11794 );
and \U$11150 ( \11982 , \11980 , \11794 );
and \U$11151 ( \11983 , \11784 , \11832 );
nor \U$11152 ( \11984 , \11982 , \11983 );
nand \U$11153 ( \11985 , \11981 , \11984 );
not \U$11154 ( \11986 , \11985 );
and \U$11155 ( \11987 , \11754 , \11821_nG31ca );
and \U$11156 ( \11988 , \11833 , \11877 );
nor \U$11157 ( \11989 , \11987 , \11988 );
not \U$11158 ( \11990 , \11989 );
and \U$11159 ( \11991 , \11986 , \11990 );
and \U$11160 ( \11992 , \11985 , \11989 );
nor \U$11161 ( \11993 , \11991 , \11992 );
not \U$11162 ( \11994 , \11993 );
or \U$11163 ( \11995 , \11979 , \11994 );
or \U$11164 ( \11996 , \11993 , \11978 );
nand \U$11165 ( \11997 , \11995 , \11996 );
not \U$11166 ( \11998 , \11997 );
xor \U$11167 ( \11999 , \11975 , \11976 );
not \U$11168 ( \12000 , \11968 );
nor \U$11169 ( \12001 , \12000 , \11970 );
xor \U$11170 ( \12002 , \11999 , \12001 );
or \U$11171 ( \12003 , \11974 , \11967 );
nand \U$11172 ( \12004 , \12003 , \11975 );
nand \U$11173 ( \12005 , \11874_nG2fb5 , \11886 );
or \U$11174 ( \12006 , \11848 , \11782_nG30bb );
nand \U$11175 ( \12007 , \12006 , \11917 );
and \U$11176 ( \12008 , \12005 , \12007 );
and \U$11177 ( \12009 , \11920 , \11782_nG30bb );
and \U$11178 ( \12010 , \11874_nG2fb5 , \11889 );
nor \U$11179 ( \12011 , \12008 , \12009 , \12010 );
and \U$11180 ( \12012 , \11846 , \11960 );
nor \U$11181 ( \12013 , \11846 , \11960 );
xor \U$11182 ( \12014 , \11960 , \11962 );
nor \U$11183 ( \12015 , \12012 , \12013 , \12014 );
and \U$11184 ( \12016 , \12015 , \11964 );
and \U$11185 ( \12017 , \11821_nG31ca , \12016 );
not \U$11186 ( \12018 , \11964 );
and \U$11187 ( \12019 , \11823 , \12018 );
or \U$11188 ( \12020 , \12015 , \11964 );
not \U$11189 ( \12021 , \12020 );
nor \U$11190 ( \12022 , \12017 , \12019 , \12021 );
or \U$11191 ( \12023 , \12011 , \12022 );
and \U$11192 ( \12024 , RIaaa2030_363, \7957 );
and \U$11193 ( \12025 , RIaaa1ce8_356, \7944 );
and \U$11194 ( \12026 , \7963 , RIaaa1dd8_358);
and \U$11195 ( \12027 , RIaaa1b80_353, \7930 );
nor \U$11196 ( \12028 , \12026 , \12027 );
and \U$11197 ( \12029 , RIaaa1b08_352, \11761 );
and \U$11198 ( \12030 , \7961 , RIaaa1f40_361);
and \U$11199 ( \12031 , RIaaa1d60_357, \7949 );
nor \U$11200 ( \12032 , \12029 , \12030 , \12031 );
and \U$11201 ( \12033 , \7928 , RIaaa1fb8_362);
and \U$11202 ( \12034 , RIaaa2198_366, \7909 );
nor \U$11203 ( \12035 , \12033 , \12034 );
nand \U$11204 ( \12036 , \12028 , \12032 , \12035 );
nor \U$11205 ( \12037 , \12024 , \12025 , \12036 );
and \U$11206 ( \12038 , \7914 , RIaaa1c70_355);
and \U$11207 ( \12039 , RIaaa20a8_364, \7959 );
nor \U$11208 ( \12040 , \12038 , \12039 );
and \U$11209 ( \12041 , \7942 , RIaaa1e50_359);
and \U$11210 ( \12042 , RIaaa1ec8_360, \7919 );
nor \U$11211 ( \12043 , \12041 , \12042 );
and \U$11212 ( \12044 , \7952 , RIaaa2120_365);
and \U$11213 ( \12045 , RIaaa1bf8_354, \7935 );
nor \U$11214 ( \12046 , \12044 , \12045 );
nand \U$11215 ( \12047 , \12037 , \12040 , \12043 , \12046 );
_DC g2ca8 ( \12048_nG2ca8 , \12047 , \11781 );
nand \U$11216 ( \12049 , \12048_nG2ca8 , \11754 );
and \U$11217 ( \12050 , \11951_nG2e94 , \11834 );
and \U$11218 ( \12051 , \11761 , RIaaa0fc8_328);
and \U$11219 ( \12052 , \7935 , RIaaa0c80_321);
and \U$11220 ( \12053 , RIaaa0cf8_322, \7957 );
nor \U$11221 ( \12054 , \12052 , \12053 );
and \U$11222 ( \12055 , \7942 , RIaaa0b18_318);
and \U$11223 ( \12056 , RIaaa0a28_316, \7944 );
nor \U$11224 ( \12057 , \12055 , \12056 );
and \U$11225 ( \12058 , \7914 , RIaaa0c08_320);
and \U$11226 ( \12059 , RIaaa1130_331, \7952 );
nor \U$11227 ( \12060 , \12058 , \12059 );
and \U$11228 ( \12061 , \7919 , RIaaa0b90_319);
and \U$11229 ( \12062 , RIaaa0d70_323, \7959 );
nor \U$11230 ( \12063 , \12061 , \12062 );
nand \U$11231 ( \12064 , \12054 , \12057 , \12060 , \12063 );
nor \U$11232 ( \12065 , \12051 , \12064 );
and \U$11233 ( \12066 , \7928 , RIaaa0e60_325);
and \U$11234 ( \12067 , RIaaa10b8_330, \7909 );
nor \U$11235 ( \12068 , \12066 , \12067 );
and \U$11236 ( \12069 , \7961 , RIaaa0de8_324);
and \U$11237 ( \12070 , RIaaa0aa0_317, \7963 );
nor \U$11238 ( \12071 , \12069 , \12070 );
and \U$11239 ( \12072 , \7949 , RIaaa0ed8_326);
and \U$11240 ( \12073 , RIaaa1040_329, \7930 );
nor \U$11241 ( \12074 , \12072 , \12073 );
nand \U$11242 ( \12075 , \12065 , \12068 , \12071 , \12074 );
_DC g2daa ( \12076_nG2daa , \12075 , \11781 );
and \U$11243 ( \12077 , \11925 , \12076_nG2daa );
nand \U$11244 ( \12078 , \11951_nG2e94 , \11827 );
or \U$11245 ( \12079 , \11795 , \12076_nG2daa );
nand \U$11246 ( \12080 , \12079 , \11831 );
and \U$11247 ( \12081 , \12078 , \12080 );
nor \U$11248 ( \12082 , \12050 , \12077 , \12081 );
or \U$11249 ( \12083 , \12049 , \12082 );
nand \U$11250 ( \12084 , \12023 , \12083 );
not \U$11251 ( \12085 , \12076_nG2daa );
nor \U$11252 ( \12086 , \11755 , \12085 );
not \U$11253 ( \12087 , \11964 );
not \U$11254 ( \12088 , \11966 );
nand \U$11255 ( \12089 , \12088 , \11958 );
not \U$11256 ( \12090 , \12089 );
or \U$11257 ( \12091 , \12087 , \12090 );
or \U$11258 ( \12092 , \12089 , \11964 );
nand \U$11259 ( \12093 , \12091 , \12092 );
xor \U$11260 ( \12094 , \12086 , \12093 );
and \U$11261 ( \12095 , \12084 , \12094 );
and \U$11262 ( \12096 , \12004 , \12095 );
and \U$11263 ( \12097 , \12002 , \12096 );
and \U$11264 ( \12098 , \11999 , \12001 );
or \U$11265 ( \12099 , \12097 , \12098 );
xor \U$11266 ( \12100 , \11914 , \11977 );
xor \U$11267 ( \12101 , \12099 , \12100 );
xor \U$11268 ( \12102 , \12004 , \12095 );
and \U$11269 ( \12103 , \12086 , \12093 );
xor \U$11270 ( \12104 , \12102 , \12103 );
xor \U$11271 ( \12105 , \8168 , \11545_nG2375 );
xor \U$11272 ( \12106 , \12105 , \11732 );
xor \U$11273 ( \12107 , \8204 , \11573_nG2307 );
xor \U$11274 ( \12108 , \12107 , \11729 );
nor \U$11275 ( \12109 , \12106 , \12108 );
or \U$11276 ( \12110 , \11962 , \12109 );
not \U$11277 ( \12111 , \12110 );
nand \U$11278 ( \12112 , \11951_nG2e94 , \11886 );
or \U$11279 ( \12113 , \11848 , \11874_nG2fb5 );
nand \U$11280 ( \12114 , \12113 , \11917 );
and \U$11281 ( \12115 , \12112 , \12114 );
and \U$11282 ( \12116 , \11920 , \11874_nG2fb5 );
and \U$11283 ( \12117 , \11951_nG2e94 , \11889 );
nor \U$11284 ( \12118 , \12115 , \12116 , \12117 );
nand \U$11285 ( \12119 , \11821_nG31ca , \12014 );
or \U$11286 ( \12120 , \11964 , \11782_nG30bb );
nand \U$11287 ( \12121 , \12120 , \12020 );
and \U$11288 ( \12122 , \12119 , \12121 );
and \U$11289 ( \12123 , \12016 , \11782_nG30bb );
not \U$11290 ( \12124 , \12014 );
nor \U$11291 ( \12125 , \12018 , \12124 );
and \U$11292 ( \12126 , \11821_nG31ca , \12125 );
nor \U$11293 ( \12127 , \12122 , \12123 , \12126 );
nor \U$11294 ( \12128 , \12118 , \12127 );
not \U$11295 ( \12129 , \12128 );
nand \U$11296 ( \12130 , \12127 , \12118 );
nand \U$11297 ( \12131 , \12129 , \12130 );
not \U$11298 ( \12132 , \12131 );
or \U$11299 ( \12133 , \12111 , \12132 );
or \U$11300 ( \12134 , \12131 , \12110 );
nand \U$11301 ( \12135 , \12133 , \12134 );
and \U$11302 ( \12136 , RIaaa1838_346, \7957 );
and \U$11303 ( \12137 , RIaaa16d0_343, \7919 );
and \U$11304 ( \12138 , \7963 , RIaaa15e0_341);
and \U$11305 ( \12139 , RIaaa1388_336, \7930 );
nor \U$11306 ( \12140 , \12138 , \12139 );
and \U$11307 ( \12141 , RIaaa1310_335, \11761 );
and \U$11308 ( \12142 , \7961 , RIaaa1748_344);
and \U$11309 ( \12143 , RIaaa1568_340, \7949 );
nor \U$11310 ( \12144 , \12141 , \12142 , \12143 );
and \U$11311 ( \12145 , \7928 , RIaaa17c0_345);
and \U$11312 ( \12146 , RIaaa19a0_349, \7909 );
nor \U$11313 ( \12147 , \12145 , \12146 );
nand \U$11314 ( \12148 , \12140 , \12144 , \12147 );
nor \U$11315 ( \12149 , \12136 , \12137 , \12148 );
and \U$11316 ( \12150 , \7952 , RIaaa1928_348);
and \U$11317 ( \12151 , RIaaa1400_337, \7935 );
nor \U$11318 ( \12152 , \12150 , \12151 );
and \U$11319 ( \12153 , \7914 , RIaaa1478_338);
and \U$11320 ( \12154 , RIaaa1658_342, \7942 );
nor \U$11321 ( \12155 , \12153 , \12154 );
and \U$11322 ( \12156 , \7959 , RIaaa18b0_347);
and \U$11323 ( \12157 , RIaaa14f0_339, \7944 );
nor \U$11324 ( \12158 , \12156 , \12157 );
nand \U$11325 ( \12159 , \12149 , \12152 , \12155 , \12158 );
_DC g2bb5 ( \12160_nG2bb5 , \12159 , \11781 );
not \U$11326 ( \12161 , \12160_nG2bb5 );
nor \U$11327 ( \12162 , \11755 , \12161 );
or \U$11328 ( \12163 , \11835 , \12085 );
not \U$11329 ( \12164 , \12048_nG2ca8 );
or \U$11330 ( \12165 , \12164 , \11829 );
or \U$11331 ( \12166 , \11826 , \12085 );
or \U$11332 ( \12167 , \11795 , \12048_nG2ca8 );
nand \U$11333 ( \12168 , \12167 , \11831 );
nand \U$11334 ( \12169 , \12166 , \12168 );
nand \U$11335 ( \12170 , \12163 , \12165 , \12169 );
xor \U$11336 ( \12171 , \12162 , \12170 );
and \U$11337 ( \12172 , \12135 , \12171 );
not \U$11338 ( \12173 , \12106 );
not \U$11339 ( \12174 , \11962 );
or \U$11340 ( \12175 , \12173 , \12174 );
or \U$11341 ( \12176 , \11962 , \12106 );
nand \U$11342 ( \12177 , \12175 , \12176 );
xor \U$11343 ( \12178 , \12108 , \12106 );
nor \U$11344 ( \12179 , \12177 , \12178 );
not \U$11345 ( \12180 , \12179 );
not \U$11346 ( \12181 , \12110 );
nor \U$11347 ( \12182 , \12180 , \12181 );
not \U$11348 ( \12183 , \12182 );
or \U$11349 ( \12184 , \12183 , \11823 );
or \U$11350 ( \12185 , \12180 , \11823 );
nand \U$11351 ( \12186 , \12185 , \12181 );
nand \U$11352 ( \12187 , \12184 , \12186 );
not \U$11353 ( \12188 , \12125 );
or \U$11354 ( \12189 , \12188 , \11783 );
not \U$11355 ( \12190 , \12016 );
or \U$11356 ( \12191 , \11896 , \12190 );
or \U$11357 ( \12192 , \12124 , \11783 );
or \U$11358 ( \12193 , \11964 , \11874_nG2fb5 );
nand \U$11359 ( \12194 , \12193 , \12020 );
nand \U$11360 ( \12195 , \12192 , \12194 );
nand \U$11361 ( \12196 , \12189 , \12191 , \12195 );
and \U$11362 ( \12197 , \12187 , \12196 );
and \U$11363 ( \12198 , \12048_nG2ca8 , \11834 );
and \U$11364 ( \12199 , \11925 , \12160_nG2bb5 );
nand \U$11365 ( \12200 , \12048_nG2ca8 , \11827 );
or \U$11366 ( \12201 , \11795 , \12160_nG2bb5 );
nand \U$11367 ( \12202 , \12201 , \11831 );
and \U$11368 ( \12203 , \12200 , \12202 );
nor \U$11369 ( \12204 , \12198 , \12199 , \12203 );
nand \U$11370 ( \12205 , \12076_nG2daa , \11886 );
or \U$11371 ( \12206 , \11848 , \11951_nG2e94 );
nand \U$11372 ( \12207 , \12206 , \11917 );
and \U$11373 ( \12208 , \12205 , \12207 );
and \U$11374 ( \12209 , \11920 , \11951_nG2e94 );
and \U$11375 ( \12210 , \12076_nG2daa , \11889 );
nor \U$11376 ( \12211 , \12208 , \12209 , \12210 );
and \U$11377 ( \12212 , \12204 , \12211 );
and \U$11378 ( \12213 , RIaaa2d50_391, \7957 );
and \U$11379 ( \12214 , RIaaa2b70_387, \7944 );
and \U$11380 ( \12215 , \7949 , RIaaa2eb8_394);
and \U$11381 ( \12216 , RIaaa3098_398, \7930 );
nor \U$11382 ( \12217 , \12215 , \12216 );
and \U$11383 ( \12218 , RIaaa3110_399, \11761 );
and \U$11384 ( \12219 , \7961 , RIaaa2e40_393);
and \U$11385 ( \12220 , RIaaa2af8_386, \7963 );
nor \U$11386 ( \12221 , \12218 , \12219 , \12220 );
and \U$11387 ( \12222 , \7928 , RIaaa2dc8_392);
and \U$11388 ( \12223 , RIaaa2f30_395, \7909 );
nor \U$11389 ( \12224 , \12222 , \12223 );
nand \U$11390 ( \12225 , \12217 , \12221 , \12224 );
nor \U$11391 ( \12226 , \12213 , \12214 , \12225 );
and \U$11392 ( \12227 , \7914 , RIaaa2c60_389);
and \U$11393 ( \12228 , RIaaa2cd8_390, \7959 );
nor \U$11394 ( \12229 , \12227 , \12228 );
and \U$11395 ( \12230 , \7942 , RIaaa2a80_385);
and \U$11396 ( \12231 , RIaaa2a08_384, \7919 );
nor \U$11397 ( \12232 , \12230 , \12231 );
and \U$11398 ( \12233 , \7952 , RIaaa2fa8_396);
and \U$11399 ( \12234 , RIaaa2be8_388, \7935 );
nor \U$11400 ( \12235 , \12233 , \12234 );
nand \U$11401 ( \12236 , \12226 , \12229 , \12232 , \12235 );
_DC g2aae ( \12237_nG2aae , \12236 , \11781 );
nand \U$11402 ( \12238 , \12237_nG2aae , \11754 );
or \U$11403 ( \12239 , \12212 , \12238 );
or \U$11404 ( \12240 , \12204 , \12211 );
nand \U$11405 ( \12241 , \12239 , \12240 );
and \U$11406 ( \12242 , \12197 , \12241 );
and \U$11407 ( \12243 , \12172 , \12242 );
and \U$11408 ( \12244 , \12130 , \12110 );
and \U$11409 ( \12245 , \12162 , \12170 );
nor \U$11410 ( \12246 , \12244 , \12245 , \12128 );
xnor \U$11411 ( \12247 , \12049 , \12082 );
not \U$11412 ( \12248 , \12247 );
xor \U$11413 ( \12249 , \12022 , \12011 );
not \U$11414 ( \12250 , \12249 );
and \U$11415 ( \12251 , \12248 , \12250 );
and \U$11416 ( \12252 , \12247 , \12249 );
nor \U$11417 ( \12253 , \12251 , \12252 );
nand \U$11418 ( \12254 , \12246 , \12253 );
xor \U$11419 ( \12255 , \12243 , \12254 );
xor \U$11420 ( \12256 , \12084 , \12094 );
and \U$11421 ( \12257 , \12255 , \12256 );
and \U$11422 ( \12258 , \12243 , \12254 );
or \U$11423 ( \12259 , \12257 , \12258 );
and \U$11424 ( \12260 , \12104 , \12259 );
and \U$11425 ( \12261 , \12102 , \12103 );
or \U$11426 ( \12262 , \12260 , \12261 );
xor \U$11427 ( \12263 , \11999 , \12001 );
xor \U$11428 ( \12264 , \12263 , \12096 );
xor \U$11429 ( \12265 , \12262 , \12264 );
and \U$11430 ( \12266 , \12160_nG2bb5 , \11834 );
and \U$11431 ( \12267 , \11925 , \12237_nG2aae );
nand \U$11432 ( \12268 , \12160_nG2bb5 , \11827 );
or \U$11433 ( \12269 , \11795 , \12237_nG2aae );
nand \U$11434 ( \12270 , \12269 , \11831 );
and \U$11435 ( \12271 , \12268 , \12270 );
nor \U$11436 ( \12272 , \12266 , \12267 , \12271 );
nand \U$11437 ( \12273 , \12048_nG2ca8 , \11886 );
or \U$11438 ( \12274 , \11848 , \12076_nG2daa );
nand \U$11439 ( \12275 , \12274 , \11917 );
and \U$11440 ( \12276 , \12273 , \12275 );
and \U$11441 ( \12277 , \11920 , \12076_nG2daa );
and \U$11442 ( \12278 , \12048_nG2ca8 , \11889 );
nor \U$11443 ( \12279 , \12276 , \12277 , \12278 );
and \U$11444 ( \12280 , \12272 , \12279 );
not \U$11445 ( \12281 , \12280 );
and \U$11446 ( \12282 , \11761 , RIaaa28a0_381);
and \U$11447 ( \12283 , \7952 , RIaaa2738_378);
and \U$11448 ( \12284 , RIaaa2300_369, \7957 );
nor \U$11449 ( \12285 , \12283 , \12284 );
and \U$11450 ( \12286 , \7942 , RIaaa2468_372);
and \U$11451 ( \12287 , RIaaa2558_374, \7944 );
nor \U$11452 ( \12288 , \12286 , \12287 );
and \U$11453 ( \12289 , \7914 , RIaaa2648_376);
and \U$11454 ( \12290 , RIaaa26c0_377, \7935 );
nor \U$11455 ( \12291 , \12289 , \12290 );
and \U$11456 ( \12292 , \7919 , RIaaa24e0_373);
and \U$11457 ( \12293 , RIaaa2378_370, \7959 );
nor \U$11458 ( \12294 , \12292 , \12293 );
nand \U$11459 ( \12295 , \12285 , \12288 , \12291 , \12294 );
nor \U$11460 ( \12296 , \12282 , \12295 );
and \U$11461 ( \12297 , \7928 , RIaaa2210_367);
and \U$11462 ( \12298 , RIaaa27b0_379, \7909 );
nor \U$11463 ( \12299 , \12297 , \12298 );
and \U$11464 ( \12300 , \7961 , RIaaa2288_368);
and \U$11465 ( \12301 , RIaaa25d0_375, \7963 );
nor \U$11466 ( \12302 , \12300 , \12301 );
and \U$11467 ( \12303 , \7949 , RIaaa23f0_371);
and \U$11468 ( \12304 , RIaaa2918_382, \7930 );
nor \U$11469 ( \12305 , \12303 , \12304 );
nand \U$11470 ( \12306 , \12296 , \12299 , \12302 , \12305 );
_DC g29cd ( \12307_nG29cd , \12306 , \11781 );
nand \U$11471 ( \12308 , \12307_nG29cd , \11754 );
not \U$11472 ( \12309 , \12308 );
and \U$11473 ( \12310 , \12281 , \12309 );
nor \U$11474 ( \12311 , \12272 , \12279 );
nor \U$11475 ( \12312 , \12310 , \12311 );
nand \U$11476 ( \12313 , \11782_nG30bb , \12179 );
or \U$11477 ( \12314 , \12110 , \11821_nG31ca );
or \U$11478 ( \12315 , \12110 , \12178 );
nand \U$11479 ( \12316 , \12314 , \12315 );
and \U$11480 ( \12317 , \12313 , \12316 );
and \U$11481 ( \12318 , \12110 , \12178 );
and \U$11482 ( \12319 , \12318 , \11821_nG31ca );
and \U$11483 ( \12320 , \11782_nG30bb , \12182 );
nor \U$11484 ( \12321 , \12317 , \12319 , \12320 );
nand \U$11485 ( \12322 , \11874_nG2fb5 , \12014 );
or \U$11486 ( \12323 , \11964 , \11951_nG2e94 );
nand \U$11487 ( \12324 , \12323 , \12020 );
and \U$11488 ( \12325 , \12322 , \12324 );
and \U$11489 ( \12326 , \12016 , \11951_nG2e94 );
and \U$11490 ( \12327 , \11874_nG2fb5 , \12125 );
nor \U$11491 ( \12328 , \12325 , \12326 , \12327 );
nand \U$11492 ( \12329 , \12321 , \12328 );
xor \U$11493 ( \12330 , \8272 , \11630_nG22ad );
xor \U$11494 ( \12331 , \12330 , \11723 );
not \U$11495 ( \12332 , \12331 );
xor \U$11496 ( \12333 , \8240 , \11602_nG2305 );
xor \U$11497 ( \12334 , \12333 , \11726 );
not \U$11498 ( \12335 , \12334 );
and \U$11499 ( \12336 , \12332 , \12335 );
or \U$11500 ( \12337 , \12108 , \12336 );
and \U$11501 ( \12338 , \12329 , \12337 );
nor \U$11502 ( \12339 , \12328 , \12321 );
nor \U$11503 ( \12340 , \12338 , \12339 );
nor \U$11504 ( \12341 , \12312 , \12340 );
xor \U$11505 ( \12342 , \12187 , \12196 );
not \U$11506 ( \12343 , \12342 );
not \U$11507 ( \12344 , \12240 );
nor \U$11508 ( \12345 , \12344 , \12212 );
not \U$11509 ( \12346 , \12345 );
not \U$11510 ( \12347 , \12238 );
and \U$11511 ( \12348 , \12346 , \12347 );
and \U$11512 ( \12349 , \12345 , \12238 );
nor \U$11513 ( \12350 , \12348 , \12349 );
nor \U$11514 ( \12351 , \12343 , \12350 );
and \U$11515 ( \12352 , \12341 , \12351 );
xor \U$11516 ( \12353 , \12135 , \12171 );
xor \U$11517 ( \12354 , \12197 , \12241 );
and \U$11518 ( \12355 , \12353 , \12354 );
xor \U$11519 ( \12356 , \12352 , \12355 );
or \U$11520 ( \12357 , \12253 , \12246 );
nand \U$11521 ( \12358 , \12357 , \12254 );
and \U$11522 ( \12359 , \12356 , \12358 );
and \U$11523 ( \12360 , \12352 , \12355 );
or \U$11524 ( \12361 , \12359 , \12360 );
not \U$11525 ( \12362 , \12249 );
nor \U$11526 ( \12363 , \12362 , \12247 );
xor \U$11527 ( \12364 , \12361 , \12363 );
xor \U$11528 ( \12365 , \12243 , \12254 );
xor \U$11529 ( \12366 , \12365 , \12256 );
and \U$11530 ( \12367 , \12364 , \12366 );
and \U$11531 ( \12368 , \12361 , \12363 );
or \U$11532 ( \12369 , \12367 , \12368 );
xor \U$11533 ( \12370 , \12102 , \12103 );
xor \U$11534 ( \12371 , \12370 , \12259 );
xor \U$11535 ( \12372 , \12369 , \12371 );
xor \U$11536 ( \12373 , \12353 , \12354 );
not \U$11537 ( \12374 , \12334 );
not \U$11538 ( \12375 , \12108 );
or \U$11539 ( \12376 , \12374 , \12375 );
or \U$11540 ( \12377 , \12108 , \12334 );
nand \U$11541 ( \12378 , \12376 , \12377 );
xor \U$11542 ( \12379 , \12332 , \12335 );
nor \U$11543 ( \12380 , \12378 , \12379 );
not \U$11544 ( \12381 , \12380 );
not \U$11545 ( \12382 , \12337 );
nor \U$11546 ( \12383 , \12381 , \12382 );
not \U$11547 ( \12384 , \12383 );
or \U$11548 ( \12385 , \12384 , \11823 );
or \U$11549 ( \12386 , \12381 , \11823 );
nand \U$11550 ( \12387 , \12386 , \12382 );
nand \U$11551 ( \12388 , \12385 , \12387 );
or \U$11552 ( \12389 , \12183 , \11896 );
not \U$11553 ( \12390 , \12318 );
or \U$11554 ( \12391 , \11783 , \12390 );
or \U$11555 ( \12392 , \12180 , \11896 );
or \U$11556 ( \12393 , \12110 , \11782_nG30bb );
nand \U$11557 ( \12394 , \12393 , \12315 );
nand \U$11558 ( \12395 , \12392 , \12394 );
nand \U$11559 ( \12396 , \12389 , \12391 , \12395 );
and \U$11560 ( \12397 , \12388 , \12396 );
nand \U$11561 ( \12398 , \12160_nG2bb5 , \11886 );
or \U$11562 ( \12399 , \11848 , \12048_nG2ca8 );
nand \U$11563 ( \12400 , \12399 , \11917 );
and \U$11564 ( \12401 , \12398 , \12400 );
and \U$11565 ( \12402 , \11920 , \12048_nG2ca8 );
and \U$11566 ( \12403 , \12160_nG2bb5 , \11889 );
nor \U$11567 ( \12404 , \12401 , \12402 , \12403 );
nand \U$11568 ( \12405 , \11951_nG2e94 , \12014 );
or \U$11569 ( \12406 , \11964 , \12076_nG2daa );
nand \U$11570 ( \12407 , \12406 , \12020 );
and \U$11571 ( \12408 , \12405 , \12407 );
and \U$11572 ( \12409 , \12016 , \12076_nG2daa );
and \U$11573 ( \12410 , \11951_nG2e94 , \12125 );
nor \U$11574 ( \12411 , \12408 , \12409 , \12410 );
xor \U$11575 ( \12412 , \12404 , \12411 );
and \U$11576 ( \12413 , \12237_nG2aae , \11834 );
and \U$11577 ( \12414 , \11925 , \12307_nG29cd );
nand \U$11578 ( \12415 , \12237_nG2aae , \11827 );
or \U$11579 ( \12416 , \11795 , \12307_nG29cd );
nand \U$11580 ( \12417 , \12416 , \11831 );
and \U$11581 ( \12418 , \12415 , \12417 );
nor \U$11582 ( \12419 , \12413 , \12414 , \12418 );
and \U$11583 ( \12420 , \12412 , \12419 );
and \U$11584 ( \12421 , \12404 , \12411 );
or \U$11585 ( \12422 , \12420 , \12421 );
not \U$11586 ( \12423 , \12422 );
and \U$11587 ( \12424 , \12397 , \12423 );
not \U$11588 ( \12425 , \12337 );
not \U$11589 ( \12426 , \12339 );
nand \U$11590 ( \12427 , \12426 , \12329 );
not \U$11591 ( \12428 , \12427 );
or \U$11592 ( \12429 , \12425 , \12428 );
or \U$11593 ( \12430 , \12427 , \12337 );
nand \U$11594 ( \12431 , \12429 , \12430 );
not \U$11595 ( \12432 , \12308 );
nor \U$11596 ( \12433 , \12280 , \12311 );
not \U$11597 ( \12434 , \12433 );
or \U$11598 ( \12435 , \12432 , \12434 );
or \U$11599 ( \12436 , \12433 , \12308 );
nand \U$11600 ( \12437 , \12435 , \12436 );
and \U$11601 ( \12438 , \12431 , \12437 );
and \U$11602 ( \12439 , \12424 , \12438 );
xor \U$11603 ( \12440 , \12373 , \12439 );
xnor \U$11604 ( \12441 , \12340 , \12312 );
not \U$11605 ( \12442 , \12350 );
not \U$11606 ( \12443 , \12342 );
and \U$11607 ( \12444 , \12442 , \12443 );
and \U$11608 ( \12445 , \12350 , \12342 );
nor \U$11609 ( \12446 , \12444 , \12445 );
nand \U$11610 ( \12447 , \12441 , \12446 );
and \U$11611 ( \12448 , \12440 , \12447 );
and \U$11612 ( \12449 , \12373 , \12439 );
or \U$11613 ( \12450 , \12448 , \12449 );
xor \U$11614 ( \12451 , \12172 , \12242 );
xor \U$11615 ( \12452 , \12450 , \12451 );
xor \U$11616 ( \12453 , \12352 , \12355 );
xor \U$11617 ( \12454 , \12453 , \12358 );
and \U$11618 ( \12455 , \12452 , \12454 );
and \U$11619 ( \12456 , \12450 , \12451 );
or \U$11620 ( \12457 , \12455 , \12456 );
xor \U$11621 ( \12458 , \12361 , \12363 );
xor \U$11622 ( \12459 , \12458 , \12366 );
xor \U$11623 ( \12460 , \12457 , \12459 );
xor \U$11624 ( \12461 , \12450 , \12451 );
xor \U$11625 ( \12462 , \12461 , \12454 );
xor \U$11626 ( \12463 , \12341 , \12351 );
xor \U$11627 ( \12464 , \12373 , \12439 );
xor \U$11628 ( \12465 , \12464 , \12447 );
and \U$11629 ( \12466 , \12463 , \12465 );
xor \U$11630 ( \12467 , \12397 , \12423 );
xor \U$11631 ( \12468 , \12431 , \12437 );
and \U$11632 ( \12469 , \12467 , \12468 );
xor \U$11633 ( \12470 , \12388 , \12396 );
not \U$11634 ( \12471 , \12470 );
xor \U$11635 ( \12472 , \12404 , \12411 );
xor \U$11636 ( \12473 , \12472 , \12419 );
nor \U$11637 ( \12474 , \12471 , \12473 );
nand \U$11638 ( \12475 , \12237_nG2aae , \11886 );
or \U$11639 ( \12476 , \11848 , \12160_nG2bb5 );
nand \U$11640 ( \12477 , \12476 , \11917 );
and \U$11641 ( \12478 , \12475 , \12477 );
and \U$11642 ( \12479 , \11920 , \12160_nG2bb5 );
and \U$11643 ( \12480 , \12237_nG2aae , \11889 );
nor \U$11644 ( \12481 , \12478 , \12479 , \12480 );
nand \U$11645 ( \12482 , \12076_nG2daa , \12014 );
or \U$11646 ( \12483 , \11964 , \12048_nG2ca8 );
nand \U$11647 ( \12484 , \12483 , \12020 );
and \U$11648 ( \12485 , \12482 , \12484 );
and \U$11649 ( \12486 , \12016 , \12048_nG2ca8 );
and \U$11650 ( \12487 , \12076_nG2daa , \12125 );
nor \U$11651 ( \12488 , \12485 , \12486 , \12487 );
xor \U$11652 ( \12489 , \12481 , \12488 );
and \U$11653 ( \12490 , \12307_nG29cd , \11834 );
and \U$11654 ( \12491 , RIaaa3ae8_420, \7957 );
and \U$11655 ( \12492 , RIaaa3ea8_428, \7944 );
and \U$11656 ( \12493 , \7963 , RIaaa4010_431);
and \U$11657 ( \12494 , RIaaa4178_434, \7930 );
nor \U$11658 ( \12495 , \12493 , \12494 );
and \U$11659 ( \12496 , RIaaa4100_433, \11761 );
and \U$11660 ( \12497 , \7961 , RIaaa3cc8_424);
and \U$11661 ( \12498 , RIaaa3f98_430, \7949 );
nor \U$11662 ( \12499 , \12496 , \12497 , \12498 );
and \U$11663 ( \12500 , \7928 , RIaaa3d40_425);
and \U$11664 ( \12501 , RIaaa3c50_423, \7909 );
nor \U$11665 ( \12502 , \12500 , \12501 );
nand \U$11666 ( \12503 , \12495 , \12499 , \12502 );
nor \U$11667 ( \12504 , \12491 , \12492 , \12503 );
and \U$11668 ( \12505 , \7914 , RIaaa3f20_429);
and \U$11669 ( \12506 , RIaaa3b60_421, \7959 );
nor \U$11670 ( \12507 , \12505 , \12506 );
and \U$11671 ( \12508 , \7942 , RIaaa39f8_418);
and \U$11672 ( \12509 , RIaaa3a70_419, \7919 );
nor \U$11673 ( \12510 , \12508 , \12509 );
and \U$11674 ( \12511 , \7952 , RIaaa3bd8_422);
and \U$11675 ( \12512 , RIaaa3e30_427, \7935 );
nor \U$11676 ( \12513 , \12511 , \12512 );
nand \U$11677 ( \12514 , \12504 , \12507 , \12510 , \12513 );
_DC g28d0 ( \12515_nG28d0 , \12514 , \11781 );
and \U$11678 ( \12516 , \11925 , \12515_nG28d0 );
nand \U$11679 ( \12517 , \12307_nG29cd , \11827 );
or \U$11680 ( \12518 , \11795 , \12515_nG28d0 );
nand \U$11681 ( \12519 , \12518 , \11831 );
and \U$11682 ( \12520 , \12517 , \12519 );
nor \U$11683 ( \12521 , \12490 , \12516 , \12520 );
and \U$11684 ( \12522 , \12489 , \12521 );
and \U$11685 ( \12523 , \12481 , \12488 );
or \U$11686 ( \12524 , \12522 , \12523 );
nand \U$11687 ( \12525 , \11782_nG30bb , \12380 );
or \U$11688 ( \12526 , \12337 , \11821_nG31ca );
or \U$11689 ( \12527 , \12337 , \12379 );
nand \U$11690 ( \12528 , \12526 , \12527 );
and \U$11691 ( \12529 , \12525 , \12528 );
and \U$11692 ( \12530 , \12337 , \12379 );
and \U$11693 ( \12531 , \12530 , \11821_nG31ca );
and \U$11694 ( \12532 , \11782_nG30bb , \12383 );
nor \U$11695 ( \12533 , \12529 , \12531 , \12532 );
xor \U$11696 ( \12534 , RIaaa91a0_605, \11687_nG223f );
xor \U$11697 ( \12535 , \12534 , \11717 );
not \U$11698 ( \12536 , \12535 );
xor \U$11699 ( \12537 , \8308 , \11658_nG22af );
xor \U$11700 ( \12538 , \12537 , \11720 );
not \U$11701 ( \12539 , \12538 );
and \U$11702 ( \12540 , \12536 , \12539 );
or \U$11703 ( \12541 , \12331 , \12540 );
not \U$11704 ( \12542 , \12541 );
xor \U$11705 ( \12543 , \12533 , \12542 );
nand \U$11706 ( \12544 , \11951_nG2e94 , \12179 );
or \U$11707 ( \12545 , \12110 , \11874_nG2fb5 );
nand \U$11708 ( \12546 , \12545 , \12315 );
and \U$11709 ( \12547 , \12544 , \12546 );
and \U$11710 ( \12548 , \12318 , \11874_nG2fb5 );
and \U$11711 ( \12549 , \11951_nG2e94 , \12182 );
nor \U$11712 ( \12550 , \12547 , \12548 , \12549 );
and \U$11713 ( \12551 , \12543 , \12550 );
and \U$11714 ( \12552 , \12533 , \12542 );
or \U$11715 ( \12553 , \12551 , \12552 );
nor \U$11716 ( \12554 , \12524 , \12553 );
and \U$11717 ( \12555 , \12474 , \12554 );
xor \U$11718 ( \12556 , \12469 , \12555 );
or \U$11719 ( \12557 , \12446 , \12441 );
nand \U$11720 ( \12558 , \12557 , \12447 );
and \U$11721 ( \12559 , \12556 , \12558 );
and \U$11722 ( \12560 , \12469 , \12555 );
or \U$11723 ( \12561 , \12559 , \12560 );
xor \U$11724 ( \12562 , \12373 , \12439 );
xor \U$11725 ( \12563 , \12562 , \12447 );
and \U$11726 ( \12564 , \12561 , \12563 );
and \U$11727 ( \12565 , \12463 , \12561 );
or \U$11728 ( \12566 , \12466 , \12564 , \12565 );
xor \U$11729 ( \12567 , \12462 , \12566 );
xor \U$11730 ( \12568 , \12373 , \12439 );
xor \U$11731 ( \12569 , \12568 , \12447 );
xor \U$11732 ( \12570 , \12463 , \12561 );
xor \U$11733 ( \12571 , \12569 , \12570 );
not \U$11734 ( \12572 , \12473 );
not \U$11735 ( \12573 , \12470 );
and \U$11736 ( \12574 , \12572 , \12573 );
and \U$11737 ( \12575 , \12473 , \12470 );
nor \U$11738 ( \12576 , \12574 , \12575 );
not \U$11739 ( \12577 , \12515_nG28d0 );
nor \U$11740 ( \12578 , \11755 , \12577 );
or \U$11741 ( \12579 , \12576 , \12578 );
xnor \U$11742 ( \12580 , \12553 , \12524 );
nand \U$11743 ( \12581 , \12579 , \12580 );
or \U$11744 ( \12582 , \12331 , \12538 );
nand \U$11745 ( \12583 , \12538 , \12331 );
nand \U$11746 ( \12584 , \12582 , \12583 );
xor \U$11747 ( \12585 , \12536 , \12539 );
nor \U$11748 ( \12586 , \12584 , \12585 );
not \U$11749 ( \12587 , \12586 );
nor \U$11750 ( \12588 , \12587 , \12542 );
not \U$11751 ( \12589 , \12588 );
or \U$11752 ( \12590 , \12589 , \11823 );
or \U$11753 ( \12591 , \12587 , \11823 );
nand \U$11754 ( \12592 , \12591 , \12542 );
nand \U$11755 ( \12593 , \12590 , \12592 );
or \U$11756 ( \12594 , \12384 , \11896 );
not \U$11757 ( \12595 , \12530 );
or \U$11758 ( \12596 , \11783 , \12595 );
or \U$11759 ( \12597 , \12381 , \11896 );
or \U$11760 ( \12598 , \12337 , \11782_nG30bb );
nand \U$11761 ( \12599 , \12598 , \12527 );
nand \U$11762 ( \12600 , \12597 , \12599 );
nand \U$11763 ( \12601 , \12594 , \12596 , \12600 );
and \U$11764 ( \12602 , \12593 , \12601 );
not \U$11765 ( \12603 , \12602 );
not \U$11766 ( \12604 , \12307_nG29cd );
or \U$11767 ( \12605 , \11890 , \12604 );
or \U$11768 ( \12606 , \11848 , \12237_nG2aae );
nand \U$11769 ( \12607 , \12606 , \11917 );
nand \U$11770 ( \12608 , \12307_nG29cd , \11886 );
and \U$11771 ( \12609 , \12607 , \12608 );
and \U$11772 ( \12610 , \12237_nG2aae , \11920 );
nor \U$11773 ( \12611 , \12609 , \12610 );
nand \U$11774 ( \12612 , \12605 , \12611 );
nand \U$11775 ( \12613 , \12076_nG2daa , \12179 );
or \U$11776 ( \12614 , \12110 , \11951_nG2e94 );
nand \U$11777 ( \12615 , \12614 , \12315 );
and \U$11778 ( \12616 , \12613 , \12615 );
and \U$11779 ( \12617 , \12318 , \11951_nG2e94 );
and \U$11780 ( \12618 , \12076_nG2daa , \12182 );
nor \U$11781 ( \12619 , \12616 , \12617 , \12618 );
nand \U$11782 ( \12620 , \12048_nG2ca8 , \12014 );
or \U$11783 ( \12621 , \11964 , \12160_nG2bb5 );
nand \U$11784 ( \12622 , \12621 , \12020 );
and \U$11785 ( \12623 , \12620 , \12622 );
and \U$11786 ( \12624 , \12016 , \12160_nG2bb5 );
and \U$11787 ( \12625 , \12048_nG2ca8 , \12125 );
nor \U$11788 ( \12626 , \12623 , \12624 , \12625 );
nand \U$11789 ( \12627 , \12619 , \12626 );
and \U$11790 ( \12628 , \12612 , \12627 );
nor \U$11791 ( \12629 , \12626 , \12619 );
nor \U$11792 ( \12630 , \12628 , \12629 );
nor \U$11793 ( \12631 , \12603 , \12630 );
xor \U$11794 ( \12632 , \12481 , \12488 );
xor \U$11795 ( \12633 , \12632 , \12521 );
xor \U$11796 ( \12634 , \12533 , \12542 );
xor \U$11797 ( \12635 , \12634 , \12550 );
nor \U$11798 ( \12636 , \12633 , \12635 );
not \U$11799 ( \12637 , \12636 );
and \U$11800 ( \12638 , RIaaa33e0_405, \7949 );
and \U$11801 ( \12639 , RIaaa36b0_411, \7909 );
and \U$11802 ( \12640 , \7930 , RIaaa35c0_409);
and \U$11803 ( \12641 , RIaaa32f0_403, \7944 );
nor \U$11804 ( \12642 , \12640 , \12641 );
and \U$11805 ( \12643 , RIaaa3548_408, \11761 );
and \U$11806 ( \12644 , \7942 , RIaaa3818_414);
and \U$11807 ( \12645 , RIaaa3908_416, \7961 );
nor \U$11808 ( \12646 , \12643 , \12644 , \12645 );
and \U$11809 ( \12647 , \7928 , RIaaa3980_417);
and \U$11810 ( \12648 , RIaaa3728_412, \7957 );
nor \U$11811 ( \12649 , \12647 , \12648 );
nand \U$11812 ( \12650 , \12642 , \12646 , \12649 );
nor \U$11813 ( \12651 , \12638 , \12639 , \12650 );
and \U$11814 ( \12652 , \7919 , RIaaa3890_415);
and \U$11815 ( \12653 , RIaaa37a0_413, \7959 );
nor \U$11816 ( \12654 , \12652 , \12653 );
and \U$11817 ( \12655 , \7914 , RIaaa3368_404);
and \U$11818 ( \12656 , RIaaa3278_402, \7935 );
nor \U$11819 ( \12657 , \12655 , \12656 );
and \U$11820 ( \12658 , \7952 , RIaaa3638_410);
and \U$11821 ( \12659 , RIaaa3458_406, \7963 );
nor \U$11822 ( \12660 , \12658 , \12659 );
nand \U$11823 ( \12661 , \12651 , \12654 , \12657 , \12660 );
_DC g27f3 ( \12662_nG27f3 , \12661 , \11781 );
nand \U$11824 ( \12663 , \12662_nG27f3 , \11754 );
nand \U$11825 ( \12664 , \12637 , \12663 );
and \U$11826 ( \12665 , \12631 , \12664 );
xor \U$11827 ( \12666 , \12581 , \12665 );
xor \U$11828 ( \12667 , \12467 , \12468 );
and \U$11829 ( \12668 , \12666 , \12667 );
and \U$11830 ( \12669 , \12581 , \12665 );
or \U$11831 ( \12670 , \12668 , \12669 );
xor \U$11832 ( \12671 , \12424 , \12438 );
xor \U$11833 ( \12672 , \12670 , \12671 );
xor \U$11834 ( \12673 , \12469 , \12555 );
xor \U$11835 ( \12674 , \12673 , \12558 );
and \U$11836 ( \12675 , \12672 , \12674 );
and \U$11837 ( \12676 , \12670 , \12671 );
or \U$11838 ( \12677 , \12675 , \12676 );
xor \U$11839 ( \12678 , \12571 , \12677 );
xor \U$11840 ( \12679 , \12670 , \12671 );
xor \U$11841 ( \12680 , \12679 , \12674 );
or \U$11842 ( \12681 , \12630 , \12602 );
and \U$11843 ( \12682 , RIaaa4808_448, \7957 );
and \U$11844 ( \12683 , RIaaa44c0_441, \7944 );
and \U$11845 ( \12684 , \7963 , RIaaa45b0_443);
and \U$11846 ( \12685 , RIaaa4358_438, \7930 );
nor \U$11847 ( \12686 , \12684 , \12685 );
and \U$11848 ( \12687 , RIaaa42e0_437, \11761 );
and \U$11849 ( \12688 , \7961 , RIaaa4718_446);
and \U$11850 ( \12689 , RIaaa4538_442, \7949 );
nor \U$11851 ( \12690 , \12687 , \12688 , \12689 );
and \U$11852 ( \12691 , \7928 , RIaaa4790_447);
and \U$11853 ( \12692 , RIaaa4970_451, \7909 );
nor \U$11854 ( \12693 , \12691 , \12692 );
nand \U$11855 ( \12694 , \12686 , \12690 , \12693 );
nor \U$11856 ( \12695 , \12682 , \12683 , \12694 );
and \U$11857 ( \12696 , \7914 , RIaaa4448_440);
and \U$11858 ( \12697 , RIaaa4880_449, \7959 );
nor \U$11859 ( \12698 , \12696 , \12697 );
and \U$11860 ( \12699 , \7942 , RIaaa4628_444);
and \U$11861 ( \12700 , RIaaa46a0_445, \7919 );
nor \U$11862 ( \12701 , \12699 , \12700 );
and \U$11863 ( \12702 , \7952 , RIaaa48f8_450);
and \U$11864 ( \12703 , RIaaa43d0_439, \7935 );
nor \U$11865 ( \12704 , \12702 , \12703 );
nand \U$11866 ( \12705 , \12695 , \12698 , \12701 , \12704 );
_DC g2723 ( \12706_nG2723 , \12705 , \11781 );
nand \U$11867 ( \12707 , \12706_nG2723 , \11754 );
and \U$11868 ( \12708 , \12515_nG28d0 , \11834 );
and \U$11869 ( \12709 , \11925 , \12662_nG27f3 );
nand \U$11870 ( \12710 , \12515_nG28d0 , \11827 );
or \U$11871 ( \12711 , \11795 , \12662_nG27f3 );
nand \U$11872 ( \12712 , \12711 , \11831 );
and \U$11873 ( \12713 , \12710 , \12712 );
nor \U$11874 ( \12714 , \12708 , \12709 , \12713 );
or \U$11875 ( \12715 , \12707 , \12714 );
nand \U$11876 ( \12716 , \12602 , \12630 );
nand \U$11877 ( \12717 , \12681 , \12715 , \12716 );
not \U$11878 ( \12718 , \12663 );
and \U$11879 ( \12719 , \12633 , \12635 );
nor \U$11880 ( \12720 , \12719 , \12636 );
not \U$11881 ( \12721 , \12720 );
or \U$11882 ( \12722 , \12718 , \12721 );
or \U$11883 ( \12723 , \12720 , \12663 );
nand \U$11884 ( \12724 , \12722 , \12723 );
and \U$11885 ( \12725 , \12717 , \12724 );
nand \U$11886 ( \12726 , \12160_nG2bb5 , \12014 );
or \U$11887 ( \12727 , \11964 , \12237_nG2aae );
nand \U$11888 ( \12728 , \12727 , \12020 );
and \U$11889 ( \12729 , \12726 , \12728 );
and \U$11890 ( \12730 , \12016 , \12237_nG2aae );
and \U$11891 ( \12731 , \12160_nG2bb5 , \12125 );
nor \U$11892 ( \12732 , \12729 , \12730 , \12731 );
nand \U$11893 ( \12733 , \12048_nG2ca8 , \12179 );
or \U$11894 ( \12734 , \12110 , \12076_nG2daa );
nand \U$11895 ( \12735 , \12734 , \12315 );
and \U$11896 ( \12736 , \12733 , \12735 );
and \U$11897 ( \12737 , \12318 , \12076_nG2daa );
and \U$11898 ( \12738 , \12048_nG2ca8 , \12182 );
nor \U$11899 ( \12739 , \12736 , \12737 , \12738 );
xor \U$11900 ( \12740 , \12732 , \12739 );
nand \U$11901 ( \12741 , \12515_nG28d0 , \11886 );
or \U$11902 ( \12742 , \11848 , \12307_nG29cd );
nand \U$11903 ( \12743 , \12742 , \11917 );
and \U$11904 ( \12744 , \12741 , \12743 );
and \U$11905 ( \12745 , \11920 , \12307_nG29cd );
and \U$11906 ( \12746 , \12515_nG28d0 , \11889 );
nor \U$11907 ( \12747 , \12744 , \12745 , \12746 );
and \U$11908 ( \12748 , \12740 , \12747 );
and \U$11909 ( \12749 , \12732 , \12739 );
or \U$11910 ( \12750 , \12748 , \12749 );
nand \U$11911 ( \12751 , \11782_nG30bb , \12586 );
or \U$11912 ( \12752 , \12541 , \11821_nG31ca );
or \U$11913 ( \12753 , \12541 , \12585 );
nand \U$11914 ( \12754 , \12752 , \12753 );
and \U$11915 ( \12755 , \12751 , \12754 );
and \U$11916 ( \12756 , \12541 , \12585 );
and \U$11917 ( \12757 , \12756 , \11821_nG31ca );
and \U$11918 ( \12758 , \11782_nG30bb , \12588 );
nor \U$11919 ( \12759 , \12755 , \12757 , \12758 );
xor \U$11920 ( \12760 , \12759 , \12536 );
nand \U$11921 ( \12761 , \11951_nG2e94 , \12380 );
or \U$11922 ( \12762 , \12337 , \11874_nG2fb5 );
nand \U$11923 ( \12763 , \12762 , \12527 );
and \U$11924 ( \12764 , \12761 , \12763 );
and \U$11925 ( \12765 , \12530 , \11874_nG2fb5 );
and \U$11926 ( \12766 , \11951_nG2e94 , \12383 );
nor \U$11927 ( \12767 , \12764 , \12765 , \12766 );
and \U$11928 ( \12768 , \12760 , \12767 );
and \U$11929 ( \12769 , \12759 , \12536 );
or \U$11930 ( \12770 , \12768 , \12769 );
nor \U$11931 ( \12771 , \12750 , \12770 );
not \U$11932 ( \12772 , \12629 );
nand \U$11933 ( \12773 , \12772 , \12627 );
not \U$11934 ( \12774 , \12773 );
not \U$11935 ( \12775 , \12612 );
or \U$11936 ( \12776 , \12774 , \12775 );
or \U$11937 ( \12777 , \12612 , \12773 );
nand \U$11938 ( \12778 , \12776 , \12777 );
xor \U$11939 ( \12779 , \12593 , \12601 );
xor \U$11940 ( \12780 , \12778 , \12779 );
xor \U$11941 ( \12781 , \12707 , \12714 );
and \U$11942 ( \12782 , \12780 , \12781 );
and \U$11943 ( \12783 , \12778 , \12779 );
or \U$11944 ( \12784 , \12782 , \12783 );
and \U$11945 ( \12785 , \12771 , \12784 );
xor \U$11946 ( \12786 , \12725 , \12785 );
not \U$11947 ( \12787 , \12580 );
xor \U$11948 ( \12788 , \12578 , \12576 );
not \U$11949 ( \12789 , \12788 );
or \U$11950 ( \12790 , \12787 , \12789 );
or \U$11951 ( \12791 , \12788 , \12580 );
nand \U$11952 ( \12792 , \12790 , \12791 );
and \U$11953 ( \12793 , \12786 , \12792 );
and \U$11954 ( \12794 , \12725 , \12785 );
or \U$11955 ( \12795 , \12793 , \12794 );
nor \U$11956 ( \12796 , \12554 , \12578 );
not \U$11957 ( \12797 , \12796 );
not \U$11958 ( \12798 , \12474 );
or \U$11959 ( \12799 , \12797 , \12798 );
or \U$11960 ( \12800 , \12474 , \12796 );
nand \U$11961 ( \12801 , \12799 , \12800 );
xor \U$11962 ( \12802 , \12795 , \12801 );
xor \U$11963 ( \12803 , \12581 , \12665 );
xor \U$11964 ( \12804 , \12803 , \12667 );
and \U$11965 ( \12805 , \12802 , \12804 );
and \U$11966 ( \12806 , \12795 , \12801 );
or \U$11967 ( \12807 , \12805 , \12806 );
xor \U$11968 ( \12808 , \12680 , \12807 );
xor \U$11969 ( \12809 , \12795 , \12801 );
xor \U$11970 ( \12810 , \12809 , \12804 );
xor \U$11971 ( \12811 , \12717 , \12724 );
xor \U$11972 ( \12812 , \12771 , \12784 );
xor \U$11973 ( \12813 , \12811 , \12812 );
nand \U$11974 ( \12814 , \12160_nG2bb5 , \12179 );
or \U$11975 ( \12815 , \12110 , \12048_nG2ca8 );
nand \U$11976 ( \12816 , \12815 , \12315 );
and \U$11977 ( \12817 , \12814 , \12816 );
and \U$11978 ( \12818 , \12318 , \12048_nG2ca8 );
and \U$11979 ( \12819 , \12160_nG2bb5 , \12182 );
nor \U$11980 ( \12820 , \12817 , \12818 , \12819 );
nand \U$11981 ( \12821 , \12076_nG2daa , \12380 );
or \U$11982 ( \12822 , \12337 , \11951_nG2e94 );
nand \U$11983 ( \12823 , \12822 , \12527 );
and \U$11984 ( \12824 , \12821 , \12823 );
and \U$11985 ( \12825 , \12530 , \11951_nG2e94 );
and \U$11986 ( \12826 , \12076_nG2daa , \12383 );
nor \U$11987 ( \12827 , \12824 , \12825 , \12826 );
xor \U$11988 ( \12828 , \12820 , \12827 );
nand \U$11989 ( \12829 , \12237_nG2aae , \12014 );
or \U$11990 ( \12830 , \11964 , \12307_nG29cd );
nand \U$11991 ( \12831 , \12830 , \12020 );
and \U$11992 ( \12832 , \12829 , \12831 );
and \U$11993 ( \12833 , \12016 , \12307_nG29cd );
and \U$11994 ( \12834 , \12237_nG2aae , \12125 );
nor \U$11995 ( \12835 , \12832 , \12833 , \12834 );
and \U$11996 ( \12836 , \12828 , \12835 );
and \U$11997 ( \12837 , \12820 , \12827 );
or \U$11998 ( \12838 , \12836 , \12837 );
nand \U$11999 ( \12839 , \11874_nG2fb5 , \12586 );
or \U$12000 ( \12840 , \12541 , \11782_nG30bb );
nand \U$12001 ( \12841 , \12840 , \12753 );
and \U$12002 ( \12842 , \12839 , \12841 );
and \U$12003 ( \12843 , \12756 , \11782_nG30bb );
and \U$12004 ( \12844 , \11874_nG2fb5 , \12588 );
nor \U$12005 ( \12845 , \12842 , \12843 , \12844 );
not \U$12006 ( \12846 , \12845 );
or \U$12007 ( \12847 , \12535 , \11821_nG31ca );
or \U$12008 ( \12848 , \8403 , \11715_nG223d );
nand \U$12009 ( \12849 , \12848 , \11716 );
nor \U$12010 ( \12850 , \12535 , \12849 );
not \U$12011 ( \12851 , \12850 );
nand \U$12012 ( \12852 , \12536 , \12851 );
nand \U$12013 ( \12853 , \12847 , \12852 );
nand \U$12014 ( \12854 , \12846 , \12853 );
xor \U$12015 ( \12855 , \12838 , \12854 );
and \U$12016 ( \12856 , \12706_nG2723 , \11834 );
and \U$12017 ( \12857 , RIaaa6860_517, \7942 );
and \U$12018 ( \12858 , RIaaa6428_508, \7914 );
and \U$12019 ( \12859 , \7963 , RIaaa6518_510);
and \U$12020 ( \12860 , RIaaa6338_506, \7930 );
nor \U$12021 ( \12861 , \12859 , \12860 );
and \U$12022 ( \12862 , RIaaa62c0_505, \11761 );
and \U$12023 ( \12863 , \7961 , RIaaa68d8_518);
and \U$12024 ( \12864 , RIaaa6590_511, \7949 );
nor \U$12025 ( \12865 , \12862 , \12863 , \12864 );
and \U$12026 ( \12866 , \7928 , RIaaa6950_519);
and \U$12027 ( \12867 , RIaaa6770_515, \7909 );
nor \U$12028 ( \12868 , \12866 , \12867 );
nand \U$12029 ( \12869 , \12861 , \12865 , \12868 );
nor \U$12030 ( \12870 , \12857 , \12858 , \12869 );
and \U$12031 ( \12871 , \7957 , RIaaa6680_513);
and \U$12032 ( \12872 , RIaaa64a0_509, \7944 );
nor \U$12033 ( \12873 , \12871 , \12872 );
and \U$12034 ( \12874 , \7935 , RIaaa63b0_507);
and \U$12035 ( \12875 , RIaaa67e8_516, \7919 );
nor \U$12036 ( \12876 , \12874 , \12875 );
and \U$12037 ( \12877 , \7952 , RIaaa66f8_514);
and \U$12038 ( \12878 , RIaaa6608_512, \7959 );
nor \U$12039 ( \12879 , \12877 , \12878 );
nand \U$12040 ( \12880 , \12870 , \12873 , \12876 , \12879 );
_DC g23c5 ( \12881_nG23c5 , \12880 , \11781 );
and \U$12041 ( \12882 , \11925 , \12881_nG23c5 );
nand \U$12042 ( \12883 , \12706_nG2723 , \11827 );
or \U$12043 ( \12884 , \11795 , \12881_nG23c5 );
nand \U$12044 ( \12885 , \12884 , \11831 );
and \U$12045 ( \12886 , \12883 , \12885 );
nor \U$12046 ( \12887 , \12856 , \12882 , \12886 );
nand \U$12047 ( \12888 , \12662_nG27f3 , \11886 );
or \U$12048 ( \12889 , \11848 , \12515_nG28d0 );
nand \U$12049 ( \12890 , \12889 , \11917 );
and \U$12050 ( \12891 , \12888 , \12890 );
and \U$12051 ( \12892 , \11920 , \12515_nG28d0 );
and \U$12052 ( \12893 , \12662_nG27f3 , \11889 );
nor \U$12053 ( \12894 , \12891 , \12892 , \12893 );
and \U$12054 ( \12895 , \12887 , \12894 );
not \U$12055 ( \12896 , \12895 );
and \U$12056 ( \12897 , \7930 , RIaaa5528_476);
and \U$12057 ( \12898 , \7952 , RIaaa57f8_482);
and \U$12058 ( \12899 , RIaaa5708_480, \7957 );
nor \U$12059 ( \12900 , \12898 , \12899 );
and \U$12060 ( \12901 , \7942 , RIaaa5618_478);
and \U$12061 ( \12902 , RIaaa52d0_471, \7944 );
nor \U$12062 ( \12903 , \12901 , \12902 );
and \U$12063 ( \12904 , \7914 , RIaaa5348_472);
and \U$12064 ( \12905 , RIaaa5258_470, \7935 );
nor \U$12065 ( \12906 , \12904 , \12905 );
and \U$12066 ( \12907 , \7919 , RIaaa5690_479);
and \U$12067 ( \12908 , RIaaa5780_481, \7959 );
nor \U$12068 ( \12909 , \12907 , \12908 );
nand \U$12069 ( \12910 , \12900 , \12903 , \12906 , \12909 );
nor \U$12070 ( \12911 , \12897 , \12910 );
and \U$12071 ( \12912 , \7961 , RIaaa5960_485);
and \U$12072 ( \12913 , RIaaa5438_474, \7963 );
nor \U$12073 ( \12914 , \12912 , \12913 );
and \U$12074 ( \12915 , \7928 , RIaaa58e8_484);
and \U$12075 ( \12916 , RIaaa5870_483, \7909 );
nor \U$12076 ( \12917 , \12915 , \12916 );
and \U$12077 ( \12918 , \11761 , RIaaa55a0_477);
and \U$12078 ( \12919 , RIaaa53c0_473, \7949 );
nor \U$12079 ( \12920 , \12918 , \12919 );
nand \U$12080 ( \12921 , \12911 , \12914 , \12917 , \12920 );
_DC g2391 ( \12922_nG2391 , \12921 , \11781 );
nand \U$12081 ( \12923 , \12922_nG2391 , \11754 );
not \U$12082 ( \12924 , \12923 );
and \U$12083 ( \12925 , \12896 , \12924 );
nor \U$12084 ( \12926 , \12887 , \12894 );
nor \U$12085 ( \12927 , \12925 , \12926 );
and \U$12086 ( \12928 , \12855 , \12927 );
and \U$12087 ( \12929 , \12838 , \12854 );
or \U$12088 ( \12930 , \12928 , \12929 );
nand \U$12089 ( \12931 , \12881_nG23c5 , \11754 );
and \U$12090 ( \12932 , \12662_nG27f3 , \11834 );
and \U$12091 ( \12933 , \11925 , \12706_nG2723 );
nand \U$12092 ( \12934 , \12662_nG27f3 , \11827 );
or \U$12093 ( \12935 , \11795 , \12706_nG2723 );
nand \U$12094 ( \12936 , \12935 , \11831 );
and \U$12095 ( \12937 , \12934 , \12936 );
nor \U$12096 ( \12938 , \12932 , \12933 , \12937 );
xor \U$12097 ( \12939 , \12931 , \12938 );
not \U$12098 ( \12940 , \12939 );
or \U$12099 ( \12941 , \12930 , \12940 );
not \U$12100 ( \12942 , \12940 );
not \U$12101 ( \12943 , \12930 );
or \U$12102 ( \12944 , \12942 , \12943 );
xor \U$12103 ( \12945 , \12778 , \12779 );
xor \U$12104 ( \12946 , \12945 , \12781 );
nand \U$12105 ( \12947 , \12944 , \12946 );
nand \U$12106 ( \12948 , \12941 , \12947 );
and \U$12107 ( \12949 , \12813 , \12948 );
and \U$12108 ( \12950 , \12811 , \12812 );
or \U$12109 ( \12951 , \12949 , \12950 );
xor \U$12110 ( \12952 , \12631 , \12664 );
xor \U$12111 ( \12953 , \12951 , \12952 );
xor \U$12112 ( \12954 , \12725 , \12785 );
xor \U$12113 ( \12955 , \12954 , \12792 );
and \U$12114 ( \12956 , \12953 , \12955 );
and \U$12115 ( \12957 , \12951 , \12952 );
or \U$12116 ( \12958 , \12956 , \12957 );
xor \U$12117 ( \12959 , \12810 , \12958 );
xor \U$12118 ( \12960 , \12951 , \12952 );
xor \U$12119 ( \12961 , \12960 , \12955 );
not \U$12120 ( \12962 , \12770 );
or \U$12121 ( \12963 , \12750 , \12962 );
not \U$12122 ( \12964 , \12750 );
or \U$12123 ( \12965 , \12770 , \12964 );
or \U$12124 ( \12966 , \12931 , \12938 );
nand \U$12125 ( \12967 , \12963 , \12965 , \12966 );
not \U$12126 ( \12968 , \12967 );
and \U$12127 ( \12969 , \12946 , \12939 );
not \U$12128 ( \12970 , \12946 );
and \U$12129 ( \12971 , \12970 , \12940 );
nor \U$12130 ( \12972 , \12969 , \12971 );
not \U$12131 ( \12973 , \12972 );
not \U$12132 ( \12974 , \12930 );
and \U$12133 ( \12975 , \12973 , \12974 );
and \U$12134 ( \12976 , \12972 , \12930 );
nor \U$12135 ( \12977 , \12975 , \12976 );
nor \U$12136 ( \12978 , \12968 , \12977 );
nand \U$12137 ( \12979 , \12307_nG29cd , \12014 );
or \U$12138 ( \12980 , \11964 , \12515_nG28d0 );
nand \U$12139 ( \12981 , \12980 , \12020 );
and \U$12140 ( \12982 , \12979 , \12981 );
and \U$12141 ( \12983 , \12016 , \12515_nG28d0 );
and \U$12142 ( \12984 , \12307_nG29cd , \12125 );
nor \U$12143 ( \12985 , \12982 , \12983 , \12984 );
nand \U$12144 ( \12986 , \12237_nG2aae , \12179 );
or \U$12145 ( \12987 , \12110 , \12160_nG2bb5 );
nand \U$12146 ( \12988 , \12987 , \12315 );
and \U$12147 ( \12989 , \12986 , \12988 );
and \U$12148 ( \12990 , \12318 , \12160_nG2bb5 );
and \U$12149 ( \12991 , \12237_nG2aae , \12182 );
nor \U$12150 ( \12992 , \12989 , \12990 , \12991 );
xor \U$12151 ( \12993 , \12985 , \12992 );
nand \U$12152 ( \12994 , \12706_nG2723 , \11886 );
or \U$12153 ( \12995 , \11848 , \12662_nG27f3 );
nand \U$12154 ( \12996 , \12995 , \11917 );
and \U$12155 ( \12997 , \12994 , \12996 );
and \U$12156 ( \12998 , \11920 , \12662_nG27f3 );
and \U$12157 ( \12999 , \12706_nG2723 , \11889 );
nor \U$12158 ( \13000 , \12997 , \12998 , \12999 );
and \U$12159 ( \13001 , \12993 , \13000 );
and \U$12160 ( \13002 , \12985 , \12992 );
or \U$12161 ( \13003 , \13001 , \13002 );
nand \U$12162 ( \13004 , \11951_nG2e94 , \12586 );
or \U$12163 ( \13005 , \12541 , \11874_nG2fb5 );
nand \U$12164 ( \13006 , \13005 , \12753 );
and \U$12165 ( \13007 , \13004 , \13006 );
and \U$12166 ( \13008 , \12756 , \11874_nG2fb5 );
and \U$12167 ( \13009 , \11951_nG2e94 , \12588 );
nor \U$12168 ( \13010 , \13007 , \13008 , \13009 );
not \U$12169 ( \13011 , \13010 );
not \U$12170 ( \13012 , \12852 );
and \U$12171 ( \13013 , \11823 , \13012 );
and \U$12172 ( \13014 , \12850 , \11783 );
and \U$12173 ( \13015 , \12535 , \12849 );
and \U$12174 ( \13016 , \11821_nG31ca , \13015 );
nor \U$12175 ( \13017 , \13013 , \13014 , \13016 );
not \U$12176 ( \13018 , \13017 );
and \U$12177 ( \13019 , \13011 , \13018 );
and \U$12178 ( \13020 , \13010 , \13017 );
nand \U$12179 ( \13021 , \12048_nG2ca8 , \12380 );
or \U$12180 ( \13022 , \12337 , \12076_nG2daa );
nand \U$12181 ( \13023 , \13022 , \12527 );
and \U$12182 ( \13024 , \13021 , \13023 );
and \U$12183 ( \13025 , \12530 , \12076_nG2daa );
and \U$12184 ( \13026 , \12048_nG2ca8 , \12383 );
nor \U$12185 ( \13027 , \13024 , \13025 , \13026 );
nor \U$12186 ( \13028 , \13020 , \13027 );
nor \U$12187 ( \13029 , \13019 , \13028 );
nor \U$12188 ( \13030 , \13003 , \13029 );
xor \U$12189 ( \13031 , \12732 , \12739 );
xor \U$12190 ( \13032 , \13031 , \12747 );
not \U$12191 ( \13033 , \13032 );
xor \U$12192 ( \13034 , \13030 , \13033 );
not \U$12193 ( \13035 , \12923 );
nor \U$12194 ( \13036 , \12895 , \12926 );
not \U$12195 ( \13037 , \13036 );
or \U$12196 ( \13038 , \13035 , \13037 );
or \U$12197 ( \13039 , \13036 , \12923 );
nand \U$12198 ( \13040 , \13038 , \13039 );
not \U$12199 ( \13041 , \13040 );
xor \U$12200 ( \13042 , \12820 , \12827 );
xor \U$12201 ( \13043 , \13042 , \12835 );
nor \U$12202 ( \13044 , \13041 , \13043 );
and \U$12203 ( \13045 , \13034 , \13044 );
and \U$12204 ( \13046 , \13030 , \13033 );
or \U$12205 ( \13047 , \13045 , \13046 );
not \U$12206 ( \13048 , \13047 );
xor \U$12207 ( \13049 , \12759 , \12536 );
xor \U$12208 ( \13050 , \13049 , \12767 );
xor \U$12209 ( \13051 , \12939 , \13050 );
xor \U$12210 ( \13052 , \12838 , \12854 );
xor \U$12211 ( \13053 , \13052 , \12927 );
and \U$12212 ( \13054 , \13051 , \13053 );
and \U$12213 ( \13055 , \12939 , \13050 );
or \U$12214 ( \13056 , \13054 , \13055 );
nand \U$12215 ( \13057 , \13048 , \13056 );
xor \U$12216 ( \13058 , \12978 , \13057 );
xor \U$12217 ( \13059 , \12811 , \12812 );
xor \U$12218 ( \13060 , \13059 , \12948 );
and \U$12219 ( \13061 , \13058 , \13060 );
and \U$12220 ( \13062 , \12978 , \13057 );
or \U$12221 ( \13063 , \13061 , \13062 );
xor \U$12222 ( \13064 , \12961 , \13063 );
xor \U$12223 ( \13065 , \12939 , \13050 );
xor \U$12224 ( \13066 , \13065 , \13053 );
not \U$12225 ( \13067 , \12845 );
not \U$12226 ( \13068 , \12853 );
and \U$12227 ( \13069 , \13067 , \13068 );
and \U$12228 ( \13070 , \12845 , \12853 );
nor \U$12229 ( \13071 , \13069 , \13070 );
nand \U$12230 ( \13072 , \12307_nG29cd , \12179 );
or \U$12231 ( \13073 , \12110 , \12237_nG2aae );
nand \U$12232 ( \13074 , \13073 , \12315 );
and \U$12233 ( \13075 , \13072 , \13074 );
and \U$12234 ( \13076 , \12318 , \12237_nG2aae );
and \U$12235 ( \13077 , \12307_nG29cd , \12182 );
nor \U$12236 ( \13078 , \13075 , \13076 , \13077 );
nand \U$12237 ( \13079 , \12160_nG2bb5 , \12380 );
or \U$12238 ( \13080 , \12337 , \12048_nG2ca8 );
nand \U$12239 ( \13081 , \13080 , \12527 );
and \U$12240 ( \13082 , \13079 , \13081 );
and \U$12241 ( \13083 , \12530 , \12048_nG2ca8 );
and \U$12242 ( \13084 , \12160_nG2bb5 , \12383 );
nor \U$12243 ( \13085 , \13082 , \13083 , \13084 );
xor \U$12244 ( \13086 , \13078 , \13085 );
nand \U$12245 ( \13087 , \12515_nG28d0 , \12014 );
or \U$12246 ( \13088 , \11964 , \12662_nG27f3 );
nand \U$12247 ( \13089 , \13088 , \12020 );
and \U$12248 ( \13090 , \13087 , \13089 );
and \U$12249 ( \13091 , \12016 , \12662_nG27f3 );
and \U$12250 ( \13092 , \12515_nG28d0 , \12125 );
nor \U$12251 ( \13093 , \13090 , \13091 , \13092 );
and \U$12252 ( \13094 , \13086 , \13093 );
and \U$12253 ( \13095 , \13078 , \13085 );
or \U$12254 ( \13096 , \13094 , \13095 );
and \U$12255 ( \13097 , \12922_nG2391 , \11834 );
and \U$12256 ( \13098 , RIaaa50f0_467, \7957 );
and \U$12257 ( \13099 , RIaaa4f88_464, \7944 );
and \U$12258 ( \13100 , \7963 , RIaaa4f10_463);
and \U$12259 ( \13101 , RIaaa4c40_457, \7930 );
nor \U$12260 ( \13102 , \13100 , \13101 );
and \U$12261 ( \13103 , RIaaa4bc8_456, \11761 );
and \U$12262 ( \13104 , \7961 , RIaaa4d30_459);
and \U$12263 ( \13105 , RIaaa4da8_460, \7949 );
nor \U$12264 ( \13106 , \13103 , \13104 , \13105 );
and \U$12265 ( \13107 , \7928 , RIaaa4cb8_458);
and \U$12266 ( \13108 , RIaaa4a60_453, \7909 );
nor \U$12267 ( \13109 , \13107 , \13108 );
nand \U$12268 ( \13110 , \13102 , \13106 , \13109 );
nor \U$12269 ( \13111 , \13098 , \13099 , \13110 );
and \U$12270 ( \13112 , \7914 , RIaaa5078_466);
and \U$12271 ( \13113 , RIaaa5168_468, \7959 );
nor \U$12272 ( \13114 , \13112 , \13113 );
and \U$12273 ( \13115 , \7942 , RIaaa4e98_462);
and \U$12274 ( \13116 , RIaaa4e20_461, \7919 );
nor \U$12275 ( \13117 , \13115 , \13116 );
and \U$12276 ( \13118 , \7952 , RIaaa49e8_452);
and \U$12277 ( \13119 , RIaaa5000_465, \7935 );
nor \U$12278 ( \13120 , \13118 , \13119 );
nand \U$12279 ( \13121 , \13111 , \13114 , \13117 , \13120 );
_DC g2354 ( \13122_nG2354 , \13121 , \11781 );
and \U$12280 ( \13123 , \11925 , \13122_nG2354 );
nand \U$12281 ( \13124 , \12922_nG2391 , \11827 );
or \U$12282 ( \13125 , \11795 , \13122_nG2354 );
nand \U$12283 ( \13126 , \13125 , \11831 );
and \U$12284 ( \13127 , \13124 , \13126 );
nor \U$12285 ( \13128 , \13097 , \13123 , \13127 );
nand \U$12286 ( \13129 , \12881_nG23c5 , \11886 );
or \U$12287 ( \13130 , \11848 , \12706_nG2723 );
nand \U$12288 ( \13131 , \13130 , \11917 );
and \U$12289 ( \13132 , \13129 , \13131 );
and \U$12290 ( \13133 , \11920 , \12706_nG2723 );
and \U$12291 ( \13134 , \12881_nG23c5 , \11889 );
nor \U$12292 ( \13135 , \13132 , \13133 , \13134 );
and \U$12293 ( \13136 , \13128 , \13135 );
not \U$12294 ( \13137 , \13136 );
and \U$12295 ( \13138 , RIaaa60e0_501, \7957 );
and \U$12296 ( \13139 , RIaaa5b40_489, \7944 );
and \U$12297 ( \13140 , \7963 , RIaaa5ac8_488);
and \U$12298 ( \13141 , RIaaa5f00_497, \7930 );
nor \U$12299 ( \13142 , \13140 , \13141 );
and \U$12300 ( \13143 , RIaaa5e88_496, \11761 );
and \U$12301 ( \13144 , \7961 , RIaaa5ff0_499);
and \U$12302 ( \13145 , RIaaa6068_500, \7949 );
nor \U$12303 ( \13146 , \13143 , \13144 , \13145 );
and \U$12304 ( \13147 , \7928 , RIaaa5f78_498);
and \U$12305 ( \13148 , RIaaa5d20_493, \7909 );
nor \U$12306 ( \13149 , \13147 , \13148 );
nand \U$12307 ( \13150 , \13142 , \13146 , \13149 );
nor \U$12308 ( \13151 , \13138 , \13139 , \13150 );
and \U$12309 ( \13152 , \7914 , RIaaa5c30_491);
and \U$12310 ( \13153 , RIaaa6158_502, \7959 );
nor \U$12311 ( \13154 , \13152 , \13153 );
and \U$12312 ( \13155 , \7942 , RIaaa59d8_486);
and \U$12313 ( \13156 , RIaaa5a50_487, \7919 );
nor \U$12314 ( \13157 , \13155 , \13156 );
and \U$12315 ( \13158 , \7952 , RIaaa5ca8_492);
and \U$12316 ( \13159 , RIaaa5bb8_490, \7935 );
nor \U$12317 ( \13160 , \13158 , \13159 );
nand \U$12318 ( \13161 , \13151 , \13154 , \13157 , \13160 );
_DC g2320 ( \13162_nG2320 , \13161 , \11781 );
nand \U$12319 ( \13163 , \13162_nG2320 , \11754 );
not \U$12320 ( \13164 , \13163 );
and \U$12321 ( \13165 , \13137 , \13164 );
nor \U$12322 ( \13166 , \13128 , \13135 );
nor \U$12323 ( \13167 , \13165 , \13166 );
nand \U$12324 ( \13168 , \13096 , \13167 );
not \U$12325 ( \13169 , \13015 );
or \U$12326 ( \13170 , \13169 , \11783 );
or \U$12327 ( \13171 , \11782_nG30bb , \12852 );
or \U$12328 ( \13172 , \11874_nG2fb5 , \12851 );
nand \U$12329 ( \13173 , \13170 , \13171 , \13172 );
or \U$12330 ( \13174 , \12589 , \12085 );
or \U$12331 ( \13175 , \12541 , \11951_nG2e94 );
nand \U$12332 ( \13176 , \13175 , \12753 );
nand \U$12333 ( \13177 , \12076_nG2daa , \12586 );
and \U$12334 ( \13178 , \13176 , \13177 );
and \U$12335 ( \13179 , \11951_nG2e94 , \12756 );
nor \U$12336 ( \13180 , \13178 , \13179 );
nand \U$12337 ( \13181 , \13174 , \13180 );
and \U$12338 ( \13182 , \13173 , \13181 );
and \U$12339 ( \13183 , \13168 , \13182 );
nor \U$12340 ( \13184 , \13167 , \13096 );
nor \U$12341 ( \13185 , \13183 , \13184 );
nand \U$12342 ( \13186 , \13071 , \13185 );
xor \U$12343 ( \13187 , \12985 , \12992 );
xor \U$12344 ( \13188 , \13187 , \13000 );
not \U$12345 ( \13189 , \13188 );
nand \U$12346 ( \13190 , \13122_nG2354 , \11754 );
and \U$12347 ( \13191 , \12881_nG23c5 , \11834 );
and \U$12348 ( \13192 , \11925 , \12922_nG2391 );
nand \U$12349 ( \13193 , \12881_nG23c5 , \11827 );
or \U$12350 ( \13194 , \11795 , \12922_nG2391 );
nand \U$12351 ( \13195 , \13194 , \11831 );
and \U$12352 ( \13196 , \13193 , \13195 );
nor \U$12353 ( \13197 , \13191 , \13192 , \13196 );
xor \U$12354 ( \13198 , \13190 , \13197 );
and \U$12355 ( \13199 , \13189 , \13198 );
and \U$12356 ( \13200 , \13186 , \13199 );
nor \U$12357 ( \13201 , \13185 , \13071 );
nor \U$12358 ( \13202 , \13200 , \13201 );
and \U$12359 ( \13203 , \13066 , \13202 );
not \U$12360 ( \13204 , \13203 );
not \U$12361 ( \13205 , \13040 );
not \U$12362 ( \13206 , \13043 );
and \U$12363 ( \13207 , \13205 , \13206 );
and \U$12364 ( \13208 , \13040 , \13043 );
nor \U$12365 ( \13209 , \13207 , \13208 );
not \U$12366 ( \13210 , \13209 );
not \U$12367 ( \13211 , \13029 );
or \U$12368 ( \13212 , \13003 , \13211 );
not \U$12369 ( \13213 , \13003 );
or \U$12370 ( \13214 , \13029 , \13213 );
or \U$12371 ( \13215 , \13190 , \13197 );
nand \U$12372 ( \13216 , \13212 , \13214 , \13215 );
nand \U$12373 ( \13217 , \13210 , \13216 );
not \U$12374 ( \13218 , \13217 );
and \U$12375 ( \13219 , \13204 , \13218 );
nor \U$12376 ( \13220 , \13066 , \13202 );
nor \U$12377 ( \13221 , \13219 , \13220 );
not \U$12378 ( \13222 , \12977 );
not \U$12379 ( \13223 , \12967 );
and \U$12380 ( \13224 , \13222 , \13223 );
and \U$12381 ( \13225 , \12977 , \12967 );
nor \U$12382 ( \13226 , \13224 , \13225 );
and \U$12383 ( \13227 , \13221 , \13226 );
not \U$12384 ( \13228 , \13227 );
not \U$12385 ( \13229 , \13047 );
not \U$12386 ( \13230 , \13056 );
or \U$12387 ( \13231 , \13229 , \13230 );
or \U$12388 ( \13232 , \13056 , \13047 );
nand \U$12389 ( \13233 , \13231 , \13232 );
not \U$12390 ( \13234 , \13233 );
and \U$12391 ( \13235 , \13228 , \13234 );
nor \U$12392 ( \13236 , \13221 , \13226 );
nor \U$12393 ( \13237 , \13235 , \13236 );
not \U$12394 ( \13238 , \13237 );
xor \U$12395 ( \13239 , \12978 , \13057 );
xor \U$12396 ( \13240 , \13239 , \13060 );
xor \U$12397 ( \13241 , \13238 , \13240 );
or \U$12398 ( \13242 , \13236 , \13227 );
not \U$12399 ( \13243 , \13242 );
not \U$12400 ( \13244 , \13233 );
and \U$12401 ( \13245 , \13243 , \13244 );
and \U$12402 ( \13246 , \13242 , \13233 );
nor \U$12403 ( \13247 , \13245 , \13246 );
not \U$12404 ( \13248 , \13216 );
not \U$12405 ( \13249 , \13209 );
or \U$12406 ( \13250 , \13248 , \13249 );
or \U$12407 ( \13251 , \13209 , \13216 );
nand \U$12408 ( \13252 , \13250 , \13251 );
not \U$12409 ( \13253 , \13010 );
xor \U$12410 ( \13254 , \13017 , \13027 );
not \U$12411 ( \13255 , \13254 );
or \U$12412 ( \13256 , \13253 , \13255 );
or \U$12413 ( \13257 , \13254 , \13010 );
nand \U$12414 ( \13258 , \13256 , \13257 );
nand \U$12415 ( \13259 , \12662_nG27f3 , \12014 );
or \U$12416 ( \13260 , \11964 , \12706_nG2723 );
nand \U$12417 ( \13261 , \13260 , \12020 );
and \U$12418 ( \13262 , \13259 , \13261 );
and \U$12419 ( \13263 , \12016 , \12706_nG2723 );
and \U$12420 ( \13264 , \12662_nG27f3 , \12125 );
nor \U$12421 ( \13265 , \13262 , \13263 , \13264 );
nand \U$12422 ( \13266 , \12515_nG28d0 , \12179 );
or \U$12423 ( \13267 , \12110 , \12307_nG29cd );
nand \U$12424 ( \13268 , \13267 , \12315 );
and \U$12425 ( \13269 , \13266 , \13268 );
and \U$12426 ( \13270 , \12318 , \12307_nG29cd );
and \U$12427 ( \13271 , \12515_nG28d0 , \12182 );
nor \U$12428 ( \13272 , \13269 , \13270 , \13271 );
xor \U$12429 ( \13273 , \13265 , \13272 );
nand \U$12430 ( \13274 , \12922_nG2391 , \11886 );
or \U$12431 ( \13275 , \11848 , \12881_nG23c5 );
nand \U$12432 ( \13276 , \13275 , \11917 );
and \U$12433 ( \13277 , \13274 , \13276 );
and \U$12434 ( \13278 , \11920 , \12881_nG23c5 );
and \U$12435 ( \13279 , \12922_nG2391 , \11889 );
nor \U$12436 ( \13280 , \13277 , \13278 , \13279 );
and \U$12437 ( \13281 , \13273 , \13280 );
and \U$12438 ( \13282 , \13265 , \13272 );
or \U$12439 ( \13283 , \13281 , \13282 );
nand \U$12440 ( \13284 , \12048_nG2ca8 , \12586 );
or \U$12441 ( \13285 , \12541 , \12076_nG2daa );
nand \U$12442 ( \13286 , \13285 , \12753 );
and \U$12443 ( \13287 , \13284 , \13286 );
and \U$12444 ( \13288 , \12756 , \12076_nG2daa );
and \U$12445 ( \13289 , \12048_nG2ca8 , \12588 );
nor \U$12446 ( \13290 , \13287 , \13288 , \13289 );
and \U$12447 ( \13291 , \11896 , \13012 );
not \U$12448 ( \13292 , \11951_nG2e94 );
and \U$12449 ( \13293 , \12850 , \13292 );
and \U$12450 ( \13294 , \11874_nG2fb5 , \13015 );
nor \U$12451 ( \13295 , \13291 , \13293 , \13294 );
xor \U$12452 ( \13296 , \13290 , \13295 );
nand \U$12453 ( \13297 , \12237_nG2aae , \12380 );
or \U$12454 ( \13298 , \12337 , \12160_nG2bb5 );
nand \U$12455 ( \13299 , \13298 , \12527 );
and \U$12456 ( \13300 , \13297 , \13299 );
and \U$12457 ( \13301 , \12530 , \12160_nG2bb5 );
and \U$12458 ( \13302 , \12237_nG2aae , \12383 );
nor \U$12459 ( \13303 , \13300 , \13301 , \13302 );
and \U$12460 ( \13304 , \13296 , \13303 );
and \U$12461 ( \13305 , \13290 , \13295 );
or \U$12462 ( \13306 , \13304 , \13305 );
nor \U$12463 ( \13307 , \13283 , \13306 );
and \U$12464 ( \13308 , \13258 , \13307 );
xor \U$12465 ( \13309 , \13252 , \13308 );
not \U$12466 ( \13310 , \13199 );
not \U$12467 ( \13311 , \13201 );
nand \U$12468 ( \13312 , \13311 , \13186 );
not \U$12469 ( \13313 , \13312 );
or \U$12470 ( \13314 , \13310 , \13313 );
or \U$12471 ( \13315 , \13312 , \13199 );
nand \U$12472 ( \13316 , \13314 , \13315 );
and \U$12473 ( \13317 , \13309 , \13316 );
and \U$12474 ( \13318 , \13252 , \13308 );
or \U$12475 ( \13319 , \13317 , \13318 );
xor \U$12476 ( \13320 , \13030 , \13033 );
xor \U$12477 ( \13321 , \13320 , \13044 );
xor \U$12478 ( \13322 , \13319 , \13321 );
not \U$12479 ( \13323 , \13217 );
nor \U$12480 ( \13324 , \13220 , \13203 );
not \U$12481 ( \13325 , \13324 );
or \U$12482 ( \13326 , \13323 , \13325 );
or \U$12483 ( \13327 , \13324 , \13217 );
nand \U$12484 ( \13328 , \13326 , \13327 );
and \U$12485 ( \13329 , \13322 , \13328 );
and \U$12486 ( \13330 , \13319 , \13321 );
or \U$12487 ( \13331 , \13329 , \13330 );
xor \U$12488 ( \13332 , \13247 , \13331 );
xor \U$12489 ( \13333 , \13319 , \13321 );
xor \U$12490 ( \13334 , \13333 , \13328 );
not \U$12491 ( \13335 , \13283 );
or \U$12492 ( \13336 , \13335 , \13306 );
not \U$12493 ( \13337 , \13306 );
or \U$12494 ( \13338 , \13337 , \13283 );
and \U$12495 ( \13339 , \7930 , RIaaa70d0_535);
and \U$12496 ( \13340 , \7952 , RIaaa6ef0_531);
and \U$12497 ( \13341 , RIaaa6d88_528, \7957 );
nor \U$12498 ( \13342 , \13340 , \13341 );
and \U$12499 ( \13343 , \7942 , RIaaa6b30_523);
and \U$12500 ( \13344 , RIaaa69c8_520, \7944 );
nor \U$12501 ( \13345 , \13343 , \13344 );
and \U$12502 ( \13346 , \7914 , RIaaa6ba8_524);
and \U$12503 ( \13347 , RIaaa6c20_525, \7935 );
nor \U$12504 ( \13348 , \13346 , \13347 );
and \U$12505 ( \13349 , \7919 , RIaaa6ab8_522);
and \U$12506 ( \13350 , RIaaa6e00_529, \7959 );
nor \U$12507 ( \13351 , \13349 , \13350 );
nand \U$12508 ( \13352 , \13342 , \13345 , \13348 , \13351 );
nor \U$12509 ( \13353 , \13339 , \13352 );
and \U$12510 ( \13354 , \7961 , RIaaa6c98_526);
and \U$12511 ( \13355 , RIaaa6a40_521, \7963 );
nor \U$12512 ( \13356 , \13354 , \13355 );
and \U$12513 ( \13357 , \7928 , RIaaa6d10_527);
and \U$12514 ( \13358 , RIaaa6f68_532, \7909 );
nor \U$12515 ( \13359 , \13357 , \13358 );
and \U$12516 ( \13360 , \11761 , RIaaa7058_534);
and \U$12517 ( \13361 , RIaaa6e78_530, \7949 );
nor \U$12518 ( \13362 , \13360 , \13361 );
nand \U$12519 ( \13363 , \13353 , \13356 , \13359 , \13362 );
_DC g22e4 ( \13364_nG22e4 , \13363 , \11781 );
nand \U$12520 ( \13365 , \13364_nG22e4 , \11754 );
and \U$12521 ( \13366 , \13122_nG2354 , \11834 );
and \U$12522 ( \13367 , \11925 , \13162_nG2320 );
nand \U$12523 ( \13368 , \13122_nG2354 , \11827 );
or \U$12524 ( \13369 , \11795 , \13162_nG2320 );
nand \U$12525 ( \13370 , \13369 , \11831 );
and \U$12526 ( \13371 , \13368 , \13370 );
nor \U$12527 ( \13372 , \13366 , \13367 , \13371 );
or \U$12528 ( \13373 , \13365 , \13372 );
nand \U$12529 ( \13374 , \13336 , \13338 , \13373 );
xor \U$12530 ( \13375 , \13173 , \13181 );
xor \U$12531 ( \13376 , \13374 , \13375 );
not \U$12532 ( \13377 , \13163 );
nor \U$12533 ( \13378 , \13136 , \13166 );
not \U$12534 ( \13379 , \13378 );
or \U$12535 ( \13380 , \13377 , \13379 );
or \U$12536 ( \13381 , \13378 , \13163 );
nand \U$12537 ( \13382 , \13380 , \13381 );
and \U$12538 ( \13383 , \13376 , \13382 );
and \U$12539 ( \13384 , \13374 , \13375 );
or \U$12540 ( \13385 , \13383 , \13384 );
xor \U$12541 ( \13386 , \13189 , \13198 );
xor \U$12542 ( \13387 , \13385 , \13386 );
xnor \U$12543 ( \13388 , \13365 , \13372 );
xor \U$12544 ( \13389 , \13265 , \13272 );
xor \U$12545 ( \13390 , \13389 , \13280 );
and \U$12546 ( \13391 , \13388 , \13390 );
not \U$12547 ( \13392 , \13391 );
xor \U$12548 ( \13393 , \13290 , \13295 );
xor \U$12549 ( \13394 , \13393 , \13303 );
not \U$12550 ( \13395 , \13394 );
and \U$12551 ( \13396 , \13392 , \13395 );
nor \U$12552 ( \13397 , \13388 , \13390 );
nor \U$12553 ( \13398 , \13396 , \13397 );
xor \U$12554 ( \13399 , \13078 , \13085 );
xor \U$12555 ( \13400 , \13399 , \13093 );
xor \U$12556 ( \13401 , \13398 , \13400 );
nand \U$12557 ( \13402 , \12662_nG27f3 , \12179 );
or \U$12558 ( \13403 , \12110 , \12515_nG28d0 );
nand \U$12559 ( \13404 , \13403 , \12315 );
and \U$12560 ( \13405 , \13402 , \13404 );
and \U$12561 ( \13406 , \12318 , \12515_nG28d0 );
and \U$12562 ( \13407 , \12662_nG27f3 , \12182 );
nor \U$12563 ( \13408 , \13405 , \13406 , \13407 );
nand \U$12564 ( \13409 , \12307_nG29cd , \12380 );
or \U$12565 ( \13410 , \12337 , \12237_nG2aae );
nand \U$12566 ( \13411 , \13410 , \12527 );
and \U$12567 ( \13412 , \13409 , \13411 );
and \U$12568 ( \13413 , \12530 , \12237_nG2aae );
and \U$12569 ( \13414 , \12307_nG29cd , \12383 );
nor \U$12570 ( \13415 , \13412 , \13413 , \13414 );
xor \U$12571 ( \13416 , \13408 , \13415 );
nand \U$12572 ( \13417 , \12706_nG2723 , \12014 );
or \U$12573 ( \13418 , \11964 , \12881_nG23c5 );
nand \U$12574 ( \13419 , \13418 , \12020 );
and \U$12575 ( \13420 , \13417 , \13419 );
and \U$12576 ( \13421 , \12016 , \12881_nG23c5 );
and \U$12577 ( \13422 , \12706_nG2723 , \12125 );
nor \U$12578 ( \13423 , \13420 , \13421 , \13422 );
and \U$12579 ( \13424 , \13416 , \13423 );
and \U$12580 ( \13425 , \13408 , \13415 );
or \U$12581 ( \13426 , \13424 , \13425 );
nand \U$12582 ( \13427 , \12160_nG2bb5 , \12586 );
or \U$12583 ( \13428 , \12541 , \12048_nG2ca8 );
nand \U$12584 ( \13429 , \13428 , \12753 );
and \U$12585 ( \13430 , \13427 , \13429 );
and \U$12586 ( \13431 , \12756 , \12048_nG2ca8 );
and \U$12587 ( \13432 , \12160_nG2bb5 , \12588 );
nor \U$12588 ( \13433 , \13430 , \13431 , \13432 );
not \U$12589 ( \13434 , \13433 );
or \U$12590 ( \13435 , \13169 , \13292 );
or \U$12591 ( \13436 , \11951_nG2e94 , \12852 );
or \U$12592 ( \13437 , \12076_nG2daa , \12851 );
nand \U$12593 ( \13438 , \13435 , \13436 , \13437 );
nand \U$12594 ( \13439 , \13434 , \13438 );
xor \U$12595 ( \13440 , \13426 , \13439 );
and \U$12596 ( \13441 , \13162_nG2320 , \11834 );
and \U$12597 ( \13442 , \11925 , \13364_nG22e4 );
nand \U$12598 ( \13443 , \13162_nG2320 , \11827 );
or \U$12599 ( \13444 , \11795 , \13364_nG22e4 );
nand \U$12600 ( \13445 , \13444 , \11831 );
and \U$12601 ( \13446 , \13443 , \13445 );
nor \U$12602 ( \13447 , \13441 , \13442 , \13446 );
nand \U$12603 ( \13448 , \13122_nG2354 , \11886 );
or \U$12604 ( \13449 , \11848 , \12922_nG2391 );
nand \U$12605 ( \13450 , \13449 , \11917 );
and \U$12606 ( \13451 , \13448 , \13450 );
and \U$12607 ( \13452 , \11920 , \12922_nG2391 );
and \U$12608 ( \13453 , \13122_nG2354 , \11889 );
nor \U$12609 ( \13454 , \13451 , \13452 , \13453 );
and \U$12610 ( \13455 , \13447 , \13454 );
not \U$12611 ( \13456 , \13455 );
and \U$12612 ( \13457 , RIaaa7850_551, \7959 );
and \U$12613 ( \13458 , RIaaa7490_543, \7944 );
and \U$12614 ( \13459 , \7963 , RIaaa7580_545);
and \U$12615 ( \13460 , RIaaa7328_540, \7930 );
nor \U$12616 ( \13461 , \13459 , \13460 );
and \U$12617 ( \13462 , RIaaa72b0_539, \11761 );
and \U$12618 ( \13463 , \7961 , RIaaa76e8_548);
and \U$12619 ( \13464 , RIaaa7508_544, \7949 );
nor \U$12620 ( \13465 , \13462 , \13463 , \13464 );
and \U$12621 ( \13466 , \7928 , RIaaa7760_549);
and \U$12622 ( \13467 , RIaaa7940_553, \7909 );
nor \U$12623 ( \13468 , \13466 , \13467 );
nand \U$12624 ( \13469 , \13461 , \13465 , \13468 );
nor \U$12625 ( \13470 , \13457 , \13458 , \13469 );
and \U$12626 ( \13471 , \7919 , RIaaa7670_547);
and \U$12627 ( \13472 , RIaaa77d8_550, \7957 );
nor \U$12628 ( \13473 , \13471 , \13472 );
and \U$12629 ( \13474 , \7914 , RIaaa7418_542);
and \U$12630 ( \13475 , RIaaa75f8_546, \7942 );
nor \U$12631 ( \13476 , \13474 , \13475 );
and \U$12632 ( \13477 , \7952 , RIaaa78c8_552);
and \U$12633 ( \13478 , RIaaa73a0_541, \7935 );
nor \U$12634 ( \13479 , \13477 , \13478 );
nand \U$12635 ( \13480 , \13470 , \13473 , \13476 , \13479 );
_DC g22ab ( \13481_nG22ab , \13480 , \11781 );
nand \U$12636 ( \13482 , \13481_nG22ab , \11754 );
not \U$12637 ( \13483 , \13482 );
and \U$12638 ( \13484 , \13456 , \13483 );
nor \U$12639 ( \13485 , \13447 , \13454 );
nor \U$12640 ( \13486 , \13484 , \13485 );
and \U$12641 ( \13487 , \13440 , \13486 );
and \U$12642 ( \13488 , \13426 , \13439 );
or \U$12643 ( \13489 , \13487 , \13488 );
and \U$12644 ( \13490 , \13401 , \13489 );
and \U$12645 ( \13491 , \13398 , \13400 );
or \U$12646 ( \13492 , \13490 , \13491 );
not \U$12647 ( \13493 , \13492 );
and \U$12648 ( \13494 , \13387 , \13493 );
and \U$12649 ( \13495 , \13385 , \13386 );
or \U$12650 ( \13496 , \13494 , \13495 );
xor \U$12651 ( \13497 , \13258 , \13307 );
not \U$12652 ( \13498 , \13182 );
not \U$12653 ( \13499 , \13184 );
nand \U$12654 ( \13500 , \13499 , \13168 );
not \U$12655 ( \13501 , \13500 );
or \U$12656 ( \13502 , \13498 , \13501 );
or \U$12657 ( \13503 , \13500 , \13182 );
nand \U$12658 ( \13504 , \13502 , \13503 );
and \U$12659 ( \13505 , \13497 , \13504 );
xor \U$12660 ( \13506 , \13496 , \13505 );
xor \U$12661 ( \13507 , \13252 , \13308 );
xor \U$12662 ( \13508 , \13507 , \13316 );
and \U$12663 ( \13509 , \13506 , \13508 );
and \U$12664 ( \13510 , \13496 , \13505 );
or \U$12665 ( \13511 , \13509 , \13510 );
xor \U$12666 ( \13512 , \13334 , \13511 );
xor \U$12667 ( \13513 , \13496 , \13505 );
xor \U$12668 ( \13514 , \13513 , \13508 );
xor \U$12669 ( \13515 , \13398 , \13400 );
xor \U$12670 ( \13516 , \13515 , \13489 );
not \U$12671 ( \13517 , \13482 );
nor \U$12672 ( \13518 , \13455 , \13485 );
not \U$12673 ( \13519 , \13518 );
or \U$12674 ( \13520 , \13517 , \13519 );
or \U$12675 ( \13521 , \13518 , \13482 );
nand \U$12676 ( \13522 , \13520 , \13521 );
not \U$12677 ( \13523 , \13522 );
xor \U$12678 ( \13524 , \13408 , \13415 );
xor \U$12679 ( \13525 , \13524 , \13423 );
nor \U$12680 ( \13526 , \13523 , \13525 );
nand \U$12681 ( \13527 , \12881_nG23c5 , \12014 );
or \U$12682 ( \13528 , \11964 , \12922_nG2391 );
nand \U$12683 ( \13529 , \13528 , \12020 );
and \U$12684 ( \13530 , \13527 , \13529 );
and \U$12685 ( \13531 , \12016 , \12922_nG2391 );
and \U$12686 ( \13532 , \12881_nG23c5 , \12125 );
nor \U$12687 ( \13533 , \13530 , \13531 , \13532 );
nand \U$12688 ( \13534 , \12706_nG2723 , \12179 );
or \U$12689 ( \13535 , \12110 , \12662_nG27f3 );
nand \U$12690 ( \13536 , \13535 , \12315 );
and \U$12691 ( \13537 , \13534 , \13536 );
and \U$12692 ( \13538 , \12318 , \12662_nG27f3 );
and \U$12693 ( \13539 , \12706_nG2723 , \12182 );
nor \U$12694 ( \13540 , \13537 , \13538 , \13539 );
xor \U$12695 ( \13541 , \13533 , \13540 );
nand \U$12696 ( \13542 , \13162_nG2320 , \11886 );
or \U$12697 ( \13543 , \11848 , \13122_nG2354 );
nand \U$12698 ( \13544 , \13543 , \11917 );
and \U$12699 ( \13545 , \13542 , \13544 );
and \U$12700 ( \13546 , \11920 , \13122_nG2354 );
and \U$12701 ( \13547 , \13162_nG2320 , \11889 );
nor \U$12702 ( \13548 , \13545 , \13546 , \13547 );
and \U$12703 ( \13549 , \13541 , \13548 );
and \U$12704 ( \13550 , \13533 , \13540 );
or \U$12705 ( \13551 , \13549 , \13550 );
nand \U$12706 ( \13552 , \12237_nG2aae , \12586 );
or \U$12707 ( \13553 , \12541 , \12160_nG2bb5 );
nand \U$12708 ( \13554 , \13553 , \12753 );
and \U$12709 ( \13555 , \13552 , \13554 );
and \U$12710 ( \13556 , \12756 , \12160_nG2bb5 );
and \U$12711 ( \13557 , \12237_nG2aae , \12588 );
nor \U$12712 ( \13558 , \13555 , \13556 , \13557 );
and \U$12713 ( \13559 , \12085 , \13012 );
and \U$12714 ( \13560 , \12850 , \12164 );
and \U$12715 ( \13561 , \12076_nG2daa , \13015 );
nor \U$12716 ( \13562 , \13559 , \13560 , \13561 );
xor \U$12717 ( \13563 , \13558 , \13562 );
nand \U$12718 ( \13564 , \12515_nG28d0 , \12380 );
or \U$12719 ( \13565 , \12337 , \12307_nG29cd );
nand \U$12720 ( \13566 , \13565 , \12527 );
and \U$12721 ( \13567 , \13564 , \13566 );
and \U$12722 ( \13568 , \12530 , \12307_nG29cd );
and \U$12723 ( \13569 , \12515_nG28d0 , \12383 );
nor \U$12724 ( \13570 , \13567 , \13568 , \13569 );
and \U$12725 ( \13571 , \13563 , \13570 );
and \U$12726 ( \13572 , \13558 , \13562 );
or \U$12727 ( \13573 , \13571 , \13572 );
nor \U$12728 ( \13574 , \13551 , \13573 );
xor \U$12729 ( \13575 , \13526 , \13574 );
not \U$12730 ( \13576 , \13394 );
nor \U$12731 ( \13577 , \13391 , \13397 );
not \U$12732 ( \13578 , \13577 );
or \U$12733 ( \13579 , \13576 , \13578 );
or \U$12734 ( \13580 , \13577 , \13394 );
nand \U$12735 ( \13581 , \13579 , \13580 );
and \U$12736 ( \13582 , \13575 , \13581 );
and \U$12737 ( \13583 , \13526 , \13574 );
or \U$12738 ( \13584 , \13582 , \13583 );
xor \U$12739 ( \13585 , \13374 , \13375 );
xor \U$12740 ( \13586 , \13585 , \13382 );
nor \U$12741 ( \13587 , \13584 , \13586 );
or \U$12742 ( \13588 , \13516 , \13587 );
nand \U$12743 ( \13589 , \13586 , \13584 );
nand \U$12744 ( \13590 , \13588 , \13589 );
xor \U$12745 ( \13591 , \13497 , \13504 );
xor \U$12746 ( \13592 , \13590 , \13591 );
xor \U$12747 ( \13593 , \13385 , \13386 );
xor \U$12748 ( \13594 , \13593 , \13493 );
and \U$12749 ( \13595 , \13592 , \13594 );
and \U$12750 ( \13596 , \13590 , \13591 );
or \U$12751 ( \13597 , \13595 , \13596 );
xor \U$12752 ( \13598 , \13514 , \13597 );
xor \U$12753 ( \13599 , \13590 , \13591 );
xor \U$12754 ( \13600 , \13599 , \13594 );
not \U$12755 ( \13601 , \13589 );
nor \U$12756 ( \13602 , \13601 , \13587 );
not \U$12757 ( \13603 , \13602 );
not \U$12758 ( \13604 , \13516 );
and \U$12759 ( \13605 , \13603 , \13604 );
and \U$12760 ( \13606 , \13602 , \13516 );
nor \U$12761 ( \13607 , \13605 , \13606 );
xor \U$12762 ( \13608 , \13533 , \13540 );
xor \U$12763 ( \13609 , \13608 , \13548 );
xor \U$12764 ( \13610 , \13558 , \13562 );
xor \U$12765 ( \13611 , \13610 , \13570 );
xor \U$12766 ( \13612 , \13609 , \13611 );
and \U$12767 ( \13613 , RIaaa87c8_584, \7957 );
and \U$12768 ( \13614 , RIaaa8408_576, \7944 );
and \U$12769 ( \13615 , \7963 , RIaaa8570_579);
and \U$12770 ( \13616 , RIaaa8318_574, \7930 );
nor \U$12771 ( \13617 , \13615 , \13616 );
and \U$12772 ( \13618 , RIaaa82a0_573, \11761 );
and \U$12773 ( \13619 , \7961 , RIaaa86d8_582);
and \U$12774 ( \13620 , RIaaa84f8_578, \7949 );
nor \U$12775 ( \13621 , \13618 , \13619 , \13620 );
and \U$12776 ( \13622 , \7928 , RIaaa8750_583);
and \U$12777 ( \13623 , RIaaa8930_587, \7909 );
nor \U$12778 ( \13624 , \13622 , \13623 );
nand \U$12779 ( \13625 , \13617 , \13621 , \13624 );
nor \U$12780 ( \13626 , \13613 , \13614 , \13625 );
and \U$12781 ( \13627 , \7914 , RIaaa8480_577);
and \U$12782 ( \13628 , RIaaa8840_585, \7959 );
nor \U$12783 ( \13629 , \13627 , \13628 );
and \U$12784 ( \13630 , \7942 , RIaaa85e8_580);
and \U$12785 ( \13631 , RIaaa8660_581, \7919 );
nor \U$12786 ( \13632 , \13630 , \13631 );
and \U$12787 ( \13633 , \7952 , RIaaa88b8_586);
and \U$12788 ( \13634 , RIaaa8390_575, \7935 );
nor \U$12789 ( \13635 , \13633 , \13634 );
nand \U$12790 ( \13636 , \13626 , \13629 , \13632 , \13635 );
_DC g2273 ( \13637_nG2273 , \13636 , \11781 );
nand \U$12791 ( \13638 , \13637_nG2273 , \11754 );
and \U$12792 ( \13639 , \13364_nG22e4 , \11834 );
and \U$12793 ( \13640 , \11925 , \13481_nG22ab );
nand \U$12794 ( \13641 , \13364_nG22e4 , \11827 );
or \U$12795 ( \13642 , \11795 , \13481_nG22ab );
nand \U$12796 ( \13643 , \13642 , \11831 );
and \U$12797 ( \13644 , \13641 , \13643 );
nor \U$12798 ( \13645 , \13639 , \13640 , \13644 );
xnor \U$12799 ( \13646 , \13638 , \13645 );
and \U$12800 ( \13647 , \13612 , \13646 );
and \U$12801 ( \13648 , \13609 , \13611 );
or \U$12802 ( \13649 , \13647 , \13648 );
not \U$12803 ( \13650 , \13433 );
not \U$12804 ( \13651 , \13438 );
and \U$12805 ( \13652 , \13650 , \13651 );
and \U$12806 ( \13653 , \13433 , \13438 );
nor \U$12807 ( \13654 , \13652 , \13653 );
xor \U$12808 ( \13655 , \13649 , \13654 );
nand \U$12809 ( \13656 , \12881_nG23c5 , \12179 );
or \U$12810 ( \13657 , \12110 , \12706_nG2723 );
nand \U$12811 ( \13658 , \13657 , \12315 );
and \U$12812 ( \13659 , \13656 , \13658 );
and \U$12813 ( \13660 , \12318 , \12706_nG2723 );
and \U$12814 ( \13661 , \12881_nG23c5 , \12182 );
nor \U$12815 ( \13662 , \13659 , \13660 , \13661 );
nand \U$12816 ( \13663 , \12662_nG27f3 , \12380 );
or \U$12817 ( \13664 , \12337 , \12515_nG28d0 );
nand \U$12818 ( \13665 , \13664 , \12527 );
and \U$12819 ( \13666 , \13663 , \13665 );
and \U$12820 ( \13667 , \12530 , \12515_nG28d0 );
and \U$12821 ( \13668 , \12662_nG27f3 , \12383 );
nor \U$12822 ( \13669 , \13666 , \13667 , \13668 );
xor \U$12823 ( \13670 , \13662 , \13669 );
nand \U$12824 ( \13671 , \12922_nG2391 , \12014 );
or \U$12825 ( \13672 , \11964 , \13122_nG2354 );
nand \U$12826 ( \13673 , \13672 , \12020 );
and \U$12827 ( \13674 , \13671 , \13673 );
and \U$12828 ( \13675 , \12016 , \13122_nG2354 );
and \U$12829 ( \13676 , \12922_nG2391 , \12125 );
nor \U$12830 ( \13677 , \13674 , \13675 , \13676 );
and \U$12831 ( \13678 , \13670 , \13677 );
and \U$12832 ( \13679 , \13662 , \13669 );
or \U$12833 ( \13680 , \13678 , \13679 );
nand \U$12834 ( \13681 , \12307_nG29cd , \12586 );
or \U$12835 ( \13682 , \12541 , \12237_nG2aae );
nand \U$12836 ( \13683 , \13682 , \12753 );
and \U$12837 ( \13684 , \13681 , \13683 );
and \U$12838 ( \13685 , \12756 , \12237_nG2aae );
and \U$12839 ( \13686 , \12307_nG29cd , \12588 );
nor \U$12840 ( \13687 , \13684 , \13685 , \13686 );
not \U$12841 ( \13688 , \13687 );
or \U$12842 ( \13689 , \13169 , \12164 );
or \U$12843 ( \13690 , \12048_nG2ca8 , \12852 );
or \U$12844 ( \13691 , \12160_nG2bb5 , \12851 );
nand \U$12845 ( \13692 , \13689 , \13690 , \13691 );
nand \U$12846 ( \13693 , \13688 , \13692 );
xor \U$12847 ( \13694 , \13680 , \13693 );
nand \U$12848 ( \13695 , \13364_nG22e4 , \11886 );
or \U$12849 ( \13696 , \11848 , \13162_nG2320 );
nand \U$12850 ( \13697 , \13696 , \11917 );
and \U$12851 ( \13698 , \13695 , \13697 );
and \U$12852 ( \13699 , \11920 , \13162_nG2320 );
and \U$12853 ( \13700 , \13364_nG22e4 , \11889 );
nor \U$12854 ( \13701 , \13698 , \13699 , \13700 );
and \U$12855 ( \13702 , RIaaa8138_570, \7959 );
and \U$12856 ( \13703 , RIaaa7c10_559, \7914 );
and \U$12857 ( \13704 , \7963 , RIaaa7b20_557);
and \U$12858 ( \13705 , RIaaa7df0_563, \7930 );
nor \U$12859 ( \13706 , \13704 , \13705 );
and \U$12860 ( \13707 , RIaaa7e68_564, \11761 );
and \U$12861 ( \13708 , \7961 , RIaaa7f58_566);
and \U$12862 ( \13709 , RIaaa8048_568, \7949 );
nor \U$12863 ( \13710 , \13707 , \13708 , \13709 );
and \U$12864 ( \13711 , \7928 , RIaaa7fd0_567);
and \U$12865 ( \13712 , RIaaa7c88_560, \7909 );
nor \U$12866 ( \13713 , \13711 , \13712 );
nand \U$12867 ( \13714 , \13706 , \13710 , \13713 );
nor \U$12868 ( \13715 , \13702 , \13703 , \13714 );
and \U$12869 ( \13716 , \7919 , RIaaa7a30_555);
and \U$12870 ( \13717 , RIaaa80c0_569, \7957 );
nor \U$12871 ( \13718 , \13716 , \13717 );
and \U$12872 ( \13719 , \7942 , RIaaa79b8_554);
and \U$12873 ( \13720 , RIaaa7d00_561, \7952 );
nor \U$12874 ( \13721 , \13719 , \13720 );
and \U$12875 ( \13722 , \7935 , RIaaa7b98_558);
and \U$12876 ( \13723 , RIaaa7aa8_556, \7944 );
nor \U$12877 ( \13724 , \13722 , \13723 );
nand \U$12878 ( \13725 , \13715 , \13718 , \13721 , \13724 );
_DC g223a ( \13726_nG223a , \13725 , \11781 );
nand \U$12879 ( \13727 , \13726_nG223a , \11754 );
xor \U$12880 ( \13728 , \13701 , \13727 );
and \U$12881 ( \13729 , \13481_nG22ab , \11834 );
and \U$12882 ( \13730 , \11925 , \13637_nG2273 );
nand \U$12883 ( \13731 , \13481_nG22ab , \11827 );
or \U$12884 ( \13732 , \11795 , \13637_nG2273 );
nand \U$12885 ( \13733 , \13732 , \11831 );
and \U$12886 ( \13734 , \13731 , \13733 );
nor \U$12887 ( \13735 , \13729 , \13730 , \13734 );
and \U$12888 ( \13736 , \13728 , \13735 );
and \U$12889 ( \13737 , \13701 , \13727 );
or \U$12890 ( \13738 , \13736 , \13737 );
and \U$12891 ( \13739 , \13694 , \13738 );
and \U$12892 ( \13740 , \13680 , \13693 );
or \U$12893 ( \13741 , \13739 , \13740 );
and \U$12894 ( \13742 , \13655 , \13741 );
and \U$12895 ( \13743 , \13649 , \13654 );
or \U$12896 ( \13744 , \13742 , \13743 );
xor \U$12897 ( \13745 , \13426 , \13439 );
xor \U$12898 ( \13746 , \13745 , \13486 );
and \U$12899 ( \13747 , \13744 , \13746 );
not \U$12900 ( \13748 , \13747 );
not \U$12901 ( \13749 , \13522 );
not \U$12902 ( \13750 , \13525 );
and \U$12903 ( \13751 , \13749 , \13750 );
and \U$12904 ( \13752 , \13522 , \13525 );
nor \U$12905 ( \13753 , \13751 , \13752 );
not \U$12906 ( \13754 , \13753 );
not \U$12907 ( \13755 , \13573 );
or \U$12908 ( \13756 , \13551 , \13755 );
not \U$12909 ( \13757 , \13551 );
or \U$12910 ( \13758 , \13573 , \13757 );
or \U$12911 ( \13759 , \13638 , \13645 );
nand \U$12912 ( \13760 , \13756 , \13758 , \13759 );
nand \U$12913 ( \13761 , \13754 , \13760 );
not \U$12914 ( \13762 , \13761 );
and \U$12915 ( \13763 , \13748 , \13762 );
nor \U$12916 ( \13764 , \13744 , \13746 );
nor \U$12917 ( \13765 , \13763 , \13764 );
nor \U$12918 ( \13766 , \13607 , \13765 );
xor \U$12919 ( \13767 , \13600 , \13766 );
and \U$12920 ( \13768 , \13607 , \13765 );
nor \U$12921 ( \13769 , \13768 , \13766 );
xor \U$12922 ( \13770 , \13526 , \13574 );
xor \U$12923 ( \13771 , \13770 , \13581 );
not \U$12924 ( \13772 , \13761 );
nor \U$12925 ( \13773 , \13764 , \13747 );
not \U$12926 ( \13774 , \13773 );
or \U$12927 ( \13775 , \13772 , \13774 );
or \U$12928 ( \13776 , \13773 , \13761 );
nand \U$12929 ( \13777 , \13775 , \13776 );
nand \U$12930 ( \13778 , \13771 , \13777 );
not \U$12931 ( \13779 , \13778 );
xor \U$12932 ( \13780 , \13769 , \13779 );
or \U$12933 ( \13781 , \13777 , \13771 );
nand \U$12934 ( \13782 , \13781 , \13778 );
not \U$12935 ( \13783 , \13753 );
not \U$12936 ( \13784 , \13760 );
and \U$12937 ( \13785 , \13783 , \13784 );
and \U$12938 ( \13786 , \13753 , \13760 );
nor \U$12939 ( \13787 , \13785 , \13786 );
xor \U$12940 ( \13788 , \13649 , \13654 );
xor \U$12941 ( \13789 , \13788 , \13741 );
and \U$12942 ( \13790 , \13787 , \13789 );
nand \U$12943 ( \13791 , \13122_nG2354 , \12014 );
or \U$12944 ( \13792 , \11964 , \13162_nG2320 );
nand \U$12945 ( \13793 , \13792 , \12020 );
and \U$12946 ( \13794 , \13791 , \13793 );
and \U$12947 ( \13795 , \12016 , \13162_nG2320 );
and \U$12948 ( \13796 , \13122_nG2354 , \12125 );
nor \U$12949 ( \13797 , \13794 , \13795 , \13796 );
nand \U$12950 ( \13798 , \12922_nG2391 , \12179 );
or \U$12951 ( \13799 , \12110 , \12881_nG23c5 );
nand \U$12952 ( \13800 , \13799 , \12315 );
and \U$12953 ( \13801 , \13798 , \13800 );
and \U$12954 ( \13802 , \12318 , \12881_nG23c5 );
and \U$12955 ( \13803 , \12922_nG2391 , \12182 );
nor \U$12956 ( \13804 , \13801 , \13802 , \13803 );
xor \U$12957 ( \13805 , \13797 , \13804 );
nand \U$12958 ( \13806 , \13481_nG22ab , \11886 );
or \U$12959 ( \13807 , \11848 , \13364_nG22e4 );
nand \U$12960 ( \13808 , \13807 , \11917 );
and \U$12961 ( \13809 , \13806 , \13808 );
and \U$12962 ( \13810 , \11920 , \13364_nG22e4 );
and \U$12963 ( \13811 , \13481_nG22ab , \11889 );
nor \U$12964 ( \13812 , \13809 , \13810 , \13811 );
and \U$12965 ( \13813 , \13805 , \13812 );
and \U$12966 ( \13814 , \13797 , \13804 );
or \U$12967 ( \13815 , \13813 , \13814 );
nand \U$12968 ( \13816 , \12515_nG28d0 , \12586 );
or \U$12969 ( \13817 , \12541 , \12307_nG29cd );
nand \U$12970 ( \13818 , \13817 , \12753 );
and \U$12971 ( \13819 , \13816 , \13818 );
and \U$12972 ( \13820 , \12756 , \12307_nG29cd );
and \U$12973 ( \13821 , \12515_nG28d0 , \12588 );
nor \U$12974 ( \13822 , \13819 , \13820 , \13821 );
and \U$12975 ( \13823 , \12161 , \13012 );
not \U$12976 ( \13824 , \12237_nG2aae );
and \U$12977 ( \13825 , \12850 , \13824 );
and \U$12978 ( \13826 , \12160_nG2bb5 , \13015 );
nor \U$12979 ( \13827 , \13823 , \13825 , \13826 );
xor \U$12980 ( \13828 , \13822 , \13827 );
nand \U$12981 ( \13829 , \12706_nG2723 , \12380 );
or \U$12982 ( \13830 , \12337 , \12662_nG27f3 );
nand \U$12983 ( \13831 , \13830 , \12527 );
and \U$12984 ( \13832 , \13829 , \13831 );
and \U$12985 ( \13833 , \12530 , \12662_nG27f3 );
and \U$12986 ( \13834 , \12706_nG2723 , \12383 );
nor \U$12987 ( \13835 , \13832 , \13833 , \13834 );
and \U$12988 ( \13836 , \13828 , \13835 );
and \U$12989 ( \13837 , \13822 , \13827 );
or \U$12990 ( \13838 , \13836 , \13837 );
xor \U$12991 ( \13839 , \13815 , \13838 );
xor \U$12992 ( \13840 , \13701 , \13727 );
xor \U$12993 ( \13841 , \13840 , \13735 );
and \U$12994 ( \13842 , \13839 , \13841 );
and \U$12995 ( \13843 , \13815 , \13838 );
or \U$12996 ( \13844 , \13842 , \13843 );
xor \U$12997 ( \13845 , \13662 , \13669 );
xor \U$12998 ( \13846 , \13845 , \13677 );
not \U$12999 ( \13847 , \13846 );
not \U$13000 ( \13848 , \13692 );
not \U$13001 ( \13849 , \13687 );
or \U$13002 ( \13850 , \13848 , \13849 );
or \U$13003 ( \13851 , \13687 , \13692 );
nand \U$13004 ( \13852 , \13850 , \13851 );
nand \U$13005 ( \13853 , \13847 , \13852 );
xor \U$13006 ( \13854 , \13844 , \13853 );
xor \U$13007 ( \13855 , \13609 , \13611 );
xor \U$13008 ( \13856 , \13855 , \13646 );
and \U$13009 ( \13857 , \13854 , \13856 );
and \U$13010 ( \13858 , \13844 , \13853 );
or \U$13011 ( \13859 , \13857 , \13858 );
xor \U$13012 ( \13860 , \13649 , \13654 );
xor \U$13013 ( \13861 , \13860 , \13741 );
and \U$13014 ( \13862 , \13859 , \13861 );
and \U$13015 ( \13863 , \13787 , \13859 );
or \U$13016 ( \13864 , \13790 , \13862 , \13863 );
xor \U$13017 ( \13865 , \13782 , \13864 );
nand \U$13018 ( \13866 , \12662_nG27f3 , \12586 );
or \U$13019 ( \13867 , \12541 , \12515_nG28d0 );
nand \U$13020 ( \13868 , \13867 , \12753 );
and \U$13021 ( \13869 , \13866 , \13868 );
and \U$13022 ( \13870 , \12756 , \12515_nG28d0 );
and \U$13023 ( \13871 , \12662_nG27f3 , \12588 );
nor \U$13024 ( \13872 , \13869 , \13870 , \13871 );
and \U$13025 ( \13873 , \13824 , \13012 );
and \U$13026 ( \13874 , \12850 , \12604 );
and \U$13027 ( \13875 , \12237_nG2aae , \13015 );
nor \U$13028 ( \13876 , \13873 , \13874 , \13875 );
xor \U$13029 ( \13877 , \13872 , \13876 );
and \U$13030 ( \13878 , \13877 , \11795 );
and \U$13031 ( \13879 , \13872 , \13876 );
or \U$13032 ( \13880 , \13878 , \13879 );
nand \U$13033 ( \13881 , \13122_nG2354 , \12179 );
or \U$13034 ( \13882 , \12110 , \12922_nG2391 );
nand \U$13035 ( \13883 , \13882 , \12315 );
and \U$13036 ( \13884 , \13881 , \13883 );
and \U$13037 ( \13885 , \12318 , \12922_nG2391 );
and \U$13038 ( \13886 , \13122_nG2354 , \12182 );
nor \U$13039 ( \13887 , \13884 , \13885 , \13886 );
nand \U$13040 ( \13888 , \12881_nG23c5 , \12380 );
or \U$13041 ( \13889 , \12337 , \12706_nG2723 );
nand \U$13042 ( \13890 , \13889 , \12527 );
and \U$13043 ( \13891 , \13888 , \13890 );
and \U$13044 ( \13892 , \12530 , \12706_nG2723 );
and \U$13045 ( \13893 , \12881_nG23c5 , \12383 );
nor \U$13046 ( \13894 , \13891 , \13892 , \13893 );
xor \U$13047 ( \13895 , \13887 , \13894 );
nand \U$13048 ( \13896 , \13162_nG2320 , \12014 );
or \U$13049 ( \13897 , \11964 , \13364_nG22e4 );
nand \U$13050 ( \13898 , \13897 , \12020 );
and \U$13051 ( \13899 , \13896 , \13898 );
and \U$13052 ( \13900 , \12016 , \13364_nG22e4 );
and \U$13053 ( \13901 , \13162_nG2320 , \12125 );
nor \U$13054 ( \13902 , \13899 , \13900 , \13901 );
and \U$13055 ( \13903 , \13895 , \13902 );
and \U$13056 ( \13904 , \13887 , \13894 );
or \U$13057 ( \13905 , \13903 , \13904 );
xor \U$13058 ( \13906 , \13880 , \13905 );
and \U$13059 ( \13907 , \13637_nG2273 , \11834 );
and \U$13060 ( \13908 , \11925 , \13726_nG223a );
nand \U$13061 ( \13909 , \13637_nG2273 , \11827 );
or \U$13062 ( \13910 , \11795 , \13726_nG223a );
nand \U$13063 ( \13911 , \13910 , \11831 );
and \U$13064 ( \13912 , \13909 , \13911 );
nor \U$13065 ( \13913 , \13907 , \13908 , \13912 );
and \U$13066 ( \13914 , \13906 , \13913 );
and \U$13067 ( \13915 , \13880 , \13905 );
or \U$13068 ( \13916 , \13914 , \13915 );
not \U$13069 ( \13917 , \13846 );
not \U$13070 ( \13918 , \13852 );
and \U$13071 ( \13919 , \13917 , \13918 );
and \U$13072 ( \13920 , \13846 , \13852 );
nor \U$13073 ( \13921 , \13919 , \13920 );
xor \U$13074 ( \13922 , \13916 , \13921 );
xor \U$13075 ( \13923 , \13815 , \13838 );
xor \U$13076 ( \13924 , \13923 , \13841 );
and \U$13077 ( \13925 , \13922 , \13924 );
and \U$13078 ( \13926 , \13916 , \13921 );
or \U$13079 ( \13927 , \13925 , \13926 );
xor \U$13080 ( \13928 , \13680 , \13693 );
xor \U$13081 ( \13929 , \13928 , \13738 );
xor \U$13082 ( \13930 , \13927 , \13929 );
xor \U$13083 ( \13931 , \13844 , \13853 );
xor \U$13084 ( \13932 , \13931 , \13856 );
and \U$13085 ( \13933 , \13930 , \13932 );
and \U$13086 ( \13934 , \13927 , \13929 );
or \U$13087 ( \13935 , \13933 , \13934 );
xor \U$13088 ( \13936 , \13649 , \13654 );
xor \U$13089 ( \13937 , \13936 , \13741 );
xor \U$13090 ( \13938 , \13787 , \13859 );
xor \U$13091 ( \13939 , \13937 , \13938 );
xor \U$13092 ( \13940 , \13935 , \13939 );
xor \U$13093 ( \13941 , \13880 , \13905 );
xor \U$13094 ( \13942 , \13941 , \13913 );
xor \U$13095 ( \13943 , \13822 , \13827 );
xor \U$13096 ( \13944 , \13943 , \13835 );
or \U$13097 ( \13945 , \13942 , \13944 );
nand \U$13098 ( \13946 , \13637_nG2273 , \11886 );
or \U$13099 ( \13947 , \11848 , \13481_nG22ab );
nand \U$13100 ( \13948 , \13947 , \11917 );
and \U$13101 ( \13949 , \13946 , \13948 );
and \U$13102 ( \13950 , \11920 , \13481_nG22ab );
and \U$13103 ( \13951 , \13637_nG2273 , \11889 );
nor \U$13104 ( \13952 , \13949 , \13950 , \13951 );
nand \U$13105 ( \13953 , \12706_nG2723 , \12586 );
or \U$13106 ( \13954 , \12541 , \12662_nG27f3 );
nand \U$13107 ( \13955 , \13954 , \12753 );
and \U$13108 ( \13956 , \13953 , \13955 );
and \U$13109 ( \13957 , \12756 , \12662_nG27f3 );
and \U$13110 ( \13958 , \12706_nG2723 , \12588 );
nor \U$13111 ( \13959 , \13956 , \13957 , \13958 );
and \U$13112 ( \13960 , \12604 , \13012 );
and \U$13113 ( \13961 , \12850 , \12577 );
and \U$13114 ( \13962 , \12307_nG29cd , \13015 );
nor \U$13115 ( \13963 , \13960 , \13961 , \13962 );
xor \U$13116 ( \13964 , \13959 , \13963 );
nand \U$13117 ( \13965 , \12922_nG2391 , \12380 );
or \U$13118 ( \13966 , \12337 , \12881_nG23c5 );
nand \U$13119 ( \13967 , \13966 , \12527 );
and \U$13120 ( \13968 , \13965 , \13967 );
and \U$13121 ( \13969 , \12530 , \12881_nG23c5 );
and \U$13122 ( \13970 , \12922_nG2391 , \12383 );
nor \U$13123 ( \13971 , \13968 , \13969 , \13970 );
and \U$13124 ( \13972 , \13964 , \13971 );
and \U$13125 ( \13973 , \13959 , \13963 );
or \U$13126 ( \13974 , \13972 , \13973 );
xor \U$13127 ( \13975 , \13952 , \13974 );
nand \U$13128 ( \13976 , \13364_nG22e4 , \12014 );
or \U$13129 ( \13977 , \11964 , \13481_nG22ab );
nand \U$13130 ( \13978 , \13977 , \12020 );
and \U$13131 ( \13979 , \13976 , \13978 );
and \U$13132 ( \13980 , \12016 , \13481_nG22ab );
and \U$13133 ( \13981 , \13364_nG22e4 , \12125 );
nor \U$13134 ( \13982 , \13979 , \13980 , \13981 );
nand \U$13135 ( \13983 , \13162_nG2320 , \12179 );
or \U$13136 ( \13984 , \12110 , \13122_nG2354 );
nand \U$13137 ( \13985 , \13984 , \12315 );
and \U$13138 ( \13986 , \13983 , \13985 );
and \U$13139 ( \13987 , \12318 , \13122_nG2354 );
and \U$13140 ( \13988 , \13162_nG2320 , \12182 );
nor \U$13141 ( \13989 , \13986 , \13987 , \13988 );
xor \U$13142 ( \13990 , \13982 , \13989 );
nand \U$13143 ( \13991 , \13726_nG223a , \11886 );
or \U$13144 ( \13992 , \11848 , \13637_nG2273 );
nand \U$13145 ( \13993 , \13992 , \11917 );
and \U$13146 ( \13994 , \13991 , \13993 );
and \U$13147 ( \13995 , \11920 , \13637_nG2273 );
and \U$13148 ( \13996 , \13726_nG223a , \11889 );
nor \U$13149 ( \13997 , \13994 , \13995 , \13996 );
and \U$13150 ( \13998 , \13990 , \13997 );
and \U$13151 ( \13999 , \13982 , \13989 );
or \U$13152 ( \14000 , \13998 , \13999 );
and \U$13153 ( \14001 , \13975 , \14000 );
and \U$13154 ( \14002 , \13952 , \13974 );
or \U$13155 ( \14003 , \14001 , \14002 );
xor \U$13156 ( \14004 , \13797 , \13804 );
xor \U$13157 ( \14005 , \14004 , \13812 );
xor \U$13158 ( \14006 , \14003 , \14005 );
xor \U$13159 ( \14007 , \13887 , \13894 );
xor \U$13160 ( \14008 , \14007 , \13902 );
xor \U$13161 ( \14009 , \13872 , \13876 );
xor \U$13162 ( \14010 , \14009 , \11795 );
and \U$13163 ( \14011 , \14008 , \14010 );
and \U$13164 ( \14012 , \11834 , \13726_nG223a );
nand \U$13165 ( \14013 , \13726_nG223a , \11827 );
and \U$13166 ( \14014 , \14013 , \11794 );
nor \U$13167 ( \14015 , \14012 , \14014 );
xor \U$13168 ( \14016 , \13872 , \13876 );
xor \U$13169 ( \14017 , \14016 , \11795 );
and \U$13170 ( \14018 , \14015 , \14017 );
and \U$13171 ( \14019 , \14008 , \14015 );
or \U$13172 ( \14020 , \14011 , \14018 , \14019 );
and \U$13173 ( \14021 , \14006 , \14020 );
and \U$13174 ( \14022 , \14003 , \14005 );
or \U$13175 ( \14023 , \14021 , \14022 );
xor \U$13176 ( \14024 , \13945 , \14023 );
xor \U$13177 ( \14025 , \13916 , \13921 );
xor \U$13178 ( \14026 , \14025 , \13924 );
and \U$13179 ( \14027 , \14024 , \14026 );
and \U$13180 ( \14028 , \13945 , \14023 );
or \U$13181 ( \14029 , \14027 , \14028 );
xor \U$13182 ( \14030 , \13927 , \13929 );
xor \U$13183 ( \14031 , \14030 , \13932 );
and \U$13184 ( \14032 , \14029 , \14031 );
nand \U$13185 ( \14033 , \13364_nG22e4 , \12179 );
or \U$13186 ( \14034 , \12110 , \13162_nG2320 );
nand \U$13187 ( \14035 , \14034 , \12315 );
and \U$13188 ( \14036 , \14033 , \14035 );
and \U$13189 ( \14037 , \12318 , \13162_nG2320 );
and \U$13190 ( \14038 , \13364_nG22e4 , \12182 );
nor \U$13191 ( \14039 , \14036 , \14037 , \14038 );
nand \U$13192 ( \14040 , \13122_nG2354 , \12380 );
or \U$13193 ( \14041 , \12337 , \12922_nG2391 );
nand \U$13194 ( \14042 , \14041 , \12527 );
and \U$13195 ( \14043 , \14040 , \14042 );
and \U$13196 ( \14044 , \12530 , \12922_nG2391 );
and \U$13197 ( \14045 , \13122_nG2354 , \12383 );
nor \U$13198 ( \14046 , \14043 , \14044 , \14045 );
xor \U$13199 ( \14047 , \14039 , \14046 );
nand \U$13200 ( \14048 , \13481_nG22ab , \12014 );
or \U$13201 ( \14049 , \11964 , \13637_nG2273 );
nand \U$13202 ( \14050 , \14049 , \12020 );
and \U$13203 ( \14051 , \14048 , \14050 );
and \U$13204 ( \14052 , \12016 , \13637_nG2273 );
and \U$13205 ( \14053 , \13481_nG22ab , \12125 );
nor \U$13206 ( \14054 , \14051 , \14052 , \14053 );
and \U$13207 ( \14055 , \14047 , \14054 );
and \U$13208 ( \14056 , \14039 , \14046 );
or \U$13209 ( \14057 , \14055 , \14056 );
nand \U$13210 ( \14058 , \12881_nG23c5 , \12586 );
or \U$13211 ( \14059 , \12541 , \12706_nG2723 );
nand \U$13212 ( \14060 , \14059 , \12753 );
and \U$13213 ( \14061 , \14058 , \14060 );
and \U$13214 ( \14062 , \12756 , \12706_nG2723 );
and \U$13215 ( \14063 , \12881_nG23c5 , \12588 );
nor \U$13216 ( \14064 , \14061 , \14062 , \14063 );
and \U$13217 ( \14065 , \12577 , \13012 );
not \U$13218 ( \14066 , \12662_nG27f3 );
and \U$13219 ( \14067 , \12850 , \14066 );
and \U$13220 ( \14068 , \12515_nG28d0 , \13015 );
nor \U$13221 ( \14069 , \14065 , \14067 , \14068 );
xor \U$13222 ( \14070 , \14064 , \14069 );
and \U$13223 ( \14071 , \14070 , \11848 );
and \U$13224 ( \14072 , \14064 , \14069 );
or \U$13225 ( \14073 , \14071 , \14072 );
xor \U$13226 ( \14074 , \14057 , \14073 );
xor \U$13227 ( \14075 , \13982 , \13989 );
xor \U$13228 ( \14076 , \14075 , \13997 );
and \U$13229 ( \14077 , \14074 , \14076 );
and \U$13230 ( \14078 , \14057 , \14073 );
or \U$13231 ( \14079 , \14077 , \14078 );
xor \U$13232 ( \14080 , \13952 , \13974 );
xor \U$13233 ( \14081 , \14080 , \14000 );
xor \U$13234 ( \14082 , \14079 , \14081 );
xor \U$13235 ( \14083 , \13872 , \13876 );
xor \U$13236 ( \14084 , \14083 , \11795 );
xor \U$13237 ( \14085 , \14008 , \14015 );
xor \U$13238 ( \14086 , \14084 , \14085 );
and \U$13239 ( \14087 , \14082 , \14086 );
and \U$13240 ( \14088 , \14079 , \14081 );
or \U$13241 ( \14089 , \14087 , \14088 );
xor \U$13242 ( \14090 , \14003 , \14005 );
xor \U$13243 ( \14091 , \14090 , \14020 );
xor \U$13244 ( \14092 , \14089 , \14091 );
xnor \U$13245 ( \14093 , \13944 , \13942 );
xor \U$13246 ( \14094 , \14092 , \14093 );
not \U$13247 ( \14095 , \14094 );
xor \U$13248 ( \14096 , \14079 , \14081 );
xor \U$13249 ( \14097 , \14096 , \14086 );
nand \U$13250 ( \14098 , \12922_nG2391 , \12586 );
or \U$13251 ( \14099 , \12541 , \12881_nG23c5 );
nand \U$13252 ( \14100 , \14099 , \12753 );
and \U$13253 ( \14101 , \14098 , \14100 );
and \U$13254 ( \14102 , \12756 , \12881_nG23c5 );
and \U$13255 ( \14103 , \12922_nG2391 , \12588 );
nor \U$13256 ( \14104 , \14101 , \14102 , \14103 );
not \U$13257 ( \14105 , \14104 );
and \U$13258 ( \14106 , \14066 , \13012 );
not \U$13259 ( \14107 , \12706_nG2723 );
and \U$13260 ( \14108 , \12850 , \14107 );
and \U$13261 ( \14109 , \12662_nG27f3 , \13015 );
nor \U$13262 ( \14110 , \14106 , \14108 , \14109 );
not \U$13263 ( \14111 , \14110 );
and \U$13264 ( \14112 , \14105 , \14111 );
and \U$13265 ( \14113 , \14104 , \14110 );
nand \U$13266 ( \14114 , \13162_nG2320 , \12380 );
or \U$13267 ( \14115 , \12337 , \13122_nG2354 );
nand \U$13268 ( \14116 , \14115 , \12527 );
and \U$13269 ( \14117 , \14114 , \14116 );
and \U$13270 ( \14118 , \12530 , \13122_nG2354 );
and \U$13271 ( \14119 , \13162_nG2320 , \12383 );
nor \U$13272 ( \14120 , \14117 , \14118 , \14119 );
nor \U$13273 ( \14121 , \14113 , \14120 );
nor \U$13274 ( \14122 , \14112 , \14121 );
xor \U$13275 ( \14123 , \14039 , \14046 );
xor \U$13276 ( \14124 , \14123 , \14054 );
and \U$13277 ( \14125 , \14122 , \14124 );
not \U$13278 ( \14126 , \13726_nG223a );
and \U$13279 ( \14127 , \14126 , \11888 );
and \U$13280 ( \14128 , \13726_nG223a , \11920 );
not \U$13281 ( \14129 , \11917 );
nor \U$13282 ( \14130 , \14127 , \14128 , \14129 );
xor \U$13283 ( \14131 , \14039 , \14046 );
xor \U$13284 ( \14132 , \14131 , \14054 );
and \U$13285 ( \14133 , \14130 , \14132 );
and \U$13286 ( \14134 , \14122 , \14130 );
or \U$13287 ( \14135 , \14125 , \14133 , \14134 );
xor \U$13288 ( \14136 , \13959 , \13963 );
xor \U$13289 ( \14137 , \14136 , \13971 );
xor \U$13290 ( \14138 , \14135 , \14137 );
xor \U$13291 ( \14139 , \14057 , \14073 );
xor \U$13292 ( \14140 , \14139 , \14076 );
and \U$13293 ( \14141 , \14138 , \14140 );
and \U$13294 ( \14142 , \14135 , \14137 );
or \U$13295 ( \14143 , \14141 , \14142 );
nor \U$13296 ( \14144 , \14097 , \14143 );
xor \U$13297 ( \14145 , \14095 , \14144 );
and \U$13298 ( \14146 , \14097 , \14143 );
nor \U$13299 ( \14147 , \14146 , \14144 );
xor \U$13300 ( \14148 , \14135 , \14137 );
xor \U$13301 ( \14149 , \14148 , \14140 );
nand \U$13302 ( \14150 , \13122_nG2354 , \12586 );
or \U$13303 ( \14151 , \12541 , \12922_nG2391 );
nand \U$13304 ( \14152 , \14151 , \12753 );
and \U$13305 ( \14153 , \14150 , \14152 );
and \U$13306 ( \14154 , \12756 , \12922_nG2391 );
and \U$13307 ( \14155 , \13122_nG2354 , \12588 );
nor \U$13308 ( \14156 , \14153 , \14154 , \14155 );
and \U$13309 ( \14157 , \14107 , \13012 );
not \U$13310 ( \14158 , \12881_nG23c5 );
and \U$13311 ( \14159 , \12850 , \14158 );
and \U$13312 ( \14160 , \12706_nG2723 , \13015 );
nor \U$13313 ( \14161 , \14157 , \14159 , \14160 );
xor \U$13314 ( \14162 , \14156 , \14161 );
and \U$13315 ( \14163 , \14162 , \11964 );
and \U$13316 ( \14164 , \14156 , \14161 );
or \U$13317 ( \14165 , \14163 , \14164 );
nand \U$13318 ( \14166 , \13481_nG22ab , \12179 );
or \U$13319 ( \14167 , \12110 , \13364_nG22e4 );
nand \U$13320 ( \14168 , \14167 , \12315 );
and \U$13321 ( \14169 , \14166 , \14168 );
and \U$13322 ( \14170 , \12318 , \13364_nG22e4 );
and \U$13323 ( \14171 , \13481_nG22ab , \12182 );
nor \U$13324 ( \14172 , \14169 , \14170 , \14171 );
xor \U$13325 ( \14173 , \14165 , \14172 );
nand \U$13326 ( \14174 , \13637_nG2273 , \12179 );
or \U$13327 ( \14175 , \12110 , \13481_nG22ab );
nand \U$13328 ( \14176 , \14175 , \12315 );
and \U$13329 ( \14177 , \14174 , \14176 );
and \U$13330 ( \14178 , \12318 , \13481_nG22ab );
and \U$13331 ( \14179 , \13637_nG2273 , \12182 );
nor \U$13332 ( \14180 , \14177 , \14178 , \14179 );
nand \U$13333 ( \14181 , \13364_nG22e4 , \12380 );
or \U$13334 ( \14182 , \12337 , \13162_nG2320 );
nand \U$13335 ( \14183 , \14182 , \12527 );
and \U$13336 ( \14184 , \14181 , \14183 );
and \U$13337 ( \14185 , \12530 , \13162_nG2320 );
and \U$13338 ( \14186 , \13364_nG22e4 , \12383 );
nor \U$13339 ( \14187 , \14184 , \14185 , \14186 );
xor \U$13340 ( \14188 , \14180 , \14187 );
and \U$13341 ( \14189 , \12125 , \13726_nG223a );
nand \U$13342 ( \14190 , \13726_nG223a , \12014 );
and \U$13343 ( \14191 , \14190 , \12018 );
nor \U$13344 ( \14192 , \14189 , \14191 );
and \U$13345 ( \14193 , \14188 , \14192 );
and \U$13346 ( \14194 , \14180 , \14187 );
or \U$13347 ( \14195 , \14193 , \14194 );
and \U$13348 ( \14196 , \14173 , \14195 );
and \U$13349 ( \14197 , \14165 , \14172 );
or \U$13350 ( \14198 , \14196 , \14197 );
xor \U$13351 ( \14199 , \14064 , \14069 );
xor \U$13352 ( \14200 , \14199 , \11848 );
nand \U$13353 ( \14201 , \14198 , \14200 );
not \U$13354 ( \14202 , \14104 );
xor \U$13355 ( \14203 , \14110 , \14120 );
not \U$13356 ( \14204 , \14203 );
or \U$13357 ( \14205 , \14202 , \14204 );
or \U$13358 ( \14206 , \14203 , \14104 );
nand \U$13359 ( \14207 , \14205 , \14206 );
not \U$13360 ( \14208 , \13637_nG2273 );
or \U$13361 ( \14209 , \12188 , \14208 );
or \U$13362 ( \14210 , \14126 , \12190 );
or \U$13363 ( \14211 , \12124 , \14208 );
or \U$13364 ( \14212 , \11964 , \13726_nG223a );
nand \U$13365 ( \14213 , \14212 , \12020 );
nand \U$13366 ( \14214 , \14211 , \14213 );
nand \U$13367 ( \14215 , \14209 , \14210 , \14214 );
and \U$13368 ( \14216 , \14207 , \14215 );
and \U$13369 ( \14217 , \14201 , \14216 );
nor \U$13370 ( \14218 , \14200 , \14198 );
nor \U$13371 ( \14219 , \14217 , \14218 );
nor \U$13372 ( \14220 , \14149 , \14219 );
xor \U$13373 ( \14221 , \14147 , \14220 );
not \U$13374 ( \14222 , \14216 );
not \U$13375 ( \14223 , \14218 );
nand \U$13376 ( \14224 , \14223 , \14201 );
not \U$13377 ( \14225 , \14224 );
or \U$13378 ( \14226 , \14222 , \14225 );
or \U$13379 ( \14227 , \14224 , \14216 );
nand \U$13380 ( \14228 , \14226 , \14227 );
xor \U$13381 ( \14229 , \14039 , \14046 );
xor \U$13382 ( \14230 , \14229 , \14054 );
xor \U$13383 ( \14231 , \14122 , \14130 );
xor \U$13384 ( \14232 , \14230 , \14231 );
not \U$13385 ( \14233 , \14232 );
xor \U$13386 ( \14234 , \14228 , \14233 );
xor \U$13387 ( \14235 , \14165 , \14172 );
xor \U$13388 ( \14236 , \14235 , \14195 );
nand \U$13389 ( \14237 , \13162_nG2320 , \12586 );
or \U$13390 ( \14238 , \12541 , \13122_nG2354 );
nand \U$13391 ( \14239 , \14238 , \12753 );
and \U$13392 ( \14240 , \14237 , \14239 );
and \U$13393 ( \14241 , \12756 , \13122_nG2354 );
and \U$13394 ( \14242 , \13162_nG2320 , \12588 );
nor \U$13395 ( \14243 , \14240 , \14241 , \14242 );
and \U$13396 ( \14244 , \14158 , \13012 );
not \U$13397 ( \14245 , \12922_nG2391 );
and \U$13398 ( \14246 , \12850 , \14245 );
and \U$13399 ( \14247 , \12881_nG23c5 , \13015 );
nor \U$13400 ( \14248 , \14244 , \14246 , \14247 );
xor \U$13401 ( \14249 , \14243 , \14248 );
nand \U$13402 ( \14250 , \13481_nG22ab , \12380 );
or \U$13403 ( \14251 , \12337 , \13364_nG22e4 );
nand \U$13404 ( \14252 , \14251 , \12527 );
and \U$13405 ( \14253 , \14250 , \14252 );
and \U$13406 ( \14254 , \12530 , \13364_nG22e4 );
and \U$13407 ( \14255 , \13481_nG22ab , \12383 );
nor \U$13408 ( \14256 , \14253 , \14254 , \14255 );
and \U$13409 ( \14257 , \14249 , \14256 );
and \U$13410 ( \14258 , \14243 , \14248 );
or \U$13411 ( \14259 , \14257 , \14258 );
xor \U$13412 ( \14260 , \14156 , \14161 );
xor \U$13413 ( \14261 , \14260 , \11964 );
and \U$13414 ( \14262 , \14259 , \14261 );
xor \U$13415 ( \14263 , \14180 , \14187 );
xor \U$13416 ( \14264 , \14263 , \14192 );
xor \U$13417 ( \14265 , \14156 , \14161 );
xor \U$13418 ( \14266 , \14265 , \11964 );
and \U$13419 ( \14267 , \14264 , \14266 );
and \U$13420 ( \14268 , \14259 , \14264 );
or \U$13421 ( \14269 , \14262 , \14267 , \14268 );
nor \U$13422 ( \14270 , \14236 , \14269 );
xor \U$13423 ( \14271 , \14207 , \14215 );
or \U$13424 ( \14272 , \14270 , \14271 );
nand \U$13425 ( \14273 , \14269 , \14236 );
nand \U$13426 ( \14274 , \14272 , \14273 );
not \U$13427 ( \14275 , \14274 );
xor \U$13428 ( \14276 , \14234 , \14275 );
not \U$13429 ( \14277 , \14273 );
nor \U$13430 ( \14278 , \14277 , \14270 );
not \U$13431 ( \14279 , \14278 );
not \U$13432 ( \14280 , \14271 );
and \U$13433 ( \14281 , \14279 , \14280 );
and \U$13434 ( \14282 , \14278 , \14271 );
nor \U$13435 ( \14283 , \14281 , \14282 );
xor \U$13436 ( \14284 , \14156 , \14161 );
xor \U$13437 ( \14285 , \14284 , \11964 );
xor \U$13438 ( \14286 , \14259 , \14264 );
xor \U$13439 ( \14287 , \14285 , \14286 );
nand \U$13440 ( \14288 , \13364_nG22e4 , \12586 );
or \U$13441 ( \14289 , \12541 , \13162_nG2320 );
nand \U$13442 ( \14290 , \14289 , \12753 );
and \U$13443 ( \14291 , \14288 , \14290 );
and \U$13444 ( \14292 , \12756 , \13162_nG2320 );
and \U$13445 ( \14293 , \13364_nG22e4 , \12588 );
nor \U$13446 ( \14294 , \14291 , \14292 , \14293 );
and \U$13447 ( \14295 , \14245 , \13012 );
not \U$13448 ( \14296 , \13122_nG2354 );
and \U$13449 ( \14297 , \12850 , \14296 );
and \U$13450 ( \14298 , \12922_nG2391 , \13015 );
nor \U$13451 ( \14299 , \14295 , \14297 , \14298 );
xor \U$13452 ( \14300 , \14294 , \14299 );
and \U$13453 ( \14301 , \14300 , \12110 );
and \U$13454 ( \14302 , \14294 , \14299 );
or \U$13455 ( \14303 , \14301 , \14302 );
nand \U$13456 ( \14304 , \13726_nG223a , \12179 );
or \U$13457 ( \14305 , \12110 , \13637_nG2273 );
nand \U$13458 ( \14306 , \14305 , \12315 );
and \U$13459 ( \14307 , \14304 , \14306 );
and \U$13460 ( \14308 , \12318 , \13637_nG2273 );
and \U$13461 ( \14309 , \13726_nG223a , \12182 );
nor \U$13462 ( \14310 , \14307 , \14308 , \14309 );
nand \U$13463 ( \14311 , \14303 , \14310 );
or \U$13464 ( \14312 , \12390 , \14126 );
or \U$13465 ( \14313 , \13726_nG223a , \12110 );
nand \U$13466 ( \14314 , \14312 , \14313 , \12315 );
not \U$13467 ( \14315 , \14314 );
nand \U$13468 ( \14316 , \13637_nG2273 , \12380 );
or \U$13469 ( \14317 , \12337 , \13481_nG22ab );
nand \U$13470 ( \14318 , \14317 , \12527 );
and \U$13471 ( \14319 , \14316 , \14318 );
and \U$13472 ( \14320 , \12530 , \13481_nG22ab );
and \U$13473 ( \14321 , \13637_nG2273 , \12383 );
nor \U$13474 ( \14322 , \14319 , \14320 , \14321 );
nor \U$13475 ( \14323 , \14315 , \14322 );
and \U$13476 ( \14324 , \14311 , \14323 );
nor \U$13477 ( \14325 , \14310 , \14303 );
nor \U$13478 ( \14326 , \14324 , \14325 );
nor \U$13479 ( \14327 , \14287 , \14326 );
xor \U$13480 ( \14328 , \14283 , \14327 );
xor \U$13481 ( \14329 , \14243 , \14248 );
xor \U$13482 ( \14330 , \14329 , \14256 );
not \U$13483 ( \14331 , \14330 );
not \U$13484 ( \14332 , \14323 );
not \U$13485 ( \14333 , \14325 );
nand \U$13486 ( \14334 , \14333 , \14311 );
not \U$13487 ( \14335 , \14334 );
or \U$13488 ( \14336 , \14332 , \14335 );
or \U$13489 ( \14337 , \14334 , \14323 );
nand \U$13490 ( \14338 , \14336 , \14337 );
xor \U$13491 ( \14339 , \14331 , \14338 );
xor \U$13492 ( \14340 , \14294 , \14299 );
xor \U$13493 ( \14341 , \14340 , \12110 );
nand \U$13494 ( \14342 , \13481_nG22ab , \12586 );
or \U$13495 ( \14343 , \12541 , \13364_nG22e4 );
nand \U$13496 ( \14344 , \14343 , \12753 );
and \U$13497 ( \14345 , \14342 , \14344 );
and \U$13498 ( \14346 , \12756 , \13364_nG22e4 );
and \U$13499 ( \14347 , \13481_nG22ab , \12588 );
nor \U$13500 ( \14348 , \14345 , \14346 , \14347 );
and \U$13501 ( \14349 , \14296 , \13012 );
not \U$13502 ( \14350 , \13162_nG2320 );
and \U$13503 ( \14351 , \12850 , \14350 );
and \U$13504 ( \14352 , \13122_nG2354 , \13015 );
nor \U$13505 ( \14353 , \14349 , \14351 , \14352 );
xor \U$13506 ( \14354 , \14348 , \14353 );
nand \U$13507 ( \14355 , \13726_nG223a , \12380 );
or \U$13508 ( \14356 , \12337 , \13637_nG2273 );
nand \U$13509 ( \14357 , \14356 , \12527 );
and \U$13510 ( \14358 , \14355 , \14357 );
and \U$13511 ( \14359 , \12530 , \13637_nG2273 );
and \U$13512 ( \14360 , \13726_nG223a , \12383 );
nor \U$13513 ( \14361 , \14358 , \14359 , \14360 );
and \U$13514 ( \14362 , \14354 , \14361 );
and \U$13515 ( \14363 , \14348 , \14353 );
or \U$13516 ( \14364 , \14362 , \14363 );
and \U$13517 ( \14365 , \14341 , \14364 );
or \U$13518 ( \14366 , \14341 , \14364 );
not \U$13519 ( \14367 , \14314 );
not \U$13520 ( \14368 , \14322 );
and \U$13521 ( \14369 , \14367 , \14368 );
and \U$13522 ( \14370 , \14314 , \14322 );
nor \U$13523 ( \14371 , \14369 , \14370 );
and \U$13524 ( \14372 , \14366 , \14371 );
nor \U$13525 ( \14373 , \14365 , \14372 );
xor \U$13526 ( \14374 , \14339 , \14373 );
xor \U$13527 ( \14375 , \14341 , \14364 );
and \U$13528 ( \14376 , \14371 , \14375 );
nor \U$13529 ( \14377 , \14371 , \14375 );
or \U$13530 ( \14378 , \14376 , \14377 );
xor \U$13531 ( \14379 , \14348 , \14353 );
xor \U$13532 ( \14380 , \14379 , \14361 );
and \U$13533 ( \14381 , \14350 , \13012 );
not \U$13534 ( \14382 , \13364_nG22e4 );
and \U$13535 ( \14383 , \12850 , \14382 );
and \U$13536 ( \14384 , \13162_nG2320 , \13015 );
nor \U$13537 ( \14385 , \14381 , \14383 , \14384 );
xor \U$13538 ( \14386 , \12337 , \14385 );
nand \U$13539 ( \14387 , \13637_nG2273 , \12586 );
or \U$13540 ( \14388 , \12541 , \13481_nG22ab );
nand \U$13541 ( \14389 , \14388 , \12753 );
and \U$13542 ( \14390 , \14387 , \14389 );
and \U$13543 ( \14391 , \12756 , \13481_nG22ab );
and \U$13544 ( \14392 , \13637_nG2273 , \12588 );
nor \U$13545 ( \14393 , \14390 , \14391 , \14392 );
and \U$13546 ( \14394 , \14386 , \14393 );
and \U$13547 ( \14395 , \12337 , \14385 );
or \U$13548 ( \14396 , \14394 , \14395 );
nor \U$13549 ( \14397 , \14380 , \14396 );
nand \U$13550 ( \14398 , \14378 , \14397 );
or \U$13551 ( \14399 , \14376 , \14377 , \14397 );
not \U$13552 ( \14400 , \14380 );
nand \U$13553 ( \14401 , \14400 , \14396 );
xor \U$13554 ( \14402 , \12337 , \14385 );
xor \U$13555 ( \14403 , \14402 , \14393 );
not \U$13556 ( \14404 , \14403 );
or \U$13557 ( \14405 , \12595 , \14126 );
or \U$13558 ( \14406 , \13726_nG223a , \12337 );
nand \U$13559 ( \14407 , \14405 , \14406 , \12527 );
nand \U$13560 ( \14408 , \14404 , \14407 );
not \U$13561 ( \14409 , \14396 );
nand \U$13562 ( \14410 , \14409 , \14380 );
and \U$13563 ( \14411 , \14401 , \14408 , \14410 );
not \U$13564 ( \14412 , \14403 );
not \U$13565 ( \14413 , \14407 );
or \U$13566 ( \14414 , \14412 , \14413 );
or \U$13567 ( \14415 , \14407 , \14403 );
nand \U$13568 ( \14416 , \14414 , \14415 );
nand \U$13569 ( \14417 , \13726_nG223a , \12586 );
or \U$13570 ( \14418 , \12541 , \13637_nG2273 );
nand \U$13571 ( \14419 , \14418 , \12753 );
and \U$13572 ( \14420 , \14417 , \14419 );
and \U$13573 ( \14421 , \12756 , \13637_nG2273 );
and \U$13574 ( \14422 , \13726_nG223a , \12588 );
nor \U$13575 ( \14423 , \14420 , \14421 , \14422 );
and \U$13576 ( \14424 , \14382 , \13012 );
not \U$13577 ( \14425 , \13481_nG22ab );
and \U$13578 ( \14426 , \12850 , \14425 );
and \U$13579 ( \14427 , \13364_nG22e4 , \13015 );
nor \U$13580 ( \14428 , \14424 , \14426 , \14427 );
nor \U$13581 ( \14429 , \14423 , \14428 );
or \U$13582 ( \14430 , \14416 , \14429 );
or \U$13583 ( \14431 , \13169 , \14425 );
or \U$13584 ( \14432 , \13481_nG22ab , \12852 );
or \U$13585 ( \14433 , \13637_nG2273 , \12851 );
nand \U$13586 ( \14434 , \14431 , \14432 , \14433 );
and \U$13587 ( \14435 , \14434 , \12542 );
not \U$13588 ( \14436 , \14435 );
and \U$13589 ( \14437 , \14423 , \14428 );
nor \U$13590 ( \14438 , \14437 , \14429 );
not \U$13591 ( \14439 , \14438 );
or \U$13592 ( \14440 , \14436 , \14439 );
or \U$13593 ( \14441 , \14438 , \14435 );
and \U$13594 ( \14442 , \12849 , \13637_nG2273 );
nor \U$13595 ( \14443 , \14442 , \12535 , \13726_nG223a );
xor \U$13596 ( \14444 , \14434 , \12542 );
or \U$13597 ( \14445 , \14443 , \14444 );
nand \U$13598 ( \14446 , \14441 , \14445 );
and \U$13599 ( \14447 , \14444 , \14443 );
not \U$13600 ( \14448 , \12756 );
and \U$13601 ( \14449 , \14448 , \13726_nG223a );
and \U$13602 ( \14450 , \14126 , \12541 );
nor \U$13603 ( \14451 , \14449 , \14450 );
not \U$13604 ( \14452 , \12753 );
nor \U$13605 ( \14453 , \14447 , \14451 , \14452 );
or \U$13606 ( \14454 , \14446 , \14453 );
nand \U$13607 ( \14455 , \14440 , \14454 );
and \U$13608 ( \14456 , \14430 , \14455 );
and \U$13609 ( \14457 , \14429 , \14416 );
nor \U$13610 ( \14458 , \14456 , \14457 );
nor \U$13611 ( \14459 , \14411 , \14458 );
and \U$13612 ( \14460 , \14401 , \14410 );
nor \U$13613 ( \14461 , \14460 , \14408 );
or \U$13614 ( \14462 , \14459 , \14461 );
nand \U$13615 ( \14463 , \14399 , \14462 );
nand \U$13616 ( \14464 , \14398 , \14463 );
and \U$13617 ( \14465 , \14374 , \14464 );
and \U$13618 ( \14466 , \14339 , \14373 );
or \U$13619 ( \14467 , \14465 , \14466 );
and \U$13620 ( \14468 , \14331 , \14338 );
xor \U$13621 ( \14469 , \14467 , \14468 );
and \U$13622 ( \14470 , \14287 , \14326 );
nor \U$13623 ( \14471 , \14470 , \14327 );
and \U$13624 ( \14472 , \14469 , \14471 );
and \U$13625 ( \14473 , \14467 , \14468 );
or \U$13626 ( \14474 , \14472 , \14473 );
and \U$13627 ( \14475 , \14328 , \14474 );
and \U$13628 ( \14476 , \14283 , \14327 );
or \U$13629 ( \14477 , \14475 , \14476 );
and \U$13630 ( \14478 , \14276 , \14477 );
and \U$13631 ( \14479 , \14234 , \14275 );
or \U$13632 ( \14480 , \14478 , \14479 );
and \U$13633 ( \14481 , \14228 , \14233 );
xor \U$13634 ( \14482 , \14480 , \14481 );
and \U$13635 ( \14483 , \14149 , \14219 );
nor \U$13636 ( \14484 , \14483 , \14220 );
and \U$13637 ( \14485 , \14482 , \14484 );
and \U$13638 ( \14486 , \14480 , \14481 );
or \U$13639 ( \14487 , \14485 , \14486 );
and \U$13640 ( \14488 , \14221 , \14487 );
and \U$13641 ( \14489 , \14147 , \14220 );
or \U$13642 ( \14490 , \14488 , \14489 );
and \U$13643 ( \14491 , \14145 , \14490 );
and \U$13644 ( \14492 , \14095 , \14144 );
or \U$13645 ( \14493 , \14491 , \14492 );
xor \U$13646 ( \14494 , \14089 , \14091 );
and \U$13647 ( \14495 , \14494 , \14093 );
and \U$13648 ( \14496 , \14089 , \14091 );
or \U$13649 ( \14497 , \14495 , \14496 );
xor \U$13650 ( \14498 , \13945 , \14023 );
xor \U$13651 ( \14499 , \14498 , \14026 );
nand \U$13652 ( \14500 , \14497 , \14499 );
and \U$13653 ( \14501 , \14493 , \14500 );
nor \U$13654 ( \14502 , \14499 , \14497 );
nor \U$13655 ( \14503 , \14501 , \14502 );
xor \U$13656 ( \14504 , \13927 , \13929 );
xor \U$13657 ( \14505 , \14504 , \13932 );
and \U$13658 ( \14506 , \14503 , \14505 );
and \U$13659 ( \14507 , \14029 , \14503 );
or \U$13660 ( \14508 , \14032 , \14506 , \14507 );
and \U$13661 ( \14509 , \13940 , \14508 );
and \U$13662 ( \14510 , \13935 , \13939 );
or \U$13663 ( \14511 , \14509 , \14510 );
and \U$13664 ( \14512 , \13865 , \14511 );
and \U$13665 ( \14513 , \13782 , \13864 );
or \U$13666 ( \14514 , \14512 , \14513 );
not \U$13667 ( \14515 , \14514 );
and \U$13668 ( \14516 , \13780 , \14515 );
and \U$13669 ( \14517 , \13769 , \13779 );
or \U$13670 ( \14518 , \14516 , \14517 );
and \U$13671 ( \14519 , \13767 , \14518 );
and \U$13672 ( \14520 , \13600 , \13766 );
or \U$13673 ( \14521 , \14519 , \14520 );
and \U$13674 ( \14522 , \13598 , \14521 );
and \U$13675 ( \14523 , \13514 , \13597 );
or \U$13676 ( \14524 , \14522 , \14523 );
and \U$13677 ( \14525 , \13512 , \14524 );
and \U$13678 ( \14526 , \13334 , \13511 );
or \U$13679 ( \14527 , \14525 , \14526 );
and \U$13680 ( \14528 , \13332 , \14527 );
and \U$13681 ( \14529 , \13247 , \13331 );
or \U$13682 ( \14530 , \14528 , \14529 );
and \U$13683 ( \14531 , \13241 , \14530 );
and \U$13684 ( \14532 , \13238 , \13240 );
or \U$13685 ( \14533 , \14531 , \14532 );
and \U$13686 ( \14534 , \13064 , \14533 );
and \U$13687 ( \14535 , \12961 , \13063 );
or \U$13688 ( \14536 , \14534 , \14535 );
and \U$13689 ( \14537 , \12959 , \14536 );
and \U$13690 ( \14538 , \12810 , \12958 );
or \U$13691 ( \14539 , \14537 , \14538 );
and \U$13692 ( \14540 , \12808 , \14539 );
and \U$13693 ( \14541 , \12680 , \12807 );
or \U$13694 ( \14542 , \14540 , \14541 );
and \U$13695 ( \14543 , \12678 , \14542 );
and \U$13696 ( \14544 , \12571 , \12677 );
or \U$13697 ( \14545 , \14543 , \14544 );
and \U$13698 ( \14546 , \12567 , \14545 );
and \U$13699 ( \14547 , \12462 , \12566 );
or \U$13700 ( \14548 , \14546 , \14547 );
and \U$13701 ( \14549 , \12460 , \14548 );
and \U$13702 ( \14550 , \12457 , \12459 );
or \U$13703 ( \14551 , \14549 , \14550 );
and \U$13704 ( \14552 , \12372 , \14551 );
and \U$13705 ( \14553 , \12369 , \12371 );
or \U$13706 ( \14554 , \14552 , \14553 );
and \U$13707 ( \14555 , \12265 , \14554 );
and \U$13708 ( \14556 , \12262 , \12264 );
or \U$13709 ( \14557 , \14555 , \14556 );
and \U$13710 ( \14558 , \12101 , \14557 );
and \U$13711 ( \14559 , \12099 , \12100 );
or \U$13712 ( \14560 , \14558 , \14559 );
not \U$13713 ( \14561 , \14560 );
or \U$13714 ( \14562 , \11998 , \14561 );
or \U$13715 ( \14563 , \14560 , \11997 );
nand \U$13716 ( \14564 , \14562 , \14563 );
buf \U$13717 ( \14565 , \11427 );
buf \U$13718 ( \14566 , \7972 );
_DC g7eb ( \14567_nG7eb , \14565 , \14566 );
not \U$13719 ( \14568 , \14567_nG7eb );
buf \U$13720 ( \14569 , \11456 );
_DC g80c ( \14570_nG80c , \14569 , \14566 );
not \U$13721 ( \14571 , \14570_nG80c );
buf \U$13722 ( \14572 , \8369 );
buf \U$13723 ( \14573 , \7972 );
_DC g906 ( \14574_nG906 , \14572 , \14573 );
not \U$13724 ( \14575 , \14574_nG906 );
not \U$13725 ( \14576 , \14575 );
buf \U$13726 ( \14577 , \11685 );
_DC g908 ( \14578_nG908 , \14577 , \14566 );
not \U$13727 ( \14579 , \14578_nG908 );
and \U$13728 ( \14580 , \14576 , \14579 );
buf \U$13729 ( \14581 , \8400 );
_DC g925 ( \14582_nG925 , \14581 , \14573 );
nor \U$13730 ( \14583 , \14580 , \14582_nG925 );
buf \U$13731 ( \14584 , \11713 );
_DC g927 ( \14585_nG927 , \14584 , \14566 );
and \U$13732 ( \14586 , \14583 , \14585_nG927 );
and \U$13733 ( \14587 , \14578_nG908 , \14575 );
nor \U$13734 ( \14588 , \14586 , \14587 );
buf \U$13735 ( \14589 , \8336 );
_DC g8e5 ( \14590_nG8e5 , \14589 , \14573 );
or \U$13736 ( \14591 , \14588 , \14590_nG8e5 );
not \U$13737 ( \14592 , \14590_nG8e5 );
not \U$13738 ( \14593 , \14588 );
or \U$13739 ( \14594 , \14592 , \14593 );
buf \U$13740 ( \14595 , \11656 );
_DC g8e7 ( \14596_nG8e7 , \14595 , \14566 );
nand \U$13741 ( \14597 , \14594 , \14596_nG8e7 );
nand \U$13742 ( \14598 , \14591 , \14597 );
buf \U$13743 ( \14599 , \11628 );
_DC g8c8 ( \14600_nG8c8 , \14599 , \14566 );
and \U$13744 ( \14601 , \14598 , \14600_nG8c8 );
not \U$13745 ( \14602 , \14598 );
not \U$13746 ( \14603 , \14600_nG8c8 );
and \U$13747 ( \14604 , \14602 , \14603 );
buf \U$13748 ( \14605 , \8300 );
_DC g8c6 ( \14606_nG8c6 , \14605 , \14573 );
nor \U$13749 ( \14607 , \14604 , \14606_nG8c6 );
nor \U$13750 ( \14608 , \14601 , \14607 );
buf \U$13751 ( \14609 , \11600 );
_DC g8a9 ( \14610_nG8a9 , \14609 , \14566 );
not \U$13752 ( \14611 , \14610_nG8a9 );
buf \U$13753 ( \14612 , \8268 );
_DC g8a7 ( \14613_nG8a7 , \14612 , \14573 );
and \U$13754 ( \14614 , \14611 , \14613_nG8a7 );
or \U$13755 ( \14615 , \14608 , \14614 );
or \U$13756 ( \14616 , \14613_nG8a7 , \14611 );
nand \U$13757 ( \14617 , \14615 , \14616 );
buf \U$13758 ( \14618 , \11571 );
_DC g88a ( \14619_nG88a , \14618 , \14566 );
and \U$13759 ( \14620 , \14617 , \14619_nG88a );
not \U$13760 ( \14621 , \14617 );
not \U$13761 ( \14622 , \14619_nG88a );
and \U$13762 ( \14623 , \14621 , \14622 );
buf \U$13763 ( \14624 , \8232 );
_DC g888 ( \14625_nG888 , \14624 , \14573 );
nor \U$13764 ( \14626 , \14623 , \14625_nG888 );
nor \U$13765 ( \14627 , \14620 , \14626 );
buf \U$13766 ( \14628 , \11543 );
_DC g86b ( \14629_nG86b , \14628 , \14566 );
not \U$13767 ( \14630 , \14629_nG86b );
buf \U$13768 ( \14631 , \8196 );
_DC g869 ( \14632_nG869 , \14631 , \14573 );
and \U$13769 ( \14633 , \14630 , \14632_nG869 );
or \U$13770 ( \14634 , \14627 , \14633 );
or \U$13771 ( \14635 , \14632_nG869 , \14630 );
nand \U$13772 ( \14636 , \14634 , \14635 );
buf \U$13773 ( \14637 , \11514 );
_DC g84c ( \14638_nG84c , \14637 , \14566 );
and \U$13774 ( \14639 , \14636 , \14638_nG84c );
not \U$13775 ( \14640 , \14636 );
not \U$13776 ( \14641 , \14638_nG84c );
and \U$13777 ( \14642 , \14640 , \14641 );
buf \U$13778 ( \14643 , \8160 );
_DC g84a ( \14644_nG84a , \14643 , \14573 );
nor \U$13779 ( \14645 , \14642 , \14644_nG84a );
nor \U$13780 ( \14646 , \14639 , \14645 );
buf \U$13781 ( \14647 , \8122 );
_DC g829 ( \14648_nG829 , \14647 , \14573 );
or \U$13782 ( \14649 , \14646 , \14648_nG829 );
not \U$13783 ( \14650 , \14648_nG829 );
not \U$13784 ( \14651 , \14646 );
or \U$13785 ( \14652 , \14650 , \14651 );
buf \U$13786 ( \14653 , \11485 );
_DC g82b ( \14654_nG82b , \14653 , \14566 );
nand \U$13787 ( \14655 , \14652 , \14654_nG82b );
nand \U$13788 ( \14656 , \14649 , \14655 );
not \U$13789 ( \14657 , \14656 );
or \U$13790 ( \14658 , \14571 , \14657 );
nor \U$13791 ( \14659 , \14656 , \14570_nG80c );
buf \U$13792 ( \14660 , \8086 );
_DC g80a ( \14661_nG80a , \14660 , \14573 );
or \U$13793 ( \14662 , \14659 , \14661_nG80a );
nand \U$13794 ( \14663 , \14658 , \14662 );
not \U$13795 ( \14664 , \14663 );
or \U$13796 ( \14665 , \14568 , \14664 );
nor \U$13797 ( \14666 , \14663 , \14567_nG7eb );
buf \U$13798 ( \14667 , \8048 );
_DC g7e9 ( \14668_nG7e9 , \14667 , \14573 );
or \U$13799 ( \14669 , \14666 , \14668_nG7e9 );
nand \U$13800 ( \14670 , \14665 , \14669 );
buf \U$13801 ( \14671 , \11399 );
_DC g7ca ( \14672_nG7ca , \14671 , \14566 );
and \U$13802 ( \14673 , \14670 , \14672_nG7ca );
not \U$13803 ( \14674 , \14670 );
not \U$13804 ( \14675 , \14672_nG7ca );
and \U$13805 ( \14676 , \14674 , \14675 );
buf \U$13806 ( \14677 , \8010 );
_DC g7c8 ( \14678_nG7c8 , \14677 , \14573 );
nor \U$13807 ( \14679 , \14676 , \14678_nG7c8 );
nor \U$13808 ( \14680 , \14673 , \14679 );
buf \U$13809 ( \14681 , \11369 );
_DC g7a9 ( \14682_nG7a9 , \14681 , \14566 );
not \U$13810 ( \14683 , \14682_nG7a9 );
buf \U$13811 ( \14684 , \7968 );
_DC g7a6 ( \14685_nG7a6 , \14684 , \14573 );
and \U$13812 ( \14686 , \14683 , \14685_nG7a6 );
or \U$13813 ( \14687 , \14680 , \14686 );
or \U$13814 ( \14688 , \14685_nG7a6 , \14683 );
nand \U$13815 ( \14689 , \14687 , \14688 );
buf \U$13816 ( \14690 , \11369 );
buf \U$13817 ( \14691 , \7972 );
_DC g62d ( \14692_nG62d , \14690 , \14691 );
nor \U$13818 ( \14693 , \7876 , RIaaa89a8_588);
nand \U$13819 ( \14694 , RIaaa9218_606, \14693 );
not \U$13820 ( \14695 , \14694 );
nand \U$13821 ( \14696 , RIaaa9290_607, \14695 );
not \U$13822 ( \14697 , \14696 );
nand \U$13823 ( \14698 , RIaaa9308_608, \14697 );
nor \U$13824 ( \14699 , \14698 , \8128 );
nand \U$13825 ( \14700 , RIaaa93f8_610, \14699 );
nor \U$13826 ( \14701 , \14700 , \8054 );
nand \U$13827 ( \14702 , RIaaa9470_611, \14701 );
not \U$13828 ( \14703 , \14702 );
nand \U$13829 ( \14704 , \14703 , RIaaa94e8_612);
not \U$13830 ( \14705 , \14704 );
not \U$13831 ( \14706 , RIaaa95d8_614);
and \U$13832 ( \14707 , \14705 , \14706 );
and \U$13833 ( \14708 , \14704 , RIaaa95d8_614);
nor \U$13834 ( \14709 , \14707 , \14708 );
nand \U$13835 ( \14710 , \14692_nG62d , \14709 );
or \U$13836 ( \14711 , \14709 , \14692_nG62d );
not \U$13837 ( \14712 , \14702 );
not \U$13838 ( \14713 , RIaaa94e8_612);
and \U$13839 ( \14714 , \14712 , \14713 );
and \U$13840 ( \14715 , \14702 , RIaaa94e8_612);
nor \U$13841 ( \14716 , \14714 , \14715 );
not \U$13842 ( \14717 , \14716 );
buf \U$13843 ( \14718 , \11399 );
_DC g64a ( \14719_nG64a , \14718 , \14691 );
not \U$13844 ( \14720 , \14719_nG64a );
and \U$13845 ( \14721 , \14717 , \14720 );
and \U$13846 ( \14722 , \14719_nG64a , \14716 );
buf \U$13847 ( \14723 , \11456 );
_DC g683 ( \14724_nG683 , \14723 , \14691 );
not \U$13848 ( \14725 , \14724_nG683 );
not \U$13849 ( \14726 , \14700 );
not \U$13850 ( \14727 , RIaaa9038_602);
and \U$13851 ( \14728 , \14726 , \14727 );
and \U$13852 ( \14729 , \14700 , RIaaa9038_602);
nor \U$13853 ( \14730 , \14728 , \14729 );
not \U$13854 ( \14731 , \14730 );
or \U$13855 ( \14732 , \14725 , \14731 );
or \U$13856 ( \14733 , \14730 , \14724_nG683 );
or \U$13857 ( \14734 , \14699 , RIaaa93f8_610);
nand \U$13858 ( \14735 , \14734 , \14700 );
buf \U$13859 ( \14736 , \11485 );
_DC g6a0 ( \14737_nG6a0 , \14736 , \14691 );
and \U$13860 ( \14738 , \14735 , \14737_nG6a0 );
buf \U$13861 ( \14739 , \11514 );
_DC g6bd ( \14740_nG6bd , \14739 , \14691 );
not \U$13862 ( \14741 , \14740_nG6bd );
not \U$13863 ( \14742 , \14698 );
not \U$13864 ( \14743 , RIaaa9380_609);
and \U$13865 ( \14744 , \14742 , \14743 );
and \U$13866 ( \14745 , \14698 , RIaaa9380_609);
nor \U$13867 ( \14746 , \14744 , \14745 );
not \U$13868 ( \14747 , \14746 );
or \U$13869 ( \14748 , \14741 , \14747 );
or \U$13870 ( \14749 , \14746 , \14740_nG6bd );
buf \U$13871 ( \14750 , \11543 );
_DC g6da ( \14751_nG6da , \14750 , \14691 );
or \U$13872 ( \14752 , \14697 , RIaaa9308_608);
nand \U$13873 ( \14753 , \14752 , \14698 );
or \U$13874 ( \14754 , \14751_nG6da , \14753 );
not \U$13875 ( \14755 , \14751_nG6da );
not \U$13876 ( \14756 , \14753 );
or \U$13877 ( \14757 , \14755 , \14756 );
buf \U$13878 ( \14758 , \11600 );
_DC g713 ( \14759_nG713 , \14758 , \14691 );
not \U$13879 ( \14760 , \14759_nG713 );
or \U$13880 ( \14761 , \14693 , RIaaa9218_606);
nand \U$13881 ( \14762 , \14761 , \14694 );
not \U$13882 ( \14763 , \14762 );
or \U$13883 ( \14764 , \14760 , \14763 );
or \U$13884 ( \14765 , \14762 , \14759_nG713 );
and \U$13885 ( \14766 , \8304 , RIaaa89a8_588);
nand \U$13886 ( \14767 , RIaaa91a0_605, \7609 );
not \U$13887 ( \14768 , \14767 );
nor \U$13888 ( \14769 , \14766 , \14768 );
buf \U$13889 ( \14770 , \11713 );
_DC g784 ( \14771_nG784 , \14770 , \14691 );
nand \U$13890 ( \14772 , \14771_nG784 , \8403 );
or \U$13891 ( \14773 , \14769 , \14772 );
not \U$13892 ( \14774 , \14772 );
not \U$13893 ( \14775 , \14769 );
or \U$13894 ( \14776 , \14774 , \14775 );
buf \U$13895 ( \14777 , \11685 );
_DC g768 ( \14778_nG768 , \14777 , \14691 );
nand \U$13896 ( \14779 , \14776 , \14778_nG768 );
nand \U$13897 ( \14780 , \14773 , \14779 );
buf \U$13898 ( \14781 , \11656 );
_DC g74b ( \14782_nG74b , \14781 , \14691 );
and \U$13899 ( \14783 , \14780 , \14782_nG74b );
and \U$13900 ( \14784 , \14767 , RIaaa9128_604);
nor \U$13901 ( \14785 , \14780 , \14782_nG74b );
nor \U$13902 ( \14786 , \14767 , RIaaa9128_604);
nor \U$13903 ( \14787 , \14784 , \14785 , \14786 );
nor \U$13904 ( \14788 , \14783 , \14787 );
and \U$13905 ( \14789 , \7875 , \7609 );
nor \U$13906 ( \14790 , \14789 , RIaaa90b0_603);
buf \U$13907 ( \14791 , \11628 );
_DC g72f ( \14792_nG72f , \14791 , \14691 );
nor \U$13908 ( \14793 , \14693 , \14790 , \14792_nG72f );
or \U$13909 ( \14794 , \14788 , \14793 );
or \U$13910 ( \14795 , \14693 , \14790 );
nand \U$13911 ( \14796 , \14795 , \14792_nG72f );
nand \U$13912 ( \14797 , \14794 , \14796 );
nand \U$13913 ( \14798 , \14765 , \14797 );
nand \U$13914 ( \14799 , \14764 , \14798 );
buf \U$13915 ( \14800 , \11571 );
_DC g6f6 ( \14801_nG6f6 , \14800 , \14691 );
or \U$13916 ( \14802 , \14799 , \14801_nG6f6 );
or \U$13917 ( \14803 , \14695 , RIaaa9290_607);
nand \U$13918 ( \14804 , \14803 , \14696 );
and \U$13919 ( \14805 , \14802 , \14804 );
and \U$13920 ( \14806 , \14801_nG6f6 , \14799 );
nor \U$13921 ( \14807 , \14805 , \14806 );
nand \U$13922 ( \14808 , \14757 , \14807 );
nand \U$13923 ( \14809 , \14749 , \14754 , \14808 );
nand \U$13924 ( \14810 , \14748 , \14809 );
or \U$13925 ( \14811 , \14738 , \14810 );
or \U$13926 ( \14812 , \14737_nG6a0 , \14735 );
nand \U$13927 ( \14813 , \14733 , \14811 , \14812 );
nand \U$13928 ( \14814 , \14732 , \14813 );
or \U$13929 ( \14815 , \14701 , RIaaa9470_611);
nand \U$13930 ( \14816 , \14815 , \14702 );
or \U$13931 ( \14817 , \14814 , \14816 );
buf \U$13932 ( \14818 , \11427 );
_DC g666 ( \14819_nG666 , \14818 , \14691 );
and \U$13933 ( \14820 , \14817 , \14819_nG666 );
and \U$13934 ( \14821 , \14816 , \14814 );
nor \U$13935 ( \14822 , \14722 , \14820 , \14821 );
nor \U$13936 ( \14823 , \14721 , \14822 );
nand \U$13937 ( \14824 , \14711 , \14823 );
nand \U$13938 ( \14825 , \14689 , \7938 , \14710 , \14824 );
nor \U$13939 ( \14826 , \14825 , \7937 );
_HMUX g3a8a_GF_PartitionCandidate ( \14827_nG3a8a , \11343 , \14564 , \14826 );
buf \U$13940 ( \14828 , \14827_nG3a8a );
xor \U$13941 ( \14829 , \8803 , \8804 );
xor \U$13942 ( \14830 , \14829 , \11336 );
xor \U$13943 ( \14831 , \12099 , \12100 );
xor \U$13944 ( \14832 , \14831 , \14557 );
_HMUX g3a4f_GF_PartitionCandidate ( \14833_nG3a4f , \14830 , \14832 , \14826 );
buf \U$13945 ( \14834 , \14833_nG3a4f );
xor \U$13946 ( \14835 , \8807 , \8972 );
xor \U$13947 ( \14836 , \14835 , \11333 );
xor \U$13948 ( \14837 , \12262 , \12264 );
xor \U$13949 ( \14838 , \14837 , \14554 );
_HMUX g3a1e_GF_PartitionCandidate ( \14839_nG3a1e , \14836 , \14838 , \14826 );
buf \U$13950 ( \14840 , \14839_nG3a1e );
xor \U$13951 ( \14841 , \8975 , \9080 );
xor \U$13952 ( \14842 , \14841 , \11330 );
xor \U$13953 ( \14843 , \12369 , \12371 );
xor \U$13954 ( \14844 , \14843 , \14551 );
_HMUX g39d7_GF_PartitionCandidate ( \14845_nG39d7 , \14842 , \14844 , \14826 );
buf \U$13955 ( \14846 , \14845_nG39d7 );
xor \U$13956 ( \14847 , \9083 , \9170 );
xor \U$13957 ( \14848 , \14847 , \11327 );
xor \U$13958 ( \14849 , \12457 , \12459 );
xor \U$13959 ( \14850 , \14849 , \14548 );
_HMUX g397e_GF_PartitionCandidate ( \14851_nG397e , \14848 , \14850 , \14826 );
buf \U$13960 ( \14852 , \14851_nG397e );
xor \U$13961 ( \14853 , \9283 , \9285 );
xor \U$13962 ( \14854 , \14853 , \11324 );
xor \U$13963 ( \14855 , \12462 , \12566 );
xor \U$13964 ( \14856 , \14855 , \14545 );
_HMUX g3917_GF_PartitionCandidate ( \14857_nG3917 , \14854 , \14856 , \14826 );
buf \U$13965 ( \14858 , \14857_nG3917 );
xor \U$13966 ( \14859 , \9290 , \9394 );
xor \U$13967 ( \14860 , \14859 , \11321 );
xor \U$13968 ( \14861 , \12571 , \12677 );
xor \U$13969 ( \14862 , \14861 , \14542 );
_HMUX g38a0_GF_PartitionCandidate ( \14863_nG38a0 , \14860 , \14862 , \14826 );
buf \U$13970 ( \14864 , \14863_nG38a0 );
xor \U$13971 ( \14865 , \9397 , \9528 );
xor \U$13972 ( \14866 , \14865 , \11318 );
xor \U$13973 ( \14867 , \12680 , \12807 );
xor \U$13974 ( \14868 , \14867 , \14539 );
_HMUX g3823_GF_PartitionCandidate ( \14869_nG3823 , \14866 , \14868 , \14826 );
buf \U$13975 ( \14870 , \14869_nG3823 );
xor \U$13976 ( \14871 , \9536 , \9703 );
xor \U$13977 ( \14872 , \14871 , \11314 );
not \U$13978 ( \14873 , \14872 );
xor \U$13979 ( \14874 , \12810 , \12958 );
xor \U$13980 ( \14875 , \14874 , \14536 );
_HMUX g378d_GF_PartitionCandidate ( \14876_nG378d , \14873 , \14875 , \14826 );
buf \U$13981 ( \14877 , \14876_nG378d );
xor \U$13982 ( \14878 , \9687 , \9692 );
xor \U$13983 ( \14879 , \14878 , \9700 );
xor \U$13984 ( \14880 , \9801 , \11309 );
xor \U$13985 ( \14881 , \14879 , \14880 );
not \U$13986 ( \14882 , \14881 );
xor \U$13987 ( \14883 , \12961 , \13063 );
xor \U$13988 ( \14884 , \14883 , \14533 );
_HMUX g36d5_GF_PartitionCandidate ( \14885_nG36d5 , \14882 , \14884 , \14826 );
buf \U$13989 ( \14886 , \14885_nG36d5 );
not \U$13990 ( \14887 , \11308 );
nand \U$13991 ( \14888 , \14887 , \11306 );
not \U$13992 ( \14889 , \14888 );
not \U$13993 ( \14890 , \11301 );
or \U$13994 ( \14891 , \14889 , \14890 );
or \U$13995 ( \14892 , \11301 , \14888 );
nand \U$13996 ( \14893 , \14891 , \14892 );
xor \U$13997 ( \14894 , \13238 , \13240 );
xor \U$13998 ( \14895 , \14894 , \14530 );
_HMUX g3621_GF_PartitionCandidate ( \14896_nG3621 , \14893 , \14895 , \14826 );
buf \U$13999 ( \14897 , \14896_nG3621 );
xor \U$14000 ( \14898 , \10058 , \10075 );
xor \U$14001 ( \14899 , \14898 , \11298 );
xor \U$14002 ( \14900 , \13247 , \13331 );
xor \U$14003 ( \14901 , \14900 , \14527 );
_HMUX g3562_GF_PartitionCandidate ( \14902_nG3562 , \14899 , \14901 , \14826 );
buf \U$14004 ( \14903 , \14902_nG3562 );
xor \U$14005 ( \14904 , \10083 , \10277 );
xor \U$14006 ( \14905 , \14904 , \11294 );
not \U$14007 ( \14906 , \14905 );
xor \U$14008 ( \14907 , \13334 , \13511 );
xor \U$14009 ( \14908 , \14907 , \14524 );
_HMUX g347c_GF_PartitionCandidate ( \14909_nG347c , \14906 , \14908 , \14826 );
buf \U$14010 ( \14910 , \14909_nG347c );
not \U$14011 ( \14911 , \11293 );
nand \U$14012 ( \14912 , \14911 , \11291 );
not \U$14013 ( \14913 , \14912 );
not \U$14014 ( \14914 , \11284 );
or \U$14015 ( \14915 , \14913 , \14914 );
or \U$14016 ( \14916 , \11284 , \14912 );
nand \U$14017 ( \14917 , \14915 , \14916 );
xor \U$14018 ( \14918 , \13514 , \13597 );
xor \U$14019 ( \14919 , \14918 , \14521 );
_HMUX g33a1_GF_PartitionCandidate ( \14920_nG33a1 , \14917 , \14919 , \14826 );
buf \U$14020 ( \14921 , \14920_nG33a1 );
xor \U$14021 ( \14922 , \10367 , \10528 );
xor \U$14022 ( \14923 , \14922 , \11281 );
xor \U$14023 ( \14924 , \13600 , \13766 );
xor \U$14024 ( \14925 , \14924 , \14518 );
_HMUX g32a4_GF_PartitionCandidate ( \14926_nG32a4 , \14923 , \14925 , \14826 );
buf \U$14025 ( \14927 , \14926_nG32a4 );
xor \U$14026 ( \14928 , \10531 , \10536 );
xor \U$14027 ( \14929 , \14928 , \11278 );
xor \U$14028 ( \14930 , \13769 , \13779 );
xor \U$14029 ( \14931 , \14930 , \14515 );
_HMUX g3195_GF_PartitionCandidate ( \14932_nG3195 , \14929 , \14931 , \14826 );
buf \U$14030 ( \14933 , \14932_nG3195 );
xor \U$14031 ( \14934 , \10539 , \10619 );
xor \U$14032 ( \14935 , \14934 , \11275 );
xor \U$14033 ( \14936 , \13782 , \13864 );
xor \U$14034 ( \14937 , \14936 , \14511 );
not \U$14035 ( \14938 , \14937 );
_HMUX g3087_GF_PartitionCandidate ( \14939_nG3087 , \14935 , \14938 , \14826 );
buf \U$14036 ( \14940 , \14939_nG3087 );
xor \U$14037 ( \14941 , \10607 , \10612 );
xor \U$14038 ( \14942 , \14941 , \10615 );
xor \U$14039 ( \14943 , \10690 , \11269 );
xor \U$14040 ( \14944 , \14942 , \14943 );
not \U$14041 ( \14945 , \14944 );
xor \U$14042 ( \14946 , \13935 , \13939 );
xor \U$14043 ( \14947 , \14946 , \14508 );
not \U$14044 ( \14948 , \14947 );
_HMUX g2f81_GF_PartitionCandidate ( \14949_nG2f81 , \14945 , \14948 , \14826 );
buf \U$14045 ( \14950 , \14949_nG2f81 );
xor \U$14046 ( \14951 , \10682 , \10684 );
xor \U$14047 ( \14952 , \14951 , \10687 );
xor \U$14048 ( \14953 , \10783 , \11264 );
xor \U$14049 ( \14954 , \14952 , \14953 );
not \U$14050 ( \14955 , \14954 );
xor \U$14051 ( \14956 , \13927 , \13929 );
xor \U$14052 ( \14957 , \14956 , \13932 );
xor \U$14053 ( \14958 , \14029 , \14503 );
xor \U$14054 ( \14959 , \14957 , \14958 );
not \U$14055 ( \14960 , \14959 );
_HMUX g2e5f_GF_PartitionCandidate ( \14961_nG2e5f , \14955 , \14960 , \14826 );
buf \U$14056 ( \14962 , \14961_nG2e5f );
not \U$14057 ( \14963 , \11254 );
not \U$14058 ( \14964 , \11263 );
nand \U$14059 ( \14965 , \14964 , \11261 );
not \U$14060 ( \14966 , \14965 );
or \U$14061 ( \14967 , \14963 , \14966 );
or \U$14062 ( \14968 , \14965 , \11254 );
nand \U$14063 ( \14969 , \14967 , \14968 );
not \U$14064 ( \14970 , \14502 );
nand \U$14065 ( \14971 , \14970 , \14500 );
not \U$14066 ( \14972 , \14971 );
not \U$14067 ( \14973 , \14493 );
or \U$14068 ( \14974 , \14972 , \14973 );
or \U$14069 ( \14975 , \14493 , \14971 );
nand \U$14070 ( \14976 , \14974 , \14975 );
_HMUX g2d75_GF_PartitionCandidate ( \14977_nG2d75 , \14969 , \14976 , \14826 );
buf \U$14071 ( \14978 , \14977_nG2d75 );
xor \U$14072 ( \14979 , \10849 , \10896 );
xor \U$14073 ( \14980 , \14979 , \11251 );
xor \U$14074 ( \14981 , \14095 , \14144 );
xor \U$14075 ( \14982 , \14981 , \14490 );
_HMUX g2c74_GF_PartitionCandidate ( \14983_nG2c74 , \14980 , \14982 , \14826 );
buf \U$14076 ( \14984 , \14983_nG2c74 );
xor \U$14077 ( \14985 , \10899 , \10969 );
xor \U$14078 ( \14986 , \14985 , \11248 );
xor \U$14079 ( \14987 , \14147 , \14220 );
xor \U$14080 ( \14988 , \14987 , \14487 );
_HMUX g2b81_GF_PartitionCandidate ( \14989_nG2b81 , \14986 , \14988 , \14826 );
buf \U$14081 ( \14990 , \14989_nG2b81 );
xor \U$14082 ( \14991 , \11241 , \11242 );
xor \U$14083 ( \14992 , \14991 , \11245 );
xor \U$14084 ( \14993 , \14480 , \14481 );
xor \U$14085 ( \14994 , \14993 , \14484 );
_HMUX g2a76_GF_PartitionCandidate ( \14995_nG2a76 , \14992 , \14994 , \14826 );
buf \U$14086 ( \14996 , \14995_nG2a76 );
xor \U$14087 ( \14997 , \10983 , \11032 );
xor \U$14088 ( \14998 , \14997 , \11238 );
xor \U$14089 ( \14999 , \14234 , \14275 );
xor \U$14090 ( \15000 , \14999 , \14477 );
_HMUX g2998_GF_PartitionCandidate ( \15001_nG2998 , \14998 , \15000 , \14826 );
buf \U$14091 ( \15002 , \15001_nG2998 );
xor \U$14092 ( \15003 , \11039 , \11083 );
xor \U$14093 ( \15004 , \15003 , \11235 );
xor \U$14094 ( \15005 , \14283 , \14327 );
xor \U$14095 ( \15006 , \15005 , \14474 );
_HMUX g2894_GF_PartitionCandidate ( \15007_nG2894 , \15004 , \15006 , \14826 );
buf \U$14096 ( \15008 , \15007_nG2894 );
xor \U$14097 ( \15009 , \11228 , \11229 );
xor \U$14098 ( \15010 , \15009 , \11232 );
xor \U$14099 ( \15011 , \14467 , \14468 );
xor \U$14100 ( \15012 , \15011 , \14471 );
_HMUX g27bf_GF_PartitionCandidate ( \15013_nG27bf , \15010 , \15012 , \14826 );
buf \U$14101 ( \15014 , \15013_nG27bf );
xor \U$14102 ( \15015 , \11098 , \11132 );
xor \U$14103 ( \15016 , \15015 , \11225 );
xor \U$14104 ( \15017 , \14339 , \14373 );
xor \U$14105 ( \15018 , \15017 , \14464 );
_HMUX g26e7_GF_PartitionCandidate ( \15019_nG26e7 , \15016 , \15018 , \14826 );
buf \U$14106 ( \15020 , \15019_nG26e7 );
endmodule

