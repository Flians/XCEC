//
// Conformal-LEC Version 20.10-d214 (03-Sep-2020)
//
module top(RI9148f90_243,RI91589e0_777,RI9158968_776,RI91588f0_775,RI9158878_774,RI9158800_773,RI9158788_772,RI9158710_771,RI9158698_770,
        RI9158620_769,RI9148810_227,RI9148090_211,RI9147910_195,RI9147190_179,RI9146a10_163,RI9146290_147,RI9145b10_131,RI9145390_115,RI9144c10_99,
        RI9144490_83,RI9143d10_67,RI9143590_51,RI90f3658_35,RI90f99b8_19,RI9138b68_3,RI91506a0_497,RI9158e18_786,RI9158da0_785,RI9158d28_784,
        RI9158cb0_783,RI9158c38_782,RI9158bc0_781,RI9158b48_780,RI9158ad0_779,RI9158a58_778,RI914ff20_481,RI914f7a0_465,RI914f020_449,RI914e8a0_433,
        RI914e120_417,RI914d9a0_401,RI914d220_385,RI914caa0_369,RI914c320_353,RI914bba0_337,RI914b420_321,RI914aca0_305,RI914a520_289,RI9149da0_273,
        RI9149620_257,RI9148f18_242,RI9148798_226,RI9148018_210,RI9147898_194,RI9147118_178,RI9146998_162,RI9146218_146,RI9145a98_130,RI9145318_114,
        RI9144b98_98,RI9144418_82,RI9143c98_66,RI9143518_50,RI90f36d0_34,RI912e758_18,RI9138be0_2,RI9150718_498,RI914ff98_482,RI914f818_466,
        RI914f098_450,RI914e918_434,RI914e198_418,RI914da18_402,RI914d298_386,RI914cb18_370,RI914c398_354,RI914bc18_338,RI914b498_322,RI914ad18_306,
        RI914a598_290,RI9149e18_274,RI9149698_258,RI9148ea0_241,RI9148720_225,RI9147fa0_209,RI9147820_193,RI91470a0_177,RI9146920_161,RI91461a0_145,
        RI9145a20_129,RI91452a0_113,RI9144b20_97,RI91443a0_81,RI9143c20_65,RI91434a0_49,RI90f3748_33,RI912e7d0_17,RI9138c58_1,RI9149008_244,
        RI9148888_228,RI9148108_212,RI9147988_196,RI9147208_180,RI9146a88_164,RI9146308_148,RI9145b88_132,RI9145408_116,RI9144c88_100,RI9144508_84,
        RI9143d88_68,RI9143608_52,RI90f35e0_36,RI90f9940_20,RI9138af0_4,RI9150790_499,RI9150010_483,RI914f890_467,RI914f110_451,RI914e990_435,
        RI914e210_419,RI914da90_403,RI914d310_387,RI914cb90_371,RI914c410_355,RI914bc90_339,RI914b510_323,RI914ad90_307,RI914a610_291,RI9149e90_275,
        RI9149710_259,RI91490f8_246,RI9148978_230,RI91481f8_214,RI9147a78_198,RI91472f8_182,RI9146b78_166,RI91463f8_150,RI9145c78_134,RI91454f8_118,
        RI9144d78_102,RI91445f8_86,RI9143e78_70,RI91436f8_54,RI90f34f0_38,RI90f9850_22,RI9138a00_6,RI9149080_245,RI9148900_229,RI9148180_213,
        RI9147a00_197,RI9147280_181,RI9146b00_165,RI9146380_149,RI9145c00_133,RI9145480_117,RI9144d00_101,RI9144580_85,RI9143e00_69,RI9143680_53,
        RI90f3568_37,RI90f98c8_21,RI9138a78_5,RI9150808_500,RI9150088_484,RI914f908_468,RI914f188_452,RI914ea08_436,RI914e288_420,RI914db08_404,
        RI914d388_388,RI914cc08_372,RI914c488_356,RI914bd08_340,RI914b588_324,RI914ae08_308,RI914a688_292,RI9149f08_276,RI9149788_260,RI9149170_247,
        RI91489f0_231,RI9148270_215,RI9147af0_199,RI9147370_183,RI9146bf0_167,RI9146470_151,RI9145cf0_135,RI9145570_119,RI9144df0_103,RI9144670_87,
        RI9143ef0_71,RI9143770_55,RI90f3478_39,RI90f97d8_23,RI9138988_7,RI9150880_501,RI9150100_485,RI914f980_469,RI914f200_453,RI914ea80_437,
        RI914e300_421,RI914db80_405,RI914d400_389,RI914cc80_373,RI914c500_357,RI914bd80_341,RI914b600_325,RI914ae80_309,RI914a700_293,RI9149f80_277,
        RI9149800_261,RI91508f8_502,RI9150178_486,RI914f9f8_470,RI914f278_454,RI914eaf8_438,RI914e378_422,RI914dbf8_406,RI914d478_390,RI914ccf8_374,
        RI914c578_358,RI914bdf8_342,RI914b678_326,RI914aef8_310,RI914a778_294,RI9149ff8_278,RI9149878_262,RI9150970_503,RI91501f0_487,RI914fa70_471,
        RI914f2f0_455,RI914eb70_439,RI914e3f0_423,RI914dc70_407,RI914d4f0_391,RI914cd70_375,RI914c5f0_359,RI914be70_343,RI914b6f0_327,RI914af70_311,
        RI914a7f0_295,RI914a070_279,RI91498f0_263,RI9149260_249,RI9148ae0_233,RI9148360_217,RI9147be0_201,RI9147460_185,RI9146ce0_169,RI9146560_153,
        RI9145de0_137,RI9145660_121,RI9144ee0_105,RI9144760_89,RI9143fe0_73,RI9143860_57,RI90f3388_41,RI90f96e8_25,RI9138898_9,RI91491e8_248,
        RI9148a68_232,RI91482e8_216,RI9147b68_200,RI91473e8_184,RI9146c68_168,RI91464e8_152,RI9145d68_136,RI91455e8_120,RI9144e68_104,RI91446e8_88,
        RI9143f68_72,RI91437e8_56,RI90f3400_40,RI90f9760_24,RI9138910_8,RI91509e8_504,RI9150268_488,RI914fae8_472,RI914f368_456,RI914ebe8_440,
        RI914e468_424,RI914dce8_408,RI914d568_392,RI914cde8_376,RI914c668_360,RI914bee8_344,RI914b768_328,RI914afe8_312,RI914a868_296,RI914a0e8_280,
        RI9149968_264,RI91492d8_250,RI9148b58_234,RI91483d8_218,RI9147c58_202,RI91474d8_186,RI9146d58_170,RI91465d8_154,RI9145e58_138,RI91456d8_122,
        RI9144f58_106,RI91447d8_90,RI9144058_74,RI91438d8_58,RI90f3310_42,RI90f9670_26,RI912eb18_10,RI9150a60_505,RI91502e0_489,RI914fb60_473,
        RI914f3e0_457,RI914ec60_441,RI914e4e0_425,RI914dd60_409,RI914d5e0_393,RI914ce60_377,RI914c6e0_361,RI914bf60_345,RI914b7e0_329,RI914b060_313,
        RI914a8e0_297,RI914a160_281,RI91499e0_265,RI91493c8_252,RI9148c48_236,RI91484c8_220,RI9147d48_204,RI91475c8_188,RI9146e48_172,RI91466c8_156,
        RI9145f48_140,RI91457c8_124,RI9145048_108,RI91448c8_92,RI9144148_76,RI91439c8_60,RI9143248_44,RI90f39a0_28,RI912ea28_12,RI9149350_251,
        RI9148bd0_235,RI9148450_219,RI9147cd0_203,RI9147550_187,RI9146dd0_171,RI9146650_155,RI9145ed0_139,RI9145750_123,RI9144fd0_107,RI9144850_91,
        RI91440d0_75,RI9143950_59,RI90f3298_43,RI90f95f8_27,RI912eaa0_11,RI9150ad8_506,RI9150358_490,RI914fbd8_474,RI914f458_458,RI914ecd8_442,
        RI914e558_426,RI914ddd8_410,RI914d658_394,RI914ced8_378,RI914c758_362,RI914bfd8_346,RI914b858_330,RI914b0d8_314,RI914a958_298,RI914a1d8_282,
        RI9149a58_266,RI9149440_253,RI9148cc0_237,RI9148540_221,RI9147dc0_205,RI9147640_189,RI9146ec0_173,RI9146740_157,RI9145fc0_141,RI9145840_125,
        RI91450c0_109,RI9144940_93,RI91441c0_77,RI9143a40_61,RI91432c0_45,RI90f3928_29,RI912e9b0_13,RI9150b50_507,RI91503d0_491,RI914fc50_475,
        RI914f4d0_459,RI914ed50_443,RI914e5d0_427,RI914de50_411,RI914d6d0_395,RI914cf50_379,RI914c7d0_363,RI914c050_347,RI914b8d0_331,RI914b150_315,
        RI914a9d0_299,RI914a250_283,RI9149ad0_267,RI9150bc8_508,RI9150448_492,RI914fcc8_476,RI914f548_460,RI914edc8_444,RI914e648_428,RI914dec8_412,
        RI914d748_396,RI914cfc8_380,RI914c848_364,RI914c0c8_348,RI914b948_332,RI914b1c8_316,RI914aa48_300,RI914a2c8_284,RI9149b48_268,RI9149530_255,
        RI9148db0_239,RI9148630_223,RI9147eb0_207,RI9147730_191,RI9146fb0_175,RI9146830_159,RI91460b0_143,RI9145930_127,RI91451b0_111,RI9144a30_95,
        RI91442b0_79,RI9143b30_63,RI91433b0_47,RI90f3838_31,RI912e8c0_15,RI91494b8_254,RI9148d38_238,RI91485b8_222,RI9147e38_206,RI91476b8_190,
        RI9146f38_174,RI91467b8_158,RI9146038_142,RI91458b8_126,RI9145138_110,RI91449b8_94,RI9144238_78,RI9143ab8_62,RI9143338_46,RI90f38b0_30,
        RI912e938_14,RI9150c40_509,RI91504c0_493,RI914fd40_477,RI914f5c0_461,RI914ee40_445,RI914e6c0_429,RI914df40_413,RI914d7c0_397,RI914d040_381,
        RI914c8c0_365,RI914c140_349,RI914b9c0_333,RI914b240_317,RI914aac0_301,RI914a340_285,RI9149bc0_269,RI91495a8_256,RI9148e28_240,RI91486a8_224,
        RI9147f28_208,RI91477a8_192,RI9147028_176,RI91468a8_160,RI9146128_144,RI91459a8_128,RI9145228_112,RI9144aa8_96,RI9144328_80,RI9143ba8_64,
        RI9143428_48,RI90f37c0_32,RI912e848_16,RI9150cb8_510,RI9150538_494,RI914fdb8_478,RI914f638_462,RI914eeb8_446,RI914e738_430,RI914dfb8_414,
        RI914d838_398,RI914d0b8_382,RI914c938_366,RI914c1b8_350,RI914ba38_334,RI914b2b8_318,RI914ab38_302,RI914a3b8_286,RI9149c38_270,RI9150d30_511,
        RI91505b0_495,RI914fe30_479,RI914f6b0_463,RI914ef30_447,RI914e7b0_431,RI914e030_415,RI914d8b0_399,RI914d130_383,RI914c9b0_367,RI914c230_351,
        RI914bab0_335,RI914b330_319,RI914abb0_303,RI914a430_287,RI9149cb0_271,RI9150da8_512,RI9150628_496,RI914fea8_480,RI914f728_464,RI914efa8_448,
        RI914e828_432,RI914e0a8_416,RI914d928_400,RI914d1a8_384,RI914ca28_368,RI914c2a8_352,RI914bb28_336,RI914b3a8_320,RI914ac28_304,RI914a4a8_288,
        RI9149d28_272,RI9157ea0_753,RI9157720_737,RI9156fa0_721,RI9156820_705,RI91560a0_689,RI9155920_673,RI91551a0_657,RI9154a20_641,RI91542a0_625,
        RI9153b20_609,RI91533a0_593,RI9152c20_577,RI91524a0_561,RI9151d20_545,RI91515a0_529,RI9150e20_513,RI9157f18_754,RI9157798_738,RI9157018_722,
        RI9156898_706,RI9156118_690,RI9155998_674,RI9155218_658,RI9154a98_642,RI9154318_626,RI9153b98_610,RI9153418_594,RI9152c98_578,RI9152518_562,
        RI9151d98_546,RI9151618_530,RI9150e98_514,RI9157f90_755,RI9157810_739,RI9157090_723,RI9156910_707,RI9156190_691,RI9155a10_675,RI9155290_659,
        RI9154b10_643,RI9154390_627,RI9153c10_611,RI9153490_595,RI9152d10_579,RI9152590_563,RI9151e10_547,RI9151690_531,RI9150f10_515,RI9158008_756,
        RI9157888_740,RI9157108_724,RI9156988_708,RI9156208_692,RI9155a88_676,RI9155308_660,RI9154b88_644,RI9154408_628,RI9153c88_612,RI9153508_596,
        RI9152d88_580,RI9152608_564,RI9151e88_548,RI9151708_532,RI9150f88_516,RI9158080_757,RI9157900_741,RI9157180_725,RI9156a00_709,RI9156280_693,
        RI9155b00_677,RI9155380_661,RI9154c00_645,RI9154480_629,RI9153d00_613,RI9153580_597,RI9152e00_581,RI9152680_565,RI9151f00_549,RI9151780_533,
        RI9151000_517,RI91580f8_758,RI9157978_742,RI91571f8_726,RI9156a78_710,RI91562f8_694,RI9155b78_678,RI91553f8_662,RI9154c78_646,RI91544f8_630,
        RI9153d78_614,RI91535f8_598,RI9152e78_582,RI91526f8_566,RI9151f78_550,RI91517f8_534,RI9151078_518,RI9158170_759,RI91579f0_743,RI9157270_727,
        RI9156af0_711,RI9156370_695,RI9155bf0_679,RI9155470_663,RI9154cf0_647,RI9154570_631,RI9153df0_615,RI9153670_599,RI9152ef0_583,RI9152770_567,
        RI9151ff0_551,RI9151870_535,RI91510f0_519,RI91581e8_760,RI9157a68_744,RI91572e8_728,RI9156b68_712,RI91563e8_696,RI9155c68_680,RI91554e8_664,
        RI9154d68_648,RI91545e8_632,RI9153e68_616,RI91536e8_600,RI9152f68_584,RI91527e8_568,RI9152068_552,RI91518e8_536,RI9151168_520,RI9158260_761,
        RI9157ae0_745,RI9157360_729,RI9156be0_713,RI9156460_697,RI9155ce0_681,RI9155560_665,RI9154de0_649,RI9154660_633,RI9153ee0_617,RI9153760_601,
        RI9152fe0_585,RI9152860_569,RI91520e0_553,RI9151960_537,RI91511e0_521,RI91582d8_762,RI9157b58_746,RI91573d8_730,RI9156c58_714,RI91564d8_698,
        RI9155d58_682,RI91555d8_666,RI9154e58_650,RI91546d8_634,RI9153f58_618,RI91537d8_602,RI9153058_586,RI91528d8_570,RI9152158_554,RI91519d8_538,
        RI9151258_522,RI9158350_763,RI9157bd0_747,RI9157450_731,RI9156cd0_715,RI9156550_699,RI9155dd0_683,RI9155650_667,RI9154ed0_651,RI9154750_635,
        RI9153fd0_619,RI9153850_603,RI91530d0_587,RI9152950_571,RI91521d0_555,RI9151a50_539,RI91512d0_523,RI91583c8_764,RI9157c48_748,RI91574c8_732,
        RI9156d48_716,RI91565c8_700,RI9155e48_684,RI91556c8_668,RI9154f48_652,RI91547c8_636,RI9154048_620,RI91538c8_604,RI9153148_588,RI91529c8_572,
        RI9152248_556,RI9151ac8_540,RI9151348_524,RI9158440_765,RI9157cc0_749,RI9157540_733,RI9156dc0_717,RI9156640_701,RI9155ec0_685,RI9155740_669,
        RI9154fc0_653,RI9154840_637,RI91540c0_621,RI9153940_605,RI91531c0_589,RI9152a40_573,RI91522c0_557,RI9151b40_541,RI91513c0_525,RI91584b8_766,
        RI9157d38_750,RI91575b8_734,RI9156e38_718,RI91566b8_702,RI9155f38_686,RI91557b8_670,RI9155038_654,RI91548b8_638,RI9154138_622,RI91539b8_606,
        RI9153238_590,RI9152ab8_574,RI9152338_558,RI9151bb8_542,RI9151438_526,RI9158530_767,RI9157db0_751,RI9157630_735,RI9156eb0_719,RI9156730_703,
        RI9155fb0_687,RI9155830_671,RI91550b0_655,RI9154930_639,RI91541b0_623,RI9153a30_607,RI91532b0_591,RI9152b30_575,RI91523b0_559,RI9151c30_543,
        RI91514b0_527,RI91585a8_768,RI9157e28_752,RI91576a8_736,RI9156f28_720,RI91567a8_704,RI9156028_688,RI91558a8_672,RI9155128_656,RI91549a8_640,
        RI9154228_624,RI9153aa8_608,RI9153328_592,RI9152ba8_576,RI9152428_560,RI9151ca8_544,RI9151528_528,R_313_9fdbc38,R_314_9fdbce0,R_315_9fdbd88,
        R_316_9fdbe30,R_317_9fdbed8,R_318_9fdbf80,R_319_9fdc028,R_31a_9fdc0d0,R_31b_9fdc178,R_31c_9fdc220,R_31d_9fdc2c8,R_31e_9fdc370,R_31f_9fdc418,
        R_320_9fdc4c0,R_321_9fdc568,R_322_9fdc610,R_323_9fdc6b8,R_324_9fdc760,R_325_9fdc808,R_326_9fdc8b0,R_327_9fdc958,R_328_9fdca00,R_329_9fdcaa8,
        R_32a_9fdcb50,R_32b_9fdcbf8,R_32c_9fdcca0,R_32d_9fdcd48);
input RI9148f90_243,RI91589e0_777,RI9158968_776,RI91588f0_775,RI9158878_774,RI9158800_773,RI9158788_772,RI9158710_771,RI9158698_770,
        RI9158620_769,RI9148810_227,RI9148090_211,RI9147910_195,RI9147190_179,RI9146a10_163,RI9146290_147,RI9145b10_131,RI9145390_115,RI9144c10_99,
        RI9144490_83,RI9143d10_67,RI9143590_51,RI90f3658_35,RI90f99b8_19,RI9138b68_3,RI91506a0_497,RI9158e18_786,RI9158da0_785,RI9158d28_784,
        RI9158cb0_783,RI9158c38_782,RI9158bc0_781,RI9158b48_780,RI9158ad0_779,RI9158a58_778,RI914ff20_481,RI914f7a0_465,RI914f020_449,RI914e8a0_433,
        RI914e120_417,RI914d9a0_401,RI914d220_385,RI914caa0_369,RI914c320_353,RI914bba0_337,RI914b420_321,RI914aca0_305,RI914a520_289,RI9149da0_273,
        RI9149620_257,RI9148f18_242,RI9148798_226,RI9148018_210,RI9147898_194,RI9147118_178,RI9146998_162,RI9146218_146,RI9145a98_130,RI9145318_114,
        RI9144b98_98,RI9144418_82,RI9143c98_66,RI9143518_50,RI90f36d0_34,RI912e758_18,RI9138be0_2,RI9150718_498,RI914ff98_482,RI914f818_466,
        RI914f098_450,RI914e918_434,RI914e198_418,RI914da18_402,RI914d298_386,RI914cb18_370,RI914c398_354,RI914bc18_338,RI914b498_322,RI914ad18_306,
        RI914a598_290,RI9149e18_274,RI9149698_258,RI9148ea0_241,RI9148720_225,RI9147fa0_209,RI9147820_193,RI91470a0_177,RI9146920_161,RI91461a0_145,
        RI9145a20_129,RI91452a0_113,RI9144b20_97,RI91443a0_81,RI9143c20_65,RI91434a0_49,RI90f3748_33,RI912e7d0_17,RI9138c58_1,RI9149008_244,
        RI9148888_228,RI9148108_212,RI9147988_196,RI9147208_180,RI9146a88_164,RI9146308_148,RI9145b88_132,RI9145408_116,RI9144c88_100,RI9144508_84,
        RI9143d88_68,RI9143608_52,RI90f35e0_36,RI90f9940_20,RI9138af0_4,RI9150790_499,RI9150010_483,RI914f890_467,RI914f110_451,RI914e990_435,
        RI914e210_419,RI914da90_403,RI914d310_387,RI914cb90_371,RI914c410_355,RI914bc90_339,RI914b510_323,RI914ad90_307,RI914a610_291,RI9149e90_275,
        RI9149710_259,RI91490f8_246,RI9148978_230,RI91481f8_214,RI9147a78_198,RI91472f8_182,RI9146b78_166,RI91463f8_150,RI9145c78_134,RI91454f8_118,
        RI9144d78_102,RI91445f8_86,RI9143e78_70,RI91436f8_54,RI90f34f0_38,RI90f9850_22,RI9138a00_6,RI9149080_245,RI9148900_229,RI9148180_213,
        RI9147a00_197,RI9147280_181,RI9146b00_165,RI9146380_149,RI9145c00_133,RI9145480_117,RI9144d00_101,RI9144580_85,RI9143e00_69,RI9143680_53,
        RI90f3568_37,RI90f98c8_21,RI9138a78_5,RI9150808_500,RI9150088_484,RI914f908_468,RI914f188_452,RI914ea08_436,RI914e288_420,RI914db08_404,
        RI914d388_388,RI914cc08_372,RI914c488_356,RI914bd08_340,RI914b588_324,RI914ae08_308,RI914a688_292,RI9149f08_276,RI9149788_260,RI9149170_247,
        RI91489f0_231,RI9148270_215,RI9147af0_199,RI9147370_183,RI9146bf0_167,RI9146470_151,RI9145cf0_135,RI9145570_119,RI9144df0_103,RI9144670_87,
        RI9143ef0_71,RI9143770_55,RI90f3478_39,RI90f97d8_23,RI9138988_7,RI9150880_501,RI9150100_485,RI914f980_469,RI914f200_453,RI914ea80_437,
        RI914e300_421,RI914db80_405,RI914d400_389,RI914cc80_373,RI914c500_357,RI914bd80_341,RI914b600_325,RI914ae80_309,RI914a700_293,RI9149f80_277,
        RI9149800_261,RI91508f8_502,RI9150178_486,RI914f9f8_470,RI914f278_454,RI914eaf8_438,RI914e378_422,RI914dbf8_406,RI914d478_390,RI914ccf8_374,
        RI914c578_358,RI914bdf8_342,RI914b678_326,RI914aef8_310,RI914a778_294,RI9149ff8_278,RI9149878_262,RI9150970_503,RI91501f0_487,RI914fa70_471,
        RI914f2f0_455,RI914eb70_439,RI914e3f0_423,RI914dc70_407,RI914d4f0_391,RI914cd70_375,RI914c5f0_359,RI914be70_343,RI914b6f0_327,RI914af70_311,
        RI914a7f0_295,RI914a070_279,RI91498f0_263,RI9149260_249,RI9148ae0_233,RI9148360_217,RI9147be0_201,RI9147460_185,RI9146ce0_169,RI9146560_153,
        RI9145de0_137,RI9145660_121,RI9144ee0_105,RI9144760_89,RI9143fe0_73,RI9143860_57,RI90f3388_41,RI90f96e8_25,RI9138898_9,RI91491e8_248,
        RI9148a68_232,RI91482e8_216,RI9147b68_200,RI91473e8_184,RI9146c68_168,RI91464e8_152,RI9145d68_136,RI91455e8_120,RI9144e68_104,RI91446e8_88,
        RI9143f68_72,RI91437e8_56,RI90f3400_40,RI90f9760_24,RI9138910_8,RI91509e8_504,RI9150268_488,RI914fae8_472,RI914f368_456,RI914ebe8_440,
        RI914e468_424,RI914dce8_408,RI914d568_392,RI914cde8_376,RI914c668_360,RI914bee8_344,RI914b768_328,RI914afe8_312,RI914a868_296,RI914a0e8_280,
        RI9149968_264,RI91492d8_250,RI9148b58_234,RI91483d8_218,RI9147c58_202,RI91474d8_186,RI9146d58_170,RI91465d8_154,RI9145e58_138,RI91456d8_122,
        RI9144f58_106,RI91447d8_90,RI9144058_74,RI91438d8_58,RI90f3310_42,RI90f9670_26,RI912eb18_10,RI9150a60_505,RI91502e0_489,RI914fb60_473,
        RI914f3e0_457,RI914ec60_441,RI914e4e0_425,RI914dd60_409,RI914d5e0_393,RI914ce60_377,RI914c6e0_361,RI914bf60_345,RI914b7e0_329,RI914b060_313,
        RI914a8e0_297,RI914a160_281,RI91499e0_265,RI91493c8_252,RI9148c48_236,RI91484c8_220,RI9147d48_204,RI91475c8_188,RI9146e48_172,RI91466c8_156,
        RI9145f48_140,RI91457c8_124,RI9145048_108,RI91448c8_92,RI9144148_76,RI91439c8_60,RI9143248_44,RI90f39a0_28,RI912ea28_12,RI9149350_251,
        RI9148bd0_235,RI9148450_219,RI9147cd0_203,RI9147550_187,RI9146dd0_171,RI9146650_155,RI9145ed0_139,RI9145750_123,RI9144fd0_107,RI9144850_91,
        RI91440d0_75,RI9143950_59,RI90f3298_43,RI90f95f8_27,RI912eaa0_11,RI9150ad8_506,RI9150358_490,RI914fbd8_474,RI914f458_458,RI914ecd8_442,
        RI914e558_426,RI914ddd8_410,RI914d658_394,RI914ced8_378,RI914c758_362,RI914bfd8_346,RI914b858_330,RI914b0d8_314,RI914a958_298,RI914a1d8_282,
        RI9149a58_266,RI9149440_253,RI9148cc0_237,RI9148540_221,RI9147dc0_205,RI9147640_189,RI9146ec0_173,RI9146740_157,RI9145fc0_141,RI9145840_125,
        RI91450c0_109,RI9144940_93,RI91441c0_77,RI9143a40_61,RI91432c0_45,RI90f3928_29,RI912e9b0_13,RI9150b50_507,RI91503d0_491,RI914fc50_475,
        RI914f4d0_459,RI914ed50_443,RI914e5d0_427,RI914de50_411,RI914d6d0_395,RI914cf50_379,RI914c7d0_363,RI914c050_347,RI914b8d0_331,RI914b150_315,
        RI914a9d0_299,RI914a250_283,RI9149ad0_267,RI9150bc8_508,RI9150448_492,RI914fcc8_476,RI914f548_460,RI914edc8_444,RI914e648_428,RI914dec8_412,
        RI914d748_396,RI914cfc8_380,RI914c848_364,RI914c0c8_348,RI914b948_332,RI914b1c8_316,RI914aa48_300,RI914a2c8_284,RI9149b48_268,RI9149530_255,
        RI9148db0_239,RI9148630_223,RI9147eb0_207,RI9147730_191,RI9146fb0_175,RI9146830_159,RI91460b0_143,RI9145930_127,RI91451b0_111,RI9144a30_95,
        RI91442b0_79,RI9143b30_63,RI91433b0_47,RI90f3838_31,RI912e8c0_15,RI91494b8_254,RI9148d38_238,RI91485b8_222,RI9147e38_206,RI91476b8_190,
        RI9146f38_174,RI91467b8_158,RI9146038_142,RI91458b8_126,RI9145138_110,RI91449b8_94,RI9144238_78,RI9143ab8_62,RI9143338_46,RI90f38b0_30,
        RI912e938_14,RI9150c40_509,RI91504c0_493,RI914fd40_477,RI914f5c0_461,RI914ee40_445,RI914e6c0_429,RI914df40_413,RI914d7c0_397,RI914d040_381,
        RI914c8c0_365,RI914c140_349,RI914b9c0_333,RI914b240_317,RI914aac0_301,RI914a340_285,RI9149bc0_269,RI91495a8_256,RI9148e28_240,RI91486a8_224,
        RI9147f28_208,RI91477a8_192,RI9147028_176,RI91468a8_160,RI9146128_144,RI91459a8_128,RI9145228_112,RI9144aa8_96,RI9144328_80,RI9143ba8_64,
        RI9143428_48,RI90f37c0_32,RI912e848_16,RI9150cb8_510,RI9150538_494,RI914fdb8_478,RI914f638_462,RI914eeb8_446,RI914e738_430,RI914dfb8_414,
        RI914d838_398,RI914d0b8_382,RI914c938_366,RI914c1b8_350,RI914ba38_334,RI914b2b8_318,RI914ab38_302,RI914a3b8_286,RI9149c38_270,RI9150d30_511,
        RI91505b0_495,RI914fe30_479,RI914f6b0_463,RI914ef30_447,RI914e7b0_431,RI914e030_415,RI914d8b0_399,RI914d130_383,RI914c9b0_367,RI914c230_351,
        RI914bab0_335,RI914b330_319,RI914abb0_303,RI914a430_287,RI9149cb0_271,RI9150da8_512,RI9150628_496,RI914fea8_480,RI914f728_464,RI914efa8_448,
        RI914e828_432,RI914e0a8_416,RI914d928_400,RI914d1a8_384,RI914ca28_368,RI914c2a8_352,RI914bb28_336,RI914b3a8_320,RI914ac28_304,RI914a4a8_288,
        RI9149d28_272,RI9157ea0_753,RI9157720_737,RI9156fa0_721,RI9156820_705,RI91560a0_689,RI9155920_673,RI91551a0_657,RI9154a20_641,RI91542a0_625,
        RI9153b20_609,RI91533a0_593,RI9152c20_577,RI91524a0_561,RI9151d20_545,RI91515a0_529,RI9150e20_513,RI9157f18_754,RI9157798_738,RI9157018_722,
        RI9156898_706,RI9156118_690,RI9155998_674,RI9155218_658,RI9154a98_642,RI9154318_626,RI9153b98_610,RI9153418_594,RI9152c98_578,RI9152518_562,
        RI9151d98_546,RI9151618_530,RI9150e98_514,RI9157f90_755,RI9157810_739,RI9157090_723,RI9156910_707,RI9156190_691,RI9155a10_675,RI9155290_659,
        RI9154b10_643,RI9154390_627,RI9153c10_611,RI9153490_595,RI9152d10_579,RI9152590_563,RI9151e10_547,RI9151690_531,RI9150f10_515,RI9158008_756,
        RI9157888_740,RI9157108_724,RI9156988_708,RI9156208_692,RI9155a88_676,RI9155308_660,RI9154b88_644,RI9154408_628,RI9153c88_612,RI9153508_596,
        RI9152d88_580,RI9152608_564,RI9151e88_548,RI9151708_532,RI9150f88_516,RI9158080_757,RI9157900_741,RI9157180_725,RI9156a00_709,RI9156280_693,
        RI9155b00_677,RI9155380_661,RI9154c00_645,RI9154480_629,RI9153d00_613,RI9153580_597,RI9152e00_581,RI9152680_565,RI9151f00_549,RI9151780_533,
        RI9151000_517,RI91580f8_758,RI9157978_742,RI91571f8_726,RI9156a78_710,RI91562f8_694,RI9155b78_678,RI91553f8_662,RI9154c78_646,RI91544f8_630,
        RI9153d78_614,RI91535f8_598,RI9152e78_582,RI91526f8_566,RI9151f78_550,RI91517f8_534,RI9151078_518,RI9158170_759,RI91579f0_743,RI9157270_727,
        RI9156af0_711,RI9156370_695,RI9155bf0_679,RI9155470_663,RI9154cf0_647,RI9154570_631,RI9153df0_615,RI9153670_599,RI9152ef0_583,RI9152770_567,
        RI9151ff0_551,RI9151870_535,RI91510f0_519,RI91581e8_760,RI9157a68_744,RI91572e8_728,RI9156b68_712,RI91563e8_696,RI9155c68_680,RI91554e8_664,
        RI9154d68_648,RI91545e8_632,RI9153e68_616,RI91536e8_600,RI9152f68_584,RI91527e8_568,RI9152068_552,RI91518e8_536,RI9151168_520,RI9158260_761,
        RI9157ae0_745,RI9157360_729,RI9156be0_713,RI9156460_697,RI9155ce0_681,RI9155560_665,RI9154de0_649,RI9154660_633,RI9153ee0_617,RI9153760_601,
        RI9152fe0_585,RI9152860_569,RI91520e0_553,RI9151960_537,RI91511e0_521,RI91582d8_762,RI9157b58_746,RI91573d8_730,RI9156c58_714,RI91564d8_698,
        RI9155d58_682,RI91555d8_666,RI9154e58_650,RI91546d8_634,RI9153f58_618,RI91537d8_602,RI9153058_586,RI91528d8_570,RI9152158_554,RI91519d8_538,
        RI9151258_522,RI9158350_763,RI9157bd0_747,RI9157450_731,RI9156cd0_715,RI9156550_699,RI9155dd0_683,RI9155650_667,RI9154ed0_651,RI9154750_635,
        RI9153fd0_619,RI9153850_603,RI91530d0_587,RI9152950_571,RI91521d0_555,RI9151a50_539,RI91512d0_523,RI91583c8_764,RI9157c48_748,RI91574c8_732,
        RI9156d48_716,RI91565c8_700,RI9155e48_684,RI91556c8_668,RI9154f48_652,RI91547c8_636,RI9154048_620,RI91538c8_604,RI9153148_588,RI91529c8_572,
        RI9152248_556,RI9151ac8_540,RI9151348_524,RI9158440_765,RI9157cc0_749,RI9157540_733,RI9156dc0_717,RI9156640_701,RI9155ec0_685,RI9155740_669,
        RI9154fc0_653,RI9154840_637,RI91540c0_621,RI9153940_605,RI91531c0_589,RI9152a40_573,RI91522c0_557,RI9151b40_541,RI91513c0_525,RI91584b8_766,
        RI9157d38_750,RI91575b8_734,RI9156e38_718,RI91566b8_702,RI9155f38_686,RI91557b8_670,RI9155038_654,RI91548b8_638,RI9154138_622,RI91539b8_606,
        RI9153238_590,RI9152ab8_574,RI9152338_558,RI9151bb8_542,RI9151438_526,RI9158530_767,RI9157db0_751,RI9157630_735,RI9156eb0_719,RI9156730_703,
        RI9155fb0_687,RI9155830_671,RI91550b0_655,RI9154930_639,RI91541b0_623,RI9153a30_607,RI91532b0_591,RI9152b30_575,RI91523b0_559,RI9151c30_543,
        RI91514b0_527,RI91585a8_768,RI9157e28_752,RI91576a8_736,RI9156f28_720,RI91567a8_704,RI9156028_688,RI91558a8_672,RI9155128_656,RI91549a8_640,
        RI9154228_624,RI9153aa8_608,RI9153328_592,RI9152ba8_576,RI9152428_560,RI9151ca8_544,RI9151528_528;
output R_313_9fdbc38,R_314_9fdbce0,R_315_9fdbd88,R_316_9fdbe30,R_317_9fdbed8,R_318_9fdbf80,R_319_9fdc028,R_31a_9fdc0d0,R_31b_9fdc178,
        R_31c_9fdc220,R_31d_9fdc2c8,R_31e_9fdc370,R_31f_9fdc418,R_320_9fdc4c0,R_321_9fdc568,R_322_9fdc610,R_323_9fdc6b8,R_324_9fdc760,R_325_9fdc808,
        R_326_9fdc8b0,R_327_9fdc958,R_328_9fdca00,R_329_9fdcaa8,R_32a_9fdcb50,R_32b_9fdcbf8,R_32c_9fdcca0,R_32d_9fdcd48;


wire \804 , \805 , \806_N$1 , \807_N$2 , \808_ZERO , \809_ONE , \810 , \811 , \812 ,
         \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 ,
         \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 ,
         \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 ,
         \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 ,
         \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 ,
         \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 ,
         \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 ,
         \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 ,
         \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 ,
         \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 ,
         \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 ,
         \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 ,
         \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 ,
         \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 ,
         \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 ,
         \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 ,
         \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 ,
         \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 ,
         \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 ,
         \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 ,
         \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 ,
         \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 ,
         \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 ,
         \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 ,
         \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 ,
         \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 ,
         \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 ,
         \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 ,
         \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 ,
         \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 ,
         \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 ,
         \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 ,
         \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 ,
         \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 ,
         \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 ,
         \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 ,
         \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 ,
         \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 ,
         \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 ,
         \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 ,
         \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 ,
         \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 ,
         \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 ,
         \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 ,
         \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 ,
         \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 ,
         \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 ,
         \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 ,
         \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 ,
         \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 ,
         \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 ,
         \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 ,
         \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 ,
         \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 ,
         \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 , \1362 ,
         \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 , \1372 ,
         \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 , \1382 ,
         \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 , \1392 ,
         \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 , \1402 ,
         \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 , \1411 , \1412 ,
         \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 , \1421 , \1422 ,
         \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 , \1431 , \1432 ,
         \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 , \1441 , \1442 ,
         \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 , \1451 , \1452 ,
         \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 , \1461 , \1462 ,
         \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 , \1471 , \1472 ,
         \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 , \1481 , \1482 ,
         \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 , \1491 , \1492 ,
         \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 , \1501 , \1502 ,
         \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 , \1511 , \1512 ,
         \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 , \1521 , \1522 ,
         \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 , \1531 , \1532 ,
         \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 , \1541 , \1542 ,
         \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 , \1551 , \1552 ,
         \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 , \1561 , \1562 ,
         \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 , \1571 , \1572 ,
         \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 , \1581 , \1582 ,
         \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 , \1591 , \1592 ,
         \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 , \1601 , \1602 ,
         \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 , \1611 , \1612 ,
         \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 , \1621 , \1622 ,
         \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 , \1631 , \1632 ,
         \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 , \1641 , \1642 ,
         \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 , \1651 , \1652 ,
         \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 , \1661 , \1662 ,
         \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 , \1671 , \1672 ,
         \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 , \1681 , \1682 ,
         \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 , \1691 , \1692 ,
         \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 , \1701 , \1702 ,
         \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 , \1711 , \1712 ,
         \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 , \1721 , \1722 ,
         \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 , \1731 , \1732 ,
         \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 , \1741 , \1742 ,
         \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 , \1751 , \1752 ,
         \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 , \1761 , \1762 ,
         \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 , \1771 , \1772 ,
         \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 , \1781 , \1782 ,
         \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 , \1791 , \1792 ,
         \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 , \1801 , \1802 ,
         \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 , \1811 , \1812 ,
         \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 , \1821 , \1822 ,
         \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 , \1831 , \1832 ,
         \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 , \1841 , \1842 ,
         \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 , \1851 , \1852 ,
         \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 , \1861 , \1862 ,
         \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 , \1871 , \1872 ,
         \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 , \1881 , \1882 ,
         \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 , \1891 , \1892 ,
         \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 , \1901 , \1902 ,
         \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 , \1911 , \1912 ,
         \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 , \1921 , \1922 ,
         \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 , \1931 , \1932 ,
         \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 , \1941 , \1942 ,
         \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 , \1951 , \1952 ,
         \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 , \1961 , \1962 ,
         \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 , \1971 , \1972 ,
         \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 , \1981 , \1982 ,
         \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 , \1991 , \1992 ,
         \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 , \2001 , \2002 ,
         \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 , \2011 , \2012 ,
         \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 , \2021 , \2022 ,
         \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 , \2031 , \2032 ,
         \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 , \2041 , \2042 ,
         \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 , \2051 , \2052 ,
         \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 , \2061 , \2062 ,
         \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 , \2071 , \2072 ,
         \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 , \2081 , \2082 ,
         \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 , \2091 , \2092 ,
         \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 , \2101 , \2102 ,
         \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 , \2111 , \2112 ,
         \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 , \2121 , \2122 ,
         \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 , \2131 , \2132 ,
         \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 , \2141 , \2142 ,
         \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 , \2151 , \2152 ,
         \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 , \2161 , \2162 ,
         \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 , \2171 , \2172 ,
         \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 , \2181 , \2182 ,
         \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 , \2191 , \2192 ,
         \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 , \2201 , \2202 ,
         \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 , \2211 , \2212 ,
         \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 , \2221 , \2222 ,
         \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 , \2231 , \2232 ,
         \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 , \2241 , \2242 ,
         \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 , \2251 , \2252 ,
         \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 , \2261 , \2262 ,
         \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 , \2271 , \2272 ,
         \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 , \2281 , \2282 ,
         \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 , \2291 , \2292 ,
         \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 , \2301 , \2302 ,
         \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 , \2311 , \2312 ,
         \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 , \2321 , \2322 ,
         \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 , \2331 , \2332 ,
         \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 , \2341 , \2342 ,
         \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 , \2351 , \2352 ,
         \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 , \2361 , \2362 ,
         \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 , \2371 , \2372 ,
         \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 , \2381 , \2382 ,
         \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 , \2391 , \2392 ,
         \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 , \2401 , \2402 ,
         \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 , \2411 , \2412 ,
         \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 , \2421 , \2422 ,
         \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 , \2431 , \2432 ,
         \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 , \2441 , \2442 ,
         \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 , \2451 , \2452 ,
         \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 , \2461 , \2462 ,
         \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 , \2471 , \2472 ,
         \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 , \2481 , \2482 ,
         \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 , \2491 , \2492 ,
         \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 , \2501 , \2502 ,
         \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 , \2511 , \2512 ,
         \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 , \2521 , \2522 ,
         \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 , \2531 , \2532 ,
         \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 , \2541 , \2542 ,
         \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 , \2551 , \2552 ,
         \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 , \2561 , \2562 ,
         \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 , \2571 , \2572 ,
         \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 , \2581 , \2582 ,
         \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 , \2591 , \2592 ,
         \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 , \2601 , \2602 ,
         \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 , \2611 , \2612 ,
         \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 , \2621 , \2622 ,
         \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 , \2631 , \2632 ,
         \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 , \2641 , \2642 ,
         \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 , \2651 , \2652 ,
         \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 , \2661 , \2662 ,
         \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 , \2671 , \2672 ,
         \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 , \2681 , \2682 ,
         \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 , \2691 , \2692 ,
         \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 , \2701 , \2702 ,
         \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 , \2711 , \2712 ,
         \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 , \2721 , \2722 ,
         \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 , \2731 , \2732 ,
         \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 , \2741 , \2742 ,
         \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 , \2751 , \2752 ,
         \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 , \2761 , \2762 ,
         \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 , \2771 , \2772 ,
         \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 , \2781 , \2782 ,
         \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 , \2791 , \2792 ,
         \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 , \2801 , \2802 ,
         \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 , \2811 , \2812 ,
         \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 , \2821 , \2822 ,
         \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 , \2831 , \2832 ,
         \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 , \2841 , \2842 ,
         \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 , \2851 , \2852 ,
         \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 , \2861 , \2862 ,
         \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 , \2871 , \2872 ,
         \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 , \2881 , \2882 ,
         \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 , \2891 , \2892 ,
         \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 , \2901 , \2902 ,
         \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 , \2911 , \2912 ,
         \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 , \2921 , \2922 ,
         \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 , \2931 , \2932 ,
         \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 , \2941 , \2942 ,
         \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 , \2951 , \2952 ,
         \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 , \2961 , \2962 ,
         \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 , \2971 , \2972 ,
         \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 , \2981 , \2982 ,
         \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 , \2991 , \2992 ,
         \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 , \3001 , \3002 ,
         \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 , \3011 , \3012 ,
         \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 , \3021 , \3022 ,
         \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 , \3031 , \3032 ,
         \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 , \3041 , \3042 ,
         \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 , \3051 , \3052 ,
         \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 , \3061 , \3062 ,
         \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 , \3071 , \3072 ,
         \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 , \3081 , \3082 ,
         \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 , \3091 , \3092 ,
         \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 , \3101 , \3102 ,
         \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 , \3111 , \3112 ,
         \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 , \3121 , \3122 ,
         \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 , \3131 , \3132 ,
         \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 , \3141 , \3142 ,
         \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 , \3151 , \3152 ,
         \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 , \3161 , \3162 ,
         \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 , \3171 , \3172 ,
         \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 , \3181 , \3182 ,
         \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 , \3191 , \3192 ,
         \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 , \3201 , \3202 ,
         \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 , \3211 , \3212 ,
         \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 , \3221 , \3222 ,
         \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 , \3231 , \3232 ,
         \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 , \3241 , \3242 ,
         \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 , \3251 , \3252 ,
         \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 , \3261 , \3262 ,
         \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 , \3271 , \3272 ,
         \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 , \3281 , \3282 ,
         \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 , \3291 , \3292 ,
         \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 , \3301 , \3302 ,
         \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 , \3311 , \3312 ,
         \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 , \3321 , \3322 ,
         \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 , \3331 , \3332 ,
         \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 , \3341 , \3342 ,
         \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 , \3351 , \3352 ,
         \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 , \3361 , \3362 ,
         \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 , \3371 , \3372 ,
         \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 , \3381 , \3382 ,
         \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 , \3391 , \3392 ,
         \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 , \3401 , \3402 ,
         \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 , \3411 , \3412 ,
         \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 , \3421 , \3422 ,
         \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 , \3431 , \3432 ,
         \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 , \3441 , \3442 ,
         \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 , \3451 , \3452 ,
         \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 , \3461 , \3462 ,
         \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 , \3471 , \3472 ,
         \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 , \3481 , \3482 ,
         \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 , \3491 , \3492 ,
         \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 , \3501 , \3502 ,
         \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 , \3511 , \3512 ,
         \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 , \3521 , \3522 ,
         \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 , \3531 , \3532 ,
         \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 , \3541 , \3542 ,
         \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 , \3551 , \3552 ,
         \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 , \3561 , \3562 ,
         \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 , \3571 , \3572 ,
         \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 , \3581 , \3582 ,
         \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 , \3591 , \3592 ,
         \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 , \3601 , \3602 ,
         \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 , \3611 , \3612 ,
         \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 , \3621 , \3622 ,
         \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 , \3631 , \3632 ,
         \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 , \3641 , \3642 ,
         \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 , \3651 , \3652 ,
         \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 , \3661 , \3662 ,
         \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 , \3671 , \3672 ,
         \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 , \3681 , \3682 ,
         \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 , \3691 , \3692 ,
         \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 , \3701 , \3702 ,
         \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 , \3711 , \3712 ,
         \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 , \3721 , \3722 ,
         \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 , \3731 , \3732 ,
         \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 , \3741 , \3742 ,
         \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 , \3751 , \3752 ,
         \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 , \3761 , \3762 ,
         \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 , \3771 , \3772 ,
         \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 , \3781 , \3782 ,
         \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 , \3791 , \3792 ,
         \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 , \3801 , \3802 ,
         \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 , \3811 , \3812 ,
         \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 , \3821 , \3822 ,
         \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 , \3831 , \3832 ,
         \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 , \3841 , \3842 ,
         \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 , \3851 , \3852 ,
         \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 , \3861 , \3862 ,
         \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 , \3871 , \3872 ,
         \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 , \3881 , \3882 ,
         \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 , \3891 , \3892 ,
         \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 , \3901 , \3902 ,
         \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 , \3911 , \3912 ,
         \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 , \3921 , \3922 ,
         \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 , \3931 , \3932 ,
         \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 , \3941 , \3942 ,
         \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 , \3951 , \3952 ,
         \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 , \3961 , \3962 ,
         \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 , \3971 , \3972 ,
         \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 , \3981 , \3982 ,
         \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 , \3991 , \3992 ,
         \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 , \4001 , \4002 ,
         \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 , \4011 , \4012 ,
         \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 , \4021 , \4022 ,
         \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 , \4031 , \4032 ,
         \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 , \4041 , \4042 ,
         \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 , \4051 , \4052 ,
         \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 , \4061 , \4062 ,
         \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 , \4071 , \4072 ,
         \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 , \4081 , \4082 ,
         \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 , \4091 , \4092 ,
         \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 , \4101 , \4102 ,
         \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 , \4111 , \4112 ,
         \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 , \4121 , \4122 ,
         \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 , \4131 , \4132 ,
         \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 , \4141 , \4142 ,
         \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 , \4151 , \4152 ,
         \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 , \4161 , \4162 ,
         \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 , \4171 , \4172 ,
         \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 , \4181 , \4182 ,
         \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 , \4191 , \4192 ,
         \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 , \4201 , \4202 ,
         \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 , \4211 , \4212 ,
         \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 , \4221 , \4222 ,
         \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 , \4231 , \4232 ,
         \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 , \4241 , \4242 ,
         \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 , \4251 , \4252 ,
         \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 , \4261 , \4262 ,
         \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 , \4271 , \4272 ,
         \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 , \4281 , \4282 ,
         \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 , \4291 , \4292 ,
         \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 , \4301 , \4302 ,
         \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 , \4311 , \4312 ,
         \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 , \4321 , \4322 ,
         \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 , \4331 , \4332 ,
         \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 , \4341 , \4342 ,
         \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 , \4351 , \4352 ,
         \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 , \4361 , \4362 ,
         \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 , \4371 , \4372 ,
         \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 , \4381 , \4382 ,
         \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 , \4391 , \4392 ,
         \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 , \4401 , \4402 ,
         \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 , \4411 , \4412 ,
         \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 , \4421 , \4422 ,
         \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 , \4431 , \4432 ,
         \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 , \4441 , \4442 ,
         \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 , \4451 , \4452 ,
         \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 , \4461 , \4462 ,
         \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 , \4471 , \4472 ,
         \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 , \4481 , \4482 ,
         \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 , \4491 , \4492 ,
         \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 , \4501 , \4502 ,
         \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 , \4511 , \4512 ,
         \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 , \4521 , \4522 ,
         \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 , \4531 , \4532 ,
         \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 , \4541 , \4542 ,
         \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 , \4551 , \4552 ,
         \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 , \4561 , \4562 ,
         \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 , \4571 , \4572 ,
         \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 , \4581 , \4582 ,
         \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 , \4591 , \4592 ,
         \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 , \4601 , \4602 ,
         \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 , \4611 , \4612 ,
         \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 , \4621 , \4622 ,
         \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 , \4631 , \4632 ,
         \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 , \4641 , \4642 ,
         \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 , \4651 , \4652 ,
         \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 , \4661 , \4662 ,
         \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 , \4671 , \4672 ,
         \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 , \4681 , \4682 ,
         \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 , \4691 , \4692 ,
         \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 , \4701 , \4702 ,
         \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 , \4711 , \4712 ,
         \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 , \4721 , \4722 ,
         \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 , \4731 , \4732 ,
         \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 , \4741 , \4742 ,
         \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 , \4751 , \4752 ,
         \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 , \4761 , \4762 ,
         \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 , \4771 , \4772 ,
         \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 , \4781 , \4782 ,
         \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 , \4791 , \4792 ,
         \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 , \4801 , \4802 ,
         \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 , \4811 , \4812 ,
         \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 , \4821 , \4822 ,
         \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 , \4831 , \4832 ,
         \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 , \4841 , \4842 ,
         \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 , \4851 , \4852 ,
         \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 , \4861 , \4862 ,
         \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 , \4871 , \4872 ,
         \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 , \4881 , \4882 ,
         \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 , \4891 , \4892 ,
         \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 , \4901 , \4902 ,
         \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 , \4911 , \4912 ,
         \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 , \4921 , \4922 ,
         \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 , \4931 , \4932 ,
         \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 , \4941 , \4942 ,
         \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 , \4951 , \4952 ,
         \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 , \4961 , \4962 ,
         \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 , \4971 , \4972 ,
         \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 , \4981 , \4982 ,
         \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 , \4991 , \4992 ,
         \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 , \5001 , \5002 ,
         \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 , \5011 , \5012 ,
         \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 , \5021 , \5022 ,
         \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 , \5031 , \5032 ,
         \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 , \5041 , \5042 ,
         \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 , \5051 , \5052 ,
         \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 , \5061 , \5062 ,
         \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 , \5071 , \5072 ,
         \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 , \5081 , \5082 ,
         \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 , \5091 , \5092 ,
         \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 , \5101 , \5102 ,
         \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 , \5111 , \5112 ,
         \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 , \5121 , \5122 ,
         \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 , \5131 , \5132 ,
         \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 , \5141 , \5142 ,
         \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 , \5151 , \5152 ,
         \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 , \5161 , \5162 ,
         \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 , \5171 , \5172 ,
         \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 , \5181 , \5182 ,
         \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 , \5191 , \5192 ,
         \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 , \5201 , \5202 ,
         \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 , \5211 , \5212 ,
         \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 , \5221 , \5222 ,
         \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 , \5231 , \5232 ,
         \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 , \5241 , \5242 ,
         \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 , \5251 , \5252 ,
         \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 , \5261 , \5262 ,
         \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 , \5271 , \5272 ,
         \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 , \5281 , \5282 ,
         \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 , \5291 , \5292 ,
         \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 , \5301 , \5302 ,
         \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 , \5311 , \5312 ,
         \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 , \5321 , \5322 ,
         \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 , \5331 , \5332 ,
         \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 , \5341 , \5342 ,
         \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 , \5351 , \5352 ,
         \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 , \5361 , \5362 ,
         \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 , \5371 , \5372 ,
         \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 , \5381 , \5382 ,
         \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 , \5391 , \5392 ,
         \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 , \5401 , \5402 ,
         \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 , \5411 , \5412 ,
         \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 , \5421 , \5422 ,
         \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 , \5431 , \5432 ,
         \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 , \5441 , \5442 ,
         \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 , \5451 , \5452 ,
         \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 , \5461 , \5462 ,
         \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 , \5471 , \5472 ,
         \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 , \5481 , \5482 ,
         \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 , \5491 , \5492 ,
         \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 , \5501 , \5502 ,
         \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 , \5511 , \5512 ,
         \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 , \5521 , \5522 ,
         \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 , \5531 , \5532 ,
         \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 , \5541 , \5542 ,
         \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 , \5551 , \5552 ,
         \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 , \5561 , \5562 ,
         \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 , \5571 , \5572 ,
         \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 , \5581 , \5582 ,
         \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 , \5591 , \5592 ,
         \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 , \5601 , \5602 ,
         \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 , \5611 , \5612 ,
         \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 , \5621 , \5622 ,
         \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 , \5631 , \5632 ,
         \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 , \5641 , \5642 ,
         \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 , \5651 , \5652 ,
         \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 , \5661 , \5662 ,
         \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 , \5671 , \5672 ,
         \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 , \5681 , \5682 ,
         \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 , \5691 , \5692 ,
         \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 , \5701 , \5702 ,
         \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 , \5711 , \5712 ,
         \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 , \5721 , \5722 ,
         \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 , \5731 , \5732 ,
         \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 , \5741 , \5742 ,
         \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 , \5751 , \5752 ,
         \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 , \5761 , \5762 ,
         \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 , \5771 , \5772 ,
         \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 , \5781 , \5782 ,
         \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 , \5791 , \5792 ,
         \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 , \5801 , \5802 ,
         \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 , \5811 , \5812 ,
         \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 , \5821 , \5822 ,
         \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 , \5831 , \5832 ,
         \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 , \5841 , \5842 ,
         \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 , \5851 , \5852 ,
         \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 , \5861 , \5862 ,
         \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 , \5871 , \5872 ,
         \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 , \5881 , \5882 ,
         \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 , \5891 , \5892 ,
         \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 , \5901 , \5902 ,
         \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 , \5911 , \5912 ,
         \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 , \5921 , \5922 ,
         \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 , \5931 , \5932 ,
         \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 , \5941 , \5942 ,
         \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 , \5951 , \5952 ,
         \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 , \5961 , \5962 ,
         \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 , \5971 , \5972 ,
         \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 , \5981 , \5982 ,
         \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 , \5991 , \5992 ,
         \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 , \6001 , \6002 ,
         \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 , \6011 , \6012 ,
         \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 , \6021 , \6022 ,
         \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 , \6031 , \6032 ,
         \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 , \6041 , \6042 ,
         \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 , \6051 , \6052 ,
         \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 , \6061 , \6062 ,
         \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 , \6071 , \6072 ,
         \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 , \6081 , \6082 ,
         \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 , \6091 , \6092 ,
         \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 , \6101 , \6102 ,
         \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 , \6111 , \6112 ,
         \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 , \6121 , \6122 ,
         \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 , \6131 , \6132 ,
         \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 , \6141 , \6142 ,
         \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 , \6151 , \6152 ,
         \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 , \6161 , \6162 ,
         \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 , \6171 , \6172 ,
         \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 , \6181 , \6182 ,
         \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 , \6191 , \6192 ,
         \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 , \6201 , \6202 ,
         \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 , \6211 , \6212 ,
         \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 , \6221 , \6222 ,
         \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 , \6231 , \6232 ,
         \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 , \6241 , \6242 ,
         \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 , \6251 , \6252 ,
         \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 , \6261 , \6262 ,
         \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 , \6271 , \6272 ,
         \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 , \6281 , \6282 ,
         \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 , \6291 , \6292 ,
         \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 , \6301 , \6302 ,
         \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 , \6311 , \6312 ,
         \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 , \6321 , \6322 ,
         \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 , \6331 , \6332 ,
         \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 , \6341 , \6342 ,
         \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 , \6351 , \6352 ,
         \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 , \6361 , \6362 ,
         \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 , \6371 , \6372 ,
         \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 , \6381 , \6382 ,
         \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 , \6391 , \6392 ,
         \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 , \6401 , \6402 ,
         \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 , \6411 , \6412 ,
         \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 , \6421 , \6422 ,
         \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 , \6431 , \6432 ,
         \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 , \6441 , \6442 ,
         \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 , \6451 , \6452 ,
         \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 , \6461 , \6462 ,
         \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 , \6471 , \6472 ,
         \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 , \6481 , \6482 ,
         \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 , \6491 , \6492 ,
         \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 , \6501 , \6502 ,
         \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 , \6511 , \6512 ,
         \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 , \6521 , \6522 ,
         \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 , \6531 , \6532 ,
         \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 , \6541 , \6542 ,
         \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 , \6551 , \6552 ,
         \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 , \6561 , \6562 ,
         \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 , \6571 , \6572 ,
         \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 , \6581 , \6582 ,
         \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 , \6591 , \6592 ,
         \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 , \6601 , \6602 ,
         \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 , \6611 , \6612 ,
         \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 , \6621 , \6622 ,
         \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 , \6631 , \6632 ,
         \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 , \6641 , \6642 ,
         \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 , \6651 , \6652 ,
         \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 , \6661 , \6662 ,
         \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 , \6671 , \6672 ,
         \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 , \6681 , \6682 ,
         \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 , \6691 , \6692 ,
         \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 , \6701 , \6702 ,
         \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 , \6711 , \6712 ,
         \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 , \6721 , \6722 ,
         \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 , \6731 , \6732 ,
         \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 , \6741 , \6742 ,
         \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 , \6751 , \6752 ,
         \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 , \6761 , \6762 ,
         \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 , \6771 , \6772 ,
         \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 , \6781 , \6782 ,
         \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 , \6791 , \6792 ,
         \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 , \6801 , \6802 ,
         \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 , \6811 , \6812 ,
         \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 , \6821 , \6822 ,
         \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 , \6831 , \6832 ,
         \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 , \6841 , \6842 ,
         \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 , \6851 , \6852 ,
         \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 , \6861 , \6862 ,
         \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 , \6871 , \6872 ,
         \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 , \6881 , \6882 ,
         \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 , \6891 , \6892 ,
         \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 , \6901 , \6902 ,
         \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 , \6911 , \6912 ,
         \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 , \6921 , \6922 ,
         \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 , \6931 , \6932 ,
         \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 , \6941 , \6942 ,
         \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 , \6951 , \6952 ,
         \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 , \6961 , \6962 ,
         \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 , \6971 , \6972 ,
         \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 , \6981 , \6982 ,
         \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 , \6991 , \6992 ,
         \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 , \7001 , \7002 ,
         \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 , \7011 , \7012 ,
         \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 , \7021 , \7022 ,
         \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 , \7031 , \7032 ,
         \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 , \7041 , \7042 ,
         \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 , \7051 , \7052 ,
         \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 , \7061 , \7062 ,
         \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 , \7071 , \7072 ,
         \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 , \7081 , \7082 ,
         \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 , \7091 , \7092 ,
         \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 , \7101 , \7102 ,
         \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 , \7111 , \7112 ,
         \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 , \7121 , \7122 ,
         \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 , \7131 , \7132 ,
         \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 , \7141 , \7142 ,
         \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 , \7151 , \7152 ,
         \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 , \7161 , \7162 ,
         \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 , \7171 , \7172 ,
         \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 , \7181 , \7182 ,
         \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 , \7191 , \7192 ,
         \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 , \7201 , \7202 ,
         \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 , \7211 , \7212 ,
         \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 , \7221 , \7222 ,
         \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 , \7231 , \7232 ,
         \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 , \7241 , \7242 ,
         \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 , \7251 , \7252 ,
         \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 , \7261 , \7262 ,
         \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 , \7271 , \7272 ,
         \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 , \7281 , \7282 ,
         \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 , \7291 , \7292 ,
         \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 , \7301 , \7302 ,
         \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 , \7311 , \7312 ,
         \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 , \7321 , \7322 ,
         \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 , \7331 , \7332 ,
         \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 , \7341 , \7342 ,
         \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 , \7351 , \7352 ,
         \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 , \7361 , \7362 ,
         \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 , \7371 , \7372 ,
         \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 , \7381 , \7382 ,
         \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 , \7391 , \7392 ,
         \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 , \7401 , \7402 ,
         \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 , \7411 , \7412 ,
         \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 , \7421 , \7422 ,
         \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 , \7431 , \7432 ,
         \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 , \7441 , \7442 ,
         \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 , \7451 , \7452 ,
         \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 , \7461 , \7462 ,
         \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 , \7471 , \7472 ,
         \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 , \7481 , \7482 ,
         \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 , \7491 , \7492 ,
         \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 , \7501 , \7502 ,
         \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 , \7511 , \7512 ,
         \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 , \7521 , \7522 ,
         \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 , \7531 , \7532 ,
         \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 , \7541 , \7542 ,
         \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 , \7551 , \7552 ,
         \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 , \7561 , \7562 ,
         \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 , \7571 , \7572 ,
         \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 , \7581 , \7582 ,
         \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 , \7591 , \7592 ,
         \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 , \7601 , \7602 ,
         \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 , \7611 , \7612 ,
         \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 , \7621 , \7622 ,
         \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 , \7631 , \7632 ,
         \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 , \7641 , \7642 ,
         \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 , \7651 , \7652 ,
         \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 , \7661 , \7662 ,
         \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 , \7671 , \7672 ,
         \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 , \7681 , \7682 ,
         \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 , \7691 , \7692 ,
         \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 , \7701 , \7702 ,
         \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 , \7711 , \7712 ,
         \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 , \7721 , \7722 ,
         \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 , \7731 , \7732 ,
         \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 , \7741 , \7742 ,
         \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 , \7751 , \7752 ,
         \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 , \7761 , \7762 ,
         \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 , \7771 , \7772 ,
         \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 , \7781 , \7782 ,
         \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 , \7791 , \7792 ,
         \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 , \7801 , \7802 ,
         \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 , \7811 , \7812 ,
         \7813 , \7814 , \7815 , \7816 , \7817 , \7818 , \7819 , \7820 , \7821 , \7822 ,
         \7823 , \7824 , \7825 , \7826 , \7827 , \7828 , \7829 , \7830 , \7831 , \7832 ,
         \7833 , \7834 , \7835 , \7836 , \7837 , \7838 , \7839 , \7840 , \7841 , \7842 ,
         \7843 , \7844 , \7845 , \7846 , \7847 , \7848 , \7849 , \7850 , \7851 , \7852 ,
         \7853 , \7854 , \7855 , \7856 , \7857 , \7858 , \7859 , \7860 , \7861 , \7862 ,
         \7863 , \7864 , \7865 , \7866 , \7867 , \7868 , \7869 , \7870 , \7871 , \7872 ,
         \7873 , \7874 , \7875 , \7876 , \7877 , \7878 , \7879 , \7880 , \7881 , \7882 ,
         \7883 , \7884 , \7885 , \7886 , \7887 , \7888 , \7889 , \7890 , \7891 , \7892 ,
         \7893 , \7894 , \7895 , \7896 , \7897 , \7898 , \7899 , \7900 , \7901 , \7902 ,
         \7903 , \7904 , \7905 , \7906 , \7907 , \7908 , \7909 , \7910 , \7911 , \7912 ,
         \7913 , \7914 , \7915 , \7916 , \7917 , \7918 , \7919 , \7920 , \7921 , \7922 ,
         \7923 , \7924 , \7925 , \7926 , \7927 , \7928 , \7929 , \7930 , \7931 , \7932 ,
         \7933 , \7934 , \7935 , \7936 , \7937 , \7938 , \7939 , \7940 , \7941 , \7942 ,
         \7943 , \7944 , \7945 , \7946 , \7947 , \7948 , \7949 , \7950 , \7951 , \7952 ,
         \7953 , \7954 , \7955 , \7956 , \7957 , \7958 , \7959 , \7960 , \7961 , \7962 ,
         \7963 , \7964 , \7965 , \7966 , \7967 , \7968 , \7969 , \7970 , \7971 , \7972 ,
         \7973 , \7974 , \7975 , \7976 , \7977 , \7978 , \7979 , \7980 , \7981 , \7982 ,
         \7983 , \7984 , \7985 , \7986 , \7987 , \7988 , \7989 , \7990 , \7991 , \7992 ,
         \7993 , \7994 , \7995 , \7996 , \7997 , \7998 , \7999 , \8000 , \8001 , \8002 ,
         \8003 , \8004 , \8005 , \8006 , \8007 , \8008 , \8009 , \8010 , \8011 , \8012 ,
         \8013 , \8014 , \8015 , \8016 , \8017 , \8018 , \8019 , \8020 , \8021 , \8022 ,
         \8023 , \8024 , \8025 , \8026 , \8027 , \8028 , \8029 , \8030 , \8031 , \8032 ,
         \8033 , \8034 , \8035 , \8036 , \8037 , \8038 , \8039 , \8040 , \8041 , \8042 ,
         \8043 , \8044 , \8045 , \8046 , \8047 , \8048 , \8049 , \8050 , \8051 , \8052 ,
         \8053 , \8054 , \8055 , \8056 , \8057 , \8058 , \8059 , \8060 , \8061 , \8062 ,
         \8063 , \8064 , \8065 , \8066 , \8067 , \8068 , \8069 , \8070 , \8071 , \8072 ,
         \8073 , \8074 , \8075 , \8076 , \8077 , \8078 , \8079 , \8080 , \8081 , \8082 ,
         \8083 , \8084 , \8085 , \8086 , \8087 , \8088 , \8089 , \8090 , \8091 , \8092 ,
         \8093 , \8094 , \8095 , \8096 , \8097 , \8098 , \8099 , \8100 , \8101 , \8102 ,
         \8103 , \8104 , \8105 , \8106 , \8107 , \8108 , \8109 , \8110 , \8111 , \8112 ,
         \8113 , \8114 , \8115 , \8116 , \8117 , \8118 , \8119 , \8120 , \8121 , \8122 ,
         \8123 , \8124 , \8125 , \8126 , \8127 , \8128 , \8129 , \8130 , \8131 , \8132 ,
         \8133 , \8134 , \8135 , \8136 , \8137 , \8138 , \8139 , \8140 , \8141 , \8142 ,
         \8143 , \8144 , \8145 , \8146 , \8147 , \8148 , \8149 , \8150 , \8151 , \8152 ,
         \8153 , \8154 , \8155 , \8156 , \8157 , \8158 , \8159 , \8160 , \8161 , \8162 ,
         \8163 , \8164 , \8165 , \8166 , \8167 , \8168 , \8169 , \8170 , \8171 , \8172 ,
         \8173 , \8174 , \8175 , \8176 , \8177 , \8178 , \8179 , \8180 , \8181 , \8182 ,
         \8183 , \8184 , \8185 , \8186 , \8187 , \8188 , \8189 , \8190 , \8191 , \8192 ,
         \8193 , \8194 , \8195 , \8196 , \8197 , \8198 , \8199 , \8200 , \8201 , \8202 ,
         \8203 , \8204 , \8205 , \8206 , \8207 , \8208 , \8209 , \8210 , \8211 , \8212 ,
         \8213 , \8214 , \8215 , \8216 , \8217 , \8218 , \8219 , \8220 , \8221 , \8222 ,
         \8223 , \8224 , \8225 , \8226 , \8227 , \8228 , \8229 , \8230 , \8231 , \8232 ,
         \8233 , \8234 , \8235 , \8236 , \8237 , \8238 , \8239 , \8240 , \8241 , \8242 ,
         \8243 , \8244 , \8245 , \8246 , \8247 , \8248 , \8249 , \8250 , \8251 , \8252 ,
         \8253 , \8254 , \8255 , \8256 , \8257 , \8258 , \8259 , \8260 , \8261 , \8262 ,
         \8263 , \8264 , \8265 , \8266 , \8267 , \8268 , \8269 , \8270 , \8271 , \8272 ,
         \8273 , \8274 , \8275 , \8276 , \8277 , \8278 , \8279 , \8280 , \8281 , \8282 ,
         \8283 , \8284 , \8285 , \8286 , \8287 , \8288 , \8289 , \8290 , \8291 , \8292 ,
         \8293 , \8294 , \8295 , \8296 , \8297 , \8298 , \8299 , \8300 , \8301 , \8302 ,
         \8303 , \8304 , \8305 , \8306 , \8307 , \8308 , \8309 , \8310 , \8311 , \8312 ,
         \8313 , \8314 , \8315 , \8316 , \8317 , \8318 , \8319 , \8320 , \8321 , \8322 ,
         \8323 , \8324 , \8325 , \8326 , \8327 , \8328 , \8329 , \8330 , \8331 , \8332 ,
         \8333 , \8334 , \8335 , \8336 , \8337 , \8338 , \8339 , \8340 , \8341 , \8342 ,
         \8343 , \8344 , \8345 , \8346 , \8347 , \8348 , \8349 , \8350 , \8351 , \8352 ,
         \8353 , \8354 , \8355 , \8356 , \8357 , \8358 , \8359 , \8360 , \8361 , \8362 ,
         \8363 , \8364 , \8365 , \8366 , \8367 , \8368 , \8369 , \8370 , \8371 , \8372 ,
         \8373 , \8374 , \8375 , \8376 , \8377 , \8378 , \8379 , \8380 , \8381 , \8382 ,
         \8383 , \8384 , \8385 , \8386 , \8387 , \8388 , \8389 , \8390 , \8391 , \8392 ,
         \8393 , \8394 , \8395 , \8396 , \8397 , \8398 , \8399 , \8400 , \8401 , \8402 ,
         \8403 , \8404 , \8405 , \8406 , \8407 , \8408 , \8409 , \8410 , \8411 , \8412 ,
         \8413 , \8414 , \8415 , \8416 , \8417 , \8418 , \8419 , \8420 , \8421 , \8422 ,
         \8423 , \8424 , \8425 , \8426 , \8427 , \8428 , \8429 , \8430 , \8431 , \8432 ,
         \8433 , \8434 , \8435 , \8436 , \8437 , \8438 , \8439 , \8440 , \8441 , \8442 ,
         \8443 , \8444 , \8445 , \8446 , \8447 , \8448 , \8449 , \8450 , \8451 , \8452 ,
         \8453 , \8454 , \8455 , \8456 , \8457 , \8458 , \8459 , \8460 , \8461 , \8462 ,
         \8463 , \8464 , \8465 , \8466 , \8467 , \8468 , \8469 , \8470 , \8471 , \8472 ,
         \8473 , \8474 , \8475 , \8476 , \8477 , \8478 , \8479 , \8480 , \8481 , \8482 ,
         \8483 , \8484 , \8485 , \8486 , \8487 , \8488 , \8489 , \8490 , \8491 , \8492 ,
         \8493 , \8494 , \8495 , \8496 , \8497 , \8498 , \8499 , \8500 , \8501 , \8502 ,
         \8503 , \8504 , \8505 , \8506 , \8507 , \8508 , \8509 , \8510 , \8511 , \8512 ,
         \8513 , \8514 , \8515 , \8516 , \8517 , \8518 , \8519 , \8520 , \8521 , \8522 ,
         \8523 , \8524 , \8525 , \8526 , \8527 , \8528 , \8529 , \8530 , \8531 , \8532 ,
         \8533 , \8534 , \8535 , \8536 , \8537 , \8538 , \8539 , \8540 , \8541 , \8542 ,
         \8543 , \8544 , \8545 , \8546 , \8547 , \8548 , \8549 , \8550 , \8551 , \8552 ,
         \8553 , \8554 , \8555 , \8556 , \8557 , \8558 , \8559 , \8560 , \8561 , \8562 ,
         \8563 , \8564 , \8565 , \8566 , \8567 , \8568 , \8569 , \8570 , \8571 , \8572 ,
         \8573 , \8574 , \8575 , \8576 , \8577 , \8578 , \8579 , \8580 , \8581 , \8582 ,
         \8583 , \8584 , \8585 , \8586 , \8587 , \8588 , \8589 , \8590 , \8591 , \8592 ,
         \8593 , \8594 , \8595 , \8596 , \8597 , \8598 , \8599 , \8600 , \8601 , \8602 ,
         \8603 , \8604 , \8605 , \8606 , \8607 , \8608 , \8609 , \8610 , \8611 , \8612 ,
         \8613 , \8614 , \8615 , \8616 , \8617 , \8618 , \8619 , \8620 , \8621 , \8622 ,
         \8623 , \8624 , \8625 , \8626 , \8627 , \8628 , \8629 , \8630 , \8631 , \8632 ,
         \8633 , \8634 , \8635 , \8636 , \8637 , \8638 , \8639 , \8640 , \8641 , \8642 ,
         \8643 , \8644 , \8645 , \8646 , \8647 , \8648 , \8649 , \8650 , \8651 , \8652 ,
         \8653 , \8654 , \8655 , \8656 , \8657 , \8658 , \8659 , \8660 , \8661 , \8662 ,
         \8663 , \8664 , \8665 , \8666 , \8667 , \8668 , \8669 , \8670 , \8671 , \8672 ,
         \8673 , \8674 , \8675 , \8676 , \8677 , \8678 , \8679 , \8680 , \8681 , \8682 ,
         \8683 , \8684 , \8685 , \8686 , \8687 , \8688 , \8689 , \8690 , \8691 , \8692 ,
         \8693 , \8694 , \8695 , \8696 , \8697 , \8698 , \8699 , \8700 , \8701 , \8702 ,
         \8703 , \8704 , \8705 , \8706 , \8707 , \8708 , \8709 , \8710 , \8711 , \8712 ,
         \8713 , \8714 , \8715 , \8716 , \8717 , \8718 , \8719 , \8720 , \8721 , \8722 ,
         \8723 , \8724 , \8725 , \8726 , \8727 , \8728 , \8729 , \8730 , \8731 , \8732 ,
         \8733 , \8734 , \8735 , \8736 , \8737 , \8738 , \8739 , \8740 , \8741 , \8742 ,
         \8743 , \8744 , \8745 , \8746 , \8747 , \8748 , \8749 , \8750 , \8751 , \8752 ,
         \8753 , \8754 , \8755 , \8756 , \8757 , \8758 , \8759 , \8760 , \8761 , \8762 ,
         \8763 , \8764 , \8765 , \8766 , \8767 , \8768 , \8769 , \8770 , \8771 , \8772 ,
         \8773 , \8774 , \8775 , \8776 , \8777 , \8778 , \8779 , \8780 , \8781 , \8782 ,
         \8783 , \8784 , \8785 , \8786 , \8787 , \8788 , \8789 , \8790 , \8791 , \8792 ,
         \8793 , \8794 , \8795 , \8796 , \8797 , \8798 , \8799 , \8800 , \8801 , \8802 ,
         \8803 , \8804 , \8805 , \8806 , \8807 , \8808 , \8809 , \8810 , \8811 , \8812 ,
         \8813 , \8814 , \8815 , \8816 , \8817 , \8818 , \8819 , \8820 , \8821 , \8822 ,
         \8823 , \8824 , \8825 , \8826 , \8827 , \8828 , \8829 , \8830 , \8831 , \8832 ,
         \8833 , \8834 , \8835 , \8836 , \8837 , \8838 , \8839 , \8840 , \8841 , \8842 ,
         \8843 , \8844 , \8845 , \8846 , \8847 , \8848 , \8849 , \8850 , \8851 , \8852 ,
         \8853 , \8854 , \8855 , \8856 , \8857 , \8858 , \8859 , \8860 , \8861 , \8862 ,
         \8863 , \8864 , \8865 , \8866 , \8867 , \8868 , \8869 , \8870 , \8871 , \8872 ,
         \8873 , \8874 , \8875 , \8876 , \8877 , \8878 , \8879 , \8880 , \8881 , \8882 ,
         \8883 , \8884 , \8885 , \8886 , \8887 , \8888 , \8889 , \8890 , \8891 , \8892 ,
         \8893 , \8894 , \8895 , \8896 , \8897 , \8898 , \8899 , \8900 , \8901 , \8902 ,
         \8903 , \8904 , \8905 , \8906 , \8907 , \8908 , \8909 , \8910 , \8911 , \8912 ,
         \8913 , \8914 , \8915 , \8916 , \8917 , \8918 , \8919 , \8920 , \8921 , \8922 ,
         \8923 , \8924 , \8925 , \8926 , \8927 , \8928 , \8929 , \8930 , \8931 , \8932 ,
         \8933 , \8934 , \8935 , \8936 , \8937 , \8938 , \8939 , \8940 , \8941 , \8942 ,
         \8943 , \8944 , \8945 , \8946 , \8947 , \8948 , \8949 , \8950 , \8951 , \8952 ,
         \8953 , \8954 , \8955 , \8956 , \8957 , \8958 , \8959 , \8960 , \8961 , \8962 ,
         \8963 , \8964 , \8965 , \8966 , \8967 , \8968 , \8969 , \8970 , \8971 , \8972 ,
         \8973 , \8974 , \8975 , \8976 , \8977 , \8978 , \8979 , \8980 , \8981 , \8982 ,
         \8983 , \8984 , \8985 , \8986 , \8987 , \8988 , \8989 , \8990 , \8991 , \8992 ,
         \8993 , \8994 , \8995 , \8996 , \8997 , \8998 , \8999 , \9000 , \9001 , \9002 ,
         \9003 , \9004 , \9005 , \9006 , \9007 , \9008 , \9009 , \9010 , \9011 , \9012 ,
         \9013 , \9014 , \9015 , \9016 , \9017 , \9018 , \9019 , \9020 , \9021 , \9022 ,
         \9023 , \9024 , \9025 , \9026 , \9027 , \9028 , \9029 , \9030 , \9031 , \9032 ,
         \9033 , \9034 , \9035 , \9036 , \9037 , \9038 , \9039 , \9040 , \9041 , \9042 ,
         \9043 , \9044 , \9045 , \9046 , \9047 , \9048 , \9049 , \9050 , \9051 , \9052 ,
         \9053 , \9054 , \9055 , \9056 , \9057 , \9058 , \9059 , \9060 , \9061 , \9062 ,
         \9063 , \9064 , \9065 , \9066 , \9067 , \9068 , \9069 , \9070 , \9071 , \9072 ,
         \9073 , \9074 , \9075 , \9076 , \9077 , \9078 , \9079 , \9080 , \9081 , \9082 ,
         \9083 , \9084 , \9085 , \9086 , \9087 , \9088 , \9089 , \9090 , \9091 , \9092 ,
         \9093 , \9094 , \9095 , \9096 , \9097 , \9098 , \9099 , \9100 , \9101 , \9102 ,
         \9103 , \9104 , \9105 , \9106 , \9107 , \9108 , \9109 , \9110 , \9111 , \9112 ,
         \9113 , \9114 , \9115 , \9116 , \9117 , \9118 , \9119 , \9120 , \9121 , \9122 ,
         \9123 , \9124 , \9125 , \9126 , \9127 , \9128 , \9129 , \9130 , \9131 , \9132 ,
         \9133 , \9134 , \9135 , \9136 , \9137 , \9138 , \9139 , \9140 , \9141 , \9142 ,
         \9143 , \9144 , \9145 , \9146 , \9147 , \9148 , \9149 , \9150 , \9151 , \9152 ,
         \9153 , \9154 , \9155 , \9156 , \9157 , \9158 , \9159 , \9160 , \9161 , \9162 ,
         \9163 , \9164 , \9165 , \9166 , \9167 , \9168 , \9169 , \9170 , \9171 , \9172 ,
         \9173 , \9174 , \9175 , \9176 , \9177 , \9178 , \9179 , \9180 , \9181 , \9182 ,
         \9183 , \9184 , \9185 , \9186 , \9187 , \9188 , \9189 , \9190 , \9191 , \9192 ,
         \9193 , \9194 , \9195 , \9196 , \9197 , \9198 , \9199 , \9200 , \9201 , \9202 ,
         \9203 , \9204 , \9205 , \9206 , \9207 , \9208 , \9209 , \9210 , \9211 , \9212 ,
         \9213 , \9214 , \9215 , \9216 , \9217 , \9218 , \9219 , \9220 , \9221 , \9222 ,
         \9223 , \9224 , \9225 , \9226 , \9227 , \9228 , \9229 , \9230 , \9231 , \9232 ,
         \9233 , \9234 , \9235 , \9236 , \9237 , \9238 , \9239 , \9240 , \9241 , \9242 ,
         \9243 , \9244 , \9245 , \9246 , \9247 , \9248 , \9249 , \9250 , \9251 , \9252 ,
         \9253 , \9254 , \9255 , \9256 , \9257 , \9258 , \9259 , \9260 , \9261 , \9262 ,
         \9263 , \9264 , \9265 , \9266 , \9267 , \9268 , \9269 , \9270 , \9271 , \9272 ,
         \9273 , \9274 , \9275 , \9276 , \9277 , \9278 , \9279 , \9280 , \9281 , \9282 ,
         \9283 , \9284 , \9285 , \9286 , \9287 , \9288 , \9289 , \9290 , \9291 , \9292 ,
         \9293 , \9294 , \9295 , \9296 , \9297 , \9298 , \9299 , \9300 , \9301 , \9302 ,
         \9303 , \9304 , \9305 , \9306 , \9307 , \9308 , \9309 , \9310 , \9311 , \9312 ,
         \9313 , \9314 , \9315 , \9316 , \9317 , \9318 , \9319 , \9320 , \9321 , \9322 ,
         \9323 , \9324 , \9325 , \9326 , \9327 , \9328 , \9329 , \9330 , \9331 , \9332 ,
         \9333 , \9334 , \9335 , \9336 , \9337 , \9338 , \9339 , \9340 , \9341 , \9342 ,
         \9343 , \9344 , \9345 , \9346 , \9347 , \9348 , \9349 , \9350 , \9351 , \9352 ,
         \9353 , \9354 , \9355 , \9356 , \9357 , \9358 , \9359 , \9360 , \9361 , \9362 ,
         \9363 , \9364 , \9365 , \9366 , \9367 , \9368 , \9369 , \9370 , \9371 , \9372 ,
         \9373 , \9374 , \9375 , \9376 , \9377 , \9378 , \9379 , \9380 , \9381 , \9382 ,
         \9383 , \9384 , \9385 , \9386 , \9387 , \9388 , \9389 , \9390 , \9391 , \9392 ,
         \9393 , \9394 , \9395 , \9396 , \9397 , \9398 , \9399 , \9400 , \9401 , \9402 ,
         \9403 , \9404 , \9405 , \9406 , \9407 , \9408 , \9409 , \9410 , \9411 , \9412 ,
         \9413 , \9414 , \9415 , \9416 , \9417 , \9418 , \9419 , \9420 , \9421 , \9422 ,
         \9423 , \9424 , \9425 , \9426 , \9427 , \9428 , \9429 , \9430 , \9431 , \9432 ,
         \9433 , \9434 , \9435 , \9436 , \9437 , \9438 , \9439 , \9440 , \9441 , \9442 ,
         \9443 , \9444 , \9445 , \9446 , \9447 , \9448 , \9449 , \9450 , \9451 , \9452 ,
         \9453 , \9454 , \9455 , \9456 , \9457 , \9458 , \9459 , \9460 , \9461 , \9462 ,
         \9463 , \9464 , \9465 , \9466 , \9467 , \9468 , \9469 , \9470 , \9471 , \9472 ,
         \9473 , \9474 , \9475 , \9476 , \9477 , \9478 , \9479 , \9480 , \9481 , \9482 ,
         \9483 , \9484 , \9485 , \9486 , \9487 , \9488 , \9489 , \9490 , \9491 , \9492 ,
         \9493 , \9494 , \9495 , \9496 , \9497 , \9498 , \9499 , \9500 , \9501 , \9502 ,
         \9503 , \9504 , \9505 , \9506 , \9507 , \9508 , \9509 , \9510 , \9511 , \9512 ,
         \9513 , \9514 , \9515 , \9516 , \9517 , \9518 , \9519 , \9520 , \9521 , \9522 ,
         \9523 , \9524 , \9525 , \9526 , \9527 , \9528 , \9529 , \9530 , \9531 , \9532 ,
         \9533 , \9534 , \9535 , \9536 , \9537 , \9538 , \9539 , \9540 , \9541 , \9542 ,
         \9543 , \9544 , \9545 , \9546 , \9547 , \9548 , \9549 , \9550 , \9551 , \9552 ,
         \9553 , \9554 , \9555 , \9556 , \9557 , \9558 , \9559 , \9560 , \9561 , \9562 ,
         \9563 , \9564 , \9565 , \9566 , \9567 , \9568 , \9569 , \9570 , \9571 , \9572 ,
         \9573 , \9574 , \9575 , \9576 , \9577 , \9578 , \9579 , \9580 , \9581 , \9582 ,
         \9583 , \9584 , \9585 , \9586 , \9587 , \9588 , \9589 , \9590 , \9591 , \9592 ,
         \9593 , \9594 , \9595 , \9596 , \9597 , \9598 , \9599 , \9600 , \9601 , \9602 ,
         \9603 , \9604 , \9605 , \9606 , \9607 , \9608 , \9609 , \9610 , \9611 , \9612 ,
         \9613 , \9614 , \9615 , \9616 , \9617 , \9618 , \9619 , \9620 , \9621 , \9622 ,
         \9623 , \9624 , \9625 , \9626 , \9627 , \9628 , \9629 , \9630 , \9631 , \9632 ,
         \9633 , \9634 , \9635 , \9636 , \9637 , \9638 , \9639 , \9640 , \9641 , \9642 ,
         \9643 , \9644 , \9645 , \9646 , \9647 , \9648 , \9649 , \9650 , \9651 , \9652 ,
         \9653 , \9654 , \9655 , \9656 , \9657 , \9658 , \9659 , \9660 , \9661 , \9662 ,
         \9663 , \9664 , \9665 , \9666 , \9667 , \9668 , \9669 , \9670 , \9671 , \9672 ,
         \9673 , \9674 , \9675 , \9676 , \9677 , \9678 , \9679 , \9680 , \9681 , \9682 ,
         \9683 , \9684 , \9685 , \9686 , \9687 , \9688 , \9689 , \9690 , \9691 , \9692 ,
         \9693 , \9694 , \9695 , \9696 , \9697 , \9698 , \9699 , \9700 , \9701 , \9702 ,
         \9703 , \9704 , \9705 , \9706 , \9707 , \9708 , \9709 , \9710 , \9711 , \9712 ,
         \9713 , \9714 , \9715 , \9716 , \9717 , \9718 , \9719 , \9720 , \9721 , \9722 ,
         \9723 , \9724 , \9725 , \9726 , \9727 , \9728 , \9729 , \9730 , \9731 , \9732 ,
         \9733 , \9734 , \9735 , \9736 , \9737 , \9738 , \9739 , \9740 , \9741 , \9742 ,
         \9743 , \9744 , \9745 , \9746 , \9747 , \9748 , \9749 , \9750 , \9751 , \9752 ,
         \9753 , \9754 , \9755 , \9756 , \9757 , \9758 , \9759 , \9760 , \9761 , \9762 ,
         \9763 , \9764 , \9765 , \9766 , \9767 , \9768 , \9769 , \9770 , \9771 , \9772 ,
         \9773 , \9774 , \9775 , \9776 , \9777 , \9778 , \9779 , \9780 , \9781 , \9782 ,
         \9783 , \9784 , \9785 , \9786 , \9787 , \9788 , \9789 , \9790 , \9791 , \9792 ,
         \9793 , \9794 , \9795 , \9796 , \9797 , \9798 , \9799 , \9800 , \9801 , \9802 ,
         \9803 , \9804 , \9805 , \9806 , \9807 , \9808 , \9809 , \9810 , \9811 , \9812 ,
         \9813 , \9814 , \9815 , \9816 , \9817 , \9818 , \9819 , \9820 , \9821 , \9822 ,
         \9823 , \9824 , \9825 , \9826 , \9827 , \9828 , \9829 , \9830 , \9831 , \9832 ,
         \9833 , \9834 , \9835 , \9836 , \9837 , \9838 , \9839 , \9840 , \9841 , \9842 ,
         \9843 , \9844 , \9845 , \9846 , \9847 , \9848 , \9849 , \9850 , \9851 , \9852 ,
         \9853 , \9854 , \9855 , \9856 , \9857 , \9858 , \9859 , \9860 , \9861 , \9862 ,
         \9863 , \9864 , \9865 , \9866 , \9867 , \9868 , \9869 , \9870 , \9871 , \9872 ,
         \9873 , \9874 , \9875 , \9876 , \9877 , \9878 , \9879 , \9880 , \9881 , \9882 ,
         \9883 , \9884 , \9885 , \9886 , \9887 , \9888 , \9889 , \9890 , \9891 , \9892 ,
         \9893 , \9894 , \9895 , \9896 , \9897 , \9898 , \9899 , \9900 , \9901 , \9902 ,
         \9903 , \9904 , \9905 , \9906 , \9907 , \9908 , \9909 , \9910 , \9911 , \9912 ,
         \9913 , \9914 , \9915 , \9916 , \9917 , \9918 , \9919 , \9920 , \9921 , \9922 ,
         \9923 , \9924 , \9925 , \9926 , \9927 , \9928 , \9929 , \9930 , \9931 , \9932 ,
         \9933 , \9934 , \9935 , \9936 , \9937 , \9938 , \9939 , \9940 , \9941 , \9942 ,
         \9943 , \9944 , \9945 , \9946 , \9947 , \9948 , \9949 , \9950 , \9951 , \9952 ,
         \9953 , \9954 , \9955 , \9956 , \9957 , \9958 , \9959 , \9960 , \9961 , \9962 ,
         \9963 , \9964 , \9965 , \9966 , \9967 , \9968 , \9969 , \9970 , \9971 , \9972 ,
         \9973 , \9974 , \9975 , \9976 , \9977 , \9978 , \9979 , \9980 , \9981 , \9982 ,
         \9983 , \9984 , \9985 , \9986 , \9987 , \9988 , \9989 , \9990 , \9991 , \9992 ,
         \9993 , \9994 , \9995 , \9996 , \9997 , \9998 , \9999 , \10000 , \10001 , \10002 ,
         \10003 , \10004 , \10005 , \10006 , \10007 , \10008 , \10009 , \10010 , \10011 , \10012 ,
         \10013 , \10014 , \10015 , \10016 , \10017 , \10018 , \10019 , \10020 , \10021 , \10022 ,
         \10023 , \10024 , \10025 , \10026 , \10027 , \10028 , \10029 , \10030 , \10031 , \10032 ,
         \10033 , \10034 , \10035 , \10036 , \10037 , \10038 , \10039 , \10040 , \10041 , \10042 ,
         \10043 , \10044 , \10045 , \10046 , \10047 , \10048 , \10049 , \10050 , \10051 , \10052 ,
         \10053 , \10054 , \10055 , \10056 , \10057 , \10058 , \10059 , \10060 , \10061 , \10062 ,
         \10063 , \10064 , \10065 , \10066 , \10067 , \10068 , \10069 , \10070 , \10071 , \10072 ,
         \10073 , \10074 , \10075 , \10076 , \10077 , \10078 , \10079 , \10080 , \10081 , \10082 ,
         \10083 , \10084 , \10085 , \10086 , \10087 , \10088 , \10089 , \10090 , \10091 , \10092 ,
         \10093 , \10094 , \10095 , \10096 , \10097 , \10098 , \10099 , \10100 , \10101 , \10102 ,
         \10103 , \10104 , \10105 , \10106 , \10107 , \10108 , \10109 , \10110 , \10111 , \10112 ,
         \10113 , \10114 , \10115 , \10116 , \10117 , \10118 , \10119 , \10120 , \10121 , \10122 ,
         \10123 , \10124 , \10125 , \10126 , \10127 , \10128 , \10129 , \10130 , \10131 , \10132 ,
         \10133 , \10134 , \10135 , \10136 , \10137 , \10138 , \10139 , \10140 , \10141 , \10142 ,
         \10143 , \10144 , \10145 , \10146 , \10147 , \10148 , \10149 , \10150 , \10151 , \10152 ,
         \10153 , \10154 , \10155 , \10156 , \10157 , \10158 , \10159 , \10160 , \10161 , \10162 ,
         \10163 , \10164 , \10165 , \10166 , \10167 , \10168 , \10169 , \10170 , \10171 , \10172 ,
         \10173 , \10174 , \10175 , \10176 , \10177 , \10178 , \10179 , \10180 , \10181 , \10182 ,
         \10183 , \10184 , \10185 , \10186 , \10187 , \10188 , \10189 , \10190 , \10191 , \10192 ,
         \10193 , \10194 , \10195 , \10196 , \10197 , \10198 , \10199 , \10200 , \10201 , \10202 ,
         \10203 , \10204 , \10205 , \10206 , \10207 , \10208 , \10209 , \10210 , \10211 , \10212 ,
         \10213 , \10214 , \10215 , \10216 , \10217 , \10218 , \10219 , \10220 , \10221 , \10222 ,
         \10223 , \10224 , \10225 , \10226 , \10227 , \10228 , \10229 , \10230 , \10231 , \10232 ,
         \10233 , \10234 , \10235 , \10236 , \10237 , \10238 , \10239 , \10240 , \10241 , \10242 ,
         \10243 , \10244 , \10245 , \10246 , \10247 , \10248 , \10249 , \10250 , \10251 , \10252 ,
         \10253 , \10254 , \10255 , \10256 , \10257 , \10258 , \10259 , \10260 , \10261 , \10262 ,
         \10263 , \10264 , \10265 , \10266 , \10267 , \10268 , \10269 , \10270 , \10271 , \10272 ,
         \10273 , \10274 , \10275 , \10276 , \10277 , \10278 , \10279 , \10280 , \10281 , \10282 ,
         \10283 , \10284 , \10285 , \10286 , \10287 , \10288 , \10289 , \10290 , \10291 , \10292 ,
         \10293 , \10294 , \10295 , \10296 , \10297 , \10298 , \10299 , \10300 , \10301 , \10302 ,
         \10303 , \10304 , \10305 , \10306 , \10307 , \10308 , \10309 , \10310 , \10311 , \10312 ,
         \10313 , \10314 , \10315 , \10316 , \10317 , \10318 , \10319 , \10320 , \10321 , \10322 ,
         \10323 , \10324 , \10325 , \10326 , \10327 , \10328 , \10329 , \10330 , \10331 , \10332 ,
         \10333 , \10334 , \10335 , \10336 , \10337 , \10338 , \10339 , \10340 , \10341 , \10342 ,
         \10343 , \10344 , \10345 , \10346 , \10347 , \10348 , \10349 , \10350 , \10351 , \10352 ,
         \10353 , \10354 , \10355 , \10356 , \10357 , \10358 , \10359 , \10360 , \10361 , \10362 ,
         \10363 , \10364 , \10365 , \10366 , \10367 , \10368 , \10369 , \10370 , \10371 , \10372 ,
         \10373 , \10374 , \10375 , \10376 , \10377 , \10378 , \10379 , \10380 , \10381 , \10382 ,
         \10383 , \10384 , \10385 , \10386 , \10387 , \10388 , \10389 , \10390 , \10391 , \10392 ,
         \10393 , \10394 , \10395 , \10396 , \10397 , \10398 , \10399 , \10400 , \10401 , \10402 ,
         \10403 , \10404 , \10405 , \10406 , \10407 , \10408 , \10409 , \10410 , \10411 , \10412 ,
         \10413 , \10414 , \10415 , \10416 , \10417 , \10418 , \10419 , \10420 , \10421 , \10422 ,
         \10423 , \10424 , \10425 , \10426 , \10427 , \10428 , \10429 , \10430 , \10431 , \10432 ,
         \10433 , \10434 , \10435 , \10436 , \10437 , \10438 , \10439 , \10440 , \10441 , \10442 ,
         \10443 , \10444 , \10445 , \10446 , \10447 , \10448 , \10449 , \10450 , \10451 , \10452 ,
         \10453 , \10454 , \10455 , \10456 , \10457 , \10458 , \10459 , \10460 , \10461 , \10462 ,
         \10463 , \10464 , \10465 , \10466 , \10467 , \10468 , \10469 , \10470 , \10471 , \10472 ,
         \10473 , \10474 , \10475 , \10476 , \10477 , \10478 , \10479 , \10480 , \10481 , \10482 ,
         \10483 , \10484 , \10485 , \10486 , \10487 , \10488 , \10489 , \10490 , \10491 , \10492 ,
         \10493 , \10494 , \10495 , \10496 , \10497 , \10498 , \10499 , \10500 , \10501 , \10502 ,
         \10503 , \10504 , \10505 , \10506 , \10507 , \10508 , \10509 , \10510 , \10511 , \10512 ,
         \10513 , \10514 , \10515 , \10516 , \10517 , \10518 , \10519 , \10520 , \10521 , \10522 ,
         \10523 , \10524 , \10525 , \10526 , \10527 , \10528 , \10529 , \10530 , \10531 , \10532 ,
         \10533 , \10534 , \10535 , \10536 , \10537 , \10538 , \10539 , \10540 , \10541 , \10542 ,
         \10543 , \10544 , \10545 , \10546 , \10547 , \10548 , \10549 , \10550 , \10551 , \10552 ,
         \10553 , \10554 , \10555 , \10556 , \10557 , \10558 , \10559 , \10560 , \10561 , \10562 ,
         \10563 , \10564 , \10565 , \10566 , \10567 , \10568 , \10569 , \10570 , \10571 , \10572 ,
         \10573 , \10574 , \10575 , \10576 , \10577 , \10578 , \10579 , \10580 , \10581 , \10582 ,
         \10583 , \10584 , \10585 , \10586 , \10587 , \10588 , \10589 , \10590 , \10591 , \10592 ,
         \10593 , \10594 , \10595 , \10596 , \10597 , \10598 , \10599 , \10600 , \10601 , \10602 ,
         \10603 , \10604 , \10605 , \10606 , \10607 , \10608 , \10609 , \10610 , \10611 , \10612 ,
         \10613 , \10614 , \10615 , \10616 , \10617 , \10618 , \10619 , \10620 , \10621 , \10622 ,
         \10623 , \10624 , \10625 , \10626 , \10627 , \10628 , \10629 , \10630 , \10631 , \10632 ,
         \10633 , \10634 , \10635 , \10636 , \10637 , \10638 , \10639 , \10640 , \10641 , \10642 ,
         \10643 , \10644 , \10645 , \10646 , \10647 , \10648 , \10649 , \10650 , \10651 , \10652 ,
         \10653 , \10654 , \10655 , \10656 , \10657 , \10658 , \10659 , \10660 , \10661 , \10662 ,
         \10663 , \10664 , \10665 , \10666 , \10667 , \10668 , \10669 , \10670 , \10671 , \10672 ,
         \10673 , \10674 , \10675 , \10676 , \10677 , \10678 , \10679 , \10680 , \10681 , \10682 ,
         \10683 , \10684 , \10685 , \10686 , \10687 , \10688 , \10689 , \10690 , \10691 , \10692 ,
         \10693 , \10694 , \10695 , \10696 , \10697 , \10698 , \10699 , \10700 , \10701 , \10702 ,
         \10703 , \10704 , \10705 , \10706 , \10707 , \10708 , \10709 , \10710 , \10711 , \10712 ,
         \10713 , \10714 , \10715 , \10716 , \10717 , \10718 , \10719 , \10720 , \10721 , \10722 ,
         \10723 , \10724 , \10725 , \10726 , \10727 , \10728 , \10729 , \10730 , \10731 , \10732 ,
         \10733 , \10734 , \10735 , \10736 , \10737 , \10738 , \10739 , \10740 , \10741 , \10742 ,
         \10743 , \10744 , \10745 , \10746 , \10747 , \10748 , \10749 , \10750 , \10751 , \10752 ,
         \10753 , \10754 , \10755 , \10756 , \10757 , \10758 , \10759 , \10760 , \10761 , \10762 ,
         \10763 , \10764 , \10765 , \10766 , \10767 , \10768 , \10769 , \10770 , \10771 , \10772 ,
         \10773 , \10774 , \10775 , \10776 , \10777 , \10778 , \10779 , \10780 , \10781 , \10782 ,
         \10783 , \10784 , \10785 , \10786 , \10787 , \10788 , \10789 , \10790 , \10791 , \10792 ,
         \10793 , \10794 , \10795 , \10796 , \10797 , \10798 , \10799 , \10800 , \10801 , \10802 ,
         \10803 , \10804 , \10805 , \10806 , \10807 , \10808 , \10809 , \10810 , \10811 , \10812 ,
         \10813 , \10814 , \10815 , \10816 , \10817 , \10818 , \10819 , \10820 , \10821 , \10822 ,
         \10823 , \10824 , \10825 , \10826 , \10827 , \10828 , \10829 , \10830 , \10831 , \10832 ,
         \10833 , \10834 , \10835 , \10836 , \10837 , \10838 , \10839 , \10840 , \10841 , \10842 ,
         \10843 , \10844 , \10845 , \10846 , \10847 , \10848 , \10849 , \10850 , \10851 , \10852 ,
         \10853 , \10854 , \10855 , \10856 , \10857 , \10858 , \10859 , \10860 , \10861 , \10862 ,
         \10863 , \10864 , \10865 , \10866 , \10867 , \10868 , \10869 , \10870 , \10871 , \10872 ,
         \10873 , \10874 , \10875 , \10876 , \10877 , \10878 , \10879 , \10880 , \10881 , \10882 ,
         \10883 , \10884 , \10885 , \10886 , \10887 , \10888 , \10889 , \10890 , \10891 , \10892 ,
         \10893 , \10894 , \10895 , \10896 , \10897 , \10898 , \10899 , \10900 , \10901 , \10902 ,
         \10903 , \10904 , \10905 , \10906 , \10907 , \10908 , \10909 , \10910 , \10911 , \10912 ,
         \10913 , \10914 , \10915 , \10916 , \10917 , \10918 , \10919 , \10920 , \10921 , \10922 ,
         \10923 , \10924 , \10925 , \10926 , \10927 , \10928 , \10929 , \10930 , \10931 , \10932 ,
         \10933 , \10934 , \10935 , \10936 , \10937 , \10938 , \10939 , \10940 ;
buf \U$labajz1181 ( R_313_9fdbc38, \10262 );
buf \U$labajz1182 ( R_314_9fdbce0, \10292 );
buf \U$labajz1183 ( R_315_9fdbd88, \10334 );
buf \U$labajz1184 ( R_316_9fdbe30, \10361 );
buf \U$labajz1185 ( R_317_9fdbed8, \10388 );
buf \U$labajz1186 ( R_318_9fdbf80, \10466 );
buf \U$labajz1187 ( R_319_9fdc028, \10504 );
buf \U$labajz1188 ( R_31a_9fdc0d0, \10520 );
buf \U$labajz1189 ( R_31b_9fdc178, \10551 );
buf \U$labajz1190 ( R_31c_9fdc220, \10579 );
buf \U$labajz1191 ( R_31d_9fdc2c8, \10606 );
buf \U$labajz1192 ( R_31e_9fdc370, \10622 );
buf \U$labajz1193 ( R_31f_9fdc418, \10663 );
buf \U$labajz1194 ( R_320_9fdc4c0, \10680 );
buf \U$labajz1195 ( R_321_9fdc568, \10706 );
buf \U$labajz1196 ( R_322_9fdc610, \10713 );
buf \U$labajz1197 ( R_323_9fdc6b8, \10752 );
buf \U$labajz1198 ( R_324_9fdc760, \10768 );
buf \U$labajz1199 ( R_325_9fdc808, \10795 );
buf \U$labajz1200 ( R_326_9fdc8b0, \10811 );
buf \U$labajz1201 ( R_327_9fdc958, \10847 );
buf \U$labajz1202 ( R_328_9fdca00, \10863 );
buf \U$labajz1203 ( R_329_9fdcaa8, \10895 );
buf \U$labajz1204 ( R_32a_9fdcb50, \10911 );
buf \U$labajz1205 ( R_32b_9fdcbf8, \10915 );
buf \U$labajz1206 ( R_32c_9fdcca0, \10931 );
buf \U$labajz1207 ( R_32d_9fdcd48, \10940 );
not \U$1 ( \810 , RI9158cb0_783);
nor \U$2 ( \811 , RI9158d28_784, RI9158da0_785);
nand \U$3 ( \812 , \810 , \811 , RI9158e18_786);
not \U$4 ( \813 , \812 );
nand \U$5 ( \814 , \813 , RI9149e90_275);
nor \U$6 ( \815 , RI9158d28_784, RI9158da0_785);
nor \U$7 ( \816 , RI9158cb0_783, RI9158e18_786);
and \U$8 ( \817 , \815 , \816 );
buf \U$9 ( \818 , \817 );
nand \U$10 ( \819 , \818 , RI9149710_259);
and \U$11 ( \820 , \814 , \819 );
not \U$12 ( \821 , RI9158cb0_783);
not \U$13 ( \822 , RI9158e18_786);
not \U$14 ( \823 , RI9158d28_784);
nand \U$15 ( \824 , \821 , \822 , \823 , RI9158da0_785);
buf \U$16 ( \825 , \824 );
not \U$17 ( \826 , \825 );
nand \U$18 ( \827 , \826 , RI914a610_291);
not \U$19 ( \828 , RI9158cb0_783);
not \U$20 ( \829 , RI9158d28_784);
nand \U$21 ( \830 , \828 , \829 , RI9158e18_786, RI9158da0_785);
not \U$22 ( \831 , \830 );
nand \U$23 ( \832 , \831 , RI914ad90_307);
and \U$24 ( \833 , \827 , \832 );
not \U$25 ( \834 , RI9158cb0_783);
not \U$26 ( \835 , RI9158da0_785);
nand \U$27 ( \836 , \834 , \822 , \835 , RI9158d28_784);
not \U$28 ( \837 , \836 );
not \U$29 ( \838 , RI914b510_323);
not \U$30 ( \839 , \838 );
and \U$31 ( \840 , \837 , \839 );
not \U$32 ( \841 , RI914bc90_339);
not \U$33 ( \842 , RI9158cb0_783);
not \U$34 ( \843 , RI9158da0_785);
nand \U$35 ( \844 , \842 , \843 , RI9158e18_786, RI9158d28_784);
nor \U$36 ( \845 , \841 , \844 );
nor \U$37 ( \846 , \840 , \845 );
not \U$38 ( \847 , RI9158cb0_783);
not \U$39 ( \848 , RI9158e18_786);
nand \U$40 ( \849 , \847 , \848 , RI9158d28_784, RI9158da0_785);
buf \U$41 ( \850 , \849 );
not \U$42 ( \851 , \850 );
not \U$43 ( \852 , RI914c410_355);
not \U$44 ( \853 , \852 );
and \U$45 ( \854 , \851 , \853 );
not \U$46 ( \855 , RI914cb90_371);
not \U$47 ( \856 , RI9158cb0_783);
nand \U$48 ( \857 , \856 , RI9158da0_785, RI9158d28_784, RI9158e18_786);
nor \U$49 ( \858 , \855 , \857 );
nor \U$50 ( \859 , \854 , \858 );
nand \U$51 ( \860 , \820 , \833 , \846 , \859 );
not \U$52 ( \861 , RI9158d28_784);
not \U$53 ( \862 , RI9158da0_785);
nand \U$54 ( \863 , \861 , \862 , \822 , RI9158cb0_783);
buf \U$55 ( \864 , \863 );
not \U$56 ( \865 , \864 );
nand \U$57 ( \866 , \865 , RI914d310_387);
not \U$58 ( \867 , RI9158d28_784);
not \U$59 ( \868 , RI9158da0_785);
nand \U$60 ( \869 , \867 , \868 , RI9158cb0_783, RI9158e18_786);
not \U$61 ( \870 , \869 );
nand \U$62 ( \871 , \870 , RI914da90_403);
and \U$63 ( \872 , \866 , \871 );
not \U$64 ( \873 , RI9158d28_784);
not \U$65 ( \874 , RI9158e18_786);
nand \U$66 ( \875 , \873 , \874 , RI9158da0_785, RI9158cb0_783);
not \U$67 ( \876 , \875 );
not \U$68 ( \877 , RI914e210_419);
not \U$69 ( \878 , \877 );
and \U$70 ( \879 , \876 , \878 );
not \U$71 ( \880 , RI914e990_435);
not \U$72 ( \881 , RI9158d28_784);
nand \U$73 ( \882 , \881 , RI9158cb0_783, RI9158e18_786, RI9158da0_785);
not \U$74 ( \883 , \882 );
not \U$75 ( \884 , \883 );
nor \U$76 ( \885 , \880 , \884 );
nor \U$77 ( \886 , \879 , \885 );
not \U$78 ( \887 , RI9158da0_785);
and \U$79 ( \888 , \822 , \887 , RI9158d28_784, RI9158cb0_783);
not \U$80 ( \889 , \888 );
not \U$81 ( \890 , \889 );
not \U$82 ( \891 , RI914f110_451);
not \U$83 ( \892 , \891 );
and \U$84 ( \893 , \890 , \892 );
not \U$85 ( \894 , RI9158da0_785);
nand \U$86 ( \895 , \894 , RI9158cb0_783, RI9158e18_786, RI9158d28_784);
not \U$87 ( \896 , \895 );
and \U$88 ( \897 , \896 , RI914f890_467);
nor \U$89 ( \898 , \893 , \897 );
not \U$90 ( \899 , RI9158e18_786);
nand \U$91 ( \900 , \899 , RI9158d28_784, RI9158da0_785, RI9158cb0_783);
not \U$92 ( \901 , \900 );
and \U$93 ( \902 , \901 , RI9150010_483);
not \U$94 ( \903 , RI9150790_499);
nand \U$95 ( \904 , RI9158d28_784, RI9158da0_785, RI9158cb0_783, RI9158e18_786);
nor \U$96 ( \905 , \903 , \904 );
nor \U$97 ( \906 , \902 , \905 );
nand \U$98 ( \907 , \872 , \886 , \898 , \906 );
nor \U$99 ( \908 , \860 , \907 );
not \U$100 ( \909 , \908 );
buf \U$101 ( \910 , \909 );
buf \U$103 ( \911 , \910 );
buf \U$104 ( \912 , \911 );
not \U$105 ( \913 , \912 );
buf \U$106 ( \914 , \913 );
buf \U$107 ( \915 , \914 );
not \U$108 ( \916 , \915 );
not \U$109 ( \917 , RI9158968_776);
nor \U$110 ( \918 , \917 , RI91588f0_775);
nor \U$111 ( \919 , RI9158878_774, RI91589e0_777);
and \U$112 ( \920 , \918 , \919 );
buf \U$113 ( \921 , \920 );
not \U$114 ( \922 , \921 );
not \U$115 ( \923 , RI90f3568_37);
or \U$116 ( \924 , \922 , \923 );
not \U$117 ( \925 , RI9158878_774);
not \U$118 ( \926 , RI91588f0_775);
nand \U$119 ( \927 , \925 , \926 , RI91589e0_777, RI9158968_776);
not \U$120 ( \928 , \927 );
not \U$121 ( \929 , \928 );
not \U$122 ( \930 , RI9143680_53);
or \U$123 ( \931 , \929 , \930 );
nand \U$124 ( \932 , \924 , \931 );
not \U$125 ( \933 , RI9145480_117);
not \U$126 ( \934 , RI9158878_774);
and \U$127 ( \935 , \934 , RI91588f0_775, RI9158968_776, RI91589e0_777);
buf \U$128 ( \936 , \935 );
not \U$129 ( \937 , \936 );
or \U$130 ( \938 , \933 , \937 );
nand \U$131 ( \939 , RI91588f0_775, RI9158968_776);
not \U$132 ( \940 , \939 );
and \U$133 ( \941 , \919 , \940 );
not \U$134 ( \942 , \941 );
not \U$135 ( \943 , \942 );
nand \U$136 ( \944 , \943 , RI9144d00_101);
nand \U$137 ( \945 , \938 , \944 );
nor \U$138 ( \946 , \932 , \945 );
not \U$139 ( \947 , RI9143e00_69);
not \U$140 ( \948 , RI91588f0_775);
nor \U$141 ( \949 , \948 , RI9158968_776);
and \U$142 ( \950 , \949 , \919 );
buf \U$143 ( \951 , \950 );
not \U$144 ( \952 , \951 );
or \U$145 ( \953 , \947 , \952 );
not \U$146 ( \954 , RI9158878_774);
not \U$147 ( \955 , RI9158968_776);
nand \U$148 ( \956 , \954 , \955 , RI91589e0_777, RI91588f0_775);
buf \U$149 ( \957 , \956 );
not \U$150 ( \958 , RI9144580_85);
or \U$151 ( \959 , \957 , \958 );
nand \U$152 ( \960 , \953 , \959 );
not \U$153 ( \961 , RI90f98c8_21);
and \U$154 ( \962 , \934 , \917 , \948 , RI91589e0_777);
buf \U$155 ( \963 , \962 );
not \U$156 ( \964 , \963 );
or \U$157 ( \965 , \961 , \964 );
nor \U$158 ( \966 , RI91588f0_775, RI9158968_776);
and \U$159 ( \967 , \966 , \919 );
buf \U$160 ( \968 , \967 );
nand \U$161 ( \969 , \968 , RI9138a78_5);
nand \U$162 ( \970 , \965 , \969 );
nor \U$163 ( \971 , \960 , \970 );
not \U$164 ( \972 , RI9145c00_133);
not \U$165 ( \973 , RI91589e0_777);
not \U$166 ( \974 , RI91588f0_775);
nand \U$167 ( \975 , \973 , \974 , \917 , RI9158878_774);
buf \U$168 ( \976 , \975 );
not \U$169 ( \977 , \976 );
not \U$170 ( \978 , \977 );
or \U$171 ( \979 , \972 , \978 );
not \U$172 ( \980 , RI91588f0_775);
not \U$173 ( \981 , RI9158968_776);
nand \U$174 ( \982 , \980 , \981 , RI9158878_774, RI91589e0_777);
buf \U$175 ( \983 , \982 );
not \U$176 ( \984 , \983 );
nand \U$177 ( \985 , \984 , RI9146380_149);
nand \U$178 ( \986 , \979 , \985 );
not \U$179 ( \987 , RI91588f0_775);
not \U$180 ( \988 , RI91589e0_777);
nand \U$181 ( \989 , \987 , \988 , RI9158968_776, RI9158878_774);
not \U$182 ( \990 , RI9146b00_165);
or \U$183 ( \991 , \989 , \990 );
not \U$184 ( \992 , RI91588f0_775);
nand \U$185 ( \993 , \992 , RI9158878_774, RI91589e0_777, RI9158968_776);
buf \U$186 ( \994 , \993 );
not \U$187 ( \995 , RI9147280_181);
or \U$188 ( \996 , \994 , \995 );
nand \U$189 ( \997 , \991 , \996 );
nor \U$190 ( \998 , \986 , \997 );
not \U$191 ( \999 , RI9147a00_197);
not \U$192 ( \1000 , RI9158968_776);
not \U$193 ( \1001 , RI91589e0_777);
nand \U$194 ( \1002 , \1000 , \1001 , RI91588f0_775, RI9158878_774);
not \U$195 ( \1003 , \1002 );
not \U$196 ( \1004 , \1003 );
or \U$197 ( \1005 , \999 , \1004 );
not \U$198 ( \1006 , RI9158968_776);
nand \U$199 ( \1007 , \1006 , RI9158878_774, RI91589e0_777, RI91588f0_775);
not \U$200 ( \1008 , \1007 );
nand \U$201 ( \1009 , RI9148180_213, \1008 );
nand \U$202 ( \1010 , \1005 , \1009 );
not \U$203 ( \1011 , RI9148900_229);
not \U$204 ( \1012 , RI91589e0_777);
and \U$205 ( \1013 , \1012 , RI91588f0_775, RI9158968_776, RI9158878_774);
buf \U$206 ( \1014 , \1013 );
not \U$207 ( \1015 , \1014 );
or \U$208 ( \1016 , \1011 , \1015 );
and \U$209 ( \1017 , RI91588f0_775, RI9158968_776, RI9158878_774, RI91589e0_777);
nand \U$210 ( \1018 , \1017 , RI9149080_245);
nand \U$211 ( \1019 , \1016 , \1018 );
nor \U$212 ( \1020 , \1010 , \1019 );
nand \U$213 ( \1021 , \946 , \971 , \998 , \1020 );
buf \U$214 ( \1022 , \1021 );
not \U$215 ( \1023 , \1022 );
buf \U$216 ( \1024 , \1023 );
buf \U$217 ( \1025 , \1024 );
not \U$218 ( \1026 , \1025 );
buf \U$219 ( \1027 , \1026 );
buf \U$220 ( \1028 , \1027 );
not \U$221 ( \1029 , \1028 );
or \U$222 ( \1030 , \916 , \1029 );
buf \U$223 ( \1031 , \1024 );
buf \U$224 ( \1032 , \911 );
nand \U$225 ( \1033 , \1031 , \1032 );
buf \U$226 ( \1034 , \1033 );
buf \U$227 ( \1035 , \1034 );
nand \U$228 ( \1036 , \1030 , \1035 );
buf \U$229 ( \1037 , \1036 );
buf \U$230 ( \1038 , \1037 );
not \U$231 ( \1039 , \1038 );
not \U$232 ( \1040 , RI914bd80_341);
not \U$233 ( \1041 , RI9158cb0_783);
not \U$234 ( \1042 , RI9158da0_785);
nand \U$235 ( \1043 , \1041 , \1042 , RI9158e18_786, RI9158d28_784);
not \U$236 ( \1044 , \1043 );
not \U$237 ( \1045 , \1044 );
or \U$238 ( \1046 , \1040 , \1045 );
not \U$239 ( \1047 , \836 );
nand \U$240 ( \1048 , \1047 , RI914b600_325);
nand \U$241 ( \1049 , \1046 , \1048 );
not \U$242 ( \1050 , RI914ae80_309);
not \U$243 ( \1051 , \831 );
or \U$244 ( \1052 , \1050 , \1051 );
not \U$245 ( \1053 , \825 );
nand \U$246 ( \1054 , \1053 , RI914a700_293);
nand \U$247 ( \1055 , \1052 , \1054 );
nor \U$248 ( \1056 , \1049 , \1055 );
not \U$249 ( \1057 , RI914d400_389);
not \U$250 ( \1058 , \864 );
not \U$251 ( \1059 , \1058 );
or \U$252 ( \1060 , \1057 , \1059 );
buf \U$253 ( \1061 , \869 );
not \U$254 ( \1062 , \1061 );
nand \U$255 ( \1063 , \1062 , RI914db80_405);
nand \U$256 ( \1064 , \1060 , \1063 );
not \U$257 ( \1065 , RI914e300_421);
not \U$258 ( \1066 , RI9158d28_784);
not \U$259 ( \1067 , RI9158e18_786);
nand \U$260 ( \1068 , \1066 , \1067 , RI9158da0_785, RI9158cb0_783);
not \U$261 ( \1069 , \1068 );
not \U$262 ( \1070 , \1069 );
or \U$263 ( \1071 , \1065 , \1070 );
nand \U$264 ( \1072 , \883 , RI914ea80_437);
nand \U$265 ( \1073 , \1071 , \1072 );
nor \U$266 ( \1074 , \1064 , \1073 );
not \U$267 ( \1075 , RI914f200_453);
not \U$268 ( \1076 , RI9158da0_785);
and \U$269 ( \1077 , \822 , \1076 , RI9158d28_784, RI9158cb0_783);
not \U$270 ( \1078 , \1077 );
or \U$271 ( \1079 , \1075 , \1078 );
buf \U$272 ( \1080 , \896 );
nand \U$273 ( \1081 , \1080 , RI914f980_469);
nand \U$274 ( \1082 , \1079 , \1081 );
not \U$275 ( \1083 , RI9150100_485);
not \U$276 ( \1084 , \901 );
or \U$277 ( \1085 , \1083 , \1084 );
nand \U$278 ( \1086 , RI9158da0_785, RI9158d28_784, RI9158cb0_783, RI9158e18_786);
not \U$279 ( \1087 , \1086 );
nand \U$280 ( \1088 , \1087 , RI9150880_501);
nand \U$281 ( \1089 , \1085 , \1088 );
nor \U$282 ( \1090 , \1082 , \1089 );
not \U$283 ( \1091 , RI914cc80_373);
not \U$284 ( \1092 , RI9158cb0_783);
nand \U$285 ( \1093 , \1092 , RI9158da0_785, RI9158d28_784, RI9158e18_786);
not \U$286 ( \1094 , \1093 );
not \U$287 ( \1095 , \1094 );
or \U$288 ( \1096 , \1091 , \1095 );
not \U$289 ( \1097 , \850 );
nand \U$290 ( \1098 , \1097 , RI914c500_357);
nand \U$291 ( \1099 , \1096 , \1098 );
not \U$292 ( \1100 , RI9149f80_277);
not \U$293 ( \1101 , \813 );
or \U$294 ( \1102 , \1100 , \1101 );
nand \U$295 ( \1103 , \818 , RI9149800_261);
nand \U$296 ( \1104 , \1102 , \1103 );
nor \U$297 ( \1105 , \1099 , \1104 );
nand \U$298 ( \1106 , \1056 , \1074 , \1090 , \1105 );
buf \U$299 ( \1107 , \1106 );
buf \U$300 ( \1108 , \1107 );
not \U$301 ( \1109 , RI914e288_420);
nor \U$302 ( \1110 , \1109 , \1068 );
not \U$303 ( \1111 , RI914ea08_436);
not \U$304 ( \1112 , \883 );
nor \U$305 ( \1113 , \1111 , \1112 );
nor \U$306 ( \1114 , \1110 , \1113 );
not \U$307 ( \1115 , \825 );
not \U$308 ( \1116 , \1115 );
not \U$309 ( \1117 , \1116 );
not \U$310 ( \1118 , RI914a688_292);
not \U$311 ( \1119 , \1118 );
and \U$312 ( \1120 , \1117 , \1119 );
not \U$313 ( \1121 , RI914ae08_308);
not \U$314 ( \1122 , \831 );
nor \U$315 ( \1123 , \1121 , \1122 );
nor \U$316 ( \1124 , \1120 , \1123 );
and \U$317 ( \1125 , \813 , RI9149f08_276);
and \U$318 ( \1126 , RI9149788_260, \818 );
nor \U$319 ( \1127 , \1125 , \1126 );
not \U$320 ( \1128 , RI9158e18_786);
nand \U$321 ( \1129 , \1128 , RI9158d28_784, RI9158da0_785, RI9158cb0_783);
not \U$322 ( \1130 , \1129 );
not \U$323 ( \1131 , RI9150088_484);
not \U$324 ( \1132 , \1131 );
and \U$325 ( \1133 , \1130 , \1132 );
not \U$326 ( \1134 , RI9150808_500);
nor \U$327 ( \1135 , \1134 , \1086 );
nor \U$328 ( \1136 , \1133 , \1135 );
nand \U$329 ( \1137 , \1114 , \1124 , \1127 , \1136 );
not \U$330 ( \1138 , RI914f188_452);
not \U$331 ( \1139 , \1077 );
nor \U$332 ( \1140 , \1138 , \1139 );
not \U$333 ( \1141 , \895 );
and \U$334 ( \1142 , \1141 , RI914f908_468);
nor \U$335 ( \1143 , \1140 , \1142 );
not \U$336 ( \1144 , \836 );
and \U$337 ( \1145 , \1144 , RI914b588_324);
and \U$338 ( \1146 , \1044 , RI914bd08_340);
nor \U$339 ( \1147 , \1145 , \1146 );
not \U$340 ( \1148 , \864 );
not \U$341 ( \1149 , RI914d388_388);
not \U$342 ( \1150 , \1149 );
and \U$343 ( \1151 , \1148 , \1150 );
not \U$344 ( \1152 , RI914db08_404);
nor \U$345 ( \1153 , \1152 , \1061 );
nor \U$346 ( \1154 , \1151 , \1153 );
not \U$347 ( \1155 , \850 );
and \U$348 ( \1156 , \1155 , RI914c488_356);
not \U$349 ( \1157 , \857 );
and \U$350 ( \1158 , \1157 , RI914cc08_372);
nor \U$351 ( \1159 , \1156 , \1158 );
nand \U$352 ( \1160 , \1143 , \1147 , \1154 , \1159 );
nor \U$353 ( \1161 , \1137 , \1160 );
not \U$354 ( \1162 , \1161 );
buf \U$355 ( \1163 , \1162 );
not \U$356 ( \1164 , \1163 );
buf \U$357 ( \1165 , \1164 );
buf \U$358 ( \1166 , \1165 );
and \U$359 ( \1167 , \1108 , \1166 );
not \U$360 ( \1168 , \1108 );
buf \U$361 ( \1169 , \1162 );
and \U$362 ( \1170 , \1168 , \1169 );
nor \U$363 ( \1171 , \1167 , \1170 );
buf \U$364 ( \1172 , \1171 );
buf \U$365 ( \1173 , \1172 );
and \U$366 ( \1174 , \1162 , \909 );
not \U$367 ( \1175 , \1162 );
buf \U$368 ( \1176 , \909 );
not \U$369 ( \1177 , \1176 );
buf \U$370 ( \1178 , \1177 );
and \U$371 ( \1179 , \1175 , \1178 );
nor \U$372 ( \1180 , \1174 , \1179 );
buf \U$373 ( \1181 , \1180 );
nand \U$374 ( \1182 , \1173 , \1181 );
buf \U$375 ( \1183 , \1182 );
buf \U$376 ( \1184 , \1183 );
not \U$377 ( \1185 , \1184 );
buf \U$378 ( \1186 , \1185 );
buf \U$381 ( \1187 , \1186 );
buf \U$382 ( \1188 , \1187 );
not \U$383 ( \1189 , \1188 );
or \U$384 ( \1190 , \1039 , \1189 );
buf \U$385 ( \1191 , \1172 );
not \U$386 ( \1192 , \1191 );
buf \U$387 ( \1193 , \1192 );
buf \U$390 ( \1194 , \1193 );
buf \U$391 ( \1195 , \1194 );
not \U$392 ( \1196 , RI9147988_196);
not \U$393 ( \1197 , \1003 );
or \U$394 ( \1198 , \1196 , \1197 );
buf \U$395 ( \1199 , \1007 );
not \U$396 ( \1200 , \1199 );
nand \U$397 ( \1201 , \1200 , RI9148108_212);
nand \U$398 ( \1202 , \1198 , \1201 );
not \U$399 ( \1203 , RI9146a88_164);
and \U$400 ( \1204 , \948 , \1012 , RI9158968_776, RI9158878_774);
not \U$401 ( \1205 , \1204 );
not \U$402 ( \1206 , \1205 );
not \U$403 ( \1207 , \1206 );
or \U$404 ( \1208 , \1203 , \1207 );
not \U$405 ( \1209 , RI9158878_774);
nand \U$406 ( \1210 , RI91589e0_777, RI9158968_776);
nor \U$407 ( \1211 , \1209 , \1210 , RI91588f0_775);
not \U$408 ( \1212 , \1211 );
not \U$409 ( \1213 , \1212 );
nand \U$410 ( \1214 , \1213 , RI9147208_180);
nand \U$411 ( \1215 , \1208 , \1214 );
nor \U$412 ( \1216 , \1202 , \1215 );
not \U$413 ( \1217 , RI9144508_84);
not \U$414 ( \1218 , \956 );
not \U$415 ( \1219 , \1218 );
or \U$416 ( \1220 , \1217 , \1219 );
nand \U$417 ( \1221 , RI9143d88_68, \951 );
nand \U$418 ( \1222 , \1220 , \1221 );
not \U$419 ( \1223 , RI9145408_116);
not \U$420 ( \1224 , \936 );
or \U$421 ( \1225 , \1223 , \1224 );
not \U$422 ( \1226 , \942 );
nand \U$423 ( \1227 , \1226 , RI9144c88_100);
nand \U$424 ( \1228 , \1225 , \1227 );
nor \U$425 ( \1229 , \1222 , \1228 );
not \U$426 ( \1230 , RI9143608_52);
not \U$427 ( \1231 , \928 );
or \U$428 ( \1232 , \1230 , \1231 );
nand \U$429 ( \1233 , \921 , RI90f35e0_36);
nand \U$430 ( \1234 , \1232 , \1233 );
not \U$431 ( \1235 , RI90f9940_20);
not \U$432 ( \1236 , \963 );
or \U$433 ( \1237 , \1235 , \1236 );
nand \U$434 ( \1238 , RI9138af0_4, \968 );
nand \U$435 ( \1239 , \1237 , \1238 );
nor \U$436 ( \1240 , \1234 , \1239 );
not \U$437 ( \1241 , RI9145b88_132);
not \U$438 ( \1242 , \977 );
or \U$439 ( \1243 , \1241 , \1242 );
not \U$440 ( \1244 , \983 );
nand \U$441 ( \1245 , \1244 , RI9146308_148);
nand \U$442 ( \1246 , \1243 , \1245 );
not \U$443 ( \1247 , RI9148888_228);
not \U$444 ( \1248 , \1014 );
or \U$445 ( \1249 , \1247 , \1248 );
not \U$446 ( \1250 , \1017 );
not \U$447 ( \1251 , \1250 );
nand \U$448 ( \1252 , \1251 , RI9149008_244);
nand \U$449 ( \1253 , \1249 , \1252 );
nor \U$450 ( \1254 , \1246 , \1253 );
nand \U$451 ( \1255 , \1216 , \1229 , \1240 , \1254 );
buf \U$452 ( \1256 , \1255 );
not \U$453 ( \1257 , \1256 );
buf \U$454 ( \1258 , \1257 );
buf \U$455 ( \1259 , \1258 );
not \U$456 ( \1260 , \1259 );
buf \U$457 ( \1261 , \1260 );
buf \U$458 ( \1262 , \1261 );
not \U$459 ( \1263 , \1262 );
buf \U$460 ( \1264 , \914 );
not \U$461 ( \1265 , \1264 );
or \U$462 ( \1266 , \1263 , \1265 );
buf \U$463 ( \1267 , \911 );
buf \U$464 ( \1268 , \1258 );
nand \U$465 ( \1269 , \1267 , \1268 );
buf \U$466 ( \1270 , \1269 );
buf \U$467 ( \1271 , \1270 );
nand \U$468 ( \1272 , \1266 , \1271 );
buf \U$469 ( \1273 , \1272 );
buf \U$470 ( \1274 , \1273 );
nand \U$471 ( \1275 , \1195 , \1274 );
buf \U$472 ( \1276 , \1275 );
buf \U$473 ( \1277 , \1276 );
nand \U$474 ( \1278 , \1190 , \1277 );
buf \U$475 ( \1279 , \1278 );
buf \U$476 ( \1280 , \1279 );
not \U$477 ( \1281 , \1280 );
not \U$478 ( \1282 , \951 );
not \U$479 ( \1283 , RI9143d10_67);
or \U$480 ( \1284 , \1282 , \1283 );
not \U$481 ( \1285 , \1218 );
not \U$482 ( \1286 , RI9144490_83);
or \U$483 ( \1287 , \1285 , \1286 );
nand \U$484 ( \1288 , \1284 , \1287 );
not \U$485 ( \1289 , RI9145390_115);
not \U$486 ( \1290 , \935 );
not \U$487 ( \1291 , \1290 );
not \U$488 ( \1292 , \1291 );
or \U$489 ( \1293 , \1289 , \1292 );
nand \U$490 ( \1294 , \943 , RI9144c10_99);
nand \U$491 ( \1295 , \1293 , \1294 );
nor \U$492 ( \1296 , \1288 , \1295 );
buf \U$493 ( \1297 , \967 );
and \U$494 ( \1298 , \1297 , RI9138b68_3);
and \U$495 ( \1299 , \963 , RI90f99b8_19);
nor \U$496 ( \1300 , \1298 , \1299 );
not \U$497 ( \1301 , \920 );
not \U$498 ( \1302 , \1301 );
nand \U$499 ( \1303 , \1302 , RI90f3658_35);
nand \U$500 ( \1304 , \928 , RI9143590_51);
and \U$501 ( \1305 , \1300 , \1303 , \1304 );
not \U$502 ( \1306 , RI9146a10_163);
or \U$503 ( \1307 , \989 , \1306 );
not \U$504 ( \1308 , RI9147190_179);
or \U$505 ( \1309 , \994 , \1308 );
nand \U$506 ( \1310 , \1307 , \1309 );
not \U$507 ( \1311 , RI9145b10_131);
not \U$508 ( \1312 , \977 );
or \U$509 ( \1313 , \1311 , \1312 );
nand \U$510 ( \1314 , \984 , RI9146290_147);
nand \U$511 ( \1315 , \1313 , \1314 );
nor \U$512 ( \1316 , \1310 , \1315 );
not \U$513 ( \1317 , RI9147910_195);
not \U$514 ( \1318 , \1003 );
or \U$515 ( \1319 , \1317 , \1318 );
nand \U$516 ( \1320 , \1008 , RI9148090_211);
nand \U$517 ( \1321 , \1319 , \1320 );
not \U$518 ( \1322 , RI9148810_227);
not \U$519 ( \1323 , \1014 );
or \U$520 ( \1324 , \1322 , \1323 );
nand \U$521 ( \1325 , \1251 , RI9148f90_243);
nand \U$522 ( \1326 , \1324 , \1325 );
nor \U$523 ( \1327 , \1321 , \1326 );
nand \U$524 ( \1328 , \1296 , \1305 , \1316 , \1327 );
buf \U$525 ( \1329 , \1328 );
not \U$526 ( \1330 , \1329 );
buf \U$527 ( \1331 , \1330 );
buf \U$528 ( \1332 , \1331 );
not \U$529 ( \1333 , \1332 );
buf \U$530 ( \1334 , \1333 );
buf \U$531 ( \1335 , \1334 );
not \U$532 ( \1336 , \1335 );
buf \U$535 ( \1337 , \1107 );
buf \U$536 ( \1338 , \1337 );
not \U$537 ( \1339 , \1338 );
buf \U$538 ( \1340 , \1339 );
buf \U$539 ( \1341 , \1340 );
not \U$540 ( \1342 , \1341 );
or \U$541 ( \1343 , \1336 , \1342 );
buf \U$542 ( \1344 , \1337 );
buf \U$543 ( \1345 , \1331 );
nand \U$544 ( \1346 , \1344 , \1345 );
buf \U$545 ( \1347 , \1346 );
buf \U$546 ( \1348 , \1347 );
nand \U$547 ( \1349 , \1343 , \1348 );
buf \U$548 ( \1350 , \1349 );
buf \U$549 ( \1351 , \1350 );
not \U$550 ( \1352 , \1351 );
not \U$551 ( \1353 , RI914a778_294);
nor \U$552 ( \1354 , \1353 , \1116 );
not \U$553 ( \1355 , RI914aef8_310);
nor \U$554 ( \1356 , \1355 , \1122 );
nor \U$555 ( \1357 , \1354 , \1356 );
not \U$556 ( \1358 , \836 );
and \U$557 ( \1359 , \1358 , RI914b678_326);
not \U$558 ( \1360 , RI914bdf8_342);
nor \U$559 ( \1361 , \1360 , \1043 );
nor \U$560 ( \1362 , \1359 , \1361 );
and \U$561 ( \1363 , \813 , RI9149ff8_278);
and \U$562 ( \1364 , \818 , RI9149878_262);
nor \U$563 ( \1365 , \1363 , \1364 );
not \U$564 ( \1366 , \850 );
not \U$565 ( \1367 , RI914c578_358);
not \U$566 ( \1368 , \1367 );
and \U$567 ( \1369 , \1366 , \1368 );
not \U$568 ( \1370 , RI914ccf8_374);
nor \U$569 ( \1371 , \1370 , \1093 );
nor \U$570 ( \1372 , \1369 , \1371 );
nand \U$571 ( \1373 , \1357 , \1362 , \1365 , \1372 );
not \U$572 ( \1374 , RI914f278_454);
nor \U$573 ( \1375 , \1374 , \1139 );
not \U$574 ( \1376 , RI914f9f8_470);
not \U$575 ( \1377 , \896 );
nor \U$576 ( \1378 , \1376 , \1377 );
nor \U$577 ( \1379 , \1375 , \1378 );
not \U$578 ( \1380 , RI914d478_390);
nor \U$579 ( \1381 , \1380 , \864 );
not \U$580 ( \1382 , RI914dbf8_406);
nor \U$581 ( \1383 , \1061 , \1382 );
nor \U$582 ( \1384 , \1381 , \1383 );
not \U$583 ( \1385 , RI914e378_422);
not \U$584 ( \1386 , \1069 );
nor \U$585 ( \1387 , \1385 , \1386 );
not \U$586 ( \1388 , RI914eaf8_438);
nor \U$587 ( \1389 , \1388 , \1112 );
nor \U$588 ( \1390 , \1387 , \1389 );
not \U$589 ( \1391 , \900 );
not \U$590 ( \1392 , RI9150178_486);
not \U$591 ( \1393 , \1392 );
and \U$592 ( \1394 , \1391 , \1393 );
not \U$593 ( \1395 , RI91508f8_502);
nor \U$594 ( \1396 , \1395 , \1086 );
nor \U$595 ( \1397 , \1394 , \1396 );
nand \U$596 ( \1398 , \1379 , \1384 , \1390 , \1397 );
nor \U$597 ( \1399 , \1373 , \1398 );
not \U$598 ( \1400 , \1399 );
buf \U$599 ( \1401 , \1400 );
nand \U$600 ( \1402 , \1115 , RI914a7f0_295);
nand \U$601 ( \1403 , \831 , RI914af70_311);
and \U$602 ( \1404 , \1402 , \1403 );
and \U$603 ( \1405 , \1144 , RI914b6f0_327);
not \U$604 ( \1406 , \844 );
and \U$605 ( \1407 , \1406 , RI914be70_343);
nor \U$606 ( \1408 , \1405 , \1407 );
not \U$607 ( \1409 , \818 );
not \U$608 ( \1410 , \1409 );
not \U$609 ( \1411 , RI91498f0_263);
not \U$610 ( \1412 , \1411 );
and \U$611 ( \1413 , \1410 , \1412 );
and \U$612 ( \1414 , \813 , RI914a070_279);
nor \U$613 ( \1415 , \1413 , \1414 );
and \U$614 ( \1416 , \1157 , RI914cd70_375);
not \U$615 ( \1417 , \850 );
and \U$616 ( \1418 , \1417 , RI914c5f0_359);
nor \U$617 ( \1419 , \1416 , \1418 );
nand \U$618 ( \1420 , \1404 , \1408 , \1415 , \1419 );
not \U$619 ( \1421 , \875 );
not \U$620 ( \1422 , RI914e3f0_423);
not \U$621 ( \1423 , \1422 );
and \U$622 ( \1424 , \1421 , \1423 );
not \U$623 ( \1425 , RI914eb70_439);
nor \U$624 ( \1426 , \1425 , \882 );
nor \U$625 ( \1427 , \1424 , \1426 );
not \U$626 ( \1428 , RI914d4f0_391);
nor \U$627 ( \1429 , \1428 , \864 );
not \U$628 ( \1430 , \870 );
not \U$629 ( \1431 , RI914dc70_407);
nor \U$630 ( \1432 , \1430 , \1431 );
nor \U$631 ( \1433 , \1429 , \1432 );
and \U$632 ( \1434 , \888 , RI914f2f0_455);
and \U$633 ( \1435 , \896 , RI914fa70_471);
nor \U$634 ( \1436 , \1434 , \1435 );
not \U$635 ( \1437 , \1129 );
and \U$636 ( \1438 , \1437 , RI91501f0_487);
not \U$637 ( \1439 , \904 );
and \U$638 ( \1440 , \1439 , RI9150970_503);
nor \U$639 ( \1441 , \1438 , \1440 );
nand \U$640 ( \1442 , \1427 , \1433 , \1436 , \1441 );
nor \U$641 ( \1443 , \1420 , \1442 );
not \U$642 ( \1444 , \1443 );
buf \U$643 ( \1445 , \1444 );
not \U$644 ( \1446 , \1445 );
buf \U$645 ( \1447 , \1446 );
buf \U$646 ( \1448 , \1447 );
and \U$647 ( \1449 , \1401 , \1448 );
not \U$648 ( \1450 , \1401 );
buf \U$649 ( \1451 , \1444 );
and \U$650 ( \1452 , \1450 , \1451 );
nor \U$651 ( \1453 , \1449 , \1452 );
buf \U$652 ( \1454 , \1453 );
buf \U$653 ( \1455 , \1454 );
buf \U$654 ( \1456 , \1400 );
buf \U$655 ( \1457 , \1107 );
and \U$656 ( \1458 , \1456 , \1457 );
not \U$657 ( \1459 , \1456 );
buf \U$658 ( \1460 , \1107 );
not \U$659 ( \1461 , \1460 );
buf \U$660 ( \1462 , \1461 );
buf \U$661 ( \1463 , \1462 );
and \U$662 ( \1464 , \1459 , \1463 );
nor \U$663 ( \1465 , \1458 , \1464 );
buf \U$664 ( \1466 , \1465 );
buf \U$665 ( \1467 , \1466 );
nand \U$666 ( \1468 , \1455 , \1467 );
buf \U$667 ( \1469 , \1468 );
buf \U$668 ( \1470 , \1469 );
not \U$669 ( \1471 , \1470 );
buf \U$670 ( \1472 , \1471 );
buf \U$671 ( \1473 , \1472 );
not \U$672 ( \1474 , \1473 );
buf \U$673 ( \1475 , \1474 );
buf \U$674 ( \1476 , \1475 );
not \U$675 ( \1477 , \1476 );
buf \U$676 ( \1478 , \1477 );
buf \U$677 ( \1479 , \1478 );
not \U$678 ( \1480 , \1479 );
or \U$679 ( \1481 , \1352 , \1480 );
buf \U$682 ( \1482 , \1454 );
buf \U$683 ( \1483 , \1482 );
not \U$684 ( \1484 , \1483 );
buf \U$685 ( \1485 , \1484 );
buf \U$686 ( \1486 , \1485 );
not \U$687 ( \1487 , RI912e758_18);
not \U$688 ( \1488 , \963 );
or \U$689 ( \1489 , \1487 , \1488 );
nand \U$690 ( \1490 , RI9138be0_2, \968 );
nand \U$691 ( \1491 , \1489 , \1490 );
not \U$692 ( \1492 , RI9143518_50);
not \U$693 ( \1493 , \928 );
or \U$694 ( \1494 , \1492 , \1493 );
not \U$695 ( \1495 , \1301 );
nand \U$696 ( \1496 , \1495 , RI90f36d0_34);
nand \U$697 ( \1497 , \1494 , \1496 );
nor \U$698 ( \1498 , \1491 , \1497 );
not \U$699 ( \1499 , RI9144418_82);
not \U$700 ( \1500 , \957 );
not \U$701 ( \1501 , \1500 );
or \U$702 ( \1502 , \1499 , \1501 );
nand \U$703 ( \1503 , RI9143c98_66, \951 );
nand \U$704 ( \1504 , \1502 , \1503 );
not \U$705 ( \1505 , RI9145318_114);
not \U$706 ( \1506 , \936 );
or \U$707 ( \1507 , \1505 , \1506 );
not \U$708 ( \1508 , \942 );
nand \U$709 ( \1509 , \1508 , RI9144b98_98);
nand \U$710 ( \1510 , \1507 , \1509 );
nor \U$711 ( \1511 , \1504 , \1510 );
not \U$712 ( \1512 , RI9146998_162);
not \U$713 ( \1513 , \1204 );
or \U$714 ( \1514 , \1512 , \1513 );
nand \U$715 ( \1515 , \1213 , RI9147118_178);
nand \U$716 ( \1516 , \1514 , \1515 );
not \U$717 ( \1517 , RI9145a98_130);
not \U$718 ( \1518 , \977 );
or \U$719 ( \1519 , \1517 , \1518 );
nand \U$720 ( \1520 , \984 , RI9146218_146);
nand \U$721 ( \1521 , \1519 , \1520 );
nor \U$722 ( \1522 , \1516 , \1521 );
not \U$723 ( \1523 , RI9147898_194);
buf \U$724 ( \1524 , \1002 );
not \U$725 ( \1525 , \1524 );
not \U$726 ( \1526 , \1525 );
or \U$727 ( \1527 , \1523 , \1526 );
nand \U$728 ( \1528 , \1008 , RI9148018_210);
nand \U$729 ( \1529 , \1527 , \1528 );
not \U$730 ( \1530 , RI9148798_226);
not \U$731 ( \1531 , \1014 );
or \U$732 ( \1532 , \1530 , \1531 );
nand \U$733 ( \1533 , \1251 , RI9148f18_242);
nand \U$734 ( \1534 , \1532 , \1533 );
nor \U$735 ( \1535 , \1529 , \1534 );
nand \U$736 ( \1536 , \1498 , \1511 , \1522 , \1535 );
buf \U$737 ( \1537 , \1536 );
not \U$738 ( \1538 , \1537 );
buf \U$739 ( \1539 , \1538 );
buf \U$740 ( \1540 , \1539 );
not \U$741 ( \1541 , \1540 );
buf \U$742 ( \1542 , \1541 );
buf \U$743 ( \1543 , \1542 );
not \U$744 ( \1544 , \1543 );
buf \U$745 ( \1545 , \1337 );
not \U$746 ( \1546 , \1545 );
buf \U$747 ( \1547 , \1546 );
buf \U$750 ( \1548 , \1547 );
buf \U$751 ( \1549 , \1548 );
not \U$752 ( \1550 , \1549 );
or \U$753 ( \1551 , \1544 , \1550 );
buf \U$754 ( \1552 , \1337 );
buf \U$755 ( \1553 , \1539 );
nand \U$756 ( \1554 , \1552 , \1553 );
buf \U$757 ( \1555 , \1554 );
buf \U$758 ( \1556 , \1555 );
nand \U$759 ( \1557 , \1551 , \1556 );
buf \U$760 ( \1558 , \1557 );
buf \U$761 ( \1559 , \1558 );
nand \U$762 ( \1560 , \1486 , \1559 );
buf \U$763 ( \1561 , \1560 );
buf \U$764 ( \1562 , \1561 );
nand \U$765 ( \1563 , \1481 , \1562 );
buf \U$766 ( \1564 , \1563 );
buf \U$767 ( \1565 , \1564 );
nand \U$768 ( \1566 , \1281 , \1565 );
buf \U$769 ( \1567 , \1566 );
buf \U$770 ( \1568 , \1567 );
not \U$771 ( \1569 , \1568 );
not \U$772 ( \1570 , RI914aca0_305);
not \U$773 ( \1571 , \831 );
or \U$774 ( \1572 , \1570 , \1571 );
nand \U$775 ( \1573 , \1053 , RI914a520_289);
nand \U$776 ( \1574 , \1572 , \1573 );
not \U$777 ( \1575 , RI914caa0_369);
not \U$778 ( \1576 , \1094 );
or \U$779 ( \1577 , \1575 , \1576 );
nand \U$780 ( \1578 , \1155 , RI914c320_353);
nand \U$781 ( \1579 , \1577 , \1578 );
nor \U$782 ( \1580 , \1574 , \1579 );
not \U$783 ( \1581 , RI914f020_449);
not \U$784 ( \1582 , \1077 );
or \U$785 ( \1583 , \1581 , \1582 );
nand \U$786 ( \1584 , \1080 , RI914f7a0_465);
nand \U$787 ( \1585 , \1583 , \1584 );
not \U$788 ( \1586 , RI914d220_385);
not \U$789 ( \1587 , \1058 );
or \U$790 ( \1588 , \1586 , \1587 );
nand \U$791 ( \1589 , \1062 , RI914d9a0_401);
nand \U$792 ( \1590 , \1588 , \1589 );
nor \U$793 ( \1591 , \1585 , \1590 );
not \U$794 ( \1592 , RI9149da0_273);
not \U$795 ( \1593 , \813 );
or \U$796 ( \1594 , \1592 , \1593 );
not \U$797 ( \1595 , \818 );
not \U$798 ( \1596 , \1595 );
nand \U$799 ( \1597 , \1596 , RI9149620_257);
nand \U$800 ( \1598 , \1594 , \1597 );
not \U$801 ( \1599 , RI914bba0_337);
not \U$802 ( \1600 , \1044 );
or \U$803 ( \1601 , \1599 , \1600 );
nand \U$804 ( \1602 , \1047 , RI914b420_321);
nand \U$805 ( \1603 , \1601 , \1602 );
nor \U$806 ( \1604 , \1598 , \1603 );
not \U$807 ( \1605 , RI914ff20_481);
not \U$808 ( \1606 , \901 );
or \U$809 ( \1607 , \1605 , \1606 );
nand \U$810 ( \1608 , \1087 , RI91506a0_497);
nand \U$811 ( \1609 , \1607 , \1608 );
not \U$812 ( \1610 , RI914e120_417);
not \U$813 ( \1611 , \1069 );
or \U$814 ( \1612 , \1610 , \1611 );
nand \U$815 ( \1613 , \883 , RI914e8a0_433);
nand \U$816 ( \1614 , \1612 , \1613 );
nor \U$817 ( \1615 , \1609 , \1614 );
nand \U$818 ( \1616 , \1580 , \1591 , \1604 , \1615 );
buf \U$819 ( \1617 , \1616 );
buf \U$821 ( \1618 , \1617 );
buf \U$824 ( \1619 , \1618 );
buf \U$825 ( \1620 , \1619 );
not \U$826 ( \1621 , RI9143860_57);
buf \U$827 ( \1622 , \927 );
not \U$828 ( \1623 , \1622 );
not \U$829 ( \1624 , \1623 );
or \U$830 ( \1625 , \1621 , \1624 );
nand \U$831 ( \1626 , \921 , RI90f3388_41);
nand \U$832 ( \1627 , \1625 , \1626 );
not \U$833 ( \1628 , RI9145660_121);
not \U$834 ( \1629 , \1291 );
or \U$835 ( \1630 , \1628 , \1629 );
nand \U$836 ( \1631 , \943 , RI9144ee0_105);
nand \U$837 ( \1632 , \1630 , \1631 );
nor \U$838 ( \1633 , \1627 , \1632 );
not \U$839 ( \1634 , RI9144760_89);
not \U$840 ( \1635 , \957 );
not \U$841 ( \1636 , \1635 );
or \U$842 ( \1637 , \1634 , \1636 );
nand \U$843 ( \1638 , \951 , RI9143fe0_73);
nand \U$844 ( \1639 , \1637 , \1638 );
not \U$845 ( \1640 , RI90f96e8_25);
not \U$846 ( \1641 , \963 );
or \U$847 ( \1642 , \1640 , \1641 );
nand \U$848 ( \1643 , \1297 , RI9138898_9);
nand \U$849 ( \1644 , \1642 , \1643 );
nor \U$850 ( \1645 , \1639 , \1644 );
not \U$851 ( \1646 , RI9146ce0_169);
not \U$852 ( \1647 , \1206 );
or \U$853 ( \1648 , \1646 , \1647 );
nand \U$854 ( \1649 , \1213 , RI9147460_185);
nand \U$855 ( \1650 , \1648 , \1649 );
not \U$856 ( \1651 , RI9145de0_137);
not \U$857 ( \1652 , \977 );
or \U$858 ( \1653 , \1651 , \1652 );
nand \U$859 ( \1654 , \1244 , RI9146560_153);
nand \U$860 ( \1655 , \1653 , \1654 );
nor \U$861 ( \1656 , \1650 , \1655 );
not \U$862 ( \1657 , RI9147be0_201);
not \U$863 ( \1658 , \1003 );
or \U$864 ( \1659 , \1657 , \1658 );
nand \U$865 ( \1660 , \1008 , RI9148360_217);
nand \U$866 ( \1661 , \1659 , \1660 );
not \U$867 ( \1662 , RI9148ae0_233);
not \U$868 ( \1663 , \1014 );
or \U$869 ( \1664 , \1662 , \1663 );
nand \U$870 ( \1665 , \1251 , RI9149260_249);
nand \U$871 ( \1666 , \1664 , \1665 );
nor \U$872 ( \1667 , \1661 , \1666 );
nand \U$873 ( \1668 , \1633 , \1645 , \1656 , \1667 );
buf \U$874 ( \1669 , \1668 );
buf \U$875 ( \1670 , \1669 );
and \U$876 ( \1671 , \1620 , \1670 );
buf \U$877 ( \1672 , \1671 );
buf \U$878 ( \1673 , \1672 );
not \U$879 ( \1674 , \1673 );
not \U$880 ( \1675 , RI9149e18_274);
not \U$881 ( \1676 , \813 );
or \U$882 ( \1677 , \1675 , \1676 );
not \U$883 ( \1678 , \818 );
not \U$884 ( \1679 , \1678 );
nand \U$885 ( \1680 , \1679 , RI9149698_258);
nand \U$886 ( \1681 , \1677 , \1680 );
not \U$887 ( \1682 , RI914ad18_306);
not \U$888 ( \1683 , \831 );
or \U$889 ( \1684 , \1682 , \1683 );
nand \U$890 ( \1685 , \1053 , RI914a598_290);
nand \U$891 ( \1686 , \1684 , \1685 );
nor \U$892 ( \1687 , \1681 , \1686 );
not \U$893 ( \1688 , RI914bc18_338);
not \U$894 ( \1689 , \1044 );
or \U$895 ( \1690 , \1688 , \1689 );
nand \U$896 ( \1691 , \1047 , RI914b498_322);
nand \U$897 ( \1692 , \1690 , \1691 );
not \U$898 ( \1693 , RI914cb18_370);
not \U$899 ( \1694 , \1094 );
or \U$900 ( \1695 , \1693 , \1694 );
not \U$901 ( \1696 , \850 );
nand \U$902 ( \1697 , \1696 , RI914c398_354);
nand \U$903 ( \1698 , \1695 , \1697 );
nor \U$904 ( \1699 , \1692 , \1698 );
not \U$905 ( \1700 , RI914d298_386);
not \U$906 ( \1701 , \1058 );
or \U$907 ( \1702 , \1700 , \1701 );
nand \U$908 ( \1703 , \1062 , RI914da18_402);
nand \U$909 ( \1704 , \1702 , \1703 );
not \U$910 ( \1705 , RI914e198_418);
not \U$911 ( \1706 , \1069 );
or \U$912 ( \1707 , \1705 , \1706 );
nand \U$913 ( \1708 , \883 , RI914e918_434);
nand \U$914 ( \1709 , \1707 , \1708 );
nor \U$915 ( \1710 , \1704 , \1709 );
not \U$916 ( \1711 , RI914f098_450);
not \U$917 ( \1712 , \1077 );
or \U$918 ( \1713 , \1711 , \1712 );
nand \U$919 ( \1714 , \1080 , RI914f818_466);
nand \U$920 ( \1715 , \1713 , \1714 );
not \U$921 ( \1716 , RI914ff98_482);
not \U$922 ( \1717 , \901 );
or \U$923 ( \1718 , \1716 , \1717 );
nand \U$924 ( \1719 , \1087 , RI9150718_498);
nand \U$925 ( \1720 , \1718 , \1719 );
nor \U$926 ( \1721 , \1715 , \1720 );
nand \U$927 ( \1722 , \1687 , \1699 , \1710 , \1721 );
buf \U$928 ( \1723 , \1722 );
buf \U$929 ( \1724 , \909 );
not \U$930 ( \1725 , \1724 );
buf \U$931 ( \1726 , \1725 );
buf \U$932 ( \1727 , \1726 );
and \U$933 ( \1728 , \1723 , \1727 );
not \U$934 ( \1729 , \1723 );
buf \U$935 ( \1730 , \909 );
and \U$936 ( \1731 , \1729 , \1730 );
nor \U$937 ( \1732 , \1728 , \1731 );
buf \U$938 ( \1733 , \1732 );
buf \U$939 ( \1734 , \1733 );
buf \U$940 ( \1735 , \1616 );
not \U$941 ( \1736 , \1735 );
buf \U$942 ( \1737 , \1736 );
buf \U$943 ( \1738 , \1737 );
not \U$944 ( \1739 , \1738 );
buf \U$945 ( \1740 , \1722 );
not \U$946 ( \1741 , \1740 );
or \U$947 ( \1742 , \1739 , \1741 );
buf \U$948 ( \1743 , \1722 );
not \U$949 ( \1744 , \1743 );
buf \U$950 ( \1745 , \1744 );
buf \U$951 ( \1746 , \1745 );
buf \U$952 ( \1747 , \1616 );
nand \U$953 ( \1748 , \1746 , \1747 );
buf \U$954 ( \1749 , \1748 );
buf \U$955 ( \1750 , \1749 );
nand \U$956 ( \1751 , \1742 , \1750 );
buf \U$957 ( \1752 , \1751 );
buf \U$958 ( \1753 , \1752 );
nand \U$959 ( \1754 , \1734 , \1753 );
buf \U$960 ( \1755 , \1754 );
buf \U$961 ( \1756 , \1755 );
not \U$962 ( \1757 , \1756 );
buf \U$963 ( \1758 , \1757 );
buf \U$964 ( \1759 , \1758 );
not \U$965 ( \1760 , \1759 );
and \U$966 ( \1761 , \1003 , RI9147b68_200);
and \U$967 ( \1762 , \1008 , RI91482e8_216);
nor \U$968 ( \1763 , \1761 , \1762 );
and \U$969 ( \1764 , \977 , RI9145d68_136);
not \U$970 ( \1765 , \983 );
and \U$971 ( \1766 , \1765 , RI91464e8_152);
nor \U$972 ( \1767 , \1764 , \1766 );
and \U$973 ( \1768 , \1206 , RI9146c68_168);
and \U$974 ( \1769 , \1213 , RI91473e8_184);
nor \U$975 ( \1770 , \1768 , \1769 );
and \U$976 ( \1771 , \1014 , RI9148a68_232);
and \U$977 ( \1772 , \1251 , RI91491e8_248);
nor \U$978 ( \1773 , \1771 , \1772 );
nand \U$979 ( \1774 , \1763 , \1767 , \1770 , \1773 );
nand \U$980 ( \1775 , \951 , RI9143f68_72);
nand \U$981 ( \1776 , \1500 , RI91446e8_88);
and \U$982 ( \1777 , \1775 , \1776 );
and \U$983 ( \1778 , \921 , RI90f3400_40);
and \U$984 ( \1779 , \928 , RI91437e8_56);
nor \U$985 ( \1780 , \1778 , \1779 );
and \U$986 ( \1781 , \1508 , RI9144e68_104);
and \U$987 ( \1782 , \936 , RI91455e8_120);
nor \U$988 ( \1783 , \1781 , \1782 );
and \U$989 ( \1784 , \963 , RI90f9760_24);
and \U$990 ( \1785 , \1297 , RI9138910_8);
nor \U$991 ( \1786 , \1784 , \1785 );
nand \U$992 ( \1787 , \1777 , \1780 , \1783 , \1786 );
nor \U$993 ( \1788 , \1774 , \1787 );
not \U$994 ( \1789 , \1788 );
buf \U$995 ( \1790 , \1789 );
not \U$996 ( \1791 , \1790 );
buf \U$997 ( \1792 , \1791 );
buf \U$998 ( \1793 , \1792 );
not \U$999 ( \1794 , \1793 );
buf \U$1000 ( \1795 , \1794 );
buf \U$1001 ( \1796 , \1795 );
not \U$1002 ( \1797 , \1796 );
buf \U$1003 ( \1798 , \1618 );
not \U$1004 ( \1799 , \1798 );
buf \U$1005 ( \1800 , \1799 );
buf \U$1006 ( \1801 , \1800 );
not \U$1007 ( \1802 , \1801 );
or \U$1008 ( \1803 , \1797 , \1802 );
buf \U$1009 ( \1804 , \1792 );
buf \U$1010 ( \1805 , \1618 );
nand \U$1011 ( \1806 , \1804 , \1805 );
buf \U$1012 ( \1807 , \1806 );
buf \U$1013 ( \1808 , \1807 );
nand \U$1014 ( \1809 , \1803 , \1808 );
buf \U$1015 ( \1810 , \1809 );
buf \U$1016 ( \1811 , \1810 );
not \U$1017 ( \1812 , \1811 );
or \U$1018 ( \1813 , \1760 , \1812 );
buf \U$1019 ( \1814 , \1618 );
not \U$1020 ( \1815 , \1814 );
buf \U$1021 ( \1816 , \1815 );
buf \U$1022 ( \1817 , \1816 );
not \U$1023 ( \1818 , \1817 );
not \U$1024 ( \1819 , \957 );
not \U$1025 ( \1820 , RI9144670_87);
not \U$1026 ( \1821 , \1820 );
and \U$1027 ( \1822 , \1819 , \1821 );
and \U$1028 ( \1823 , \951 , RI9143ef0_71);
nor \U$1029 ( \1824 , \1822 , \1823 );
not \U$1030 ( \1825 , \1622 );
not \U$1031 ( \1826 , RI9143770_55);
not \U$1032 ( \1827 , \1826 );
and \U$1033 ( \1828 , \1825 , \1827 );
not \U$1034 ( \1829 , RI90f3478_39);
nor \U$1035 ( \1830 , \1829 , \1301 );
nor \U$1036 ( \1831 , \1828 , \1830 );
and \U$1037 ( \1832 , \936 , RI9145570_119);
and \U$1038 ( \1833 , \1508 , RI9144df0_103);
nor \U$1039 ( \1834 , \1832 , \1833 );
nand \U$1040 ( \1835 , \963 , RI90f97d8_23);
nand \U$1041 ( \1836 , \1297 , RI9138988_7);
and \U$1042 ( \1837 , \1835 , \1836 );
nand \U$1043 ( \1838 , \1824 , \1831 , \1834 , \1837 );
not \U$1044 ( \1839 , RI9146bf0_167);
nor \U$1045 ( \1840 , \1839 , \989 );
not \U$1046 ( \1841 , RI9147370_183);
nor \U$1047 ( \1842 , \1841 , \994 );
nor \U$1048 ( \1843 , \1840 , \1842 );
not \U$1049 ( \1844 , RI9147af0_199);
nor \U$1050 ( \1845 , \1844 , \1524 );
not \U$1051 ( \1846 , RI9148270_215);
not \U$1052 ( \1847 , \1008 );
nor \U$1053 ( \1848 , \1846 , \1847 );
nor \U$1054 ( \1849 , \1845 , \1848 );
not \U$1055 ( \1850 , RI9145cf0_135);
nor \U$1056 ( \1851 , \1850 , \976 );
not \U$1057 ( \1852 , RI9146470_151);
nor \U$1058 ( \1853 , \1852 , \983 );
nor \U$1059 ( \1854 , \1851 , \1853 );
and \U$1060 ( \1855 , \1014 , RI91489f0_231);
not \U$1061 ( \1856 , RI9149170_247);
nand \U$1062 ( \1857 , RI91588f0_775, RI9158968_776, RI9158878_774, RI91589e0_777);
nor \U$1063 ( \1858 , \1856 , \1857 );
nor \U$1064 ( \1859 , \1855 , \1858 );
nand \U$1065 ( \1860 , \1843 , \1849 , \1854 , \1859 );
nor \U$1066 ( \1861 , \1838 , \1860 );
not \U$1067 ( \1862 , \1861 );
buf \U$1068 ( \1863 , \1862 );
not \U$1069 ( \1864 , \1863 );
buf \U$1070 ( \1865 , \1864 );
buf \U$1071 ( \1866 , \1865 );
not \U$1072 ( \1867 , \1866 );
buf \U$1073 ( \1868 , \1867 );
buf \U$1074 ( \1869 , \1868 );
not \U$1075 ( \1870 , \1869 );
or \U$1076 ( \1871 , \1818 , \1870 );
buf \U$1077 ( \1872 , \1865 );
buf \U$1078 ( \1873 , \1618 );
nand \U$1079 ( \1874 , \1872 , \1873 );
buf \U$1080 ( \1875 , \1874 );
buf \U$1081 ( \1876 , \1875 );
nand \U$1082 ( \1877 , \1871 , \1876 );
buf \U$1083 ( \1878 , \1877 );
buf \U$1084 ( \1879 , \1878 );
buf \U$1085 ( \1880 , \1733 );
not \U$1086 ( \1881 , \1880 );
buf \U$1087 ( \1882 , \1881 );
buf \U$1088 ( \1883 , \1882 );
nand \U$1089 ( \1884 , \1879 , \1883 );
buf \U$1090 ( \1885 , \1884 );
buf \U$1091 ( \1886 , \1885 );
nand \U$1092 ( \1887 , \1813 , \1886 );
buf \U$1093 ( \1888 , \1887 );
buf \U$1094 ( \1889 , \1888 );
not \U$1095 ( \1890 , \1889 );
or \U$1096 ( \1891 , \1674 , \1890 );
or \U$1097 ( \1892 , \1672 , \1888 );
and \U$1098 ( \1893 , \1340 , \1261 );
not \U$1099 ( \1894 , \1340 );
and \U$1100 ( \1895 , \1894 , \1258 );
or \U$1101 ( \1896 , \1893 , \1895 );
buf \U$1102 ( \1897 , \1896 );
not \U$1103 ( \1898 , \1897 );
buf \U$1104 ( \1899 , \1478 );
not \U$1105 ( \1900 , \1899 );
or \U$1106 ( \1901 , \1898 , \1900 );
buf \U$1107 ( \1902 , \1482 );
not \U$1108 ( \1903 , \1902 );
buf \U$1109 ( \1904 , \1903 );
buf \U$1110 ( \1905 , \1904 );
buf \U$1111 ( \1906 , \1350 );
nand \U$1112 ( \1907 , \1905 , \1906 );
buf \U$1113 ( \1908 , \1907 );
buf \U$1114 ( \1909 , \1908 );
nand \U$1115 ( \1910 , \1901 , \1909 );
buf \U$1116 ( \1911 , \1910 );
nand \U$1117 ( \1912 , \1892 , \1911 );
buf \U$1118 ( \1913 , \1912 );
nand \U$1119 ( \1914 , \1891 , \1913 );
buf \U$1120 ( \1915 , \1914 );
buf \U$1121 ( \1916 , \1915 );
not \U$1122 ( \1917 , \1916 );
or \U$1123 ( \1918 , \1569 , \1917 );
buf \U$1124 ( \1919 , \1564 );
not \U$1125 ( \1920 , \1919 );
buf \U$1126 ( \1921 , \1279 );
nand \U$1127 ( \1922 , \1920 , \1921 );
buf \U$1128 ( \1923 , \1922 );
buf \U$1129 ( \1924 , \1923 );
nand \U$1130 ( \1925 , \1918 , \1924 );
buf \U$1131 ( \1926 , \1925 );
buf \U$1132 ( \1927 , \1926 );
buf \U$1133 ( \1928 , \1619 );
buf \U$1134 ( \1929 , \1789 );
not \U$1135 ( \1930 , \1929 );
buf \U$1136 ( \1931 , \1930 );
buf \U$1137 ( \1932 , \1931 );
not \U$1138 ( \1933 , \1932 );
buf \U$1139 ( \1934 , \1933 );
buf \U$1140 ( \1935 , \1934 );
and \U$1141 ( \1936 , \1928 , \1935 );
buf \U$1142 ( \1937 , \1936 );
buf \U$1143 ( \1938 , \1937 );
buf \U$1144 ( \1939 , \1878 );
not \U$1145 ( \1940 , \1939 );
buf \U$1146 ( \1941 , \1758 );
not \U$1147 ( \1942 , \1941 );
buf \U$1148 ( \1943 , \1942 );
buf \U$1149 ( \1944 , \1943 );
not \U$1150 ( \1945 , \1944 );
buf \U$1151 ( \1946 , \1945 );
buf \U$1152 ( \1947 , \1946 );
not \U$1153 ( \1948 , \1947 );
or \U$1154 ( \1949 , \1940 , \1948 );
buf \U$1157 ( \1950 , \1882 );
buf \U$1158 ( \1951 , \1950 );
nand \U$1159 ( \1952 , \951 , RI9143e78_70);
nand \U$1160 ( \1953 , \1218 , RI91445f8_86);
nand \U$1161 ( \1954 , \1014 , RI9148978_230);
nand \U$1162 ( \1955 , \1251 , RI91490f8_246);
and \U$1163 ( \1956 , \1952 , \1953 , \1954 , \1955 );
not \U$1164 ( \1957 , RI9147a78_198);
not \U$1165 ( \1958 , \1003 );
or \U$1166 ( \1959 , \1957 , \1958 );
nand \U$1167 ( \1960 , \1200 , RI91481f8_214);
nand \U$1168 ( \1961 , \1959 , \1960 );
not \U$1169 ( \1962 , RI91454f8_118);
not \U$1170 ( \1963 , \1291 );
or \U$1171 ( \1964 , \1962 , \1963 );
nand \U$1172 ( \1965 , \1226 , RI9144d78_102);
nand \U$1173 ( \1966 , \1964 , \1965 );
nor \U$1174 ( \1967 , \1961 , \1966 );
not \U$1175 ( \1968 , RI91436f8_54);
not \U$1176 ( \1969 , \928 );
or \U$1177 ( \1970 , \1968 , \1969 );
nand \U$1178 ( \1971 , \1495 , RI90f34f0_38);
nand \U$1179 ( \1972 , \1970 , \1971 );
not \U$1180 ( \1973 , RI90f9850_22);
not \U$1181 ( \1974 , \963 );
or \U$1182 ( \1975 , \1973 , \1974 );
nand \U$1183 ( \1976 , \968 , RI9138a00_6);
nand \U$1184 ( \1977 , \1975 , \1976 );
nor \U$1185 ( \1978 , \1972 , \1977 );
not \U$1186 ( \1979 , RI9145c78_134);
not \U$1187 ( \1980 , \977 );
or \U$1188 ( \1981 , \1979 , \1980 );
nand \U$1189 ( \1982 , \1244 , RI91463f8_150);
nand \U$1190 ( \1983 , \1981 , \1982 );
not \U$1191 ( \1984 , RI9146b78_166);
not \U$1192 ( \1985 , \1204 );
or \U$1193 ( \1986 , \1984 , \1985 );
nand \U$1194 ( \1987 , \1211 , RI91472f8_182);
nand \U$1195 ( \1988 , \1986 , \1987 );
nor \U$1196 ( \1989 , \1983 , \1988 );
nand \U$1197 ( \1990 , \1956 , \1967 , \1978 , \1989 );
buf \U$1198 ( \1991 , \1990 );
not \U$1199 ( \1992 , \1991 );
buf \U$1200 ( \1993 , \1619 );
not \U$1201 ( \1994 , \1993 );
buf \U$1202 ( \1995 , \1994 );
buf \U$1203 ( \1996 , \1995 );
not \U$1204 ( \1997 , \1996 );
or \U$1205 ( \1998 , \1992 , \1997 );
not \U$1206 ( \1999 , \1990 );
buf \U$1207 ( \2000 , \1999 );
buf \U$1208 ( \2001 , \1619 );
nand \U$1209 ( \2002 , \2000 , \2001 );
buf \U$1210 ( \2003 , \2002 );
buf \U$1211 ( \2004 , \2003 );
nand \U$1212 ( \2005 , \1998 , \2004 );
buf \U$1213 ( \2006 , \2005 );
buf \U$1214 ( \2007 , \2006 );
nand \U$1215 ( \2008 , \1951 , \2007 );
buf \U$1216 ( \2009 , \2008 );
buf \U$1217 ( \2010 , \2009 );
nand \U$1218 ( \2011 , \1949 , \2010 );
buf \U$1219 ( \2012 , \2011 );
buf \U$1220 ( \2013 , \2012 );
xor \U$1221 ( \2014 , \1938 , \2013 );
not \U$1222 ( \2015 , RI90f3748_33);
or \U$1223 ( \2016 , \922 , \2015 );
not \U$1224 ( \2017 , \1622 );
nand \U$1225 ( \2018 , \2017 , RI91434a0_49);
nand \U$1226 ( \2019 , \2016 , \2018 );
not \U$1227 ( \2020 , RI91452a0_113);
not \U$1228 ( \2021 , \1291 );
or \U$1229 ( \2022 , \2020 , \2021 );
nand \U$1230 ( \2023 , \943 , RI9144b20_97);
nand \U$1231 ( \2024 , \2022 , \2023 );
nor \U$1232 ( \2025 , \2019 , \2024 );
not \U$1233 ( \2026 , RI912e7d0_17);
not \U$1234 ( \2027 , \963 );
or \U$1235 ( \2028 , \2026 , \2027 );
nand \U$1236 ( \2029 , \968 , RI9138c58_1);
nand \U$1237 ( \2030 , \2028 , \2029 );
not \U$1238 ( \2031 , \951 );
not \U$1239 ( \2032 , RI9143c20_65);
or \U$1240 ( \2033 , \2031 , \2032 );
not \U$1241 ( \2034 , RI91443a0_81);
or \U$1242 ( \2035 , \1285 , \2034 );
nand \U$1243 ( \2036 , \2033 , \2035 );
nor \U$1244 ( \2037 , \2030 , \2036 );
not \U$1245 ( \2038 , RI9145a20_129);
not \U$1246 ( \2039 , \977 );
or \U$1247 ( \2040 , \2038 , \2039 );
nand \U$1248 ( \2041 , \984 , RI91461a0_145);
nand \U$1249 ( \2042 , \2040 , \2041 );
not \U$1250 ( \2043 , RI9146920_161);
or \U$1251 ( \2044 , \989 , \2043 );
not \U$1252 ( \2045 , RI91470a0_177);
or \U$1253 ( \2046 , \994 , \2045 );
nand \U$1254 ( \2047 , \2044 , \2046 );
nor \U$1255 ( \2048 , \2042 , \2047 );
not \U$1256 ( \2049 , RI9147820_193);
not \U$1257 ( \2050 , \1525 );
or \U$1258 ( \2051 , \2049 , \2050 );
not \U$1259 ( \2052 , \1199 );
nand \U$1260 ( \2053 , \2052 , RI9147fa0_209);
nand \U$1261 ( \2054 , \2051 , \2053 );
not \U$1262 ( \2055 , RI9148720_225);
not \U$1263 ( \2056 , \1014 );
or \U$1264 ( \2057 , \2055 , \2056 );
nand \U$1265 ( \2058 , \1251 , RI9148ea0_241);
nand \U$1266 ( \2059 , \2057 , \2058 );
nor \U$1267 ( \2060 , \2054 , \2059 );
nand \U$1268 ( \2061 , \2025 , \2037 , \2048 , \2060 );
buf \U$1269 ( \2062 , \2061 );
buf \U$1271 ( \2063 , \2062 );
buf \U$1272 ( \2064 , \2063 );
not \U$1273 ( \2065 , \2064 );
buf \U$1274 ( \2066 , \1444 );
buf \U$1276 ( \2067 , \2066 );
buf \U$1279 ( \2068 , \2067 );
buf \U$1280 ( \2069 , \2068 );
not \U$1281 ( \2070 , \2069 );
buf \U$1282 ( \2071 , \2070 );
buf \U$1283 ( \2072 , \2071 );
not \U$1284 ( \2073 , \2072 );
or \U$1285 ( \2074 , \2065 , \2073 );
buf \U$1286 ( \2075 , \2068 );
buf \U$1287 ( \2076 , \2063 );
not \U$1288 ( \2077 , \2076 );
buf \U$1289 ( \2078 , \2077 );
buf \U$1290 ( \2079 , \2078 );
nand \U$1291 ( \2080 , \2075 , \2079 );
buf \U$1292 ( \2081 , \2080 );
buf \U$1293 ( \2082 , \2081 );
nand \U$1294 ( \2083 , \2074 , \2082 );
buf \U$1295 ( \2084 , \2083 );
buf \U$1296 ( \2085 , \2084 );
not \U$1297 ( \2086 , \2085 );
not \U$1298 ( \2087 , RI914ce60_377);
not \U$1299 ( \2088 , \1094 );
or \U$1300 ( \2089 , \2087 , \2088 );
nand \U$1301 ( \2090 , RI914c6e0_361, \1097 );
nand \U$1302 ( \2091 , \2089 , \2090 );
not \U$1303 ( \2092 , RI914a160_281);
not \U$1304 ( \2093 , \813 );
or \U$1305 ( \2094 , \2092 , \2093 );
nand \U$1306 ( \2095 , \818 , RI91499e0_265);
nand \U$1307 ( \2096 , \2094 , \2095 );
nor \U$1308 ( \2097 , \2091 , \2096 );
not \U$1309 ( \2098 , RI914e4e0_425);
not \U$1310 ( \2099 , \1069 );
or \U$1311 ( \2100 , \2098 , \2099 );
nand \U$1312 ( \2101 , \883 , RI914ec60_441);
nand \U$1313 ( \2102 , \2100 , \2101 );
not \U$1314 ( \2103 , RI914d5e0_393);
not \U$1315 ( \2104 , \865 );
or \U$1316 ( \2105 , \2103 , \2104 );
nand \U$1317 ( \2106 , \1062 , RI914dd60_409);
nand \U$1318 ( \2107 , \2105 , \2106 );
nor \U$1319 ( \2108 , \2102 , \2107 );
not \U$1320 ( \2109 , RI914f3e0_457);
not \U$1321 ( \2110 , \1077 );
or \U$1322 ( \2111 , \2109 , \2110 );
nand \U$1323 ( \2112 , \1080 , RI914fb60_473);
nand \U$1324 ( \2113 , \2111 , \2112 );
not \U$1325 ( \2114 , RI91502e0_489);
not \U$1326 ( \2115 , \901 );
or \U$1327 ( \2116 , \2114 , \2115 );
nand \U$1328 ( \2117 , \1087 , RI9150a60_505);
nand \U$1329 ( \2118 , \2116 , \2117 );
nor \U$1330 ( \2119 , \2113 , \2118 );
not \U$1331 ( \2120 , RI914b060_313);
not \U$1332 ( \2121 , \831 );
or \U$1333 ( \2122 , \2120 , \2121 );
nand \U$1334 ( \2123 , \1053 , RI914a8e0_297);
nand \U$1335 ( \2124 , \2122 , \2123 );
not \U$1336 ( \2125 , RI914bf60_345);
not \U$1337 ( \2126 , \1044 );
or \U$1338 ( \2127 , \2125 , \2126 );
nand \U$1339 ( \2128 , \1358 , RI914b7e0_329);
nand \U$1340 ( \2129 , \2127 , \2128 );
nor \U$1341 ( \2130 , \2124 , \2129 );
nand \U$1342 ( \2131 , \2097 , \2108 , \2119 , \2130 );
buf \U$1343 ( \2132 , \2131 );
and \U$1344 ( \2133 , \813 , RI914a0e8_280);
not \U$1345 ( \2134 , RI9149968_264);
nor \U$1346 ( \2135 , \2134 , \1595 );
nor \U$1347 ( \2136 , \2133 , \2135 );
nand \U$1348 ( \2137 , \1358 , RI914b768_328);
nand \U$1349 ( \2138 , \1406 , RI914bee8_344);
and \U$1350 ( \2139 , \2137 , \2138 );
not \U$1351 ( \2140 , \825 );
nand \U$1352 ( \2141 , \2140 , RI914a868_296);
nand \U$1353 ( \2142 , \831 , RI914afe8_312);
and \U$1354 ( \2143 , \2141 , \2142 );
and \U$1355 ( \2144 , \1155 , RI914c668_360);
and \U$1356 ( \2145 , \1157 , RI914cde8_376);
nor \U$1357 ( \2146 , \2144 , \2145 );
nand \U$1358 ( \2147 , \2136 , \2139 , \2143 , \2146 );
not \U$1359 ( \2148 , \1068 );
not \U$1360 ( \2149 , RI914e468_424);
not \U$1361 ( \2150 , \2149 );
and \U$1362 ( \2151 , \2148 , \2150 );
not \U$1363 ( \2152 , RI914ebe8_440);
nor \U$1364 ( \2153 , \2152 , \884 );
nor \U$1365 ( \2154 , \2151 , \2153 );
not \U$1366 ( \2155 , RI914d568_392);
nor \U$1367 ( \2156 , \2155 , \864 );
not \U$1368 ( \2157 , RI914dce8_408);
nor \U$1369 ( \2158 , \2157 , \1430 );
nor \U$1370 ( \2159 , \2156 , \2158 );
and \U$1371 ( \2160 , \888 , RI914f368_456);
and \U$1372 ( \2161 , \1141 , RI914fae8_472);
nor \U$1373 ( \2162 , \2160 , \2161 );
and \U$1374 ( \2163 , \1437 , RI9150268_488);
and \U$1375 ( \2164 , \1439 , RI91509e8_504);
nor \U$1376 ( \2165 , \2163 , \2164 );
nand \U$1377 ( \2166 , \2154 , \2159 , \2162 , \2165 );
nor \U$1378 ( \2167 , \2147 , \2166 );
not \U$1379 ( \2168 , \2167 );
buf \U$1380 ( \2169 , \2168 );
not \U$1381 ( \2170 , \2169 );
buf \U$1382 ( \2171 , \2170 );
buf \U$1383 ( \2172 , \2171 );
and \U$1384 ( \2173 , \2132 , \2172 );
not \U$1385 ( \2174 , \2132 );
buf \U$1386 ( \2175 , \2168 );
and \U$1387 ( \2176 , \2174 , \2175 );
nor \U$1388 ( \2177 , \2173 , \2176 );
buf \U$1389 ( \2178 , \2177 );
buf \U$1390 ( \2179 , \2178 );
buf \U$1391 ( \2180 , \1447 );
not \U$1392 ( \2181 , \2180 );
buf \U$1393 ( \2182 , \2168 );
not \U$1394 ( \2183 , \2182 );
or \U$1395 ( \2184 , \2181 , \2183 );
buf \U$1396 ( \2185 , \2168 );
not \U$1397 ( \2186 , \2185 );
buf \U$1398 ( \2187 , \2186 );
buf \U$1399 ( \2188 , \2187 );
buf \U$1400 ( \2189 , \1444 );
nand \U$1401 ( \2190 , \2188 , \2189 );
buf \U$1402 ( \2191 , \2190 );
buf \U$1403 ( \2192 , \2191 );
nand \U$1404 ( \2193 , \2184 , \2192 );
buf \U$1405 ( \2194 , \2193 );
buf \U$1406 ( \2195 , \2194 );
nand \U$1407 ( \2196 , \2179 , \2195 );
buf \U$1408 ( \2197 , \2196 );
buf \U$1409 ( \2198 , \2197 );
not \U$1410 ( \2199 , \2198 );
buf \U$1411 ( \2200 , \2199 );
buf \U$1414 ( \2201 , \2200 );
buf \U$1415 ( \2202 , \2201 );
not \U$1416 ( \2203 , \2202 );
or \U$1417 ( \2204 , \2086 , \2203 );
buf \U$1418 ( \2205 , \2067 );
buf \U$1419 ( \2206 , \2178 );
not \U$1420 ( \2207 , \2206 );
buf \U$1421 ( \2208 , \2207 );
buf \U$1422 ( \2209 , \2208 );
not \U$1423 ( \2210 , \2209 );
buf \U$1424 ( \2211 , \2210 );
buf \U$1425 ( \2212 , \2211 );
not \U$1426 ( \2213 , \2212 );
buf \U$1427 ( \2214 , \2213 );
buf \U$1428 ( \2215 , \2214 );
nand \U$1429 ( \2216 , \2205 , \2215 );
buf \U$1430 ( \2217 , \2216 );
buf \U$1431 ( \2218 , \2217 );
nand \U$1432 ( \2219 , \2204 , \2218 );
buf \U$1433 ( \2220 , \2219 );
buf \U$1434 ( \2221 , \2220 );
and \U$1435 ( \2222 , \2014 , \2221 );
and \U$1436 ( \2223 , \1938 , \2013 );
or \U$1437 ( \2224 , \2222 , \2223 );
buf \U$1438 ( \2225 , \2224 );
buf \U$1439 ( \2226 , \2225 );
buf \U$1440 ( \2227 , \1619 );
buf \U$1441 ( \2228 , \1868 );
and \U$1442 ( \2229 , \2227 , \2228 );
buf \U$1443 ( \2230 , \2229 );
buf \U$1444 ( \2231 , \2230 );
buf \U$1445 ( \2232 , \1564 );
xor \U$1446 ( \2233 , \2231 , \2232 );
buf \U$1447 ( \2234 , \1273 );
not \U$1448 ( \2235 , \2234 );
buf \U$1449 ( \2236 , \1187 );
not \U$1450 ( \2237 , \2236 );
or \U$1451 ( \2238 , \2235 , \2237 );
buf \U$1452 ( \2239 , \1194 );
buf \U$1453 ( \2240 , \1334 );
buf \U$1454 ( \2241 , \911 );
and \U$1455 ( \2242 , \2240 , \2241 );
not \U$1456 ( \2243 , \2240 );
buf \U$1457 ( \2244 , \914 );
and \U$1458 ( \2245 , \2243 , \2244 );
nor \U$1459 ( \2246 , \2242 , \2245 );
buf \U$1460 ( \2247 , \2246 );
buf \U$1461 ( \2248 , \2247 );
nand \U$1462 ( \2249 , \2239 , \2248 );
buf \U$1463 ( \2250 , \2249 );
buf \U$1464 ( \2251 , \2250 );
nand \U$1465 ( \2252 , \2238 , \2251 );
buf \U$1466 ( \2253 , \2252 );
buf \U$1467 ( \2254 , \2253 );
xor \U$1468 ( \2255 , \2233 , \2254 );
buf \U$1469 ( \2256 , \2255 );
buf \U$1470 ( \2257 , \2256 );
xor \U$1471 ( \2258 , \2226 , \2257 );
buf \U$1472 ( \2259 , \1558 );
not \U$1473 ( \2260 , \2259 );
buf \U$1476 ( \2261 , \1478 );
buf \U$1477 ( \2262 , \2261 );
not \U$1478 ( \2263 , \2262 );
or \U$1479 ( \2264 , \2260 , \2263 );
buf \U$1480 ( \2265 , \1485 );
buf \U$1481 ( \2266 , \2063 );
not \U$1482 ( \2267 , \2266 );
buf \U$1483 ( \2268 , \1548 );
not \U$1484 ( \2269 , \2268 );
or \U$1485 ( \2270 , \2267 , \2269 );
buf \U$1486 ( \2271 , \1107 );
not \U$1487 ( \2272 , \2271 );
buf \U$1488 ( \2273 , \2272 );
buf \U$1489 ( \2274 , \2273 );
not \U$1490 ( \2275 , \2274 );
buf \U$1491 ( \2276 , \2275 );
buf \U$1492 ( \2277 , \2276 );
buf \U$1493 ( \2278 , \2063 );
not \U$1494 ( \2279 , \2278 );
buf \U$1495 ( \2280 , \2279 );
buf \U$1496 ( \2281 , \2280 );
nand \U$1497 ( \2282 , \2277 , \2281 );
buf \U$1498 ( \2283 , \2282 );
buf \U$1499 ( \2284 , \2283 );
nand \U$1500 ( \2285 , \2270 , \2284 );
buf \U$1501 ( \2286 , \2285 );
buf \U$1502 ( \2287 , \2286 );
nand \U$1503 ( \2288 , \2265 , \2287 );
buf \U$1504 ( \2289 , \2288 );
buf \U$1505 ( \2290 , \2289 );
nand \U$1506 ( \2291 , \2264 , \2290 );
buf \U$1507 ( \2292 , \2291 );
buf \U$1508 ( \2293 , \2292 );
buf \U$1509 ( \2294 , \2006 );
not \U$1510 ( \2295 , \2294 );
buf \U$1513 ( \2296 , \1946 );
buf \U$1514 ( \2297 , \2296 );
not \U$1515 ( \2298 , \2297 );
or \U$1516 ( \2299 , \2295 , \2298 );
buf \U$1517 ( \2300 , \1950 );
buf \U$1518 ( \2301 , \1027 );
buf \U$1519 ( \2302 , \1619 );
xor \U$1520 ( \2303 , \2301 , \2302 );
buf \U$1521 ( \2304 , \2303 );
buf \U$1522 ( \2305 , \2304 );
nand \U$1523 ( \2306 , \2300 , \2305 );
buf \U$1524 ( \2307 , \2306 );
buf \U$1525 ( \2308 , \2307 );
nand \U$1526 ( \2309 , \2299 , \2308 );
buf \U$1527 ( \2310 , \2309 );
buf \U$1528 ( \2311 , \2310 );
xor \U$1529 ( \2312 , \2293 , \2311 );
buf \U$1530 ( \2313 , \2211 );
not \U$1531 ( \2314 , \2313 );
buf \U$1532 ( \2315 , \2201 );
not \U$1533 ( \2316 , \2315 );
buf \U$1534 ( \2317 , \2316 );
buf \U$1535 ( \2318 , \2317 );
not \U$1536 ( \2319 , \2318 );
or \U$1537 ( \2320 , \2314 , \2319 );
buf \U$1538 ( \2321 , \2067 );
nand \U$1539 ( \2322 , \2320 , \2321 );
buf \U$1540 ( \2323 , \2322 );
buf \U$1541 ( \2324 , \2323 );
xor \U$1542 ( \2325 , \2312 , \2324 );
buf \U$1543 ( \2326 , \2325 );
buf \U$1544 ( \2327 , \2326 );
xor \U$1545 ( \2328 , \2258 , \2327 );
buf \U$1546 ( \2329 , \2328 );
buf \U$1547 ( \2330 , \2329 );
xor \U$1548 ( \2331 , \1927 , \2330 );
xor \U$1549 ( \2332 , \1938 , \2013 );
xor \U$1550 ( \2333 , \2332 , \2221 );
buf \U$1551 ( \2334 , \2333 );
buf \U$1552 ( \2335 , \2334 );
not \U$1553 ( \2336 , \2335 );
buf \U$1554 ( \2337 , \1915 );
not \U$1555 ( \2338 , \2337 );
buf \U$1556 ( \2339 , \1564 );
buf \U$1557 ( \2340 , \1279 );
xor \U$1558 ( \2341 , \2339 , \2340 );
buf \U$1559 ( \2342 , \2341 );
buf \U$1560 ( \2343 , \2342 );
not \U$1561 ( \2344 , \2343 );
and \U$1562 ( \2345 , \2338 , \2344 );
buf \U$1563 ( \2346 , \1915 );
buf \U$1564 ( \2347 , \2342 );
and \U$1565 ( \2348 , \2346 , \2347 );
nor \U$1566 ( \2349 , \2345 , \2348 );
buf \U$1567 ( \2350 , \2349 );
buf \U$1568 ( \2351 , \2350 );
not \U$1569 ( \2352 , \2351 );
buf \U$1570 ( \2353 , \2352 );
buf \U$1571 ( \2354 , \2353 );
not \U$1572 ( \2355 , \2354 );
or \U$1573 ( \2356 , \2336 , \2355 );
buf \U$1574 ( \2357 , \2353 );
buf \U$1575 ( \2358 , \2334 );
or \U$1576 ( \2359 , \2357 , \2358 );
not \U$1577 ( \2360 , RI914a1d8_282);
not \U$1578 ( \2361 , \813 );
or \U$1579 ( \2362 , \2360 , \2361 );
nand \U$1580 ( \2363 , \1596 , RI9149a58_266);
nand \U$1581 ( \2364 , \2362 , \2363 );
not \U$1582 ( \2365 , RI914b0d8_314);
not \U$1583 ( \2366 , \831 );
or \U$1584 ( \2367 , \2365 , \2366 );
nand \U$1585 ( \2368 , \1053 , RI914a958_298);
nand \U$1586 ( \2369 , \2367 , \2368 );
nor \U$1587 ( \2370 , \2364 , \2369 );
not \U$1588 ( \2371 , RI914bfd8_346);
not \U$1589 ( \2372 , \1044 );
or \U$1590 ( \2373 , \2371 , \2372 );
nand \U$1591 ( \2374 , \1047 , RI914b858_330);
nand \U$1592 ( \2375 , \2373 , \2374 );
not \U$1593 ( \2376 , RI914ced8_378);
not \U$1594 ( \2377 , \1094 );
or \U$1595 ( \2378 , \2376 , \2377 );
nand \U$1596 ( \2379 , \1696 , RI914c758_362);
nand \U$1597 ( \2380 , \2378 , \2379 );
nor \U$1598 ( \2381 , \2375 , \2380 );
not \U$1599 ( \2382 , RI914f458_458);
not \U$1600 ( \2383 , \1077 );
or \U$1601 ( \2384 , \2382 , \2383 );
nand \U$1602 ( \2385 , \1080 , RI914fbd8_474);
nand \U$1603 ( \2386 , \2384 , \2385 );
not \U$1604 ( \2387 , RI914d658_394);
not \U$1605 ( \2388 , \1058 );
or \U$1606 ( \2389 , \2387 , \2388 );
nand \U$1607 ( \2390 , \1062 , RI914ddd8_410);
nand \U$1608 ( \2391 , \2389 , \2390 );
nor \U$1609 ( \2392 , \2386 , \2391 );
not \U$1610 ( \2393 , RI914e558_426);
not \U$1611 ( \2394 , \1069 );
or \U$1612 ( \2395 , \2393 , \2394 );
nand \U$1613 ( \2396 , \883 , RI914ecd8_442);
nand \U$1614 ( \2397 , \2395 , \2396 );
not \U$1615 ( \2398 , RI9150358_490);
not \U$1616 ( \2399 , \901 );
or \U$1617 ( \2400 , \2398 , \2399 );
nand \U$1618 ( \2401 , \1087 , RI9150ad8_506);
nand \U$1619 ( \2402 , \2400 , \2401 );
nor \U$1620 ( \2403 , \2397 , \2402 );
nand \U$1621 ( \2404 , \2370 , \2381 , \2392 , \2403 );
buf \U$1622 ( \2405 , \2404 );
not \U$1623 ( \2406 , \2405 );
buf \U$1624 ( \2407 , \2406 );
buf \U$1625 ( \2408 , \2407 );
not \U$1626 ( \2409 , \2408 );
buf \U$1627 ( \2410 , \2131 );
not \U$1628 ( \2411 , \2410 );
buf \U$1629 ( \2412 , \2411 );
buf \U$1630 ( \2413 , \2412 );
not \U$1631 ( \2414 , \2413 );
buf \U$1632 ( \2415 , \2414 );
buf \U$1633 ( \2416 , \2415 );
not \U$1634 ( \2417 , \2416 );
or \U$1635 ( \2418 , \2409 , \2417 );
buf \U$1636 ( \2419 , \2412 );
buf \U$1637 ( \2420 , \2404 );
nand \U$1638 ( \2421 , \2419 , \2420 );
buf \U$1639 ( \2422 , \2421 );
buf \U$1640 ( \2423 , \2422 );
nand \U$1641 ( \2424 , \2418 , \2423 );
buf \U$1642 ( \2425 , \2424 );
buf \U$1643 ( \2426 , \2425 );
and \U$1644 ( \2427 , \1358 , RI914b8d0_331);
and \U$1645 ( \2428 , \1406 , RI914c050_347);
nor \U$1646 ( \2429 , \2427 , \2428 );
and \U$1647 ( \2430 , \826 , RI914a9d0_299);
and \U$1648 ( \2431 , \831 , RI914b150_315);
nor \U$1649 ( \2432 , \2430 , \2431 );
nand \U$1650 ( \2433 , \813 , RI914a250_283);
nand \U$1651 ( \2434 , \818 , RI9149ad0_267);
and \U$1652 ( \2435 , \2433 , \2434 );
and \U$1653 ( \2436 , \1417 , RI914c7d0_363);
and \U$1654 ( \2437 , \1157 , RI914cf50_379);
nor \U$1655 ( \2438 , \2436 , \2437 );
nand \U$1656 ( \2439 , \2429 , \2432 , \2435 , \2438 );
not \U$1657 ( \2440 , \864 );
not \U$1658 ( \2441 , RI914d6d0_395);
not \U$1659 ( \2442 , \2441 );
and \U$1660 ( \2443 , \2440 , \2442 );
not \U$1661 ( \2444 , RI914de50_411);
nor \U$1662 ( \2445 , \2444 , \1061 );
nor \U$1663 ( \2446 , \2443 , \2445 );
not \U$1664 ( \2447 , \889 );
not \U$1665 ( \2448 , RI914f4d0_459);
not \U$1666 ( \2449 , \2448 );
and \U$1667 ( \2450 , \2447 , \2449 );
not \U$1668 ( \2451 , RI914fc50_475);
nor \U$1669 ( \2452 , \2451 , \1377 );
nor \U$1670 ( \2453 , \2450 , \2452 );
and \U$1671 ( \2454 , \1069 , RI914e5d0_427);
and \U$1672 ( \2455 , \883 , RI914ed50_443);
nor \U$1673 ( \2456 , \2454 , \2455 );
and \U$1674 ( \2457 , \1437 , RI91503d0_491);
and \U$1675 ( \2458 , \1087 , RI9150b50_507);
nor \U$1676 ( \2459 , \2457 , \2458 );
nand \U$1677 ( \2460 , \2446 , \2453 , \2456 , \2459 );
nor \U$1678 ( \2461 , \2439 , \2460 );
not \U$1679 ( \2462 , \2461 );
xor \U$1680 ( \2463 , \2462 , \2404 );
buf \U$1681 ( \2464 , \2463 );
not \U$1682 ( \2465 , \2464 );
buf \U$1683 ( \2466 , \2465 );
buf \U$1684 ( \2467 , \2466 );
nand \U$1685 ( \2468 , \2426 , \2467 );
buf \U$1686 ( \2469 , \2468 );
buf \U$1689 ( \2470 , \2469 );
buf \U$1690 ( \2471 , \2470 );
buf \U$1691 ( \2472 , \2463 );
buf \U$1693 ( \2473 , \2472 );
buf \U$1694 ( \2474 , \2473 );
not \U$1695 ( \2475 , \2474 );
buf \U$1696 ( \2476 , \2475 );
buf \U$1697 ( \2477 , \2476 );
and \U$1698 ( \2478 , \2471 , \2477 );
buf \U$1701 ( \2479 , \2412 );
buf \U$1702 ( \2480 , \2479 );
nor \U$1703 ( \2481 , \2478 , \2480 );
buf \U$1704 ( \2482 , \2481 );
buf \U$1705 ( \2483 , \2482 );
buf \U$1706 ( \2484 , \1542 );
not \U$1707 ( \2485 , \2484 );
buf \U$1708 ( \2486 , \2067 );
not \U$1709 ( \2487 , \2486 );
buf \U$1710 ( \2488 , \2487 );
buf \U$1711 ( \2489 , \2488 );
not \U$1712 ( \2490 , \2489 );
or \U$1713 ( \2491 , \2485 , \2490 );
buf \U$1714 ( \2492 , \2068 );
buf \U$1715 ( \2493 , \1539 );
nand \U$1716 ( \2494 , \2492 , \2493 );
buf \U$1717 ( \2495 , \2494 );
buf \U$1718 ( \2496 , \2495 );
nand \U$1719 ( \2497 , \2491 , \2496 );
buf \U$1720 ( \2498 , \2497 );
buf \U$1721 ( \2499 , \2498 );
not \U$1722 ( \2500 , \2499 );
buf \U$1726 ( \2501 , \2197 );
not \U$1727 ( \2502 , \2501 );
buf \U$1728 ( \2503 , \2502 );
buf \U$1729 ( \2504 , \2503 );
not \U$1730 ( \2505 , \2504 );
or \U$1731 ( \2506 , \2500 , \2505 );
buf \U$1732 ( \2507 , \2214 );
buf \U$1733 ( \2508 , \2084 );
nand \U$1734 ( \2509 , \2507 , \2508 );
buf \U$1735 ( \2510 , \2509 );
buf \U$1736 ( \2511 , \2510 );
nand \U$1737 ( \2512 , \2506 , \2511 );
buf \U$1738 ( \2513 , \2512 );
buf \U$1739 ( \2514 , \2513 );
not \U$1740 ( \2515 , \2514 );
buf \U$1741 ( \2516 , \2515 );
buf \U$1742 ( \2517 , \2516 );
nand \U$1743 ( \2518 , \2483 , \2517 );
buf \U$1744 ( \2519 , \2518 );
buf \U$1745 ( \2520 , \2519 );
buf \U$1746 ( \2521 , \1990 );
and \U$1747 ( \2522 , \2521 , \914 );
not \U$1748 ( \2523 , \2521 );
and \U$1749 ( \2524 , \2523 , \911 );
or \U$1750 ( \2525 , \2522 , \2524 );
buf \U$1751 ( \2526 , \2525 );
not \U$1752 ( \2527 , \2526 );
buf \U$1753 ( \2528 , \1187 );
not \U$1754 ( \2529 , \2528 );
or \U$1755 ( \2530 , \2527 , \2529 );
buf \U$1756 ( \2531 , \1194 );
buf \U$1757 ( \2532 , \1037 );
nand \U$1758 ( \2533 , \2531 , \2532 );
buf \U$1759 ( \2534 , \2533 );
buf \U$1760 ( \2535 , \2534 );
nand \U$1761 ( \2536 , \2530 , \2535 );
buf \U$1762 ( \2537 , \2536 );
buf \U$1763 ( \2538 , \2537 );
and \U$1764 ( \2539 , \2520 , \2538 );
buf \U$1765 ( \2540 , \2482 );
not \U$1766 ( \2541 , \2540 );
buf \U$1767 ( \2542 , \2541 );
buf \U$1768 ( \2543 , \2542 );
buf \U$1769 ( \2544 , \2513 );
and \U$1770 ( \2545 , \2543 , \2544 );
buf \U$1771 ( \2546 , \2545 );
buf \U$1772 ( \2547 , \2546 );
nor \U$1773 ( \2548 , \2539 , \2547 );
buf \U$1774 ( \2549 , \2548 );
buf \U$1775 ( \2550 , \2549 );
not \U$1776 ( \2551 , \2550 );
buf \U$1777 ( \2552 , \2551 );
buf \U$1778 ( \2553 , \2552 );
nand \U$1779 ( \2554 , \2359 , \2553 );
buf \U$1780 ( \2555 , \2554 );
buf \U$1781 ( \2556 , \2555 );
nand \U$1782 ( \2557 , \2356 , \2556 );
buf \U$1783 ( \2558 , \2557 );
buf \U$1784 ( \2559 , \2558 );
xnor \U$1785 ( \2560 , \2331 , \2559 );
buf \U$1786 ( \2561 , \2560 );
buf \U$1787 ( \2562 , \2561 );
buf \U$1788 ( \2563 , \1328 );
not \U$1789 ( \2564 , \2563 );
buf \U$1790 ( \2565 , \2564 );
buf \U$1791 ( \2566 , \2565 );
not \U$1792 ( \2567 , \2566 );
buf \U$1793 ( \2568 , \2567 );
buf \U$1794 ( \2569 , \2568 );
not \U$1795 ( \2570 , \2569 );
buf \U$1796 ( \2571 , \2488 );
not \U$1797 ( \2572 , \2571 );
or \U$1798 ( \2573 , \2570 , \2572 );
buf \U$1799 ( \2574 , \2068 );
buf \U$1800 ( \2575 , \2565 );
nand \U$1801 ( \2576 , \2574 , \2575 );
buf \U$1802 ( \2577 , \2576 );
buf \U$1803 ( \2578 , \2577 );
nand \U$1804 ( \2579 , \2573 , \2578 );
buf \U$1805 ( \2580 , \2579 );
buf \U$1806 ( \2581 , \2580 );
not \U$1807 ( \2582 , \2581 );
buf \U$1808 ( \2583 , \2201 );
not \U$1809 ( \2584 , \2583 );
or \U$1810 ( \2585 , \2582 , \2584 );
buf \U$1811 ( \2586 , \2498 );
buf \U$1812 ( \2587 , \2214 );
nand \U$1813 ( \2588 , \2586 , \2587 );
buf \U$1814 ( \2589 , \2588 );
buf \U$1815 ( \2590 , \2589 );
nand \U$1816 ( \2591 , \2585 , \2590 );
buf \U$1817 ( \2592 , \2591 );
buf \U$1818 ( \2593 , \2592 );
not \U$1819 ( \2594 , \2593 );
buf \U$1820 ( \2595 , \2594 );
buf \U$1821 ( \2596 , \2595 );
buf \U$1822 ( \2597 , \1672 );
buf \U$1823 ( \2598 , \1888 );
xor \U$1824 ( \2599 , \2597 , \2598 );
buf \U$1825 ( \2600 , \1911 );
xnor \U$1826 ( \2601 , \2599 , \2600 );
buf \U$1827 ( \2602 , \2601 );
buf \U$1828 ( \2603 , \2602 );
xor \U$1829 ( \2604 , \2596 , \2603 );
and \U$1830 ( \2605 , \1669 , \1800 );
not \U$1831 ( \2606 , \1669 );
and \U$1832 ( \2607 , \2606 , \1618 );
or \U$1833 ( \2608 , \2605 , \2607 );
buf \U$1834 ( \2609 , \2608 );
not \U$1835 ( \2610 , \2609 );
buf \U$1836 ( \2611 , \1946 );
not \U$1837 ( \2612 , \2611 );
or \U$1838 ( \2613 , \2610 , \2612 );
buf \U$1839 ( \2614 , \1950 );
buf \U$1840 ( \2615 , \1810 );
nand \U$1841 ( \2616 , \2614 , \2615 );
buf \U$1842 ( \2617 , \2616 );
buf \U$1843 ( \2618 , \2617 );
nand \U$1844 ( \2619 , \2613 , \2618 );
buf \U$1845 ( \2620 , \2619 );
buf \U$1846 ( \2621 , \2620 );
not \U$1847 ( \2622 , \2621 );
buf \U$1848 ( \2623 , \2622 );
buf \U$1849 ( \2624 , \2623 );
buf \U$1850 ( \2625 , \2063 );
not \U$1851 ( \2626 , \2625 );
buf \U$1854 ( \2627 , \2479 );
buf \U$1855 ( \2628 , \2627 );
not \U$1856 ( \2629 , \2628 );
or \U$1857 ( \2630 , \2626 , \2629 );
buf \U$1858 ( \2631 , \2479 );
not \U$1859 ( \2632 , \2631 );
buf \U$1860 ( \2633 , \2632 );
buf \U$1861 ( \2634 , \2633 );
buf \U$1862 ( \2635 , \2280 );
nand \U$1863 ( \2636 , \2634 , \2635 );
buf \U$1864 ( \2637 , \2636 );
buf \U$1865 ( \2638 , \2637 );
nand \U$1866 ( \2639 , \2630 , \2638 );
buf \U$1867 ( \2640 , \2639 );
buf \U$1868 ( \2641 , \2640 );
not \U$1869 ( \2642 , \2641 );
buf \U$1870 ( \2643 , \2470 );
not \U$1871 ( \2644 , \2643 );
buf \U$1872 ( \2645 , \2644 );
buf \U$1873 ( \2646 , \2645 );
not \U$1874 ( \2647 , \2646 );
or \U$1875 ( \2648 , \2642 , \2647 );
buf \U$1876 ( \2649 , \2479 );
not \U$1877 ( \2650 , \2649 );
buf \U$1878 ( \2651 , \2473 );
nand \U$1879 ( \2652 , \2650 , \2651 );
buf \U$1880 ( \2653 , \2652 );
buf \U$1881 ( \2654 , \2653 );
nand \U$1882 ( \2655 , \2648 , \2654 );
buf \U$1883 ( \2656 , \2655 );
buf \U$1884 ( \2657 , \2656 );
not \U$1885 ( \2658 , \2657 );
buf \U$1886 ( \2659 , \2658 );
buf \U$1887 ( \2660 , \2659 );
and \U$1888 ( \2661 , \2624 , \2660 );
buf \U$1889 ( \2662 , \1187 );
buf \U$1890 ( \2663 , \1868 );
not \U$1891 ( \2664 , \2663 );
buf \U$1892 ( \2665 , \1178 );
not \U$1893 ( \2666 , \2665 );
or \U$1894 ( \2667 , \2664 , \2666 );
buf \U$1895 ( \2668 , \1862 );
not \U$1896 ( \2669 , \2668 );
buf \U$1897 ( \2670 , \2669 );
buf \U$1898 ( \2671 , \2670 );
buf \U$1899 ( \2672 , \911 );
nand \U$1900 ( \2673 , \2671 , \2672 );
buf \U$1901 ( \2674 , \2673 );
buf \U$1902 ( \2675 , \2674 );
nand \U$1903 ( \2676 , \2667 , \2675 );
buf \U$1904 ( \2677 , \2676 );
buf \U$1905 ( \2678 , \2677 );
and \U$1906 ( \2679 , \2662 , \2678 );
buf \U$1907 ( \2680 , \1194 );
buf \U$1908 ( \2681 , \2525 );
and \U$1909 ( \2682 , \2680 , \2681 );
nor \U$1910 ( \2683 , \2679 , \2682 );
buf \U$1911 ( \2684 , \2683 );
buf \U$1912 ( \2685 , \2684 );
nor \U$1913 ( \2686 , \2661 , \2685 );
buf \U$1914 ( \2687 , \2686 );
buf \U$1915 ( \2688 , \2687 );
buf \U$1916 ( \2689 , \2659 );
buf \U$1917 ( \2690 , \2623 );
nor \U$1918 ( \2691 , \2689 , \2690 );
buf \U$1919 ( \2692 , \2691 );
buf \U$1920 ( \2693 , \2692 );
nor \U$1921 ( \2694 , \2688 , \2693 );
buf \U$1922 ( \2695 , \2694 );
buf \U$1923 ( \2696 , \2695 );
and \U$1924 ( \2697 , \2604 , \2696 );
and \U$1925 ( \2698 , \2596 , \2603 );
or \U$1926 ( \2699 , \2697 , \2698 );
buf \U$1927 ( \2700 , \2699 );
buf \U$1928 ( \2701 , \2700 );
xor \U$1929 ( \2702 , \2549 , \2334 );
xnor \U$1930 ( \2703 , \2702 , \2350 );
buf \U$1931 ( \2704 , \2703 );
xor \U$1932 ( \2705 , \2701 , \2704 );
buf \U$1933 ( \2706 , \2516 );
not \U$1934 ( \2707 , \2706 );
buf \U$1935 ( \2708 , \2542 );
not \U$1936 ( \2709 , \2708 );
or \U$1937 ( \2710 , \2707 , \2709 );
buf \U$1938 ( \2711 , \2513 );
buf \U$1939 ( \2712 , \2482 );
nand \U$1940 ( \2713 , \2711 , \2712 );
buf \U$1941 ( \2714 , \2713 );
buf \U$1942 ( \2715 , \2714 );
nand \U$1943 ( \2716 , \2710 , \2715 );
buf \U$1944 ( \2717 , \2716 );
buf \U$1945 ( \2718 , \2717 );
buf \U$1946 ( \2719 , \2537 );
xor \U$1947 ( \2720 , \2718 , \2719 );
buf \U$1948 ( \2721 , \2720 );
buf \U$1949 ( \2722 , \2721 );
not \U$1950 ( \2723 , \2722 );
buf \U$1951 ( \2724 , \2723 );
buf \U$1952 ( \2725 , \2724 );
not \U$1953 ( \2726 , \2725 );
nand \U$1954 ( \2727 , \951 , RI9144058_74);
nand \U$1955 ( \2728 , \1500 , RI91447d8_90);
and \U$1956 ( \2729 , \2727 , \2728 );
and \U$1957 ( \2730 , \1495 , RI90f3310_42);
and \U$1958 ( \2731 , \928 , RI91438d8_58);
nor \U$1959 ( \2732 , \2730 , \2731 );
and \U$1960 ( \2733 , \1508 , RI9144f58_106);
and \U$1961 ( \2734 , \1291 , RI91456d8_122);
nor \U$1962 ( \2735 , \2733 , \2734 );
and \U$1963 ( \2736 , \963 , RI90f9670_26);
and \U$1964 ( \2737 , \1297 , RI912eb18_10);
nor \U$1965 ( \2738 , \2736 , \2737 );
nand \U$1966 ( \2739 , \2729 , \2732 , \2735 , \2738 );
and \U$1967 ( \2740 , \1204 , RI9146d58_170);
and \U$1968 ( \2741 , \1213 , RI91474d8_186);
nor \U$1969 ( \2742 , \2740 , \2741 );
and \U$1970 ( \2743 , \1525 , RI9147c58_202);
and \U$1971 ( \2744 , \1008 , RI91483d8_218);
nor \U$1972 ( \2745 , \2743 , \2744 );
not \U$1973 ( \2746 , \976 );
not \U$1974 ( \2747 , RI9145e58_138);
not \U$1975 ( \2748 , \2747 );
and \U$1976 ( \2749 , \2746 , \2748 );
not \U$1977 ( \2750 , RI91465d8_154);
nor \U$1978 ( \2751 , \2750 , \983 );
nor \U$1979 ( \2752 , \2749 , \2751 );
and \U$1980 ( \2753 , \1014 , RI9148b58_234);
and \U$1981 ( \2754 , \1017 , RI91492d8_250);
nor \U$1982 ( \2755 , \2753 , \2754 );
nand \U$1983 ( \2756 , \2742 , \2745 , \2752 , \2755 );
nor \U$1984 ( \2757 , \2739 , \2756 );
not \U$1985 ( \2758 , \2757 );
buf \U$1986 ( \2759 , \2758 );
buf \U$1987 ( \2760 , \1619 );
nand \U$1988 ( \2761 , \2759 , \2760 );
buf \U$1989 ( \2762 , \2761 );
buf \U$1990 ( \2763 , \2762 );
buf \U$1991 ( \2764 , \2592 );
xor \U$1992 ( \2765 , \2763 , \2764 );
buf \U$1993 ( \2766 , \2261 );
buf \U$1994 ( \2767 , \1027 );
not \U$1995 ( \2768 , \2767 );
buf \U$1996 ( \2769 , \2273 );
not \U$1997 ( \2770 , \2769 );
or \U$1998 ( \2771 , \2768 , \2770 );
buf \U$1999 ( \2772 , \1024 );
buf \U$2000 ( \2773 , \1337 );
nand \U$2001 ( \2774 , \2772 , \2773 );
buf \U$2002 ( \2775 , \2774 );
buf \U$2003 ( \2776 , \2775 );
nand \U$2004 ( \2777 , \2771 , \2776 );
buf \U$2005 ( \2778 , \2777 );
buf \U$2006 ( \2779 , \2778 );
and \U$2007 ( \2780 , \2766 , \2779 );
buf \U$2008 ( \2781 , \1485 );
buf \U$2009 ( \2782 , \1896 );
and \U$2010 ( \2783 , \2781 , \2782 );
nor \U$2011 ( \2784 , \2780 , \2783 );
buf \U$2012 ( \2785 , \2784 );
buf \U$2013 ( \2786 , \2785 );
and \U$2014 ( \2787 , \2765 , \2786 );
and \U$2015 ( \2788 , \2763 , \2764 );
or \U$2016 ( \2789 , \2787 , \2788 );
buf \U$2017 ( \2790 , \2789 );
buf \U$2018 ( \2791 , \2790 );
not \U$2019 ( \2792 , \2791 );
and \U$2020 ( \2793 , \2726 , \2792 );
xor \U$2021 ( \2794 , \2596 , \2603 );
xor \U$2022 ( \2795 , \2794 , \2696 );
buf \U$2023 ( \2796 , \2795 );
not \U$2024 ( \2797 , \2796 );
buf \U$2025 ( \2798 , \2797 );
buf \U$2026 ( \2799 , \2724 );
buf \U$2027 ( \2800 , \2790 );
nand \U$2028 ( \2801 , \2799 , \2800 );
buf \U$2029 ( \2802 , \2801 );
buf \U$2030 ( \2803 , \2802 );
and \U$2031 ( \2804 , \2798 , \2803 );
nor \U$2032 ( \2805 , \2793 , \2804 );
buf \U$2033 ( \2806 , \2805 );
buf \U$2034 ( \2807 , \2806 );
and \U$2035 ( \2808 , \2705 , \2807 );
and \U$2036 ( \2809 , \2701 , \2704 );
or \U$2037 ( \2810 , \2808 , \2809 );
buf \U$2038 ( \2811 , \2810 );
buf \U$2039 ( \2812 , \2811 );
nand \U$2040 ( \2813 , \2562 , \2812 );
buf \U$2041 ( \2814 , \2813 );
buf \U$2042 ( \2815 , \2814 );
xor \U$2043 ( \2816 , \2701 , \2704 );
xor \U$2044 ( \2817 , \2816 , \2807 );
buf \U$2045 ( \2818 , \2817 );
buf \U$2046 ( \2819 , \2818 );
buf \U$2047 ( \2820 , \2790 );
not \U$2048 ( \2821 , \2820 );
buf \U$2049 ( \2822 , \2721 );
not \U$2050 ( \2823 , \2822 );
or \U$2051 ( \2824 , \2821 , \2823 );
buf \U$2052 ( \2825 , \2721 );
buf \U$2053 ( \2826 , \2790 );
or \U$2054 ( \2827 , \2825 , \2826 );
nand \U$2055 ( \2828 , \2824 , \2827 );
buf \U$2056 ( \2829 , \2828 );
not \U$2057 ( \2830 , \2829 );
buf \U$2058 ( \2831 , \2830 );
not \U$2059 ( \2832 , \2831 );
not \U$2060 ( \2833 , \2796 );
buf \U$2061 ( \2834 , \2833 );
not \U$2062 ( \2835 , \2834 );
or \U$2063 ( \2836 , \2832 , \2835 );
buf \U$2064 ( \2837 , \2796 );
buf \U$2065 ( \2838 , \2829 );
nand \U$2066 ( \2839 , \2837 , \2838 );
buf \U$2067 ( \2840 , \2839 );
buf \U$2068 ( \2841 , \2840 );
nand \U$2069 ( \2842 , \2836 , \2841 );
buf \U$2070 ( \2843 , \2842 );
not \U$2071 ( \2844 , \2843 );
buf \U$2072 ( \2845 , \2844 );
buf \U$2073 ( \2846 , \2758 );
not \U$2074 ( \2847 , \2846 );
buf \U$2075 ( \2848 , \1800 );
not \U$2076 ( \2849 , \2848 );
or \U$2077 ( \2850 , \2847 , \2849 );
buf \U$2078 ( \2851 , \2758 );
not \U$2079 ( \2852 , \2851 );
buf \U$2080 ( \2853 , \2852 );
buf \U$2081 ( \2854 , \2853 );
buf \U$2082 ( \2855 , \1618 );
nand \U$2083 ( \2856 , \2854 , \2855 );
buf \U$2084 ( \2857 , \2856 );
buf \U$2085 ( \2858 , \2857 );
nand \U$2086 ( \2859 , \2850 , \2858 );
buf \U$2087 ( \2860 , \2859 );
buf \U$2088 ( \2861 , \2860 );
not \U$2089 ( \2862 , \2861 );
buf \U$2090 ( \2863 , \1758 );
not \U$2091 ( \2864 , \2863 );
or \U$2092 ( \2865 , \2862 , \2864 );
buf \U$2093 ( \2866 , \2608 );
buf \U$2094 ( \2867 , \1882 );
nand \U$2095 ( \2868 , \2866 , \2867 );
buf \U$2096 ( \2869 , \2868 );
buf \U$2097 ( \2870 , \2869 );
nand \U$2098 ( \2871 , \2865 , \2870 );
buf \U$2099 ( \2872 , \2871 );
buf \U$2100 ( \2873 , \2872 );
buf \U$2101 ( \2874 , \1261 );
not \U$2102 ( \2875 , \2874 );
buf \U$2103 ( \2876 , \1444 );
not \U$2104 ( \2877 , \2876 );
buf \U$2105 ( \2878 , \2877 );
buf \U$2106 ( \2879 , \2878 );
not \U$2107 ( \2880 , \2879 );
or \U$2108 ( \2881 , \2875 , \2880 );
buf \U$2109 ( \2882 , \2878 );
not \U$2110 ( \2883 , \2882 );
buf \U$2111 ( \2884 , \2883 );
buf \U$2112 ( \2885 , \2884 );
buf \U$2113 ( \2886 , \1258 );
nand \U$2114 ( \2887 , \2885 , \2886 );
buf \U$2115 ( \2888 , \2887 );
buf \U$2116 ( \2889 , \2888 );
nand \U$2117 ( \2890 , \2881 , \2889 );
buf \U$2118 ( \2891 , \2890 );
buf \U$2119 ( \2892 , \2891 );
not \U$2120 ( \2893 , \2892 );
buf \U$2121 ( \2894 , \2200 );
not \U$2122 ( \2895 , \2894 );
or \U$2123 ( \2896 , \2893 , \2895 );
buf \U$2126 ( \2897 , \2208 );
buf \U$2127 ( \2898 , \2897 );
buf \U$2128 ( \2899 , \2580 );
nand \U$2129 ( \2900 , \2898 , \2899 );
buf \U$2130 ( \2901 , \2900 );
buf \U$2131 ( \2902 , \2901 );
nand \U$2132 ( \2903 , \2896 , \2902 );
buf \U$2133 ( \2904 , \2903 );
buf \U$2134 ( \2905 , \2904 );
xor \U$2135 ( \2906 , \2873 , \2905 );
buf \U$2136 ( \2907 , \1934 );
not \U$2137 ( \2908 , \2907 );
buf \U$2138 ( \2909 , \914 );
not \U$2139 ( \2910 , \2909 );
or \U$2140 ( \2911 , \2908 , \2910 );
buf \U$2141 ( \2912 , \1931 );
buf \U$2142 ( \2913 , \911 );
nand \U$2143 ( \2914 , \2912 , \2913 );
buf \U$2144 ( \2915 , \2914 );
buf \U$2145 ( \2916 , \2915 );
nand \U$2146 ( \2917 , \2911 , \2916 );
buf \U$2147 ( \2918 , \2917 );
buf \U$2148 ( \2919 , \2918 );
not \U$2149 ( \2920 , \2919 );
buf \U$2150 ( \2921 , \1186 );
not \U$2151 ( \2922 , \2921 );
or \U$2152 ( \2923 , \2920 , \2922 );
buf \U$2153 ( \2924 , \2677 );
buf \U$2154 ( \2925 , \1194 );
nand \U$2155 ( \2926 , \2924 , \2925 );
buf \U$2156 ( \2927 , \2926 );
buf \U$2157 ( \2928 , \2927 );
nand \U$2158 ( \2929 , \2923 , \2928 );
buf \U$2159 ( \2930 , \2929 );
buf \U$2160 ( \2931 , \2930 );
and \U$2161 ( \2932 , \2906 , \2931 );
and \U$2162 ( \2933 , \2873 , \2905 );
or \U$2163 ( \2934 , \2932 , \2933 );
buf \U$2164 ( \2935 , \2934 );
buf \U$2165 ( \2936 , \2935 );
buf \U$2166 ( \2937 , \2521 );
not \U$2167 ( \2938 , \2937 );
buf \U$2168 ( \2939 , \2273 );
not \U$2169 ( \2940 , \2939 );
or \U$2170 ( \2941 , \2938 , \2940 );
buf \U$2171 ( \2942 , \1337 );
buf \U$2172 ( \2943 , \1999 );
nand \U$2173 ( \2944 , \2942 , \2943 );
buf \U$2174 ( \2945 , \2944 );
buf \U$2175 ( \2946 , \2945 );
nand \U$2176 ( \2947 , \2941 , \2946 );
buf \U$2177 ( \2948 , \2947 );
buf \U$2178 ( \2949 , \2948 );
not \U$2179 ( \2950 , \2949 );
buf \U$2180 ( \2951 , \1478 );
not \U$2181 ( \2952 , \2951 );
or \U$2182 ( \2953 , \2950 , \2952 );
buf \U$2183 ( \2954 , \1485 );
buf \U$2184 ( \2955 , \2778 );
nand \U$2185 ( \2956 , \2954 , \2955 );
buf \U$2186 ( \2957 , \2956 );
buf \U$2187 ( \2958 , \2957 );
nand \U$2188 ( \2959 , \2953 , \2958 );
buf \U$2189 ( \2960 , \2959 );
buf \U$2190 ( \2961 , \2960 );
not \U$2191 ( \2962 , \2961 );
buf \U$2192 ( \2963 , \2962 );
buf \U$2193 ( \2964 , \2963 );
not \U$2194 ( \2965 , \2964 );
buf \U$2195 ( \2966 , \1542 );
not \U$2196 ( \2967 , \2966 );
buf \U$2197 ( \2968 , \2627 );
not \U$2198 ( \2969 , \2968 );
or \U$2199 ( \2970 , \2967 , \2969 );
buf \U$2200 ( \2971 , \2479 );
not \U$2201 ( \2972 , \2971 );
buf \U$2202 ( \2973 , \1539 );
nand \U$2203 ( \2974 , \2972 , \2973 );
buf \U$2204 ( \2975 , \2974 );
buf \U$2205 ( \2976 , \2975 );
nand \U$2206 ( \2977 , \2970 , \2976 );
buf \U$2207 ( \2978 , \2977 );
buf \U$2208 ( \2979 , \2978 );
not \U$2209 ( \2980 , \2979 );
buf \U$2210 ( \2981 , \2470 );
not \U$2211 ( \2982 , \2981 );
buf \U$2212 ( \2983 , \2982 );
buf \U$2213 ( \2984 , \2983 );
not \U$2214 ( \2985 , \2984 );
or \U$2215 ( \2986 , \2980 , \2985 );
buf \U$2216 ( \2987 , \2473 );
buf \U$2217 ( \2988 , \2640 );
nand \U$2218 ( \2989 , \2987 , \2988 );
buf \U$2219 ( \2990 , \2989 );
buf \U$2220 ( \2991 , \2990 );
nand \U$2221 ( \2992 , \2986 , \2991 );
buf \U$2222 ( \2993 , \2992 );
buf \U$2223 ( \2994 , \2993 );
not \U$2224 ( \2995 , \2994 );
buf \U$2225 ( \2996 , \2995 );
buf \U$2226 ( \2997 , \2996 );
not \U$2227 ( \2998 , \2997 );
or \U$2228 ( \2999 , \2965 , \2998 );
not \U$2229 ( \3000 , RI914c140_349);
not \U$2230 ( \3001 , \1044 );
or \U$2231 ( \3002 , \3000 , \3001 );
nand \U$2232 ( \3003 , \1144 , RI914b9c0_333);
nand \U$2233 ( \3004 , \3002 , \3003 );
not \U$2234 ( \3005 , RI914d040_381);
not \U$2235 ( \3006 , \1094 );
or \U$2236 ( \3007 , \3005 , \3006 );
nand \U$2237 ( \3008 , \1097 , RI914c8c0_365);
nand \U$2238 ( \3009 , \3007 , \3008 );
nor \U$2239 ( \3010 , \3004 , \3009 );
not \U$2240 ( \3011 , RI914b240_317);
not \U$2241 ( \3012 , \831 );
or \U$2242 ( \3013 , \3011 , \3012 );
nand \U$2243 ( \3014 , \1115 , RI914aac0_301);
nand \U$2244 ( \3015 , \3013 , \3014 );
not \U$2245 ( \3016 , RI914a340_285);
not \U$2246 ( \3017 , \813 );
or \U$2247 ( \3018 , \3016 , \3017 );
nand \U$2248 ( \3019 , \818 , RI9149bc0_269);
nand \U$2249 ( \3020 , \3018 , \3019 );
nor \U$2250 ( \3021 , \3015 , \3020 );
not \U$2251 ( \3022 , RI914e6c0_429);
not \U$2252 ( \3023 , \1069 );
or \U$2253 ( \3024 , \3022 , \3023 );
nand \U$2254 ( \3025 , \883 , RI914ee40_445);
nand \U$2255 ( \3026 , \3024 , \3025 );
not \U$2256 ( \3027 , RI914d7c0_397);
not \U$2257 ( \3028 , \865 );
or \U$2258 ( \3029 , \3027 , \3028 );
nand \U$2259 ( \3030 , \870 , RI914df40_413);
nand \U$2260 ( \3031 , \3029 , \3030 );
nor \U$2261 ( \3032 , \3026 , \3031 );
not \U$2262 ( \3033 , RI914f5c0_461);
not \U$2263 ( \3034 , \888 );
or \U$2264 ( \3035 , \3033 , \3034 );
nand \U$2265 ( \3036 , \1141 , RI914fd40_477);
nand \U$2266 ( \3037 , \3035 , \3036 );
not \U$2267 ( \3038 , RI91504c0_493);
not \U$2268 ( \3039 , \1437 );
or \U$2269 ( \3040 , \3038 , \3039 );
nand \U$2270 ( \3041 , \1439 , RI9150c40_509);
nand \U$2271 ( \3042 , \3040 , \3041 );
nor \U$2272 ( \3043 , \3037 , \3042 );
nand \U$2273 ( \3044 , \3010 , \3021 , \3032 , \3043 );
not \U$2274 ( \3045 , RI914cfc8_380);
not \U$2275 ( \3046 , \1094 );
or \U$2276 ( \3047 , \3045 , \3046 );
nand \U$2277 ( \3048 , \1097 , RI914c848_364);
nand \U$2278 ( \3049 , \3047 , \3048 );
not \U$2279 ( \3050 , RI914c0c8_348);
not \U$2280 ( \3051 , \1044 );
or \U$2281 ( \3052 , \3050 , \3051 );
nand \U$2282 ( \3053 , \1144 , RI914b948_332);
nand \U$2283 ( \3054 , \3052 , \3053 );
nor \U$2284 ( \3055 , \3049 , \3054 );
not \U$2285 ( \3056 , RI914a2c8_284);
not \U$2286 ( \3057 , \813 );
or \U$2287 ( \3058 , \3056 , \3057 );
nand \U$2288 ( \3059 , \818 , RI9149b48_268);
nand \U$2289 ( \3060 , \3058 , \3059 );
not \U$2290 ( \3061 , RI914b1c8_316);
not \U$2291 ( \3062 , \831 );
or \U$2292 ( \3063 , \3061 , \3062 );
nand \U$2293 ( \3064 , \1115 , RI914aa48_300);
nand \U$2294 ( \3065 , \3063 , \3064 );
nor \U$2295 ( \3066 , \3060 , \3065 );
not \U$2296 ( \3067 , RI914d748_396);
not \U$2297 ( \3068 , \865 );
or \U$2298 ( \3069 , \3067 , \3068 );
not \U$2299 ( \3070 , \869 );
nand \U$2300 ( \3071 , \3070 , RI914dec8_412);
nand \U$2301 ( \3072 , \3069 , \3071 );
not \U$2302 ( \3073 , RI914e648_428);
not \U$2303 ( \3074 , \1069 );
or \U$2304 ( \3075 , \3073 , \3074 );
nand \U$2305 ( \3076 , \883 , RI914edc8_444);
nand \U$2306 ( \3077 , \3075 , \3076 );
nor \U$2307 ( \3078 , \3072 , \3077 );
not \U$2308 ( \3079 , RI914f548_460);
not \U$2309 ( \3080 , \888 );
or \U$2310 ( \3081 , \3079 , \3080 );
nand \U$2311 ( \3082 , \1141 , RI914fcc8_476);
nand \U$2312 ( \3083 , \3081 , \3082 );
not \U$2313 ( \3084 , RI9150448_492);
not \U$2314 ( \3085 , \1437 );
or \U$2315 ( \3086 , \3084 , \3085 );
nand \U$2316 ( \3087 , \1439 , RI9150bc8_508);
nand \U$2317 ( \3088 , \3086 , \3087 );
nor \U$2318 ( \3089 , \3083 , \3088 );
nand \U$2319 ( \3090 , \3055 , \3066 , \3078 , \3089 );
xnor \U$2320 ( \3091 , \3044 , \3090 );
buf \U$2321 ( \3092 , \3091 );
not \U$2322 ( \3093 , \3092 );
buf \U$2323 ( \3094 , \3093 );
buf \U$2326 ( \3095 , \3094 );
buf \U$2327 ( \3096 , \3095 );
not \U$2328 ( \3097 , \3096 );
buf \U$2329 ( \3098 , \3097 );
buf \U$2330 ( \3099 , \3098 );
not \U$2331 ( \3100 , \3099 );
buf \U$2332 ( \3101 , \3091 );
nand \U$2333 ( \3102 , \3055 , \3066 , \3078 , \3089 );
buf \U$2334 ( \3103 , \3102 );
not \U$2335 ( \3104 , \3103 );
buf \U$2336 ( \3105 , \2462 );
not \U$2337 ( \3106 , \3105 );
buf \U$2338 ( \3107 , \3106 );
buf \U$2339 ( \3108 , \3107 );
not \U$2340 ( \3109 , \3108 );
or \U$2341 ( \3110 , \3104 , \3109 );
buf \U$2342 ( \3111 , \3107 );
not \U$2343 ( \3112 , \3111 );
buf \U$2344 ( \3113 , \3102 );
not \U$2345 ( \3114 , \3113 );
buf \U$2346 ( \3115 , \3114 );
buf \U$2347 ( \3116 , \3115 );
nand \U$2348 ( \3117 , \3112 , \3116 );
buf \U$2349 ( \3118 , \3117 );
buf \U$2350 ( \3119 , \3118 );
nand \U$2351 ( \3120 , \3110 , \3119 );
buf \U$2352 ( \3121 , \3120 );
buf \U$2353 ( \3122 , \3121 );
nand \U$2354 ( \3123 , \3101 , \3122 );
buf \U$2355 ( \3124 , \3123 );
buf \U$2356 ( \3125 , \3124 );
not \U$2357 ( \3126 , \3125 );
or \U$2358 ( \3127 , \3100 , \3126 );
buf \U$2359 ( \3128 , \2462 );
not \U$2360 ( \3129 , \3128 );
buf \U$2361 ( \3130 , \3129 );
buf \U$2362 ( \3131 , \3130 );
not \U$2363 ( \3132 , \3131 );
buf \U$2364 ( \3133 , \3132 );
buf \U$2367 ( \3134 , \3133 );
buf \U$2368 ( \3135 , \3134 );
nand \U$2369 ( \3136 , \3127 , \3135 );
buf \U$2370 ( \3137 , \3136 );
buf \U$2371 ( \3138 , \3137 );
nand \U$2372 ( \3139 , \2999 , \3138 );
buf \U$2373 ( \3140 , \3139 );
buf \U$2374 ( \3141 , \3140 );
buf \U$2375 ( \3142 , \2996 );
not \U$2376 ( \3143 , \3142 );
buf \U$2377 ( \3144 , \2960 );
nand \U$2378 ( \3145 , \3143 , \3144 );
buf \U$2379 ( \3146 , \3145 );
buf \U$2380 ( \3147 , \3146 );
nand \U$2381 ( \3148 , \3141 , \3147 );
buf \U$2382 ( \3149 , \3148 );
buf \U$2383 ( \3150 , \3149 );
xor \U$2384 ( \3151 , \2936 , \3150 );
buf \U$2385 ( \3152 , \2684 );
not \U$2386 ( \3153 , \3152 );
buf \U$2387 ( \3154 , \3153 );
buf \U$2388 ( \3155 , \3154 );
not \U$2389 ( \3156 , \3155 );
buf \U$2390 ( \3157 , \2656 );
buf \U$2391 ( \3158 , \2623 );
and \U$2392 ( \3159 , \3157 , \3158 );
not \U$2393 ( \3160 , \3157 );
buf \U$2394 ( \3161 , \2620 );
and \U$2395 ( \3162 , \3160 , \3161 );
nor \U$2396 ( \3163 , \3159 , \3162 );
buf \U$2397 ( \3164 , \3163 );
buf \U$2398 ( \3165 , \3164 );
not \U$2399 ( \3166 , \3165 );
or \U$2400 ( \3167 , \3156 , \3166 );
buf \U$2401 ( \3168 , \3164 );
buf \U$2402 ( \3169 , \3154 );
or \U$2403 ( \3170 , \3168 , \3169 );
nand \U$2404 ( \3171 , \3167 , \3170 );
buf \U$2405 ( \3172 , \3171 );
buf \U$2406 ( \3173 , \3172 );
and \U$2407 ( \3174 , \3151 , \3173 );
and \U$2408 ( \3175 , \2936 , \3150 );
or \U$2409 ( \3176 , \3174 , \3175 );
buf \U$2410 ( \3177 , \3176 );
buf \U$2411 ( \3178 , \3177 );
not \U$2412 ( \3179 , \3178 );
buf \U$2413 ( \3180 , \3179 );
buf \U$2414 ( \3181 , \3180 );
nand \U$2415 ( \3182 , \2845 , \3181 );
buf \U$2416 ( \3183 , \3182 );
buf \U$2417 ( \3184 , \3183 );
not \U$2418 ( \3185 , RI9145ed0_139);
nor \U$2419 ( \3186 , \3185 , \976 );
not \U$2420 ( \3187 , RI9146650_155);
nor \U$2421 ( \3188 , \3187 , \983 );
nor \U$2422 ( \3189 , \3186 , \3188 );
not \U$2423 ( \3190 , RI9146dd0_171);
nor \U$2424 ( \3191 , \3190 , \989 );
not \U$2425 ( \3192 , RI9147550_187);
nor \U$2426 ( \3193 , \3192 , \994 );
nor \U$2427 ( \3194 , \3191 , \3193 );
nand \U$2428 ( \3195 , \3189 , \3194 );
not \U$2429 ( \3196 , RI9147cd0_203);
nor \U$2430 ( \3197 , \3196 , \1524 );
not \U$2431 ( \3198 , RI9148450_219);
nor \U$2432 ( \3199 , \3198 , \1199 );
nor \U$2433 ( \3200 , \3197 , \3199 );
and \U$2434 ( \3201 , \1014 , RI9148bd0_235);
not \U$2435 ( \3202 , RI9149350_251);
nor \U$2436 ( \3203 , \3202 , \1857 );
nor \U$2437 ( \3204 , \3201 , \3203 );
nand \U$2438 ( \3205 , \3200 , \3204 );
nor \U$2439 ( \3206 , \3195 , \3205 );
not \U$2440 ( \3207 , RI9144850_91);
nor \U$2441 ( \3208 , \3207 , \957 );
not \U$2442 ( \3209 , \3208 );
not \U$2443 ( \3210 , \2031 );
nand \U$2444 ( \3211 , \3210 , RI91440d0_75);
and \U$2445 ( \3212 , \963 , RI90f95f8_27);
and \U$2446 ( \3213 , \968 , RI912eaa0_11);
nor \U$2447 ( \3214 , \3212 , \3213 );
nand \U$2448 ( \3215 , \3209 , \3211 , \3214 );
nand \U$2449 ( \3216 , \1302 , RI90f3298_43);
nand \U$2450 ( \3217 , \928 , RI9143950_59);
nand \U$2451 ( \3218 , \1291 , RI9145750_123);
nand \U$2452 ( \3219 , \943 , RI9144fd0_107);
nand \U$2453 ( \3220 , \3216 , \3217 , \3218 , \3219 );
nor \U$2454 ( \3221 , \3215 , \3220 );
nand \U$2455 ( \3222 , \3206 , \3221 );
buf \U$2456 ( \3223 , \3222 );
buf \U$2457 ( \3224 , \3223 );
not \U$2458 ( \3225 , \3224 );
buf \U$2459 ( \3226 , \1995 );
nor \U$2460 ( \3227 , \3225 , \3226 );
buf \U$2461 ( \3228 , \3227 );
buf \U$2462 ( \3229 , \3228 );
not \U$2463 ( \3230 , \3229 );
buf \U$2464 ( \3231 , \2061 );
not \U$2465 ( \3232 , \3231 );
buf \U$2466 ( \3233 , \3130 );
not \U$2467 ( \3234 , \3233 );
or \U$2468 ( \3235 , \3232 , \3234 );
buf \U$2469 ( \3236 , \2061 );
not \U$2470 ( \3237 , \3236 );
buf \U$2471 ( \3238 , \3133 );
nand \U$2472 ( \3239 , \3237 , \3238 );
buf \U$2473 ( \3240 , \3239 );
buf \U$2474 ( \3241 , \3240 );
nand \U$2475 ( \3242 , \3235 , \3241 );
buf \U$2476 ( \3243 , \3242 );
buf \U$2477 ( \3244 , \3243 );
not \U$2478 ( \3245 , \3244 );
buf \U$2479 ( \3246 , \3121 );
buf \U$2480 ( \3247 , \3091 );
nand \U$2481 ( \3248 , \3246 , \3247 );
buf \U$2482 ( \3249 , \3248 );
not \U$2483 ( \3250 , \3249 );
buf \U$2484 ( \3251 , \3250 );
not \U$2485 ( \3252 , \3251 );
or \U$2486 ( \3253 , \3245 , \3252 );
buf \U$2487 ( \3254 , \3095 );
buf \U$2488 ( \3255 , \3134 );
nand \U$2489 ( \3256 , \3254 , \3255 );
buf \U$2490 ( \3257 , \3256 );
buf \U$2491 ( \3258 , \3257 );
nand \U$2492 ( \3259 , \3253 , \3258 );
buf \U$2493 ( \3260 , \3259 );
buf \U$2494 ( \3261 , \3260 );
not \U$2495 ( \3262 , \3261 );
buf \U$2496 ( \3263 , \3262 );
buf \U$2497 ( \3264 , \3263 );
nand \U$2498 ( \3265 , \3230 , \3264 );
buf \U$2499 ( \3266 , \3265 );
buf \U$2500 ( \3267 , \3266 );
not \U$2501 ( \3268 , \3267 );
buf \U$2502 ( \3269 , \2568 );
not \U$2503 ( \3270 , \3269 );
buf \U$2504 ( \3271 , \2479 );
not \U$2505 ( \3272 , \3271 );
or \U$2506 ( \3273 , \3270 , \3272 );
buf \U$2507 ( \3274 , \2479 );
not \U$2508 ( \3275 , \3274 );
buf \U$2509 ( \3276 , \3275 );
buf \U$2510 ( \3277 , \3276 );
buf \U$2511 ( \3278 , \1331 );
nand \U$2512 ( \3279 , \3277 , \3278 );
buf \U$2513 ( \3280 , \3279 );
buf \U$2514 ( \3281 , \3280 );
nand \U$2515 ( \3282 , \3273 , \3281 );
buf \U$2516 ( \3283 , \3282 );
buf \U$2517 ( \3284 , \3283 );
not \U$2518 ( \3285 , \3284 );
buf \U$2519 ( \3286 , \2469 );
not \U$2520 ( \3287 , \3286 );
buf \U$2521 ( \3288 , \3287 );
buf \U$2522 ( \3289 , \3288 );
not \U$2523 ( \3290 , \3289 );
or \U$2524 ( \3291 , \3285 , \3290 );
buf \U$2525 ( \3292 , \2473 );
buf \U$2526 ( \3293 , \2978 );
nand \U$2527 ( \3294 , \3292 , \3293 );
buf \U$2528 ( \3295 , \3294 );
buf \U$2529 ( \3296 , \3295 );
nand \U$2530 ( \3297 , \3291 , \3296 );
buf \U$2531 ( \3298 , \3297 );
buf \U$2532 ( \3299 , \1337 );
not \U$2533 ( \3300 , \3299 );
buf \U$2534 ( \3301 , \2670 );
not \U$2535 ( \3302 , \3301 );
and \U$2536 ( \3303 , \3300 , \3302 );
buf \U$2537 ( \3304 , \1337 );
buf \U$2538 ( \3305 , \1865 );
and \U$2539 ( \3306 , \3304 , \3305 );
nor \U$2540 ( \3307 , \3303 , \3306 );
buf \U$2541 ( \3308 , \3307 );
buf \U$2542 ( \3309 , \3308 );
not \U$2543 ( \3310 , \3309 );
buf \U$2544 ( \3311 , \3310 );
buf \U$2545 ( \3312 , \3311 );
not \U$2546 ( \3313 , \3312 );
buf \U$2547 ( \3314 , \1472 );
not \U$2548 ( \3315 , \3314 );
or \U$2549 ( \3316 , \3313 , \3315 );
buf \U$2550 ( \3317 , \1485 );
buf \U$2551 ( \3318 , \2948 );
nand \U$2552 ( \3319 , \3317 , \3318 );
buf \U$2553 ( \3320 , \3319 );
buf \U$2554 ( \3321 , \3320 );
nand \U$2555 ( \3322 , \3316 , \3321 );
buf \U$2556 ( \3323 , \3322 );
or \U$2557 ( \3324 , \3298 , \3323 );
and \U$2558 ( \3325 , \1669 , \1178 );
not \U$2559 ( \3326 , \1669 );
buf \U$2560 ( \3327 , \1178 );
not \U$2561 ( \3328 , \3327 );
buf \U$2562 ( \3329 , \3328 );
and \U$2563 ( \3330 , \3326 , \3329 );
or \U$2564 ( \3331 , \3325 , \3330 );
buf \U$2565 ( \3332 , \3331 );
not \U$2566 ( \3333 , \3332 );
buf \U$2567 ( \3334 , \1187 );
not \U$2568 ( \3335 , \3334 );
or \U$2569 ( \3336 , \3333 , \3335 );
buf \U$2570 ( \3337 , \1194 );
buf \U$2571 ( \3338 , \2918 );
nand \U$2572 ( \3339 , \3337 , \3338 );
buf \U$2573 ( \3340 , \3339 );
buf \U$2574 ( \3341 , \3340 );
nand \U$2575 ( \3342 , \3336 , \3341 );
buf \U$2576 ( \3343 , \3342 );
nand \U$2577 ( \3344 , \3324 , \3343 );
buf \U$2578 ( \3345 , \3323 );
buf \U$2579 ( \3346 , \3298 );
nand \U$2580 ( \3347 , \3345 , \3346 );
buf \U$2581 ( \3348 , \3347 );
nand \U$2582 ( \3349 , \3344 , \3348 );
buf \U$2583 ( \3350 , \3349 );
not \U$2584 ( \3351 , \3350 );
or \U$2585 ( \3352 , \3268 , \3351 );
buf \U$2586 ( \3353 , \3260 );
buf \U$2587 ( \3354 , \3228 );
nand \U$2588 ( \3355 , \3353 , \3354 );
buf \U$2589 ( \3356 , \3355 );
buf \U$2590 ( \3357 , \3356 );
nand \U$2591 ( \3358 , \3352 , \3357 );
buf \U$2592 ( \3359 , \3358 );
buf \U$2593 ( \3360 , \3359 );
not \U$2594 ( \3361 , \3360 );
xor \U$2595 ( \3362 , \2763 , \2764 );
xor \U$2596 ( \3363 , \3362 , \2786 );
buf \U$2597 ( \3364 , \3363 );
buf \U$2598 ( \3365 , \3364 );
nand \U$2599 ( \3366 , \3361 , \3365 );
buf \U$2600 ( \3367 , \3366 );
buf \U$2601 ( \3368 , \3367 );
not \U$2602 ( \3369 , \3368 );
buf \U$2603 ( \3370 , \3137 );
not \U$2604 ( \3371 , \3370 );
buf \U$2605 ( \3372 , \2996 );
not \U$2606 ( \3373 , \3372 );
or \U$2607 ( \3374 , \3371 , \3373 );
buf \U$2608 ( \3375 , \3137 );
not \U$2609 ( \3376 , \3375 );
buf \U$2610 ( \3377 , \2993 );
nand \U$2611 ( \3378 , \3376 , \3377 );
buf \U$2612 ( \3379 , \3378 );
buf \U$2613 ( \3380 , \3379 );
nand \U$2614 ( \3381 , \3374 , \3380 );
buf \U$2615 ( \3382 , \3381 );
buf \U$2616 ( \3383 , \3382 );
buf \U$2617 ( \3384 , \2963 );
and \U$2618 ( \3385 , \3383 , \3384 );
not \U$2619 ( \3386 , \3383 );
buf \U$2620 ( \3387 , \2960 );
and \U$2621 ( \3388 , \3386 , \3387 );
nor \U$2622 ( \3389 , \3385 , \3388 );
buf \U$2623 ( \3390 , \3389 );
buf \U$2624 ( \3391 , \3390 );
not \U$2625 ( \3392 , \2214 );
not \U$2626 ( \3393 , \2891 );
or \U$2627 ( \3394 , \3392 , \3393 );
buf \U$2628 ( \3395 , \1021 );
buf \U$2629 ( \3396 , \2488 );
and \U$2630 ( \3397 , \3395 , \3396 );
not \U$2631 ( \3398 , \3395 );
buf \U$2632 ( \3399 , \2067 );
and \U$2633 ( \3400 , \3398 , \3399 );
nor \U$2634 ( \3401 , \3397 , \3400 );
buf \U$2635 ( \3402 , \3401 );
not \U$2636 ( \3403 , \3402 );
nand \U$2637 ( \3404 , \3403 , \2200 );
nand \U$2638 ( \3405 , \3394 , \3404 );
buf \U$2639 ( \3406 , \3405 );
not \U$2640 ( \3407 , \3406 );
buf \U$2641 ( \3408 , \1619 );
and \U$2642 ( \3409 , \1525 , RI9147d48_204);
and \U$2643 ( \3410 , \1200 , RI91484c8_220);
nor \U$2644 ( \3411 , \3409 , \3410 );
not \U$2645 ( \3412 , RI9145f48_140);
nor \U$2646 ( \3413 , \3412 , \976 );
not \U$2647 ( \3414 , RI91466c8_156);
nor \U$2648 ( \3415 , \3414 , \983 );
nor \U$2649 ( \3416 , \3413 , \3415 );
nand \U$2650 ( \3417 , \3411 , \3416 );
nand \U$2651 ( \3418 , \1014 , RI9148c48_236);
nand \U$2652 ( \3419 , \1213 , RI91475c8_188);
nand \U$2653 ( \3420 , \1206 , RI9146e48_172);
nand \U$2654 ( \3421 , \1017 , RI91493c8_252);
nand \U$2655 ( \3422 , \3418 , \3419 , \3420 , \3421 );
nor \U$2656 ( \3423 , \3417 , \3422 );
not \U$2657 ( \3424 , RI9144148_76);
nor \U$2658 ( \3425 , \3424 , \2031 );
not \U$2659 ( \3426 , RI91448c8_92);
nor \U$2660 ( \3427 , \3426 , \957 );
nor \U$2661 ( \3428 , \3425 , \3427 );
not \U$2662 ( \3429 , \929 );
not \U$2663 ( \3430 , RI91439c8_60);
not \U$2664 ( \3431 , \3430 );
and \U$2665 ( \3432 , \3429 , \3431 );
not \U$2666 ( \3433 , RI9143248_44);
nor \U$2667 ( \3434 , \3433 , \1301 );
nor \U$2668 ( \3435 , \3432 , \3434 );
nand \U$2669 ( \3436 , \3428 , \3435 );
nand \U$2670 ( \3437 , \1508 , RI9145048_108);
nand \U$2671 ( \3438 , \968 , RI912ea28_12);
nand \U$2672 ( \3439 , \1291 , RI91457c8_124);
nand \U$2673 ( \3440 , \963 , RI90f39a0_28);
nand \U$2674 ( \3441 , \3437 , \3438 , \3439 , \3440 );
nor \U$2675 ( \3442 , \3436 , \3441 );
nand \U$2676 ( \3443 , \3423 , \3442 );
buf \U$2677 ( \3444 , \3443 );
buf \U$2678 ( \3445 , \3444 );
and \U$2679 ( \3446 , \3408 , \3445 );
buf \U$2680 ( \3447 , \3446 );
buf \U$2681 ( \3448 , \3447 );
not \U$2682 ( \3449 , \3448 );
buf \U$2683 ( \3450 , \3449 );
buf \U$2684 ( \3451 , \3450 );
nand \U$2685 ( \3452 , \3407 , \3451 );
buf \U$2686 ( \3453 , \3452 );
buf \U$2687 ( \3454 , \3453 );
buf \U$2688 ( \3455 , \1618 );
not \U$2689 ( \3456 , \3455 );
buf \U$2690 ( \3457 , \3223 );
not \U$2691 ( \3458 , \3457 );
buf \U$2692 ( \3459 , \3458 );
buf \U$2693 ( \3460 , \3459 );
not \U$2694 ( \3461 , \3460 );
or \U$2695 ( \3462 , \3456 , \3461 );
buf \U$2696 ( \3463 , \1618 );
not \U$2697 ( \3464 , \3463 );
buf \U$2698 ( \3465 , \3464 );
buf \U$2699 ( \3466 , \3465 );
buf \U$2700 ( \3467 , \3223 );
nand \U$2701 ( \3468 , \3466 , \3467 );
buf \U$2702 ( \3469 , \3468 );
buf \U$2703 ( \3470 , \3469 );
nand \U$2704 ( \3471 , \3462 , \3470 );
buf \U$2705 ( \3472 , \3471 );
buf \U$2706 ( \3473 , \3472 );
not \U$2707 ( \3474 , \3473 );
buf \U$2708 ( \3475 , \1946 );
not \U$2709 ( \3476 , \3475 );
or \U$2710 ( \3477 , \3474 , \3476 );
buf \U$2711 ( \3478 , \1950 );
buf \U$2712 ( \3479 , \2860 );
nand \U$2713 ( \3480 , \3478 , \3479 );
buf \U$2714 ( \3481 , \3480 );
buf \U$2715 ( \3482 , \3481 );
nand \U$2716 ( \3483 , \3477 , \3482 );
buf \U$2717 ( \3484 , \3483 );
buf \U$2718 ( \3485 , \3484 );
and \U$2719 ( \3486 , \3454 , \3485 );
buf \U$2720 ( \3487 , \3405 );
buf \U$2721 ( \3488 , \3447 );
and \U$2722 ( \3489 , \3487 , \3488 );
buf \U$2723 ( \3490 , \3489 );
buf \U$2724 ( \3491 , \3490 );
nor \U$2725 ( \3492 , \3486 , \3491 );
buf \U$2726 ( \3493 , \3492 );
buf \U$2727 ( \3494 , \3493 );
buf \U$2728 ( \3495 , \3494 );
nand \U$2729 ( \3496 , \3391 , \3495 );
buf \U$2730 ( \3497 , \3496 );
buf \U$2731 ( \3498 , \3497 );
xor \U$2732 ( \3499 , \2873 , \2905 );
xor \U$2733 ( \3500 , \3499 , \2931 );
buf \U$2734 ( \3501 , \3500 );
buf \U$2738 ( \3502 , \3501 );
and \U$2739 ( \3503 , \3498 , \3502 );
buf \U$2740 ( \3504 , \3390 );
buf \U$2741 ( \3505 , \3494 );
nor \U$2742 ( \3506 , \3504 , \3505 );
buf \U$2743 ( \3507 , \3506 );
buf \U$2744 ( \3508 , \3507 );
nor \U$2745 ( \3509 , \3503 , \3508 );
buf \U$2746 ( \3510 , \3509 );
not \U$2747 ( \3511 , \3510 );
buf \U$2748 ( \3512 , \3511 );
not \U$2749 ( \3513 , \3512 );
or \U$2750 ( \3514 , \3369 , \3513 );
buf \U$2751 ( \3515 , \3364 );
not \U$2752 ( \3516 , \3515 );
buf \U$2753 ( \3517 , \3359 );
nand \U$2754 ( \3518 , \3516 , \3517 );
buf \U$2755 ( \3519 , \3518 );
buf \U$2756 ( \3520 , \3519 );
nand \U$2757 ( \3521 , \3514 , \3520 );
buf \U$2758 ( \3522 , \3521 );
buf \U$2759 ( \3523 , \3522 );
and \U$2760 ( \3524 , \3184 , \3523 );
buf \U$2761 ( \3525 , \2844 );
buf \U$2762 ( \3526 , \3180 );
nor \U$2763 ( \3527 , \3525 , \3526 );
buf \U$2764 ( \3528 , \3527 );
buf \U$2765 ( \3529 , \3528 );
nor \U$2766 ( \3530 , \3524 , \3529 );
buf \U$2767 ( \3531 , \3530 );
buf \U$2768 ( \3532 , \3531 );
nand \U$2769 ( \3533 , \2819 , \3532 );
buf \U$2770 ( \3534 , \3533 );
buf \U$2771 ( \3535 , \3534 );
nand \U$2772 ( \3536 , \2815 , \3535 );
buf \U$2773 ( \3537 , \3536 );
buf \U$2774 ( \3538 , \3537 );
or \U$2775 ( \3539 , \2329 , \1926 );
nand \U$2776 ( \3540 , \3539 , \2558 );
buf \U$2777 ( \3541 , \3540 );
buf \U$2778 ( \3542 , \2329 );
buf \U$2779 ( \3543 , \1926 );
nand \U$2780 ( \3544 , \3542 , \3543 );
buf \U$2781 ( \3545 , \3544 );
buf \U$2782 ( \3546 , \3545 );
nand \U$2783 ( \3547 , \3541 , \3546 );
buf \U$2784 ( \3548 , \3547 );
buf \U$2785 ( \3549 , \3548 );
xor \U$2786 ( \3550 , \2231 , \2232 );
and \U$2787 ( \3551 , \3550 , \2254 );
and \U$2788 ( \3552 , \2231 , \2232 );
or \U$2789 ( \3553 , \3551 , \3552 );
buf \U$2790 ( \3554 , \3553 );
buf \U$2791 ( \3555 , \3554 );
xor \U$2792 ( \3556 , \2226 , \2257 );
and \U$2793 ( \3557 , \3556 , \2327 );
and \U$2794 ( \3558 , \2226 , \2257 );
or \U$2795 ( \3559 , \3557 , \3558 );
buf \U$2796 ( \3560 , \3559 );
buf \U$2797 ( \3561 , \3560 );
xor \U$2798 ( \3562 , \3555 , \3561 );
buf \U$2799 ( \3563 , \2261 );
not \U$2800 ( \3564 , \3563 );
buf \U$2801 ( \3565 , \3564 );
buf \U$2802 ( \3566 , \3565 );
buf \U$2803 ( \3567 , \2286 );
not \U$2804 ( \3568 , \3567 );
buf \U$2805 ( \3569 , \3568 );
buf \U$2806 ( \3570 , \3569 );
or \U$2807 ( \3571 , \3566 , \3570 );
buf \U$2808 ( \3572 , \1485 );
not \U$2809 ( \3573 , \3572 );
buf \U$2810 ( \3574 , \3573 );
buf \U$2811 ( \3575 , \3574 );
buf \U$2812 ( \3576 , \1548 );
or \U$2813 ( \3577 , \3575 , \3576 );
nand \U$2814 ( \3578 , \3571 , \3577 );
buf \U$2815 ( \3579 , \3578 );
buf \U$2816 ( \3580 , \3579 );
not \U$2817 ( \3581 , \3580 );
buf \U$2818 ( \3582 , \3581 );
buf \U$2819 ( \3583 , \3582 );
buf \U$2820 ( \3584 , \1619 );
buf \U$2821 ( \3585 , \1990 );
and \U$2822 ( \3586 , \3584 , \3585 );
buf \U$2823 ( \3587 , \3586 );
buf \U$2824 ( \3588 , \3587 );
buf \U$2825 ( \3589 , \2304 );
not \U$2826 ( \3590 , \3589 );
buf \U$2827 ( \3591 , \2296 );
not \U$2828 ( \3592 , \3591 );
or \U$2829 ( \3593 , \3590 , \3592 );
buf \U$2830 ( \3594 , \1950 );
buf \U$2831 ( \3595 , \1261 );
buf \U$2832 ( \3596 , \1619 );
xor \U$2833 ( \3597 , \3595 , \3596 );
buf \U$2834 ( \3598 , \3597 );
buf \U$2835 ( \3599 , \3598 );
nand \U$2836 ( \3600 , \3594 , \3599 );
buf \U$2837 ( \3601 , \3600 );
buf \U$2838 ( \3602 , \3601 );
nand \U$2839 ( \3603 , \3593 , \3602 );
buf \U$2840 ( \3604 , \3603 );
buf \U$2841 ( \3605 , \3604 );
xor \U$2842 ( \3606 , \3588 , \3605 );
buf \U$2843 ( \3607 , \2247 );
not \U$2844 ( \3608 , \3607 );
buf \U$2845 ( \3609 , \1187 );
not \U$2846 ( \3610 , \3609 );
or \U$2847 ( \3611 , \3608 , \3610 );
buf \U$2848 ( \3612 , \1194 );
buf \U$2849 ( \3613 , \1542 );
buf \U$2850 ( \3614 , \911 );
and \U$2851 ( \3615 , \3613 , \3614 );
not \U$2852 ( \3616 , \3613 );
buf \U$2853 ( \3617 , \914 );
and \U$2854 ( \3618 , \3616 , \3617 );
nor \U$2855 ( \3619 , \3615 , \3618 );
buf \U$2856 ( \3620 , \3619 );
buf \U$2857 ( \3621 , \3620 );
nand \U$2858 ( \3622 , \3612 , \3621 );
buf \U$2859 ( \3623 , \3622 );
buf \U$2860 ( \3624 , \3623 );
nand \U$2861 ( \3625 , \3611 , \3624 );
buf \U$2862 ( \3626 , \3625 );
buf \U$2863 ( \3627 , \3626 );
xor \U$2864 ( \3628 , \3606 , \3627 );
buf \U$2865 ( \3629 , \3628 );
buf \U$2866 ( \3630 , \3629 );
xor \U$2867 ( \3631 , \3583 , \3630 );
xor \U$2868 ( \3632 , \2293 , \2311 );
and \U$2869 ( \3633 , \3632 , \2324 );
and \U$2870 ( \3634 , \2293 , \2311 );
or \U$2871 ( \3635 , \3633 , \3634 );
buf \U$2872 ( \3636 , \3635 );
buf \U$2873 ( \3637 , \3636 );
xor \U$2874 ( \3638 , \3631 , \3637 );
buf \U$2875 ( \3639 , \3638 );
buf \U$2876 ( \3640 , \3639 );
xor \U$2877 ( \3641 , \3562 , \3640 );
buf \U$2878 ( \3642 , \3641 );
buf \U$2879 ( \3643 , \3642 );
nor \U$2880 ( \3644 , \3549 , \3643 );
buf \U$2881 ( \3645 , \3644 );
buf \U$2882 ( \3646 , \3645 );
nor \U$2883 ( \3647 , \3538 , \3646 );
buf \U$2884 ( \3648 , \3647 );
buf \U$2885 ( \3649 , \3648 );
and \U$2886 ( \3650 , \2301 , \2302 );
buf \U$2887 ( \3651 , \3650 );
buf \U$2888 ( \3652 , \3651 );
buf \U$2889 ( \3653 , \3574 );
not \U$2890 ( \3654 , \3653 );
buf \U$2891 ( \3655 , \3565 );
not \U$2892 ( \3656 , \3655 );
or \U$2893 ( \3657 , \3654 , \3656 );
buf \U$2894 ( \3658 , \1548 );
not \U$2895 ( \3659 , \3658 );
buf \U$2896 ( \3660 , \3659 );
buf \U$2897 ( \3661 , \3660 );
nand \U$2898 ( \3662 , \3657 , \3661 );
buf \U$2899 ( \3663 , \3662 );
buf \U$2900 ( \3664 , \3663 );
xor \U$2901 ( \3665 , \3652 , \3664 );
buf \U$2902 ( \3666 , \1187 );
not \U$2903 ( \3667 , \3666 );
buf \U$2904 ( \3668 , \3667 );
buf \U$2905 ( \3669 , \3668 );
buf \U$2906 ( \3670 , \3620 );
not \U$2907 ( \3671 , \3670 );
buf \U$2908 ( \3672 , \3671 );
buf \U$2909 ( \3673 , \3672 );
or \U$2910 ( \3674 , \3669 , \3673 );
buf \U$2911 ( \3675 , \911 );
buf \U$2912 ( \3676 , \2280 );
or \U$2913 ( \3677 , \3675 , \3676 );
buf \U$2914 ( \3678 , \914 );
buf \U$2915 ( \3679 , \2063 );
or \U$2916 ( \3680 , \3678 , \3679 );
nand \U$2917 ( \3681 , \3677 , \3680 );
buf \U$2918 ( \3682 , \3681 );
buf \U$2919 ( \3683 , \3682 );
not \U$2920 ( \3684 , \3683 );
buf \U$2921 ( \3685 , \3684 );
buf \U$2922 ( \3686 , \3685 );
buf \U$2923 ( \3687 , \1194 );
not \U$2924 ( \3688 , \3687 );
buf \U$2925 ( \3689 , \3688 );
buf \U$2926 ( \3690 , \3689 );
or \U$2927 ( \3691 , \3686 , \3690 );
nand \U$2928 ( \3692 , \3674 , \3691 );
buf \U$2929 ( \3693 , \3692 );
buf \U$2930 ( \3694 , \3693 );
xor \U$2931 ( \3695 , \3665 , \3694 );
buf \U$2932 ( \3696 , \3695 );
buf \U$2933 ( \3697 , \3696 );
buf \U$2934 ( \3698 , \3579 );
buf \U$2935 ( \3699 , \2296 );
not \U$2936 ( \3700 , \3699 );
buf \U$2937 ( \3701 , \3700 );
buf \U$2938 ( \3702 , \3701 );
buf \U$2939 ( \3703 , \3598 );
not \U$2940 ( \3704 , \3703 );
buf \U$2941 ( \3705 , \3704 );
buf \U$2942 ( \3706 , \3705 );
or \U$2943 ( \3707 , \3702 , \3706 );
buf \U$2944 ( \3708 , \1950 );
not \U$2945 ( \3709 , \3708 );
buf \U$2946 ( \3710 , \3709 );
buf \U$2947 ( \3711 , \3710 );
buf \U$2948 ( \3712 , \1995 );
buf \U$2949 ( \3713 , \1334 );
and \U$2950 ( \3714 , \3712 , \3713 );
buf \U$2951 ( \3715 , \1619 );
buf \U$2952 ( \3716 , \1331 );
and \U$2953 ( \3717 , \3715 , \3716 );
nor \U$2954 ( \3718 , \3714 , \3717 );
buf \U$2955 ( \3719 , \3718 );
buf \U$2956 ( \3720 , \3719 );
or \U$2957 ( \3721 , \3711 , \3720 );
nand \U$2958 ( \3722 , \3707 , \3721 );
buf \U$2959 ( \3723 , \3722 );
buf \U$2960 ( \3724 , \3723 );
xor \U$2961 ( \3725 , \3698 , \3724 );
xor \U$2962 ( \3726 , \3588 , \3605 );
and \U$2963 ( \3727 , \3726 , \3627 );
and \U$2964 ( \3728 , \3588 , \3605 );
or \U$2965 ( \3729 , \3727 , \3728 );
buf \U$2966 ( \3730 , \3729 );
buf \U$2967 ( \3731 , \3730 );
xor \U$2968 ( \3732 , \3725 , \3731 );
buf \U$2969 ( \3733 , \3732 );
buf \U$2970 ( \3734 , \3733 );
xor \U$2971 ( \3735 , \3697 , \3734 );
xor \U$2972 ( \3736 , \3583 , \3630 );
and \U$2973 ( \3737 , \3736 , \3637 );
and \U$2974 ( \3738 , \3583 , \3630 );
or \U$2975 ( \3739 , \3737 , \3738 );
buf \U$2976 ( \3740 , \3739 );
buf \U$2977 ( \3741 , \3740 );
xor \U$2978 ( \3742 , \3735 , \3741 );
buf \U$2979 ( \3743 , \3742 );
buf \U$2980 ( \3744 , \3743 );
xor \U$2981 ( \3745 , \3555 , \3561 );
and \U$2982 ( \3746 , \3745 , \3640 );
and \U$2983 ( \3747 , \3555 , \3561 );
or \U$2984 ( \3748 , \3746 , \3747 );
buf \U$2985 ( \3749 , \3748 );
buf \U$2986 ( \3750 , \3749 );
or \U$2987 ( \3751 , \3744 , \3750 );
buf \U$2988 ( \3752 , \3751 );
buf \U$2989 ( \3753 , \3752 );
and \U$2990 ( \3754 , \3649 , \3753 );
buf \U$2991 ( \3755 , \3754 );
buf \U$2992 ( \3756 , \3755 );
xor \U$2993 ( \3757 , \3652 , \3664 );
and \U$2994 ( \3758 , \3757 , \3694 );
and \U$2995 ( \3759 , \3652 , \3664 );
or \U$2996 ( \3760 , \3758 , \3759 );
buf \U$2997 ( \3761 , \3760 );
buf \U$2998 ( \3762 , \3761 );
buf \U$2999 ( \3763 , \3701 );
buf \U$3000 ( \3764 , \3719 );
or \U$3001 ( \3765 , \3763 , \3764 );
buf \U$3002 ( \3766 , \1995 );
buf \U$3003 ( \3767 , \1542 );
and \U$3004 ( \3768 , \3766 , \3767 );
buf \U$3005 ( \3769 , \1619 );
buf \U$3006 ( \3770 , \1539 );
and \U$3007 ( \3771 , \3769 , \3770 );
nor \U$3008 ( \3772 , \3768 , \3771 );
buf \U$3009 ( \3773 , \3772 );
buf \U$3010 ( \3774 , \3773 );
buf \U$3011 ( \3775 , \3710 );
or \U$3012 ( \3776 , \3774 , \3775 );
nand \U$3013 ( \3777 , \3765 , \3776 );
buf \U$3014 ( \3778 , \3777 );
buf \U$3015 ( \3779 , \3778 );
and \U$3016 ( \3780 , \3595 , \3596 );
buf \U$3017 ( \3781 , \3780 );
buf \U$3018 ( \3782 , \3781 );
xor \U$3019 ( \3783 , \3779 , \3782 );
buf \U$3020 ( \3784 , \1187 );
buf \U$3021 ( \3785 , \3682 );
and \U$3022 ( \3786 , \3784 , \3785 );
buf \U$3023 ( \3787 , \1194 );
buf \U$3024 ( \3788 , \911 );
and \U$3025 ( \3789 , \3787 , \3788 );
nor \U$3026 ( \3790 , \3786 , \3789 );
buf \U$3027 ( \3791 , \3790 );
buf \U$3028 ( \3792 , \3791 );
xor \U$3029 ( \3793 , \3783 , \3792 );
buf \U$3030 ( \3794 , \3793 );
buf \U$3031 ( \3795 , \3794 );
xor \U$3032 ( \3796 , \3762 , \3795 );
xor \U$3033 ( \3797 , \3698 , \3724 );
and \U$3034 ( \3798 , \3797 , \3731 );
and \U$3035 ( \3799 , \3698 , \3724 );
or \U$3036 ( \3800 , \3798 , \3799 );
buf \U$3037 ( \3801 , \3800 );
buf \U$3038 ( \3802 , \3801 );
xor \U$3039 ( \3803 , \3796 , \3802 );
buf \U$3040 ( \3804 , \3803 );
buf \U$3041 ( \3805 , \3804 );
xor \U$3042 ( \3806 , \3697 , \3734 );
and \U$3043 ( \3807 , \3806 , \3741 );
and \U$3044 ( \3808 , \3697 , \3734 );
or \U$3045 ( \3809 , \3807 , \3808 );
buf \U$3046 ( \3810 , \3809 );
buf \U$3047 ( \3811 , \3810 );
nor \U$3048 ( \3812 , \3805 , \3811 );
buf \U$3049 ( \3813 , \3812 );
buf \U$3050 ( \3814 , \3813 );
not \U$3051 ( \3815 , \3814 );
buf \U$3052 ( \3816 , \3815 );
buf \U$3053 ( \3817 , \3816 );
and \U$3054 ( \3818 , \3756 , \3817 );
buf \U$3055 ( \3819 , \3818 );
buf \U$3056 ( \3820 , \3819 );
xor \U$3057 ( \3821 , \3779 , \3782 );
and \U$3058 ( \3822 , \3821 , \3792 );
and \U$3059 ( \3823 , \3779 , \3782 );
or \U$3060 ( \3824 , \3822 , \3823 );
buf \U$3061 ( \3825 , \3824 );
buf \U$3062 ( \3826 , \3825 );
buf \U$3063 ( \3827 , \3791 );
not \U$3064 ( \3828 , \3827 );
buf \U$3065 ( \3829 , \3828 );
buf \U$3066 ( \3830 , \3829 );
xor \U$3067 ( \3831 , \3826 , \3830 );
buf \U$3068 ( \3832 , \3701 );
buf \U$3069 ( \3833 , \3773 );
or \U$3070 ( \3834 , \3832 , \3833 );
buf \U$3071 ( \3835 , \3710 );
buf \U$3072 ( \3836 , \1995 );
buf \U$3073 ( \3837 , \2063 );
and \U$3074 ( \3838 , \3836 , \3837 );
buf \U$3075 ( \3839 , \1619 );
buf \U$3076 ( \3840 , \2280 );
and \U$3077 ( \3841 , \3839 , \3840 );
nor \U$3078 ( \3842 , \3838 , \3841 );
buf \U$3079 ( \3843 , \3842 );
buf \U$3080 ( \3844 , \3843 );
or \U$3081 ( \3845 , \3835 , \3844 );
nand \U$3082 ( \3846 , \3834 , \3845 );
buf \U$3083 ( \3847 , \3846 );
buf \U$3084 ( \3848 , \3847 );
buf \U$3085 ( \3849 , \1995 );
buf \U$3086 ( \3850 , \1331 );
nor \U$3087 ( \3851 , \3849 , \3850 );
buf \U$3088 ( \3852 , \3851 );
buf \U$3089 ( \3853 , \3852 );
xor \U$3090 ( \3854 , \3848 , \3853 );
buf \U$3091 ( \3855 , \3689 );
not \U$3092 ( \3856 , \3855 );
buf \U$3093 ( \3857 , \3668 );
not \U$3094 ( \3858 , \3857 );
or \U$3095 ( \3859 , \3856 , \3858 );
buf \U$3096 ( \3860 , \911 );
nand \U$3097 ( \3861 , \3859 , \3860 );
buf \U$3098 ( \3862 , \3861 );
buf \U$3099 ( \3863 , \3862 );
xor \U$3100 ( \3864 , \3854 , \3863 );
buf \U$3101 ( \3865 , \3864 );
buf \U$3102 ( \3866 , \3865 );
xor \U$3103 ( \3867 , \3831 , \3866 );
buf \U$3104 ( \3868 , \3867 );
buf \U$3105 ( \3869 , \3868 );
xor \U$3106 ( \3870 , \3762 , \3795 );
and \U$3107 ( \3871 , \3870 , \3802 );
and \U$3108 ( \3872 , \3762 , \3795 );
or \U$3109 ( \3873 , \3871 , \3872 );
buf \U$3110 ( \3874 , \3873 );
buf \U$3111 ( \3875 , \3874 );
or \U$3112 ( \3876 , \3869 , \3875 );
buf \U$3113 ( \3877 , \3876 );
buf \U$3114 ( \3878 , \3877 );
nand \U$3115 ( \3879 , \3820 , \3878 );
buf \U$3116 ( \3880 , \3879 );
buf \U$3117 ( \3881 , \3880 );
xor \U$3118 ( \3882 , \3826 , \3830 );
and \U$3119 ( \3883 , \3882 , \3866 );
and \U$3120 ( \3884 , \3826 , \3830 );
or \U$3121 ( \3885 , \3883 , \3884 );
buf \U$3122 ( \3886 , \3885 );
buf \U$3123 ( \3887 , \3886 );
buf \U$3124 ( \3888 , \3701 );
buf \U$3125 ( \3889 , \3843 );
or \U$3126 ( \3890 , \3888 , \3889 );
buf \U$3127 ( \3891 , \3710 );
buf \U$3128 ( \3892 , \1995 );
or \U$3129 ( \3893 , \3891 , \3892 );
nand \U$3130 ( \3894 , \3890 , \3893 );
buf \U$3131 ( \3895 , \3894 );
buf \U$3132 ( \3896 , \3895 );
buf \U$3133 ( \3897 , \1619 );
buf \U$3134 ( \3898 , \1542 );
nand \U$3135 ( \3899 , \3897 , \3898 );
buf \U$3136 ( \3900 , \3899 );
buf \U$3137 ( \3901 , \3900 );
xor \U$3138 ( \3902 , \3896 , \3901 );
xor \U$3139 ( \3903 , \3848 , \3853 );
and \U$3140 ( \3904 , \3903 , \3863 );
and \U$3141 ( \3905 , \3848 , \3853 );
or \U$3142 ( \3906 , \3904 , \3905 );
buf \U$3143 ( \3907 , \3906 );
buf \U$3144 ( \3908 , \3907 );
xor \U$3145 ( \3909 , \3902 , \3908 );
buf \U$3146 ( \3910 , \3909 );
buf \U$3147 ( \3911 , \3910 );
nor \U$3148 ( \3912 , \3887 , \3911 );
buf \U$3149 ( \3913 , \3912 );
buf \U$3150 ( \3914 , \3913 );
nor \U$3151 ( \3915 , \3881 , \3914 );
buf \U$3152 ( \3916 , \3915 );
buf \U$3153 ( \3917 , \3916 );
not \U$3154 ( \3918 , \3917 );
buf \U$3155 ( \3919 , \3177 );
buf \U$3156 ( \3920 , \2843 );
xor \U$3157 ( \3921 , \3919 , \3920 );
buf \U$3158 ( \3922 , \3522 );
xor \U$3159 ( \3923 , \3921 , \3922 );
buf \U$3160 ( \3924 , \3923 );
buf \U$3161 ( \3925 , \3924 );
xor \U$3162 ( \3926 , \2936 , \3150 );
xor \U$3163 ( \3927 , \3926 , \3173 );
buf \U$3164 ( \3928 , \3927 );
buf \U$3165 ( \3929 , \3928 );
buf \U$3166 ( \3930 , \3359 );
not \U$3167 ( \3931 , \3930 );
buf \U$3168 ( \3932 , \3364 );
not \U$3169 ( \3933 , \3932 );
or \U$3170 ( \3934 , \3931 , \3933 );
buf \U$3171 ( \3935 , \3359 );
buf \U$3172 ( \3936 , \3364 );
or \U$3173 ( \3937 , \3935 , \3936 );
nand \U$3174 ( \3938 , \3934 , \3937 );
buf \U$3175 ( \3939 , \3938 );
buf \U$3176 ( \3940 , \3939 );
not \U$3177 ( \3941 , \3940 );
buf \U$3178 ( \3942 , \3941 );
buf \U$3179 ( \3943 , \3942 );
not \U$3180 ( \3944 , \3943 );
buf \U$3181 ( \3945 , \3511 );
not \U$3182 ( \3946 , \3945 );
or \U$3183 ( \3947 , \3944 , \3946 );
buf \U$3184 ( \3948 , \3510 );
buf \U$3185 ( \3949 , \3939 );
nand \U$3186 ( \3950 , \3948 , \3949 );
buf \U$3187 ( \3951 , \3950 );
buf \U$3188 ( \3952 , \3951 );
nand \U$3189 ( \3953 , \3947 , \3952 );
buf \U$3190 ( \3954 , \3953 );
buf \U$3191 ( \3955 , \3954 );
xor \U$3192 ( \3956 , \3929 , \3955 );
buf \U$3193 ( \3957 , \3493 );
not \U$3194 ( \3958 , \3957 );
buf \U$3195 ( \3959 , \3501 );
not \U$3196 ( \3960 , \3959 );
or \U$3197 ( \3961 , \3958 , \3960 );
buf \U$3198 ( \3962 , \3493 );
buf \U$3199 ( \3963 , \3501 );
or \U$3200 ( \3964 , \3962 , \3963 );
nand \U$3201 ( \3965 , \3961 , \3964 );
buf \U$3202 ( \3966 , \3965 );
buf \U$3203 ( \3967 , \3966 );
buf \U$3204 ( \3968 , \3390 );
not \U$3205 ( \3969 , \3968 );
buf \U$3206 ( \3970 , \3969 );
buf \U$3207 ( \3971 , \3970 );
and \U$3208 ( \3972 , \3967 , \3971 );
not \U$3209 ( \3973 , \3967 );
buf \U$3210 ( \3974 , \3390 );
and \U$3211 ( \3975 , \3973 , \3974 );
nor \U$3212 ( \3976 , \3972 , \3975 );
buf \U$3213 ( \3977 , \3976 );
not \U$3214 ( \3978 , \3977 );
buf \U$3215 ( \3979 , \3228 );
not \U$3216 ( \3980 , \3979 );
buf \U$3217 ( \3981 , \3263 );
not \U$3218 ( \3982 , \3981 );
or \U$3219 ( \3983 , \3980 , \3982 );
buf \U$3220 ( \3984 , \3263 );
buf \U$3221 ( \3985 , \3228 );
or \U$3222 ( \3986 , \3984 , \3985 );
nand \U$3223 ( \3987 , \3983 , \3986 );
buf \U$3224 ( \3988 , \3987 );
xnor \U$3225 ( \3989 , \3349 , \3988 );
buf \U$3226 ( \3990 , \3989 );
not \U$3227 ( \3991 , \3990 );
buf \U$3228 ( \3992 , \3991 );
not \U$3229 ( \3993 , \3992 );
or \U$3230 ( \3994 , \3978 , \3993 );
buf \U$3231 ( \3995 , \3992 );
buf \U$3232 ( \3996 , \3977 );
or \U$3233 ( \3997 , \3995 , \3996 );
buf \U$3234 ( \3998 , \3260 );
not \U$3235 ( \3999 , \3998 );
buf \U$3236 ( \4000 , \1816 );
not \U$3237 ( \4001 , \4000 );
nand \U$3238 ( \4002 , \1291 , RI9145840_125);
not \U$3239 ( \4003 , \1524 );
nand \U$3240 ( \4004 , \4003 , RI9147dc0_205);
nand \U$3241 ( \4005 , \1008 , RI9148540_221);
nand \U$3242 ( \4006 , \943 , RI91450c0_109);
nand \U$3243 ( \4007 , \4002 , \4004 , \4005 , \4006 );
nand \U$3244 ( \4008 , \977 , RI9145fc0_141);
nand \U$3245 ( \4009 , \1014 , RI9148cc0_237);
nand \U$3246 ( \4010 , \1244 , RI9146740_157);
not \U$3247 ( \4011 , \1250 );
nand \U$3248 ( \4012 , \4011 , RI9149440_253);
nand \U$3249 ( \4013 , \4008 , \4009 , \4010 , \4012 );
nor \U$3250 ( \4014 , \4007 , \4013 );
nand \U$3251 ( \4015 , \951 , RI91441c0_77);
nand \U$3252 ( \4016 , \1218 , RI9144940_93);
nand \U$3253 ( \4017 , \1206 , RI9146ec0_173);
nand \U$3254 ( \4018 , \1213 , RI9147640_189);
nand \U$3255 ( \4019 , \4015 , \4016 , \4017 , \4018 );
nand \U$3256 ( \4020 , \963 , RI90f3928_29);
nand \U$3257 ( \4021 , \1302 , RI91432c0_45);
nand \U$3258 ( \4022 , \928 , RI9143a40_61);
nand \U$3259 ( \4023 , RI912e9b0_13, \968 );
nand \U$3260 ( \4024 , \4020 , \4021 , \4022 , \4023 );
nor \U$3261 ( \4025 , \4019 , \4024 );
nand \U$3262 ( \4026 , \4014 , \4025 );
buf \U$3263 ( \4027 , \4026 );
not \U$3264 ( \4028 , \4027 );
buf \U$3265 ( \4029 , \4028 );
buf \U$3266 ( \4030 , \4029 );
not \U$3267 ( \4031 , \4030 );
buf \U$3268 ( \4032 , \4031 );
buf \U$3269 ( \4033 , \4032 );
nand \U$3270 ( \4034 , \4001 , \4033 );
buf \U$3271 ( \4035 , \4034 );
buf \U$3272 ( \4036 , \4035 );
buf \U$3273 ( \4037 , \1107 );
not \U$3274 ( \4038 , \4037 );
buf \U$3275 ( \4039 , \1792 );
not \U$3276 ( \4040 , \4039 );
and \U$3277 ( \4041 , \4038 , \4040 );
buf \U$3278 ( \4042 , \1931 );
buf \U$3279 ( \4043 , \1337 );
and \U$3280 ( \4044 , \4042 , \4043 );
nor \U$3281 ( \4045 , \4041 , \4044 );
buf \U$3282 ( \4046 , \4045 );
buf \U$3283 ( \4047 , \4046 );
not \U$3284 ( \4048 , \4047 );
buf \U$3285 ( \4049 , \1469 );
not \U$3286 ( \4050 , \4049 );
and \U$3287 ( \4051 , \4048 , \4050 );
buf \U$3288 ( \4052 , \3308 );
buf \U$3289 ( \4053 , \1482 );
nor \U$3290 ( \4054 , \4052 , \4053 );
buf \U$3291 ( \4055 , \4054 );
buf \U$3292 ( \4056 , \4055 );
nor \U$3293 ( \4057 , \4051 , \4056 );
buf \U$3294 ( \4058 , \4057 );
buf \U$3295 ( \4059 , \4058 );
xor \U$3296 ( \4060 , \4036 , \4059 );
buf \U$3297 ( \4061 , \3288 );
not \U$3298 ( \4062 , \4061 );
buf \U$3299 ( \4063 , \1261 );
not \U$3300 ( \4064 , \4063 );
buf \U$3301 ( \4065 , \2479 );
not \U$3302 ( \4066 , \4065 );
or \U$3303 ( \4067 , \4064 , \4066 );
buf \U$3304 ( \4068 , \2479 );
not \U$3305 ( \4069 , \4068 );
buf \U$3306 ( \4070 , \4069 );
buf \U$3307 ( \4071 , \4070 );
buf \U$3308 ( \4072 , \1258 );
nand \U$3309 ( \4073 , \4071 , \4072 );
buf \U$3310 ( \4074 , \4073 );
buf \U$3311 ( \4075 , \4074 );
nand \U$3312 ( \4076 , \4067 , \4075 );
buf \U$3313 ( \4077 , \4076 );
buf \U$3314 ( \4078 , \4077 );
not \U$3315 ( \4079 , \4078 );
or \U$3316 ( \4080 , \4062 , \4079 );
buf \U$3317 ( \4081 , \3283 );
buf \U$3318 ( \4082 , \2473 );
nand \U$3319 ( \4083 , \4081 , \4082 );
buf \U$3320 ( \4084 , \4083 );
buf \U$3321 ( \4085 , \4084 );
nand \U$3322 ( \4086 , \4080 , \4085 );
buf \U$3323 ( \4087 , \4086 );
not \U$3324 ( \4088 , \4087 );
buf \U$3325 ( \4089 , \4088 );
and \U$3326 ( \4090 , \4060 , \4089 );
and \U$3327 ( \4091 , \4036 , \4059 );
or \U$3328 ( \4092 , \4090 , \4091 );
buf \U$3329 ( \4093 , \4092 );
buf \U$3330 ( \4094 , \4093 );
not \U$3331 ( \4095 , \4094 );
or \U$3332 ( \4096 , \3999 , \4095 );
and \U$3333 ( \4097 , \1536 , \3130 );
not \U$3334 ( \4098 , \1536 );
buf \U$3335 ( \4099 , \2462 );
buf \U$3337 ( \4100 , \4099 );
and \U$3338 ( \4101 , \4098 , \4100 );
or \U$3339 ( \4102 , \4097 , \4101 );
buf \U$3340 ( \4103 , \4102 );
buf \U$3341 ( \4104 , \3121 );
nand \U$3342 ( \4105 , \4103 , \4104 );
buf \U$3343 ( \4106 , \4105 );
buf \U$3344 ( \4107 , \4106 );
buf \U$3345 ( \4108 , \3094 );
or \U$3346 ( \4109 , \4107 , \4108 );
buf \U$3347 ( \4110 , \3243 );
buf \U$3348 ( \4111 , \3094 );
nand \U$3349 ( \4112 , \4110 , \4111 );
buf \U$3350 ( \4113 , \4112 );
buf \U$3351 ( \4114 , \4113 );
nand \U$3352 ( \4115 , \4109 , \4114 );
buf \U$3353 ( \4116 , \4115 );
buf \U$3354 ( \4117 , \4116 );
not \U$3355 ( \4118 , \4117 );
buf \U$3356 ( \4119 , \3402 );
not \U$3357 ( \4120 , \4119 );
buf \U$3358 ( \4121 , \2178 );
not \U$3359 ( \4122 , \4121 );
and \U$3360 ( \4123 , \4120 , \4122 );
buf \U$3361 ( \4124 , \2211 );
buf \U$3362 ( \4125 , \2194 );
not \U$3363 ( \4126 , \4125 );
buf \U$3364 ( \4127 , \4126 );
buf \U$3365 ( \4128 , \4127 );
buf \U$3366 ( \4129 , \1990 );
buf \U$3367 ( \4130 , \2878 );
and \U$3368 ( \4131 , \4129 , \4130 );
not \U$3369 ( \4132 , \4129 );
buf \U$3370 ( \4133 , \2067 );
and \U$3371 ( \4134 , \4132 , \4133 );
nor \U$3372 ( \4135 , \4131 , \4134 );
buf \U$3373 ( \4136 , \4135 );
buf \U$3374 ( \4137 , \4136 );
nor \U$3375 ( \4138 , \4128 , \4137 );
buf \U$3376 ( \4139 , \4138 );
buf \U$3377 ( \4140 , \4139 );
and \U$3378 ( \4141 , \4124 , \4140 );
nor \U$3379 ( \4142 , \4123 , \4141 );
buf \U$3380 ( \4143 , \4142 );
not \U$3381 ( \4144 , \4143 );
buf \U$3382 ( \4145 , \4144 );
not \U$3383 ( \4146 , \4145 );
or \U$3384 ( \4147 , \4118 , \4146 );
buf \U$3385 ( \4148 , \4143 );
not \U$3386 ( \4149 , \4148 );
buf \U$3387 ( \4150 , \4116 );
not \U$3388 ( \4151 , \4150 );
buf \U$3389 ( \4152 , \4151 );
buf \U$3390 ( \4153 , \4152 );
not \U$3391 ( \4154 , \4153 );
or \U$3392 ( \4155 , \4149 , \4154 );
not \U$3393 ( \4156 , RI914b330_319);
not \U$3394 ( \4157 , \831 );
or \U$3395 ( \4158 , \4156 , \4157 );
nand \U$3396 ( \4159 , \826 , RI914abb0_303);
nand \U$3397 ( \4160 , \4158 , \4159 );
not \U$3398 ( \4161 , RI914a430_287);
not \U$3399 ( \4162 , \813 );
or \U$3400 ( \4163 , \4161 , \4162 );
nand \U$3401 ( \4164 , \818 , RI9149cb0_271);
nand \U$3402 ( \4165 , \4163 , \4164 );
nor \U$3403 ( \4166 , \4160 , \4165 );
not \U$3404 ( \4167 , RI914c230_351);
not \U$3405 ( \4168 , \1044 );
or \U$3406 ( \4169 , \4167 , \4168 );
nand \U$3407 ( \4170 , \1144 , RI914bab0_335);
nand \U$3408 ( \4171 , \4169 , \4170 );
not \U$3409 ( \4172 , RI914d130_383);
not \U$3410 ( \4173 , \1094 );
or \U$3411 ( \4174 , \4172 , \4173 );
nand \U$3412 ( \4175 , \1155 , RI914c9b0_367);
nand \U$3413 ( \4176 , \4174 , \4175 );
nor \U$3414 ( \4177 , \4171 , \4176 );
not \U$3415 ( \4178 , RI914e7b0_431);
not \U$3416 ( \4179 , \1069 );
or \U$3417 ( \4180 , \4178 , \4179 );
nand \U$3418 ( \4181 , \883 , RI914ef30_447);
nand \U$3419 ( \4182 , \4180 , \4181 );
not \U$3420 ( \4183 , RI914d8b0_399);
not \U$3421 ( \4184 , \865 );
or \U$3422 ( \4185 , \4183 , \4184 );
nand \U$3423 ( \4186 , \870 , RI914e030_415);
nand \U$3424 ( \4187 , \4185 , \4186 );
nor \U$3425 ( \4188 , \4182 , \4187 );
not \U$3426 ( \4189 , RI914f6b0_463);
not \U$3427 ( \4190 , \1077 );
or \U$3428 ( \4191 , \4189 , \4190 );
nand \U$3429 ( \4192 , \1141 , RI914fe30_479);
nand \U$3430 ( \4193 , \4191 , \4192 );
not \U$3431 ( \4194 , RI91505b0_495);
not \U$3432 ( \4195 , \901 );
or \U$3433 ( \4196 , \4194 , \4195 );
and \U$3434 ( \4197 , RI9158d28_784, RI9158da0_785, RI9158cb0_783);
nand \U$3435 ( \4198 , \4197 , RI9158e18_786, RI9150d30_511);
nand \U$3436 ( \4199 , \4196 , \4198 );
nor \U$3437 ( \4200 , \4193 , \4199 );
nand \U$3438 ( \4201 , \4166 , \4177 , \4188 , \4200 );
buf \U$3439 ( \4202 , \4201 );
buf \U$3440 ( \4203 , \4202 );
nand \U$3441 ( \4204 , \826 , RI914ab38_302);
nand \U$3442 ( \4205 , \831 , RI914b2b8_318);
and \U$3443 ( \4206 , \4204 , \4205 );
and \U$3444 ( \4207 , \813 , RI914a3b8_286);
not \U$3445 ( \4208 , RI9149c38_270);
nor \U$3446 ( \4209 , \4208 , \1678 );
nor \U$3447 ( \4210 , \4207 , \4209 );
nand \U$3448 ( \4211 , \1358 , RI914ba38_334);
nand \U$3449 ( \4212 , \1406 , RI914c1b8_350);
and \U$3450 ( \4213 , \4211 , \4212 );
and \U$3451 ( \4214 , \1696 , RI914c938_366);
and \U$3452 ( \4215 , \1094 , RI914d0b8_382);
nor \U$3453 ( \4216 , \4214 , \4215 );
nand \U$3454 ( \4217 , \4206 , \4210 , \4213 , \4216 );
not \U$3455 ( \4218 , \1386 );
not \U$3456 ( \4219 , RI914e738_430);
not \U$3457 ( \4220 , \4219 );
and \U$3458 ( \4221 , \4218 , \4220 );
not \U$3459 ( \4222 , RI914eeb8_446);
nor \U$3460 ( \4223 , \4222 , \884 );
nor \U$3461 ( \4224 , \4221 , \4223 );
not \U$3462 ( \4225 , RI914d838_398);
nor \U$3463 ( \4226 , \4225 , \864 );
not \U$3464 ( \4227 , RI914dfb8_414);
nor \U$3465 ( \4228 , \4227 , \1061 );
nor \U$3466 ( \4229 , \4226 , \4228 );
and \U$3467 ( \4230 , \1077 , RI914f638_462);
and \U$3468 ( \4231 , \1141 , RI914fdb8_478);
nor \U$3469 ( \4232 , \4230 , \4231 );
and \U$3470 ( \4233 , \901 , RI9150538_494);
and \U$3471 ( \4234 , \1439 , RI9150cb8_510);
nor \U$3472 ( \4235 , \4233 , \4234 );
nand \U$3473 ( \4236 , \4224 , \4229 , \4232 , \4235 );
nor \U$3474 ( \4237 , \4217 , \4236 );
not \U$3475 ( \4238 , \4237 );
buf \U$3476 ( \4239 , \4238 );
not \U$3477 ( \4240 , \4239 );
buf \U$3478 ( \4241 , \4240 );
buf \U$3479 ( \4242 , \4241 );
and \U$3480 ( \4243 , \4203 , \4242 );
not \U$3481 ( \4244 , \4203 );
buf \U$3482 ( \4245 , \4238 );
and \U$3483 ( \4246 , \4244 , \4245 );
nor \U$3484 ( \4247 , \4243 , \4246 );
buf \U$3485 ( \4248 , \4247 );
buf \U$3486 ( \4249 , \4248 );
not \U$3487 ( \4250 , \4249 );
buf \U$3488 ( \4251 , \3044 );
buf \U$3490 ( \4252 , \4251 );
buf \U$3491 ( \4253 , \4252 );
not \U$3492 ( \4254 , \4253 );
buf \U$3493 ( \4255 , \4254 );
buf \U$3494 ( \4256 , \4255 );
not \U$3495 ( \4257 , \4256 );
buf \U$3496 ( \4258 , \4241 );
not \U$3497 ( \4259 , \4258 );
buf \U$3498 ( \4260 , \4259 );
buf \U$3499 ( \4261 , \4260 );
not \U$3500 ( \4262 , \4261 );
or \U$3501 ( \4263 , \4257 , \4262 );
buf \U$3502 ( \4264 , \4252 );
buf \U$3503 ( \4265 , \4241 );
nand \U$3504 ( \4266 , \4264 , \4265 );
buf \U$3505 ( \4267 , \4266 );
buf \U$3506 ( \4268 , \4267 );
nand \U$3507 ( \4269 , \4263 , \4268 );
buf \U$3508 ( \4270 , \4269 );
buf \U$3509 ( \4271 , \4270 );
buf \U$3510 ( \4272 , \4248 );
nand \U$3511 ( \4273 , \4271 , \4272 );
buf \U$3512 ( \4274 , \4273 );
buf \U$3513 ( \4275 , \4274 );
not \U$3514 ( \4276 , \4275 );
or \U$3515 ( \4277 , \4250 , \4276 );
buf \U$3518 ( \4278 , \4252 );
buf \U$3519 ( \4279 , \4278 );
not \U$3520 ( \4280 , \4279 );
buf \U$3521 ( \4281 , \4280 );
buf \U$3524 ( \4282 , \4281 );
buf \U$3525 ( \4283 , \4282 );
not \U$3526 ( \4284 , \4283 );
buf \U$3527 ( \4285 , \4284 );
buf \U$3528 ( \4286 , \4285 );
nand \U$3529 ( \4287 , \4277 , \4286 );
buf \U$3530 ( \4288 , \4287 );
buf \U$3531 ( \4289 , \4288 );
nand \U$3532 ( \4290 , \4155 , \4289 );
buf \U$3533 ( \4291 , \4290 );
buf \U$3534 ( \4292 , \4291 );
nand \U$3535 ( \4293 , \4147 , \4292 );
buf \U$3536 ( \4294 , \4293 );
buf \U$3540 ( \4295 , \4294 );
nand \U$3541 ( \4296 , \4096 , \4295 );
buf \U$3542 ( \4297 , \4296 );
buf \U$3543 ( \4298 , \4297 );
not \U$3544 ( \4299 , \4093 );
nand \U$3545 ( \4300 , \4299 , \3263 );
buf \U$3546 ( \4301 , \4300 );
nand \U$3547 ( \4302 , \4298 , \4301 );
buf \U$3548 ( \4303 , \4302 );
buf \U$3549 ( \4304 , \4303 );
nand \U$3550 ( \4305 , \3997 , \4304 );
buf \U$3551 ( \4306 , \4305 );
nand \U$3552 ( \4307 , \3994 , \4306 );
buf \U$3553 ( \4308 , \4307 );
and \U$3554 ( \4309 , \3956 , \4308 );
and \U$3555 ( \4310 , \3929 , \3955 );
or \U$3556 ( \4311 , \4309 , \4310 );
buf \U$3557 ( \4312 , \4311 );
buf \U$3558 ( \4313 , \4312 );
nand \U$3559 ( \4314 , \3925 , \4313 );
buf \U$3560 ( \4315 , \4314 );
buf \U$3561 ( \4316 , \4315 );
xor \U$3562 ( \4317 , \3929 , \3955 );
xor \U$3563 ( \4318 , \4317 , \4308 );
buf \U$3564 ( \4319 , \4318 );
buf \U$3565 ( \4320 , \4319 );
buf \U$3566 ( \4321 , \4303 );
not \U$3567 ( \4322 , \4321 );
buf \U$3568 ( \4323 , \3989 );
not \U$3569 ( \4324 , \4323 );
and \U$3570 ( \4325 , \4322 , \4324 );
buf \U$3571 ( \4326 , \4303 );
buf \U$3572 ( \4327 , \3989 );
and \U$3573 ( \4328 , \4326 , \4327 );
nor \U$3574 ( \4329 , \4325 , \4328 );
buf \U$3575 ( \4330 , \4329 );
buf \U$3576 ( \4331 , \4330 );
not \U$3577 ( \4332 , \4331 );
buf \U$3578 ( \4333 , \3977 );
not \U$3579 ( \4334 , \4333 );
or \U$3580 ( \4335 , \4332 , \4334 );
buf \U$3581 ( \4336 , \4330 );
buf \U$3582 ( \4337 , \3977 );
or \U$3583 ( \4338 , \4336 , \4337 );
nand \U$3584 ( \4339 , \4335 , \4338 );
buf \U$3585 ( \4340 , \4339 );
not \U$3586 ( \4341 , \4340 );
buf \U$3587 ( \4342 , \3298 );
buf \U$3588 ( \4343 , \3323 );
and \U$3589 ( \4344 , \4342 , \4343 );
not \U$3590 ( \4345 , \4342 );
buf \U$3591 ( \4346 , \3323 );
not \U$3592 ( \4347 , \4346 );
buf \U$3593 ( \4348 , \4347 );
buf \U$3594 ( \4349 , \4348 );
and \U$3595 ( \4350 , \4345 , \4349 );
nor \U$3596 ( \4351 , \4344 , \4350 );
buf \U$3597 ( \4352 , \4351 );
buf \U$3598 ( \4353 , \4352 );
not \U$3599 ( \4354 , \3331 );
not \U$3600 ( \4355 , \1187 );
or \U$3601 ( \4356 , \4354 , \4355 );
nand \U$3602 ( \4357 , \4356 , \3340 );
buf \U$3603 ( \4358 , \4357 );
and \U$3604 ( \4359 , \4353 , \4358 );
not \U$3605 ( \4360 , \4353 );
buf \U$3606 ( \4361 , \4357 );
not \U$3607 ( \4362 , \4361 );
buf \U$3608 ( \4363 , \4362 );
buf \U$3609 ( \4364 , \4363 );
and \U$3610 ( \4365 , \4360 , \4364 );
nor \U$3611 ( \4366 , \4359 , \4365 );
buf \U$3612 ( \4367 , \4366 );
buf \U$3613 ( \4368 , \4367 );
buf \U$3614 ( \4369 , \3450 );
buf \U$3615 ( \4370 , \3484 );
xor \U$3616 ( \4371 , \4369 , \4370 );
buf \U$3617 ( \4372 , \3405 );
xnor \U$3618 ( \4373 , \4371 , \4372 );
buf \U$3619 ( \4374 , \4373 );
buf \U$3620 ( \4375 , \4374 );
xor \U$3621 ( \4376 , \4368 , \4375 );
buf \U$3622 ( \4377 , \1618 );
not \U$3623 ( \4378 , \4377 );
buf \U$3624 ( \4379 , \3444 );
not \U$3625 ( \4380 , \4379 );
buf \U$3626 ( \4381 , \4380 );
buf \U$3627 ( \4382 , \4381 );
not \U$3628 ( \4383 , \4382 );
or \U$3629 ( \4384 , \4378 , \4383 );
buf \U$3630 ( \4385 , \3465 );
buf \U$3631 ( \4386 , \3444 );
nand \U$3632 ( \4387 , \4385 , \4386 );
buf \U$3633 ( \4388 , \4387 );
buf \U$3634 ( \4389 , \4388 );
nand \U$3635 ( \4390 , \4384 , \4389 );
buf \U$3636 ( \4391 , \4390 );
buf \U$3637 ( \4392 , \4391 );
not \U$3638 ( \4393 , \4392 );
buf \U$3639 ( \4394 , \1758 );
not \U$3640 ( \4395 , \4394 );
or \U$3641 ( \4396 , \4393 , \4395 );
buf \U$3642 ( \4397 , \3472 );
buf \U$3643 ( \4398 , \1882 );
nand \U$3644 ( \4399 , \4397 , \4398 );
buf \U$3645 ( \4400 , \4399 );
buf \U$3646 ( \4401 , \4400 );
nand \U$3647 ( \4402 , \4396 , \4401 );
buf \U$3648 ( \4403 , \4402 );
buf \U$3649 ( \4404 , \4403 );
not \U$3650 ( \4405 , \4404 );
buf \U$3651 ( \4406 , \1178 );
not \U$3652 ( \4407 , \4406 );
buf \U$3653 ( \4408 , \2758 );
not \U$3654 ( \4409 , \4408 );
or \U$3655 ( \4410 , \4407 , \4409 );
buf \U$3656 ( \4411 , \3329 );
buf \U$3657 ( \4412 , \2853 );
nand \U$3658 ( \4413 , \4411 , \4412 );
buf \U$3659 ( \4414 , \4413 );
buf \U$3660 ( \4415 , \4414 );
nand \U$3661 ( \4416 , \4410 , \4415 );
buf \U$3662 ( \4417 , \4416 );
buf \U$3663 ( \4418 , \4417 );
not \U$3664 ( \4419 , \4418 );
buf \U$3665 ( \4420 , \1186 );
not \U$3666 ( \4421 , \4420 );
or \U$3667 ( \4422 , \4419 , \4421 );
buf \U$3668 ( \4423 , \3331 );
buf \U$3669 ( \4424 , \1194 );
nand \U$3670 ( \4425 , \4423 , \4424 );
buf \U$3671 ( \4426 , \4425 );
buf \U$3672 ( \4427 , \4426 );
nand \U$3673 ( \4428 , \4422 , \4427 );
buf \U$3674 ( \4429 , \4428 );
buf \U$3675 ( \4430 , \4429 );
not \U$3676 ( \4431 , \4430 );
buf \U$3677 ( \4432 , \4431 );
buf \U$3678 ( \4433 , \4432 );
nand \U$3679 ( \4434 , \4405 , \4433 );
buf \U$3680 ( \4435 , \4434 );
buf \U$3681 ( \4436 , \4435 );
not \U$3682 ( \4437 , \4436 );
buf \U$3683 ( \4438 , \3223 );
not \U$3684 ( \4439 , \4438 );
buf \U$3685 ( \4440 , \914 );
not \U$3686 ( \4441 , \4440 );
or \U$3687 ( \4442 , \4439 , \4441 );
buf \U$3688 ( \4443 , \3459 );
buf \U$3689 ( \4444 , \3329 );
nand \U$3690 ( \4445 , \4443 , \4444 );
buf \U$3691 ( \4446 , \4445 );
buf \U$3692 ( \4447 , \4446 );
nand \U$3693 ( \4448 , \4442 , \4447 );
buf \U$3694 ( \4449 , \4448 );
buf \U$3695 ( \4450 , \4449 );
not \U$3696 ( \4451 , \4450 );
buf \U$3697 ( \4452 , \1186 );
not \U$3698 ( \4453 , \4452 );
or \U$3699 ( \4454 , \4451 , \4453 );
buf \U$3700 ( \4455 , \4417 );
buf \U$3701 ( \4456 , \1194 );
nand \U$3702 ( \4457 , \4455 , \4456 );
buf \U$3703 ( \4458 , \4457 );
buf \U$3704 ( \4459 , \4458 );
nand \U$3705 ( \4460 , \4454 , \4459 );
buf \U$3706 ( \4461 , \4460 );
buf \U$3707 ( \4462 , \4461 );
buf \U$3708 ( \4463 , \1027 );
not \U$3709 ( \4464 , \4463 );
buf \U$3710 ( \4465 , \2627 );
not \U$3711 ( \4466 , \4465 );
or \U$3712 ( \4467 , \4464 , \4466 );
buf \U$3713 ( \4468 , \2633 );
buf \U$3714 ( \4469 , \1024 );
nand \U$3715 ( \4470 , \4468 , \4469 );
buf \U$3716 ( \4471 , \4470 );
buf \U$3717 ( \4472 , \4471 );
nand \U$3718 ( \4473 , \4467 , \4472 );
buf \U$3719 ( \4474 , \4473 );
buf \U$3720 ( \4475 , \4474 );
not \U$3721 ( \4476 , \4475 );
buf \U$3722 ( \4477 , \3288 );
not \U$3723 ( \4478 , \4477 );
or \U$3724 ( \4479 , \4476 , \4478 );
buf \U$3725 ( \4480 , \2473 );
buf \U$3726 ( \4481 , \4077 );
nand \U$3727 ( \4482 , \4480 , \4481 );
buf \U$3728 ( \4483 , \4482 );
buf \U$3729 ( \4484 , \4483 );
nand \U$3730 ( \4485 , \4479 , \4484 );
buf \U$3731 ( \4486 , \4485 );
buf \U$3732 ( \4487 , \4486 );
and \U$3733 ( \4488 , \4462 , \4487 );
buf \U$3734 ( \4489 , \4488 );
buf \U$3735 ( \4490 , \4489 );
not \U$3736 ( \4491 , \4490 );
or \U$3737 ( \4492 , \4437 , \4491 );
buf \U$3738 ( \4493 , \4432 );
not \U$3739 ( \4494 , \4493 );
buf \U$3740 ( \4495 , \4403 );
nand \U$3741 ( \4496 , \4494 , \4495 );
buf \U$3742 ( \4497 , \4496 );
buf \U$3743 ( \4498 , \4497 );
nand \U$3744 ( \4499 , \4492 , \4498 );
buf \U$3745 ( \4500 , \4499 );
buf \U$3746 ( \4501 , \4500 );
and \U$3747 ( \4502 , \4376 , \4501 );
and \U$3748 ( \4503 , \4368 , \4375 );
or \U$3749 ( \4504 , \4502 , \4503 );
buf \U$3750 ( \4505 , \4504 );
buf \U$3751 ( \4506 , \4505 );
not \U$3752 ( \4507 , \4506 );
or \U$3753 ( \4508 , \4341 , \4507 );
buf \U$3754 ( \4509 , \4506 );
buf \U$3755 ( \4510 , \4340 );
or \U$3756 ( \4511 , \4509 , \4510 );
buf \U$3757 ( \4512 , \1334 );
not \U$3758 ( \4513 , \4512 );
buf \U$3759 ( \4514 , \4100 );
not \U$3760 ( \4515 , \4514 );
buf \U$3761 ( \4516 , \4515 );
buf \U$3762 ( \4517 , \4516 );
not \U$3763 ( \4518 , \4517 );
or \U$3764 ( \4519 , \4513 , \4518 );
buf \U$3765 ( \4520 , \3134 );
buf \U$3766 ( \4521 , \2565 );
nand \U$3767 ( \4522 , \4520 , \4521 );
buf \U$3768 ( \4523 , \4522 );
buf \U$3769 ( \4524 , \4523 );
nand \U$3770 ( \4525 , \4519 , \4524 );
buf \U$3771 ( \4526 , \4525 );
buf \U$3772 ( \4527 , \4526 );
not \U$3773 ( \4528 , \4527 );
buf \U$3774 ( \4529 , \3250 );
not \U$3775 ( \4530 , \4529 );
or \U$3776 ( \4531 , \4528 , \4530 );
buf \U$3777 ( \4532 , \3095 );
buf \U$3778 ( \4533 , \4102 );
nand \U$3779 ( \4534 , \4532 , \4533 );
buf \U$3780 ( \4535 , \4534 );
buf \U$3781 ( \4536 , \4535 );
nand \U$3782 ( \4537 , \4531 , \4536 );
buf \U$3783 ( \4538 , \4537 );
buf \U$3784 ( \4539 , \4538 );
not \U$3785 ( \4540 , \4539 );
buf \U$3786 ( \4541 , \4274 );
not \U$3787 ( \4542 , \4541 );
buf \U$3788 ( \4543 , \4542 );
buf \U$3789 ( \4544 , \4543 );
not \U$3790 ( \4545 , \4544 );
buf \U$3791 ( \4546 , \2063 );
not \U$3792 ( \4547 , \4546 );
buf \U$3793 ( \4548 , \4278 );
not \U$3794 ( \4549 , \4548 );
buf \U$3795 ( \4550 , \4549 );
buf \U$3796 ( \4551 , \4550 );
not \U$3797 ( \4552 , \4551 );
or \U$3798 ( \4553 , \4547 , \4552 );
buf \U$3799 ( \4554 , \4278 );
buf \U$3800 ( \4555 , \2280 );
nand \U$3801 ( \4556 , \4554 , \4555 );
buf \U$3802 ( \4557 , \4556 );
buf \U$3803 ( \4558 , \4557 );
nand \U$3804 ( \4559 , \4553 , \4558 );
buf \U$3805 ( \4560 , \4559 );
buf \U$3806 ( \4561 , \4560 );
not \U$3807 ( \4562 , \4561 );
or \U$3808 ( \4563 , \4545 , \4562 );
buf \U$3809 ( \4564 , \4550 );
not \U$3810 ( \4565 , \4564 );
buf \U$3811 ( \4566 , \4238 );
not \U$3812 ( \4567 , \4566 );
buf \U$3813 ( \4568 , \4567 );
buf \U$3814 ( \4569 , \4568 );
not \U$3815 ( \4570 , \4569 );
buf \U$3816 ( \4571 , \4202 );
not \U$3817 ( \4572 , \4571 );
or \U$3818 ( \4573 , \4570 , \4572 );
not \U$3819 ( \4574 , \4202 );
buf \U$3820 ( \4575 , \4574 );
buf \U$3821 ( \4576 , \4238 );
nand \U$3822 ( \4577 , \4575 , \4576 );
buf \U$3823 ( \4578 , \4577 );
buf \U$3824 ( \4579 , \4578 );
nand \U$3825 ( \4580 , \4573 , \4579 );
buf \U$3826 ( \4581 , \4580 );
buf \U$3827 ( \4582 , \4581 );
nand \U$3828 ( \4583 , \4565 , \4582 );
buf \U$3829 ( \4584 , \4583 );
buf \U$3830 ( \4585 , \4584 );
nand \U$3831 ( \4586 , \4563 , \4585 );
buf \U$3832 ( \4587 , \4586 );
buf \U$3833 ( \4588 , \4587 );
not \U$3834 ( \4589 , \4588 );
buf \U$3835 ( \4590 , \4589 );
buf \U$3836 ( \4591 , \4590 );
nand \U$3837 ( \4592 , \4540 , \4591 );
buf \U$3838 ( \4593 , \4592 );
buf \U$3839 ( \4594 , \4593 );
not \U$3840 ( \4595 , \4594 );
buf \U$3841 ( \4596 , \4595 );
buf \U$3842 ( \4597 , \4596 );
not \U$3843 ( \4598 , \4597 );
buf \U$3844 ( \4599 , \1862 );
not \U$3845 ( \4600 , \4599 );
buf \U$3846 ( \4601 , \2488 );
not \U$3847 ( \4602 , \4601 );
or \U$3848 ( \4603 , \4600 , \4602 );
buf \U$3849 ( \4604 , \2670 );
buf \U$3850 ( \4605 , \2067 );
nand \U$3851 ( \4606 , \4604 , \4605 );
buf \U$3852 ( \4607 , \4606 );
buf \U$3853 ( \4608 , \4607 );
nand \U$3854 ( \4609 , \4603 , \4608 );
buf \U$3855 ( \4610 , \4609 );
buf \U$3856 ( \4611 , \4610 );
not \U$3857 ( \4612 , \4611 );
buf \U$3858 ( \4613 , \2197 );
not \U$3859 ( \4614 , \4613 );
buf \U$3860 ( \4615 , \4614 );
buf \U$3861 ( \4616 , \4615 );
not \U$3862 ( \4617 , \4616 );
or \U$3863 ( \4618 , \4612 , \4617 );
not \U$3864 ( \4619 , \4136 );
nand \U$3865 ( \4620 , \4619 , \2208 );
buf \U$3866 ( \4621 , \4620 );
nand \U$3867 ( \4622 , \4618 , \4621 );
buf \U$3868 ( \4623 , \4622 );
buf \U$3869 ( \4624 , \4623 );
not \U$3870 ( \4625 , \4624 );
buf \U$3871 ( \4626 , \1618 );
not \U$3872 ( \4627 , RI9144238_78);
or \U$3873 ( \4628 , \952 , \4627 );
not \U$3874 ( \4629 , RI91449b8_94);
or \U$3875 ( \4630 , \957 , \4629 );
nand \U$3876 ( \4631 , \4628 , \4630 );
not \U$3877 ( \4632 , RI91458b8_126);
not \U$3878 ( \4633 , \936 );
or \U$3879 ( \4634 , \4632 , \4633 );
nand \U$3880 ( \4635 , \1226 , RI9145138_110);
nand \U$3881 ( \4636 , \4634 , \4635 );
nor \U$3882 ( \4637 , \4631 , \4636 );
not \U$3883 ( \4638 , RI9146f38_174);
not \U$3884 ( \4639 , \1206 );
or \U$3885 ( \4640 , \4638 , \4639 );
nand \U$3886 ( \4641 , \1213 , RI91476b8_190);
nand \U$3887 ( \4642 , \4640 , \4641 );
not \U$3888 ( \4643 , RI9146038_142);
not \U$3889 ( \4644 , \976 );
not \U$3890 ( \4645 , \4644 );
or \U$3891 ( \4646 , \4643 , \4645 );
nand \U$3892 ( \4647 , \1244 , RI91467b8_158);
nand \U$3893 ( \4648 , \4646 , \4647 );
nor \U$3894 ( \4649 , \4642 , \4648 );
not \U$3895 ( \4650 , RI9143338_46);
or \U$3896 ( \4651 , \922 , \4650 );
not \U$3897 ( \4652 , RI9143ab8_62);
or \U$3898 ( \4653 , \1622 , \4652 );
nand \U$3899 ( \4654 , \4651 , \4653 );
not \U$3900 ( \4655 , RI90f38b0_30);
not \U$3901 ( \4656 , \963 );
or \U$3902 ( \4657 , \4655 , \4656 );
nand \U$3903 ( \4658 , RI912e938_14, \968 );
nand \U$3904 ( \4659 , \4657 , \4658 );
nor \U$3905 ( \4660 , \4654 , \4659 );
not \U$3906 ( \4661 , RI9148d38_238);
not \U$3907 ( \4662 , \1014 );
or \U$3908 ( \4663 , \4661 , \4662 );
nand \U$3909 ( \4664 , \1251 , RI91494b8_254);
nand \U$3910 ( \4665 , \4663 , \4664 );
not \U$3911 ( \4666 , RI9147e38_206);
not \U$3912 ( \4667 , \1003 );
or \U$3913 ( \4668 , \4666 , \4667 );
nand \U$3914 ( \4669 , \1008 , RI91485b8_222);
nand \U$3915 ( \4670 , \4668 , \4669 );
nor \U$3916 ( \4671 , \4665 , \4670 );
nand \U$3917 ( \4672 , \4637 , \4649 , \4660 , \4671 );
buf \U$3918 ( \4673 , \4672 );
not \U$3919 ( \4674 , \4673 );
buf \U$3920 ( \4675 , \4674 );
buf \U$3921 ( \4676 , \4675 );
not \U$3922 ( \4677 , \4676 );
buf \U$3923 ( \4678 , \4677 );
buf \U$3924 ( \4679 , \4678 );
and \U$3925 ( \4680 , \4626 , \4679 );
buf \U$3926 ( \4681 , \4680 );
buf \U$3927 ( \4682 , \4681 );
not \U$3928 ( \4683 , \4682 );
buf \U$3929 ( \4684 , \4683 );
buf \U$3930 ( \4685 , \4684 );
nand \U$3931 ( \4686 , \4625 , \4685 );
buf \U$3932 ( \4687 , \4686 );
buf \U$3933 ( \4688 , \4687 );
buf \U$3934 ( \4689 , \1107 );
not \U$3935 ( \4690 , \4689 );
buf \U$3936 ( \4691 , \4690 );
and \U$3937 ( \4692 , \1669 , \4691 );
not \U$3938 ( \4693 , \1669 );
and \U$3939 ( \4694 , \4693 , \1337 );
or \U$3940 ( \4695 , \4692 , \4694 );
buf \U$3941 ( \4696 , \4695 );
not \U$3942 ( \4697 , \4696 );
buf \U$3943 ( \4698 , \1472 );
not \U$3944 ( \4699 , \4698 );
or \U$3945 ( \4700 , \4697 , \4699 );
buf \U$3946 ( \4701 , \4046 );
not \U$3947 ( \4702 , \4701 );
buf \U$3948 ( \4703 , \1904 );
nand \U$3949 ( \4704 , \4702 , \4703 );
buf \U$3950 ( \4705 , \4704 );
buf \U$3951 ( \4706 , \4705 );
nand \U$3952 ( \4707 , \4700 , \4706 );
buf \U$3953 ( \4708 , \4707 );
buf \U$3954 ( \4709 , \4708 );
and \U$3955 ( \4710 , \4688 , \4709 );
buf \U$3956 ( \4711 , \4623 );
buf \U$3957 ( \4712 , \4681 );
and \U$3958 ( \4713 , \4711 , \4712 );
buf \U$3959 ( \4714 , \4713 );
buf \U$3960 ( \4715 , \4714 );
nor \U$3961 ( \4716 , \4710 , \4715 );
buf \U$3962 ( \4717 , \4716 );
buf \U$3963 ( \4718 , \4717 );
not \U$3964 ( \4719 , \4718 );
or \U$3965 ( \4720 , \4598 , \4719 );
buf \U$3966 ( \4721 , \4116 );
buf \U$3967 ( \4722 , \4144 );
xor \U$3968 ( \4723 , \4721 , \4722 );
buf \U$3969 ( \4724 , \4288 );
xor \U$3970 ( \4725 , \4723 , \4724 );
buf \U$3971 ( \4726 , \4725 );
buf \U$3972 ( \4727 , \4726 );
nand \U$3973 ( \4728 , \4720 , \4727 );
buf \U$3974 ( \4729 , \4728 );
buf \U$3975 ( \4730 , \4729 );
buf \U$3976 ( \4731 , \4596 );
not \U$3977 ( \4732 , \4731 );
buf \U$3978 ( \4733 , \4717 );
not \U$3979 ( \4734 , \4733 );
buf \U$3980 ( \4735 , \4734 );
buf \U$3981 ( \4736 , \4735 );
nand \U$3982 ( \4737 , \4732 , \4736 );
buf \U$3983 ( \4738 , \4737 );
buf \U$3984 ( \4739 , \4738 );
nand \U$3985 ( \4740 , \4730 , \4739 );
buf \U$3986 ( \4741 , \4740 );
buf \U$3987 ( \4742 , \4741 );
not \U$3988 ( \4743 , \4742 );
buf \U$3989 ( \4744 , \4743 );
buf \U$3990 ( \4745 , \4744 );
buf \U$3991 ( \4746 , \3260 );
buf \U$3992 ( \4747 , \4294 );
xor \U$3993 ( \4748 , \4746 , \4747 );
buf \U$3994 ( \4749 , \4093 );
xnor \U$3995 ( \4750 , \4748 , \4749 );
buf \U$3996 ( \4751 , \4750 );
buf \U$3997 ( \4752 , \4751 );
nand \U$3998 ( \4753 , \4745 , \4752 );
buf \U$3999 ( \4754 , \4753 );
buf \U$4000 ( \4755 , \4754 );
not \U$4001 ( \4756 , \4755 );
xor \U$4002 ( \4757 , \4036 , \4059 );
xor \U$4003 ( \4758 , \4757 , \4089 );
buf \U$4004 ( \4759 , \4758 );
buf \U$4005 ( \4760 , \4759 );
not \U$4006 ( \4761 , \4760 );
xor \U$4007 ( \4762 , \4403 , \4432 );
xor \U$4008 ( \4763 , \4762 , \4489 );
buf \U$4009 ( \4764 , \4763 );
not \U$4010 ( \4765 , \4764 );
or \U$4011 ( \4766 , \4761 , \4765 );
buf \U$4012 ( \4767 , \4026 );
buf \U$4014 ( \4768 , \4767 );
buf \U$4015 ( \4769 , \4768 );
not \U$4016 ( \4770 , \4769 );
buf \U$4017 ( \4771 , \1800 );
not \U$4018 ( \4772 , \4771 );
or \U$4019 ( \4773 , \4770 , \4772 );
buf \U$4020 ( \4774 , \4029 );
buf \U$4021 ( \4775 , \1618 );
nand \U$4022 ( \4776 , \4774 , \4775 );
buf \U$4023 ( \4777 , \4776 );
buf \U$4024 ( \4778 , \4777 );
nand \U$4025 ( \4779 , \4773 , \4778 );
buf \U$4026 ( \4780 , \4779 );
buf \U$4027 ( \4781 , \4780 );
not \U$4028 ( \4782 , \4781 );
buf \U$4029 ( \4783 , \1946 );
not \U$4030 ( \4784 , \4783 );
or \U$4031 ( \4785 , \4782 , \4784 );
buf \U$4032 ( \4786 , \4391 );
buf \U$4033 ( \4787 , \1950 );
nand \U$4034 ( \4788 , \4786 , \4787 );
buf \U$4035 ( \4789 , \4788 );
buf \U$4036 ( \4790 , \4789 );
nand \U$4037 ( \4791 , \4785 , \4790 );
buf \U$4038 ( \4792 , \4791 );
buf \U$4039 ( \4793 , \4792 );
buf \U$4040 ( \4794 , \4201 );
not \U$4041 ( \4795 , \4794 );
not \U$4042 ( \4796 , \4795 );
buf \U$4043 ( \4797 , \2488 );
not \U$4044 ( \4798 , \4797 );
buf \U$4045 ( \4799 , \1795 );
not \U$4046 ( \4800 , \4799 );
or \U$4047 ( \4801 , \4798 , \4800 );
buf \U$4048 ( \4802 , \2068 );
buf \U$4049 ( \4803 , \1931 );
nand \U$4050 ( \4804 , \4802 , \4803 );
buf \U$4051 ( \4805 , \4804 );
buf \U$4052 ( \4806 , \4805 );
nand \U$4053 ( \4807 , \4801 , \4806 );
buf \U$4054 ( \4808 , \4807 );
nand \U$4055 ( \4809 , \2200 , \4808 );
not \U$4056 ( \4810 , \4809 );
not \U$4057 ( \4811 , \4610 );
buf \U$4058 ( \4812 , \2897 );
not \U$4059 ( \4813 , \4812 );
buf \U$4060 ( \4814 , \4813 );
nor \U$4061 ( \4815 , \4811 , \4814 );
nor \U$4062 ( \4816 , \4810 , \4815 );
nand \U$4063 ( \4817 , \4796 , \4816 );
buf \U$4064 ( \4818 , \4817 );
xor \U$4065 ( \4819 , \4793 , \4818 );
buf \U$4066 ( \4820 , \1618 );
and \U$4067 ( \4821 , \1525 , RI9147eb0_207);
and \U$4068 ( \4822 , \1200 , RI9148630_223);
nor \U$4069 ( \4823 , \4821 , \4822 );
not \U$4070 ( \4824 , RI91460b0_143);
nor \U$4071 ( \4825 , \4824 , \976 );
not \U$4072 ( \4826 , RI9146830_159);
nor \U$4073 ( \4827 , \4826 , \983 );
nor \U$4074 ( \4828 , \4825 , \4827 );
nand \U$4075 ( \4829 , \4823 , \4828 );
nand \U$4076 ( \4830 , \1204 , RI9146fb0_175);
nand \U$4077 ( \4831 , \1213 , RI9147730_191);
nand \U$4078 ( \4832 , \1014 , RI9148db0_239);
nand \U$4079 ( \4833 , \1017 , RI9149530_255);
nand \U$4080 ( \4834 , \4830 , \4831 , \4832 , \4833 );
nor \U$4081 ( \4835 , \4829 , \4834 );
nand \U$4082 ( \4836 , \921 , RI91433b0_47);
nand \U$4083 ( \4837 , \928 , RI9143b30_63);
nand \U$4084 ( \4838 , \1291 , RI9145930_127);
nand \U$4085 ( \4839 , \1508 , RI91451b0_111);
nand \U$4086 ( \4840 , \4836 , \4837 , \4838 , \4839 );
nand \U$4087 ( \4841 , \963 , RI90f3838_31);
nand \U$4088 ( \4842 , \1297 , RI912e8c0_15);
nand \U$4089 ( \4843 , \951 , RI91442b0_79);
nand \U$4090 ( \4844 , \1218 , RI9144a30_95);
nand \U$4091 ( \4845 , \4841 , \4842 , \4843 , \4844 );
nor \U$4092 ( \4846 , \4840 , \4845 );
nand \U$4093 ( \4847 , \4835 , \4846 );
buf \U$4094 ( \4848 , \4847 );
buf \U$4095 ( \4849 , \4848 );
and \U$4096 ( \4850 , \4820 , \4849 );
buf \U$4097 ( \4851 , \4850 );
buf \U$4098 ( \4852 , \4851 );
not \U$4099 ( \4853 , \4852 );
buf \U$4100 ( \4854 , \4672 );
buf \U$4102 ( \4855 , \4854 );
buf \U$4103 ( \4856 , \4855 );
not \U$4104 ( \4857 , \4856 );
buf \U$4105 ( \4858 , \3465 );
not \U$4106 ( \4859 , \4858 );
or \U$4107 ( \4860 , \4857 , \4859 );
buf \U$4108 ( \4861 , \4855 );
not \U$4109 ( \4862 , \4861 );
buf \U$4110 ( \4863 , \4862 );
buf \U$4111 ( \4864 , \4863 );
buf \U$4112 ( \4865 , \1618 );
nand \U$4113 ( \4866 , \4864 , \4865 );
buf \U$4114 ( \4867 , \4866 );
buf \U$4115 ( \4868 , \4867 );
nand \U$4116 ( \4869 , \4860 , \4868 );
buf \U$4117 ( \4870 , \4869 );
buf \U$4118 ( \4871 , \4870 );
not \U$4119 ( \4872 , \4871 );
buf \U$4120 ( \4873 , \1758 );
not \U$4121 ( \4874 , \4873 );
or \U$4122 ( \4875 , \4872 , \4874 );
buf \U$4123 ( \4876 , \4780 );
buf \U$4124 ( \4877 , \1882 );
nand \U$4125 ( \4878 , \4876 , \4877 );
buf \U$4126 ( \4879 , \4878 );
buf \U$4127 ( \4880 , \4879 );
nand \U$4128 ( \4881 , \4875 , \4880 );
buf \U$4129 ( \4882 , \4881 );
buf \U$4130 ( \4883 , \4882 );
not \U$4131 ( \4884 , \4883 );
or \U$4132 ( \4885 , \4853 , \4884 );
or \U$4133 ( \4886 , \4851 , \4882 );
buf \U$4134 ( \4887 , \2521 );
not \U$4135 ( \4888 , \4887 );
buf \U$4136 ( \4889 , \2627 );
not \U$4137 ( \4890 , \4889 );
or \U$4138 ( \4891 , \4888 , \4890 );
buf \U$4139 ( \4892 , \4070 );
buf \U$4140 ( \4893 , \1999 );
nand \U$4141 ( \4894 , \4892 , \4893 );
buf \U$4142 ( \4895 , \4894 );
buf \U$4143 ( \4896 , \4895 );
nand \U$4144 ( \4897 , \4891 , \4896 );
buf \U$4145 ( \4898 , \4897 );
buf \U$4146 ( \4899 , \4898 );
not \U$4147 ( \4900 , \4899 );
buf \U$4148 ( \4901 , \2983 );
not \U$4149 ( \4902 , \4901 );
or \U$4150 ( \4903 , \4900 , \4902 );
buf \U$4151 ( \4904 , \4474 );
buf \U$4152 ( \4905 , \2473 );
nand \U$4153 ( \4906 , \4904 , \4905 );
buf \U$4154 ( \4907 , \4906 );
buf \U$4155 ( \4908 , \4907 );
nand \U$4156 ( \4909 , \4903 , \4908 );
buf \U$4157 ( \4910 , \4909 );
nand \U$4158 ( \4911 , \4886 , \4910 );
buf \U$4159 ( \4912 , \4911 );
nand \U$4160 ( \4913 , \4885 , \4912 );
buf \U$4161 ( \4914 , \4913 );
buf \U$4162 ( \4915 , \4914 );
and \U$4163 ( \4916 , \4819 , \4915 );
and \U$4164 ( \4917 , \4793 , \4818 );
or \U$4165 ( \4918 , \4916 , \4917 );
buf \U$4166 ( \4919 , \4918 );
buf \U$4167 ( \4920 , \4919 );
nand \U$4168 ( \4921 , \4766 , \4920 );
buf \U$4169 ( \4922 , \4921 );
buf \U$4170 ( \4923 , \4922 );
buf \U$4171 ( \4924 , \4759 );
not \U$4172 ( \4925 , \4924 );
buf \U$4173 ( \4926 , \4763 );
not \U$4174 ( \4927 , \4926 );
buf \U$4175 ( \4928 , \4927 );
buf \U$4176 ( \4929 , \4928 );
nand \U$4177 ( \4930 , \4925 , \4929 );
buf \U$4178 ( \4931 , \4930 );
buf \U$4179 ( \4932 , \4931 );
nand \U$4180 ( \4933 , \4923 , \4932 );
buf \U$4181 ( \4934 , \4933 );
buf \U$4182 ( \4935 , \4934 );
not \U$4183 ( \4936 , \4935 );
or \U$4184 ( \4937 , \4756 , \4936 );
buf \U$4185 ( \4938 , \4751 );
buf \U$4186 ( \4939 , \4744 );
or \U$4187 ( \4940 , \4938 , \4939 );
buf \U$4188 ( \4941 , \4940 );
buf \U$4189 ( \4942 , \4941 );
nand \U$4190 ( \4943 , \4937 , \4942 );
buf \U$4191 ( \4944 , \4943 );
buf \U$4192 ( \4945 , \4944 );
nand \U$4193 ( \4946 , \4511 , \4945 );
buf \U$4194 ( \4947 , \4946 );
nand \U$4195 ( \4948 , \4508 , \4947 );
buf \U$4196 ( \4949 , \4948 );
nand \U$4197 ( \4950 , \4320 , \4949 );
buf \U$4198 ( \4951 , \4950 );
buf \U$4199 ( \4952 , \4951 );
nand \U$4200 ( \4953 , \4316 , \4952 );
buf \U$4201 ( \4954 , \4953 );
buf \U$4202 ( \4955 , \4954 );
not \U$4203 ( \4956 , \4955 );
buf \U$4204 ( \4957 , \4956 );
buf \U$4205 ( \4958 , \4957 );
buf \U$4206 ( \4959 , \4759 );
buf \U$4207 ( \4960 , \4919 );
xor \U$4208 ( \4961 , \4959 , \4960 );
buf \U$4209 ( \4962 , \4928 );
xnor \U$4210 ( \4963 , \4961 , \4962 );
buf \U$4211 ( \4964 , \4963 );
buf \U$4212 ( \4965 , \4964 );
buf \U$4213 ( \4966 , \4851 );
buf \U$4214 ( \4967 , \4882 );
xor \U$4215 ( \4968 , \4966 , \4967 );
buf \U$4216 ( \4969 , \4910 );
xnor \U$4217 ( \4970 , \4968 , \4969 );
buf \U$4218 ( \4971 , \4970 );
buf \U$4219 ( \4972 , \4971 );
not \U$4220 ( \4973 , \4972 );
buf \U$4221 ( \4974 , \4973 );
not \U$4222 ( \4975 , \4974 );
not \U$4223 ( \4976 , \4816 );
nand \U$4224 ( \4977 , \4976 , \4795 );
nand \U$4225 ( \4978 , \4977 , \4817 );
not \U$4226 ( \4979 , \4978 );
or \U$4227 ( \4980 , \4975 , \4979 );
not \U$4228 ( \4981 , \4971 );
buf \U$4229 ( \4982 , \4978 );
not \U$4230 ( \4983 , \4982 );
buf \U$4231 ( \4984 , \4983 );
not \U$4232 ( \4985 , \4984 );
or \U$4233 ( \4986 , \4981 , \4985 );
buf \U$4234 ( \4987 , \1618 );
not \U$4235 ( \4988 , \4987 );
buf \U$4236 ( \4989 , \4848 );
not \U$4237 ( \4990 , \4989 );
buf \U$4238 ( \4991 , \4990 );
buf \U$4239 ( \4992 , \4991 );
not \U$4240 ( \4993 , \4992 );
or \U$4241 ( \4994 , \4988 , \4993 );
buf \U$4242 ( \4995 , \1816 );
buf \U$4243 ( \4996 , \4848 );
nand \U$4244 ( \4997 , \4995 , \4996 );
buf \U$4245 ( \4998 , \4997 );
buf \U$4246 ( \4999 , \4998 );
nand \U$4247 ( \5000 , \4994 , \4999 );
buf \U$4248 ( \5001 , \5000 );
buf \U$4249 ( \5002 , \5001 );
not \U$4250 ( \5003 , \5002 );
buf \U$4251 ( \5004 , \1758 );
not \U$4252 ( \5005 , \5004 );
or \U$4253 ( \5006 , \5003 , \5005 );
buf \U$4254 ( \5007 , \4870 );
buf \U$4255 ( \5008 , \1882 );
nand \U$4256 ( \5009 , \5007 , \5008 );
buf \U$4257 ( \5010 , \5009 );
buf \U$4258 ( \5011 , \5010 );
nand \U$4259 ( \5012 , \5006 , \5011 );
buf \U$4260 ( \5013 , \5012 );
buf \U$4261 ( \5014 , \5013 );
buf \U$4262 ( \5015 , \2670 );
not \U$4263 ( \5016 , \5015 );
buf \U$4264 ( \5017 , \5016 );
buf \U$4265 ( \5018 , \5017 );
not \U$4266 ( \5019 , \5018 );
buf \U$4267 ( \5020 , \2479 );
not \U$4268 ( \5021 , \5020 );
or \U$4269 ( \5022 , \5019 , \5021 );
buf \U$4270 ( \5023 , \3276 );
buf \U$4271 ( \5024 , \2670 );
nand \U$4272 ( \5025 , \5023 , \5024 );
buf \U$4273 ( \5026 , \5025 );
buf \U$4274 ( \5027 , \5026 );
nand \U$4275 ( \5028 , \5022 , \5027 );
buf \U$4276 ( \5029 , \5028 );
buf \U$4277 ( \5030 , \5029 );
not \U$4278 ( \5031 , \5030 );
buf \U$4279 ( \5032 , \3288 );
not \U$4280 ( \5033 , \5032 );
or \U$4281 ( \5034 , \5031 , \5033 );
buf \U$4282 ( \5035 , \4898 );
buf \U$4283 ( \5036 , \2473 );
nand \U$4284 ( \5037 , \5035 , \5036 );
buf \U$4285 ( \5038 , \5037 );
buf \U$4286 ( \5039 , \5038 );
nand \U$4287 ( \5040 , \5034 , \5039 );
buf \U$4288 ( \5041 , \5040 );
buf \U$4289 ( \5042 , \5041 );
xor \U$4290 ( \5043 , \5014 , \5042 );
buf \U$4291 ( \5044 , \4543 );
not \U$4292 ( \5045 , \5044 );
buf \U$4293 ( \5046 , \5045 );
buf \U$4294 ( \5047 , \5046 );
buf \U$4295 ( \5048 , \1334 );
not \U$4296 ( \5049 , \5048 );
buf \U$4297 ( \5050 , \4550 );
not \U$4298 ( \5051 , \5050 );
or \U$4299 ( \5052 , \5049 , \5051 );
buf \U$4300 ( \5053 , \4278 );
buf \U$4301 ( \5054 , \1331 );
nand \U$4302 ( \5055 , \5053 , \5054 );
buf \U$4303 ( \5056 , \5055 );
buf \U$4304 ( \5057 , \5056 );
nand \U$4305 ( \5058 , \5052 , \5057 );
buf \U$4306 ( \5059 , \5058 );
buf \U$4307 ( \5060 , \5059 );
not \U$4308 ( \5061 , \5060 );
buf \U$4309 ( \5062 , \5061 );
buf \U$4310 ( \5063 , \5062 );
or \U$4311 ( \5064 , \5047 , \5063 );
buf \U$4314 ( \5065 , \4248 );
buf \U$4315 ( \5066 , \5065 );
buf \U$4316 ( \5067 , \1542 );
not \U$4317 ( \5068 , \5067 );
buf \U$4318 ( \5069 , \4281 );
not \U$4319 ( \5070 , \5069 );
or \U$4320 ( \5071 , \5068 , \5070 );
buf \U$4321 ( \5072 , \4278 );
buf \U$4322 ( \5073 , \1539 );
nand \U$4323 ( \5074 , \5072 , \5073 );
buf \U$4324 ( \5075 , \5074 );
buf \U$4325 ( \5076 , \5075 );
nand \U$4326 ( \5077 , \5071 , \5076 );
buf \U$4327 ( \5078 , \5077 );
buf \U$4328 ( \5079 , \5078 );
not \U$4329 ( \5080 , \5079 );
buf \U$4330 ( \5081 , \5080 );
buf \U$4331 ( \5082 , \5081 );
or \U$4332 ( \5083 , \5066 , \5082 );
nand \U$4333 ( \5084 , \5064 , \5083 );
buf \U$4334 ( \5085 , \5084 );
buf \U$4335 ( \5086 , \5085 );
and \U$4336 ( \5087 , \5043 , \5086 );
and \U$4337 ( \5088 , \5014 , \5042 );
or \U$4338 ( \5089 , \5087 , \5088 );
buf \U$4339 ( \5090 , \5089 );
nand \U$4340 ( \5091 , \4986 , \5090 );
nand \U$4341 ( \5092 , \4980 , \5091 );
buf \U$4342 ( \5093 , \5092 );
buf \U$4344 ( \5094 , \5093 );
buf \U$4345 ( \5095 , \5094 );
not \U$4346 ( \5096 , \5095 );
xor \U$4347 ( \5097 , \4462 , \4487 );
buf \U$4348 ( \5098 , \5097 );
buf \U$4349 ( \5099 , \5098 );
buf \U$4350 ( \5100 , \2758 );
not \U$4351 ( \5101 , \5100 );
buf \U$4352 ( \5102 , \4691 );
not \U$4353 ( \5103 , \5102 );
or \U$4354 ( \5104 , \5101 , \5103 );
buf \U$4355 ( \5105 , \2853 );
buf \U$4356 ( \5106 , \1337 );
nand \U$4357 ( \5107 , \5105 , \5106 );
buf \U$4358 ( \5108 , \5107 );
buf \U$4359 ( \5109 , \5108 );
nand \U$4360 ( \5110 , \5104 , \5109 );
buf \U$4361 ( \5111 , \5110 );
buf \U$4362 ( \5112 , \5111 );
not \U$4363 ( \5113 , \5112 );
buf \U$4364 ( \5114 , \1472 );
not \U$4365 ( \5115 , \5114 );
or \U$4366 ( \5116 , \5113 , \5115 );
buf \U$4367 ( \5117 , \1482 );
not \U$4368 ( \5118 , \5117 );
buf \U$4369 ( \5119 , \4695 );
nand \U$4370 ( \5120 , \5118 , \5119 );
buf \U$4371 ( \5121 , \5120 );
buf \U$4372 ( \5122 , \5121 );
nand \U$4373 ( \5123 , \5116 , \5122 );
buf \U$4374 ( \5124 , \5123 );
buf \U$4377 ( \5125 , \5124 );
buf \U$4378 ( \5126 , \5125 );
buf \U$4379 ( \5127 , \1255 );
buf \U$4381 ( \5128 , \5127 );
buf \U$4382 ( \5129 , \5128 );
not \U$4383 ( \5130 , \5129 );
buf \U$4384 ( \5131 , \4516 );
not \U$4385 ( \5132 , \5131 );
or \U$4386 ( \5133 , \5130 , \5132 );
buf \U$4387 ( \5134 , \3134 );
buf \U$4388 ( \5135 , \1258 );
nand \U$4389 ( \5136 , \5134 , \5135 );
buf \U$4390 ( \5137 , \5136 );
buf \U$4391 ( \5138 , \5137 );
nand \U$4392 ( \5139 , \5133 , \5138 );
buf \U$4393 ( \5140 , \5139 );
buf \U$4394 ( \5141 , \5140 );
not \U$4395 ( \5142 , \5141 );
not \U$4396 ( \5143 , \3249 );
buf \U$4397 ( \5144 , \5143 );
not \U$4398 ( \5145 , \5144 );
or \U$4399 ( \5146 , \5142 , \5145 );
buf \U$4400 ( \5147 , \3095 );
buf \U$4401 ( \5148 , \4526 );
nand \U$4402 ( \5149 , \5147 , \5148 );
buf \U$4403 ( \5150 , \5149 );
buf \U$4404 ( \5151 , \5150 );
nand \U$4405 ( \5152 , \5146 , \5151 );
buf \U$4406 ( \5153 , \5152 );
buf \U$4407 ( \5154 , \5153 );
nor \U$4408 ( \5155 , \5126 , \5154 );
buf \U$4409 ( \5156 , \5155 );
buf \U$4410 ( \5157 , \5156 );
buf \U$4411 ( \5158 , \5078 );
not \U$4412 ( \5159 , \5158 );
buf \U$4413 ( \5160 , \4543 );
not \U$4414 ( \5161 , \5160 );
or \U$4415 ( \5162 , \5159 , \5161 );
buf \U$4416 ( \5163 , \4560 );
buf \U$4417 ( \5164 , \4581 );
nand \U$4418 ( \5165 , \5163 , \5164 );
buf \U$4419 ( \5166 , \5165 );
buf \U$4420 ( \5167 , \5166 );
nand \U$4421 ( \5168 , \5162 , \5167 );
buf \U$4422 ( \5169 , \5168 );
buf \U$4423 ( \5170 , \5169 );
not \U$4424 ( \5171 , \5170 );
buf \U$4425 ( \5172 , \5171 );
buf \U$4426 ( \5173 , \5172 );
or \U$4427 ( \5174 , \5157 , \5173 );
buf \U$4428 ( \5175 , \5125 );
buf \U$4429 ( \5176 , \5153 );
nand \U$4430 ( \5177 , \5175 , \5176 );
buf \U$4431 ( \5178 , \5177 );
buf \U$4432 ( \5179 , \5178 );
nand \U$4433 ( \5180 , \5174 , \5179 );
buf \U$4434 ( \5181 , \5180 );
buf \U$4435 ( \5182 , \5181 );
xor \U$4436 ( \5183 , \5099 , \5182 );
buf \U$4437 ( \5184 , \4538 );
not \U$4438 ( \5185 , \5184 );
buf \U$4439 ( \5186 , \4590 );
nor \U$4440 ( \5187 , \5185 , \5186 );
buf \U$4441 ( \5188 , \5187 );
buf \U$4442 ( \5189 , \5188 );
not \U$4443 ( \5190 , \5189 );
buf \U$4444 ( \5191 , \4593 );
nand \U$4445 ( \5192 , \5190 , \5191 );
buf \U$4446 ( \5193 , \5192 );
buf \U$4447 ( \5194 , \5193 );
xor \U$4448 ( \5195 , \5183 , \5194 );
buf \U$4449 ( \5196 , \5195 );
buf \U$4450 ( \5197 , \5196 );
not \U$4451 ( \5198 , \5197 );
or \U$4452 ( \5199 , \5096 , \5198 );
buf \U$4453 ( \5200 , \5094 );
buf \U$4454 ( \5201 , \5196 );
or \U$4455 ( \5202 , \5200 , \5201 );
buf \U$4456 ( \5203 , \5124 );
buf \U$4457 ( \5204 , \5153 );
xor \U$4458 ( \5205 , \5203 , \5204 );
buf \U$4459 ( \5206 , \5172 );
xor \U$4460 ( \5207 , \5205 , \5206 );
buf \U$4461 ( \5208 , \5207 );
not \U$4462 ( \5209 , \5208 );
buf \U$4463 ( \5210 , \3223 );
not \U$4464 ( \5211 , \5210 );
buf \U$4465 ( \5212 , \1547 );
not \U$4466 ( \5213 , \5212 );
or \U$4467 ( \5214 , \5211 , \5213 );
buf \U$4468 ( \5215 , \3459 );
buf \U$4469 ( \5216 , \1337 );
nand \U$4470 ( \5217 , \5215 , \5216 );
buf \U$4471 ( \5218 , \5217 );
buf \U$4472 ( \5219 , \5218 );
nand \U$4473 ( \5220 , \5214 , \5219 );
buf \U$4474 ( \5221 , \5220 );
buf \U$4475 ( \5222 , \5221 );
not \U$4476 ( \5223 , \5222 );
buf \U$4477 ( \5224 , \1472 );
not \U$4478 ( \5225 , \5224 );
or \U$4479 ( \5226 , \5223 , \5225 );
buf \U$4480 ( \5227 , \1482 );
not \U$4481 ( \5228 , \5227 );
buf \U$4482 ( \5229 , \5111 );
nand \U$4483 ( \5230 , \5228 , \5229 );
buf \U$4484 ( \5231 , \5230 );
buf \U$4485 ( \5232 , \5231 );
nand \U$4486 ( \5233 , \5226 , \5232 );
buf \U$4487 ( \5234 , \5233 );
buf \U$4488 ( \5235 , \5234 );
buf \U$4489 ( \5236 , \914 );
not \U$4490 ( \5237 , \5236 );
buf \U$4491 ( \5238 , \4768 );
not \U$4492 ( \5239 , \5238 );
or \U$4493 ( \5240 , \5237 , \5239 );
buf \U$4494 ( \5241 , \4768 );
not \U$4495 ( \5242 , \5241 );
buf \U$4496 ( \5243 , \5242 );
buf \U$4497 ( \5244 , \5243 );
buf \U$4498 ( \5245 , \911 );
nand \U$4499 ( \5246 , \5244 , \5245 );
buf \U$4500 ( \5247 , \5246 );
buf \U$4501 ( \5248 , \5247 );
nand \U$4502 ( \5249 , \5240 , \5248 );
buf \U$4503 ( \5250 , \5249 );
buf \U$4504 ( \5251 , \5250 );
not \U$4505 ( \5252 , \5251 );
buf \U$4506 ( \5253 , \1186 );
not \U$4507 ( \5254 , \5253 );
or \U$4508 ( \5255 , \5252 , \5254 );
buf \U$4509 ( \5256 , \1178 );
not \U$4510 ( \5257 , \5256 );
buf \U$4511 ( \5258 , \3444 );
not \U$4512 ( \5259 , \5258 );
or \U$4513 ( \5260 , \5257 , \5259 );
buf \U$4514 ( \5261 , \4381 );
buf \U$4515 ( \5262 , \911 );
nand \U$4516 ( \5263 , \5261 , \5262 );
buf \U$4517 ( \5264 , \5263 );
buf \U$4518 ( \5265 , \5264 );
nand \U$4519 ( \5266 , \5260 , \5265 );
buf \U$4520 ( \5267 , \5266 );
buf \U$4521 ( \5268 , \5267 );
buf \U$4522 ( \5269 , \1194 );
nand \U$4523 ( \5270 , \5268 , \5269 );
buf \U$4524 ( \5271 , \5270 );
buf \U$4525 ( \5272 , \5271 );
nand \U$4526 ( \5273 , \5255 , \5272 );
buf \U$4527 ( \5274 , \5273 );
buf \U$4528 ( \5275 , \5274 );
xor \U$4529 ( \5276 , \5235 , \5275 );
nand \U$4530 ( \5277 , \1218 , RI9144aa8_96);
nand \U$4531 ( \5278 , RI9144328_80, \950 );
and \U$4532 ( \5279 , \5277 , \5278 );
and \U$4533 ( \5280 , \920 , RI9143428_48);
not \U$4534 ( \5281 , RI9143ba8_64);
nor \U$4535 ( \5282 , \5281 , \927 );
nor \U$4536 ( \5283 , \5280 , \5282 );
nand \U$4537 ( \5284 , \941 , RI9145228_112);
nand \U$4538 ( \5285 , \935 , RI91459a8_128);
and \U$4539 ( \5286 , \5284 , \5285 );
nor \U$4540 ( \5287 , RI9158968_776, RI9158878_774, RI91588f0_775);
and \U$4541 ( \5288 , RI91589e0_777, RI90f37c0_32);
not \U$4542 ( \5289 , RI91589e0_777);
and \U$4543 ( \5290 , \5289 , RI912e848_16);
or \U$4544 ( \5291 , \5288 , \5290 );
nand \U$4545 ( \5292 , \5287 , \5291 );
nand \U$4546 ( \5293 , \5279 , \5283 , \5286 , \5292 );
not \U$4547 ( \5294 , \975 );
nand \U$4548 ( \5295 , \5294 , RI9146128_144);
not \U$4549 ( \5296 , \982 );
nand \U$4550 ( \5297 , \5296 , RI91468a8_160);
and \U$4551 ( \5298 , \5295 , \5297 );
not \U$4552 ( \5299 , \989 );
not \U$4553 ( \5300 , RI9147028_176);
not \U$4554 ( \5301 , \5300 );
and \U$4555 ( \5302 , \5299 , \5301 );
not \U$4556 ( \5303 , RI91477a8_192);
nor \U$4557 ( \5304 , \5303 , \993 );
nor \U$4558 ( \5305 , \5302 , \5304 );
not \U$4559 ( \5306 , \1002 );
not \U$4560 ( \5307 , RI9147f28_208);
not \U$4561 ( \5308 , \5307 );
and \U$4562 ( \5309 , \5306 , \5308 );
not \U$4563 ( \5310 , RI91486a8_224);
nor \U$4564 ( \5311 , \5310 , \1007 );
nor \U$4565 ( \5312 , \5309 , \5311 );
and \U$4566 ( \5313 , \1013 , RI9148e28_240);
not \U$4567 ( \5314 , RI91495a8_256);
nor \U$4568 ( \5315 , \5314 , \1857 );
nor \U$4569 ( \5316 , \5313 , \5315 );
nand \U$4570 ( \5317 , \5298 , \5305 , \5312 , \5316 );
nor \U$4571 ( \5318 , \5293 , \5317 );
not \U$4572 ( \5319 , \5318 );
buf \U$4573 ( \5320 , \5319 );
buf \U$4575 ( \5321 , \5320 );
buf \U$4576 ( \5322 , \5321 );
buf \U$4577 ( \5323 , \1619 );
nand \U$4578 ( \5324 , \5322 , \5323 );
buf \U$4579 ( \5325 , \5324 );
buf \U$4580 ( \5326 , \5325 );
not \U$4581 ( \5327 , \5326 );
buf \U$4582 ( \5328 , \2063 );
not \U$4583 ( \5329 , \5328 );
not \U$4584 ( \5330 , \4794 );
buf \U$4585 ( \5331 , \5330 );
not \U$4586 ( \5332 , \5331 );
or \U$4587 ( \5333 , \5329 , \5332 );
buf \U$4588 ( \5334 , \4202 );
buf \U$4589 ( \5335 , \5334 );
buf \U$4590 ( \5336 , \2078 );
nand \U$4591 ( \5337 , \5335 , \5336 );
buf \U$4592 ( \5338 , \5337 );
buf \U$4593 ( \5339 , \5338 );
nand \U$4594 ( \5340 , \5333 , \5339 );
buf \U$4595 ( \5341 , \5340 );
buf \U$4596 ( \5342 , \5341 );
not \U$4597 ( \5343 , \5342 );
not \U$4598 ( \5344 , RI914b3a8_320);
nor \U$4599 ( \5345 , \5344 , \1122 );
not \U$4600 ( \5346 , RI914ac28_304);
nor \U$4601 ( \5347 , \5346 , \825 );
nor \U$4602 ( \5348 , \5345 , \5347 );
and \U$4603 ( \5349 , \813 , RI914a4a8_288);
and \U$4604 ( \5350 , \1679 , RI9149d28_272);
nor \U$4605 ( \5351 , \5349 , \5350 );
nand \U$4606 ( \5352 , \5348 , \5351 );
and \U$4607 ( \5353 , \1047 , RI914bb28_336);
not \U$4608 ( \5354 , RI914c2a8_352);
nor \U$4609 ( \5355 , \5354 , \1043 );
nor \U$4610 ( \5356 , \5353 , \5355 );
and \U$4611 ( \5357 , \1094 , RI914d1a8_384);
not \U$4612 ( \5358 , RI914ca28_368);
nor \U$4613 ( \5359 , \5358 , \850 );
nor \U$4614 ( \5360 , \5357 , \5359 );
nand \U$4615 ( \5361 , \5356 , \5360 );
nor \U$4616 ( \5362 , \5352 , \5361 );
and \U$4617 ( \5363 , \901 , RI9150628_496);
and \U$4618 ( \5364 , \1087 , RI9150da8_512);
nor \U$4619 ( \5365 , \5363 , \5364 );
not \U$4620 ( \5366 , RI914f728_464);
nor \U$4621 ( \5367 , \5366 , \1139 );
and \U$4622 ( \5368 , \1080 , RI914fea8_480);
nor \U$4623 ( \5369 , \5367 , \5368 );
nand \U$4624 ( \5370 , \5365 , \5369 );
and \U$4625 ( \5371 , \1062 , RI914e0a8_416);
not \U$4626 ( \5372 , RI914d928_400);
nor \U$4627 ( \5373 , \5372 , \864 );
nor \U$4628 ( \5374 , \5371 , \5373 );
not \U$4629 ( \5375 , RI914e828_432);
nor \U$4630 ( \5376 , \5375 , \1386 );
not \U$4631 ( \5377 , RI914efa8_448);
nor \U$4632 ( \5378 , \5377 , \884 );
nor \U$4633 ( \5379 , \5376 , \5378 );
nand \U$4634 ( \5380 , \5374 , \5379 );
nor \U$4635 ( \5381 , \5370 , \5380 );
nand \U$4636 ( \5382 , \5362 , \5381 );
buf \U$4637 ( \5383 , \5382 );
not \U$4638 ( \5384 , \5383 );
buf \U$4639 ( \5385 , \4794 );
nand \U$4640 ( \5386 , \5384 , \5385 );
buf \U$4641 ( \5387 , \5386 );
buf \U$4644 ( \5388 , \5387 );
buf \U$4645 ( \5389 , \5388 );
not \U$4646 ( \5390 , \5389 );
buf \U$4647 ( \5391 , \5390 );
buf \U$4648 ( \5392 , \5391 );
not \U$4649 ( \5393 , \5392 );
or \U$4650 ( \5394 , \5343 , \5393 );
buf \U$4651 ( \5395 , \4794 );
buf \U$4652 ( \5396 , \5382 );
buf \U$4654 ( \5397 , \5396 );
buf \U$4657 ( \5398 , \5397 );
buf \U$4658 ( \5399 , \5398 );
nand \U$4659 ( \5400 , \5395 , \5399 );
buf \U$4660 ( \5401 , \5400 );
buf \U$4661 ( \5402 , \5401 );
nand \U$4662 ( \5403 , \5394 , \5402 );
buf \U$4663 ( \5404 , \5403 );
buf \U$4664 ( \5405 , \5404 );
not \U$4665 ( \5406 , \5405 );
or \U$4666 ( \5407 , \5327 , \5406 );
buf \U$4667 ( \5408 , \5404 );
buf \U$4668 ( \5409 , \5325 );
or \U$4669 ( \5410 , \5408 , \5409 );
nand \U$4670 ( \5411 , \5407 , \5410 );
buf \U$4671 ( \5412 , \5411 );
buf \U$4672 ( \5413 , \5412 );
and \U$4673 ( \5414 , \5276 , \5413 );
and \U$4674 ( \5415 , \5235 , \5275 );
or \U$4675 ( \5416 , \5414 , \5415 );
buf \U$4676 ( \5417 , \5416 );
buf \U$4677 ( \5418 , \5417 );
not \U$4678 ( \5419 , \5418 );
buf \U$4679 ( \5420 , \5419 );
not \U$4680 ( \5421 , \5420 );
or \U$4681 ( \5422 , \5209 , \5421 );
not \U$4682 ( \5423 , RI9154a20_641);
nor \U$4683 ( \5424 , \5423 , \976 );
not \U$4684 ( \5425 , RI91551a0_657);
nor \U$4685 ( \5426 , \5425 , \983 );
nor \U$4686 ( \5427 , \5424 , \5426 );
not \U$4687 ( \5428 , \1205 );
and \U$4688 ( \5429 , \5428 , RI9155920_673);
buf \U$4689 ( \5430 , \1213 );
and \U$4690 ( \5431 , \5430 , RI91560a0_689);
nor \U$4691 ( \5432 , \5429 , \5431 );
nand \U$4692 ( \5433 , \5427 , \5432 );
not \U$4693 ( \5434 , \1524 );
and \U$4694 ( \5435 , \5434 , RI9156820_705);
and \U$4695 ( \5436 , \2052 , RI9156fa0_721);
nor \U$4696 ( \5437 , \5435 , \5436 );
and \U$4697 ( \5438 , \1014 , RI9157720_737);
not \U$4698 ( \5439 , \1250 );
and \U$4699 ( \5440 , \5439 , RI9157ea0_753);
nor \U$4700 ( \5441 , \5438 , \5440 );
nand \U$4701 ( \5442 , \5437 , \5441 );
nor \U$4702 ( \5443 , \5433 , \5442 );
not \U$4703 ( \5444 , \929 );
not \U$4704 ( \5445 , RI91524a0_561);
not \U$4705 ( \5446 , \5445 );
and \U$4706 ( \5447 , \5444 , \5446 );
not \U$4707 ( \5448 , RI9151d20_545);
nor \U$4708 ( \5449 , \5448 , \922 );
nor \U$4709 ( \5450 , \5447 , \5449 );
buf \U$4710 ( \5451 , \943 );
and \U$4711 ( \5452 , \5451 , RI9153b20_609);
buf \U$4712 ( \5453 , \1291 );
and \U$4713 ( \5454 , \5453 , RI91542a0_625);
nor \U$4714 ( \5455 , \5452 , \5454 );
nand \U$4715 ( \5456 , \5450 , \5455 );
and \U$4716 ( \5457 , \1635 , RI91533a0_593);
not \U$4717 ( \5458 , RI9152c20_577);
nor \U$4718 ( \5459 , \5458 , \1282 );
nor \U$4719 ( \5460 , \5457 , \5459 );
and \U$4720 ( \5461 , \963 , RI91515a0_529);
not \U$4721 ( \5462 , RI9150e20_513);
buf \U$4722 ( \5463 , \968 );
not \U$4723 ( \5464 , \5463 );
nor \U$4724 ( \5465 , \5462 , \5464 );
nor \U$4725 ( \5466 , \5461 , \5465 );
nand \U$4726 ( \5467 , \5460 , \5466 );
nor \U$4727 ( \5468 , \5456 , \5467 );
nand \U$4728 ( \5469 , \5443 , \5468 );
buf \U$4729 ( \5470 , \5469 );
buf \U$4730 ( \5471 , \5319 );
buf \U$4732 ( \5472 , \5471 );
buf \U$4733 ( \5473 , \5472 );
not \U$4734 ( \5474 , \5473 );
buf \U$4735 ( \5475 , \5474 );
buf \U$4736 ( \5476 , \5475 );
buf \U$4737 ( \5477 , \1745 );
nand \U$4738 ( \5478 , \5476 , \5477 );
buf \U$4739 ( \5479 , \5478 );
buf \U$4740 ( \5480 , \5479 );
buf \U$4741 ( \5481 , \3329 );
and \U$4742 ( \5482 , \5480 , \5481 );
buf \U$4743 ( \5483 , \1745 );
not \U$4744 ( \5484 , \5483 );
buf \U$4745 ( \5485 , \5484 );
buf \U$4746 ( \5486 , \5485 );
not \U$4747 ( \5487 , \5486 );
buf \U$4748 ( \5488 , \5472 );
not \U$4749 ( \5489 , \5488 );
or \U$4750 ( \5490 , \5487 , \5489 );
buf \U$4751 ( \5491 , \1737 );
not \U$4752 ( \5492 , \5491 );
buf \U$4753 ( \5493 , \5492 );
buf \U$4754 ( \5494 , \5493 );
nand \U$4755 ( \5495 , \5490 , \5494 );
buf \U$4756 ( \5496 , \5495 );
buf \U$4757 ( \5497 , \5496 );
nor \U$4758 ( \5498 , \5482 , \5497 );
buf \U$4759 ( \5499 , \5498 );
buf \U$4760 ( \5500 , \5499 );
xor \U$4761 ( \5501 , \5470 , \5500 );
buf \U$4762 ( \5502 , \5501 );
buf \U$4763 ( \5503 , \5502 );
buf \U$4764 ( \5504 , \5387 );
not \U$4765 ( \5505 , \5504 );
buf \U$4766 ( \5506 , \5505 );
buf \U$4767 ( \5507 , \5506 );
not \U$4768 ( \5508 , \5507 );
buf \U$4769 ( \5509 , \1542 );
not \U$4770 ( \5510 , \5509 );
buf \U$4771 ( \5511 , \4795 );
not \U$4772 ( \5512 , \5511 );
or \U$4773 ( \5513 , \5510 , \5512 );
buf \U$4774 ( \5514 , \4794 );
buf \U$4775 ( \5515 , \1539 );
nand \U$4776 ( \5516 , \5514 , \5515 );
buf \U$4777 ( \5517 , \5516 );
buf \U$4778 ( \5518 , \5517 );
nand \U$4779 ( \5519 , \5513 , \5518 );
buf \U$4780 ( \5520 , \5519 );
buf \U$4781 ( \5521 , \5520 );
not \U$4782 ( \5522 , \5521 );
or \U$4783 ( \5523 , \5508 , \5522 );
buf \U$4784 ( \5524 , \5341 );
buf \U$4785 ( \5525 , \5398 );
nand \U$4786 ( \5526 , \5524 , \5525 );
buf \U$4787 ( \5527 , \5526 );
buf \U$4788 ( \5528 , \5527 );
nand \U$4789 ( \5529 , \5523 , \5528 );
buf \U$4790 ( \5530 , \5529 );
buf \U$4791 ( \5531 , \5530 );
or \U$4792 ( \5532 , \5503 , \5531 );
buf \U$4793 ( \5533 , \1795 );
not \U$4794 ( \5534 , \5533 );
buf \U$4795 ( \5535 , \2479 );
not \U$4796 ( \5536 , \5535 );
or \U$4797 ( \5537 , \5534 , \5536 );
buf \U$4798 ( \5538 , \1792 );
buf \U$4799 ( \5539 , \4070 );
nand \U$4800 ( \5540 , \5538 , \5539 );
buf \U$4801 ( \5541 , \5540 );
buf \U$4802 ( \5542 , \5541 );
nand \U$4803 ( \5543 , \5537 , \5542 );
buf \U$4804 ( \5544 , \5543 );
buf \U$4805 ( \5545 , \5544 );
not \U$4806 ( \5546 , \5545 );
buf \U$4807 ( \5547 , \3288 );
not \U$4808 ( \5548 , \5547 );
or \U$4809 ( \5549 , \5546 , \5548 );
buf \U$4810 ( \5550 , \5029 );
buf \U$4811 ( \5551 , \2473 );
nand \U$4812 ( \5552 , \5550 , \5551 );
buf \U$4813 ( \5553 , \5552 );
buf \U$4814 ( \5554 , \5553 );
nand \U$4815 ( \5555 , \5549 , \5554 );
buf \U$4816 ( \5556 , \5555 );
buf \U$4817 ( \5557 , \5556 );
nand \U$4818 ( \5558 , \5532 , \5557 );
buf \U$4819 ( \5559 , \5558 );
buf \U$4820 ( \5560 , \5559 );
buf \U$4821 ( \5561 , \5502 );
buf \U$4822 ( \5562 , \5530 );
nand \U$4823 ( \5563 , \5561 , \5562 );
buf \U$4824 ( \5564 , \5563 );
buf \U$4825 ( \5565 , \5564 );
nand \U$4826 ( \5566 , \5560 , \5565 );
buf \U$4827 ( \5567 , \5566 );
buf \U$4828 ( \5568 , \5567 );
buf \U$4829 ( \5569 , \1618 );
not \U$4830 ( \5570 , \5569 );
buf \U$4831 ( \5571 , \5321 );
not \U$4832 ( \5572 , \5571 );
buf \U$4833 ( \5573 , \5572 );
buf \U$4834 ( \5574 , \5573 );
not \U$4835 ( \5575 , \5574 );
or \U$4836 ( \5576 , \5570 , \5575 );
buf \U$4837 ( \5577 , \5321 );
buf \U$4838 ( \5578 , \3465 );
nand \U$4839 ( \5579 , \5577 , \5578 );
buf \U$4840 ( \5580 , \5579 );
buf \U$4841 ( \5581 , \5580 );
nand \U$4842 ( \5582 , \5576 , \5581 );
buf \U$4843 ( \5583 , \5582 );
buf \U$4844 ( \5584 , \5583 );
not \U$4845 ( \5585 , \5584 );
buf \U$4846 ( \5586 , \1758 );
not \U$4847 ( \5587 , \5586 );
or \U$4848 ( \5588 , \5585 , \5587 );
buf \U$4849 ( \5589 , \5001 );
buf \U$4850 ( \5590 , \1882 );
nand \U$4851 ( \5591 , \5589 , \5590 );
buf \U$4852 ( \5592 , \5591 );
buf \U$4853 ( \5593 , \5592 );
nand \U$4854 ( \5594 , \5588 , \5593 );
buf \U$4855 ( \5595 , \5594 );
buf \U$4856 ( \5596 , \5595 );
not \U$4857 ( \5597 , \5596 );
buf \U$4858 ( \5598 , \2521 );
not \U$4859 ( \5599 , \5598 );
buf \U$4860 ( \5600 , \4516 );
not \U$4861 ( \5601 , \5600 );
or \U$4862 ( \5602 , \5599 , \5601 );
buf \U$4865 ( \5603 , \4100 );
buf \U$4866 ( \5604 , \5603 );
buf \U$4867 ( \5605 , \1999 );
nand \U$4868 ( \5606 , \5604 , \5605 );
buf \U$4869 ( \5607 , \5606 );
buf \U$4870 ( \5608 , \5607 );
nand \U$4871 ( \5609 , \5602 , \5608 );
buf \U$4872 ( \5610 , \5609 );
buf \U$4873 ( \5611 , \5610 );
not \U$4874 ( \5612 , \5611 );
buf \U$4875 ( \5613 , \3124 );
not \U$4876 ( \5614 , \5613 );
buf \U$4877 ( \5615 , \5614 );
buf \U$4878 ( \5616 , \5615 );
not \U$4879 ( \5617 , \5616 );
or \U$4880 ( \5618 , \5612 , \5617 );
buf \U$4881 ( \5619 , \1024 );
not \U$4882 ( \5620 , \5619 );
buf \U$4883 ( \5621 , \5620 );
buf \U$4884 ( \5622 , \5621 );
not \U$4885 ( \5623 , \5622 );
buf \U$4886 ( \5624 , \4516 );
not \U$4887 ( \5625 , \5624 );
or \U$4888 ( \5626 , \5623 , \5625 );
buf \U$4889 ( \5627 , \5603 );
buf \U$4890 ( \5628 , \1024 );
nand \U$4891 ( \5629 , \5627 , \5628 );
buf \U$4892 ( \5630 , \5629 );
buf \U$4893 ( \5631 , \5630 );
nand \U$4894 ( \5632 , \5626 , \5631 );
buf \U$4895 ( \5633 , \5632 );
buf \U$4896 ( \5634 , \5633 );
buf \U$4897 ( \5635 , \3095 );
nand \U$4898 ( \5636 , \5634 , \5635 );
buf \U$4899 ( \5637 , \5636 );
buf \U$4900 ( \5638 , \5637 );
nand \U$4901 ( \5639 , \5618 , \5638 );
buf \U$4902 ( \5640 , \5639 );
buf \U$4903 ( \5641 , \5640 );
not \U$4904 ( \5642 , \5641 );
or \U$4905 ( \5643 , \5597 , \5642 );
buf \U$4906 ( \5644 , \5640 );
buf \U$4907 ( \5645 , \5595 );
or \U$4908 ( \5646 , \5644 , \5645 );
buf \U$4909 ( \5647 , \1178 );
not \U$4910 ( \5648 , \5647 );
buf \U$4911 ( \5649 , \4678 );
not \U$4912 ( \5650 , \5649 );
or \U$4913 ( \5651 , \5648 , \5650 );
buf \U$4914 ( \5652 , \4863 );
buf \U$4915 ( \5653 , \911 );
nand \U$4916 ( \5654 , \5652 , \5653 );
buf \U$4917 ( \5655 , \5654 );
buf \U$4918 ( \5656 , \5655 );
nand \U$4919 ( \5657 , \5651 , \5656 );
buf \U$4920 ( \5658 , \5657 );
buf \U$4921 ( \5659 , \5658 );
not \U$4922 ( \5660 , \5659 );
buf \U$4923 ( \5661 , \1186 );
not \U$4924 ( \5662 , \5661 );
or \U$4925 ( \5663 , \5660 , \5662 );
buf \U$4926 ( \5664 , \5250 );
buf \U$4927 ( \5665 , \1194 );
nand \U$4928 ( \5666 , \5664 , \5665 );
buf \U$4929 ( \5667 , \5666 );
buf \U$4930 ( \5668 , \5667 );
nand \U$4931 ( \5669 , \5663 , \5668 );
buf \U$4932 ( \5670 , \5669 );
buf \U$4933 ( \5671 , \5670 );
nand \U$4934 ( \5672 , \5646 , \5671 );
buf \U$4935 ( \5673 , \5672 );
buf \U$4936 ( \5674 , \5673 );
nand \U$4937 ( \5675 , \5643 , \5674 );
buf \U$4938 ( \5676 , \5675 );
buf \U$4939 ( \5677 , \5676 );
xor \U$4940 ( \5678 , \5568 , \5677 );
buf \U$4941 ( \5679 , \2758 );
not \U$4942 ( \5680 , \5679 );
buf \U$4943 ( \5681 , \2488 );
not \U$4944 ( \5682 , \5681 );
or \U$4945 ( \5683 , \5680 , \5682 );
buf \U$4946 ( \5684 , \2068 );
buf \U$4947 ( \5685 , \2853 );
nand \U$4948 ( \5686 , \5684 , \5685 );
buf \U$4949 ( \5687 , \5686 );
buf \U$4950 ( \5688 , \5687 );
nand \U$4951 ( \5689 , \5683 , \5688 );
buf \U$4952 ( \5690 , \5689 );
buf \U$4953 ( \5691 , \5690 );
not \U$4954 ( \5692 , \5691 );
buf \U$4955 ( \5693 , \2200 );
not \U$4956 ( \5694 , \5693 );
or \U$4957 ( \5695 , \5692 , \5694 );
buf \U$4958 ( \5696 , \2214 );
and \U$4959 ( \5697 , \1669 , \2488 );
not \U$4960 ( \5698 , \1669 );
and \U$4961 ( \5699 , \5698 , \2068 );
or \U$4962 ( \5700 , \5697 , \5699 );
buf \U$4963 ( \5701 , \5700 );
nand \U$4964 ( \5702 , \5696 , \5701 );
buf \U$4965 ( \5703 , \5702 );
buf \U$4966 ( \5704 , \5703 );
nand \U$4967 ( \5705 , \5695 , \5704 );
buf \U$4968 ( \5706 , \5705 );
not \U$4969 ( \5707 , \5706 );
buf \U$4970 ( \5708 , \3444 );
not \U$4971 ( \5709 , \5708 );
buf \U$4972 ( \5710 , \2273 );
not \U$4973 ( \5711 , \5710 );
or \U$4974 ( \5712 , \5709 , \5711 );
buf \U$4975 ( \5713 , \1337 );
buf \U$4976 ( \5714 , \4381 );
nand \U$4977 ( \5715 , \5713 , \5714 );
buf \U$4978 ( \5716 , \5715 );
buf \U$4979 ( \5717 , \5716 );
nand \U$4980 ( \5718 , \5712 , \5717 );
buf \U$4981 ( \5719 , \5718 );
buf \U$4982 ( \5720 , \5719 );
not \U$4983 ( \5721 , \5720 );
buf \U$4984 ( \5722 , \1472 );
not \U$4985 ( \5723 , \5722 );
or \U$4986 ( \5724 , \5721 , \5723 );
buf \U$4987 ( \5725 , \5221 );
buf \U$4988 ( \5726 , \1904 );
nand \U$4989 ( \5727 , \5725 , \5726 );
buf \U$4990 ( \5728 , \5727 );
buf \U$4991 ( \5729 , \5728 );
nand \U$4992 ( \5730 , \5724 , \5729 );
buf \U$4993 ( \5731 , \5730 );
not \U$4994 ( \5732 , \5731 );
or \U$4995 ( \5733 , \5707 , \5732 );
buf \U$4996 ( \5734 , \5731 );
not \U$4997 ( \5735 , \5734 );
buf \U$4998 ( \5736 , \5735 );
not \U$4999 ( \5737 , \5736 );
buf \U$5000 ( \5738 , \5706 );
not \U$5001 ( \5739 , \5738 );
buf \U$5002 ( \5740 , \5739 );
not \U$5003 ( \5741 , \5740 );
or \U$5004 ( \5742 , \5737 , \5741 );
buf \U$5005 ( \5743 , \5128 );
not \U$5006 ( \5744 , \5743 );
buf \U$5007 ( \5745 , \4281 );
not \U$5008 ( \5746 , \5745 );
or \U$5009 ( \5747 , \5744 , \5746 );
buf \U$5010 ( \5748 , \4278 );
buf \U$5011 ( \5749 , \1258 );
nand \U$5012 ( \5750 , \5748 , \5749 );
buf \U$5013 ( \5751 , \5750 );
buf \U$5014 ( \5752 , \5751 );
nand \U$5015 ( \5753 , \5747 , \5752 );
buf \U$5016 ( \5754 , \5753 );
buf \U$5017 ( \5755 , \5754 );
not \U$5018 ( \5756 , \5755 );
buf \U$5019 ( \5757 , \4543 );
not \U$5020 ( \5758 , \5757 );
or \U$5021 ( \5759 , \5756 , \5758 );
buf \U$5022 ( \5760 , \4581 );
buf \U$5023 ( \5761 , \5059 );
nand \U$5024 ( \5762 , \5760 , \5761 );
buf \U$5025 ( \5763 , \5762 );
buf \U$5026 ( \5764 , \5763 );
nand \U$5027 ( \5765 , \5759 , \5764 );
buf \U$5028 ( \5766 , \5765 );
nand \U$5029 ( \5767 , \5742 , \5766 );
nand \U$5030 ( \5768 , \5733 , \5767 );
buf \U$5031 ( \5769 , \5768 );
and \U$5032 ( \5770 , \5678 , \5769 );
and \U$5033 ( \5771 , \5568 , \5677 );
or \U$5034 ( \5772 , \5770 , \5771 );
buf \U$5035 ( \5773 , \5772 );
nand \U$5036 ( \5774 , \5422 , \5773 );
buf \U$5037 ( \5775 , \5208 );
buf \U$5038 ( \5776 , \5420 );
or \U$5039 ( \5777 , \5775 , \5776 );
buf \U$5040 ( \5778 , \5777 );
nand \U$5041 ( \5779 , \5774 , \5778 );
buf \U$5042 ( \5780 , \5779 );
nand \U$5043 ( \5781 , \5202 , \5780 );
buf \U$5044 ( \5782 , \5781 );
buf \U$5045 ( \5783 , \5782 );
nand \U$5046 ( \5784 , \5199 , \5783 );
buf \U$5047 ( \5785 , \5784 );
buf \U$5048 ( \5786 , \5785 );
xor \U$5049 ( \5787 , \4965 , \5786 );
buf \U$5050 ( \5788 , \4593 );
buf \U$5051 ( \5789 , \4735 );
xor \U$5052 ( \5790 , \5788 , \5789 );
buf \U$5053 ( \5791 , \4726 );
xnor \U$5054 ( \5792 , \5790 , \5791 );
buf \U$5055 ( \5793 , \5792 );
buf \U$5056 ( \5794 , \5793 );
not \U$5057 ( \5795 , \5794 );
buf \U$5058 ( \5796 , \5795 );
buf \U$5059 ( \5797 , \5796 );
not \U$5060 ( \5798 , \5797 );
xor \U$5061 ( \5799 , \5099 , \5182 );
and \U$5062 ( \5800 , \5799 , \5194 );
and \U$5063 ( \5801 , \5099 , \5182 );
or \U$5064 ( \5802 , \5800 , \5801 );
buf \U$5065 ( \5803 , \5802 );
not \U$5066 ( \5804 , \5803 );
buf \U$5067 ( \5805 , \5804 );
not \U$5068 ( \5806 , \5805 );
or \U$5069 ( \5807 , \5798 , \5806 );
buf \U$5070 ( \5808 , \5793 );
buf \U$5071 ( \5809 , \5803 );
nand \U$5072 ( \5810 , \5808 , \5809 );
buf \U$5073 ( \5811 , \5810 );
buf \U$5074 ( \5812 , \5811 );
nand \U$5075 ( \5813 , \5807 , \5812 );
buf \U$5076 ( \5814 , \5813 );
buf \U$5077 ( \5815 , \5814 );
and \U$5078 ( \5816 , \4623 , \4681 );
not \U$5079 ( \5817 , \4623 );
and \U$5080 ( \5818 , \5817 , \4684 );
nor \U$5081 ( \5819 , \5816 , \5818 );
xor \U$5082 ( \5820 , \5819 , \4708 );
buf \U$5083 ( \5821 , \5820 );
not \U$5084 ( \5822 , \5821 );
xor \U$5085 ( \5823 , \4793 , \4818 );
xor \U$5086 ( \5824 , \5823 , \4915 );
buf \U$5087 ( \5825 , \5824 );
buf \U$5088 ( \5826 , \5825 );
not \U$5089 ( \5827 , \5826 );
or \U$5090 ( \5828 , \5822 , \5827 );
buf \U$5091 ( \5829 , \5825 );
buf \U$5092 ( \5830 , \5820 );
or \U$5093 ( \5831 , \5829 , \5830 );
buf \U$5094 ( \5832 , \1186 );
not \U$5095 ( \5833 , \5832 );
buf \U$5096 ( \5834 , \5267 );
not \U$5097 ( \5835 , \5834 );
or \U$5098 ( \5836 , \5833 , \5835 );
buf \U$5099 ( \5837 , \1194 );
buf \U$5100 ( \5838 , \4449 );
nand \U$5101 ( \5839 , \5837 , \5838 );
buf \U$5102 ( \5840 , \5839 );
buf \U$5103 ( \5841 , \5840 );
nand \U$5104 ( \5842 , \5836 , \5841 );
buf \U$5105 ( \5843 , \5842 );
buf \U$5106 ( \5844 , \5843 );
not \U$5107 ( \5845 , \5844 );
buf \U$5108 ( \5846 , \5325 );
not \U$5109 ( \5847 , \5846 );
buf \U$5112 ( \5848 , \5404 );
buf \U$5113 ( \5849 , \5848 );
nand \U$5114 ( \5850 , \5847 , \5849 );
buf \U$5115 ( \5851 , \5850 );
buf \U$5116 ( \5852 , \5851 );
nand \U$5117 ( \5853 , \5845 , \5852 );
buf \U$5118 ( \5854 , \5853 );
buf \U$5119 ( \5855 , \5854 );
not \U$5120 ( \5856 , \5855 );
and \U$5121 ( \5857 , \5470 , \5500 );
buf \U$5122 ( \5858 , \5857 );
buf \U$5123 ( \5859 , \5858 );
buf \U$5124 ( \5860 , \5700 );
not \U$5125 ( \5861 , \5860 );
buf \U$5126 ( \5862 , \2200 );
not \U$5127 ( \5863 , \5862 );
or \U$5128 ( \5864 , \5861 , \5863 );
buf \U$5129 ( \5865 , \2897 );
buf \U$5130 ( \5866 , \4808 );
nand \U$5131 ( \5867 , \5865 , \5866 );
buf \U$5132 ( \5868 , \5867 );
buf \U$5133 ( \5869 , \5868 );
nand \U$5134 ( \5870 , \5864 , \5869 );
buf \U$5135 ( \5871 , \5870 );
buf \U$5136 ( \5872 , \5871 );
xor \U$5137 ( \5873 , \5859 , \5872 );
buf \U$5138 ( \5874 , \5633 );
not \U$5139 ( \5875 , \5874 );
buf \U$5140 ( \5876 , \5615 );
not \U$5141 ( \5877 , \5876 );
or \U$5142 ( \5878 , \5875 , \5877 );
buf \U$5143 ( \5879 , \3095 );
buf \U$5144 ( \5880 , \5140 );
nand \U$5145 ( \5881 , \5879 , \5880 );
buf \U$5146 ( \5882 , \5881 );
buf \U$5147 ( \5883 , \5882 );
nand \U$5148 ( \5884 , \5878 , \5883 );
buf \U$5149 ( \5885 , \5884 );
buf \U$5150 ( \5886 , \5885 );
and \U$5151 ( \5887 , \5873 , \5886 );
and \U$5152 ( \5888 , \5859 , \5872 );
or \U$5153 ( \5889 , \5887 , \5888 );
buf \U$5154 ( \5890 , \5889 );
buf \U$5155 ( \5891 , \5890 );
not \U$5156 ( \5892 , \5891 );
or \U$5157 ( \5893 , \5856 , \5892 );
buf \U$5158 ( \5894 , \5851 );
not \U$5159 ( \5895 , \5894 );
buf \U$5160 ( \5896 , \5843 );
nand \U$5161 ( \5897 , \5895 , \5896 );
buf \U$5162 ( \5898 , \5897 );
buf \U$5163 ( \5899 , \5898 );
nand \U$5164 ( \5900 , \5893 , \5899 );
buf \U$5165 ( \5901 , \5900 );
buf \U$5166 ( \5902 , \5901 );
nand \U$5167 ( \5903 , \5831 , \5902 );
buf \U$5168 ( \5904 , \5903 );
buf \U$5169 ( \5905 , \5904 );
nand \U$5170 ( \5906 , \5828 , \5905 );
buf \U$5171 ( \5907 , \5906 );
buf \U$5172 ( \5908 , \5907 );
not \U$5173 ( \5909 , \5908 );
buf \U$5174 ( \5910 , \5909 );
buf \U$5175 ( \5911 , \5910 );
and \U$5176 ( \5912 , \5815 , \5911 );
not \U$5177 ( \5913 , \5815 );
buf \U$5178 ( \5914 , \5907 );
and \U$5179 ( \5915 , \5913 , \5914 );
nor \U$5180 ( \5916 , \5912 , \5915 );
buf \U$5181 ( \5917 , \5916 );
not \U$5182 ( \5918 , \5917 );
buf \U$5183 ( \5919 , \5918 );
xnor \U$5184 ( \5920 , \5787 , \5919 );
buf \U$5185 ( \5921 , \5920 );
buf \U$5186 ( \5922 , \5921 );
buf \U$5187 ( \5923 , \5820 );
buf \U$5188 ( \5924 , \5901 );
xor \U$5189 ( \5925 , \5923 , \5924 );
buf \U$5190 ( \5926 , \5825 );
xnor \U$5191 ( \5927 , \5925 , \5926 );
buf \U$5192 ( \5928 , \5927 );
buf \U$5193 ( \5929 , \5928 );
buf \U$5194 ( \5930 , \5325 );
not \U$5195 ( \5931 , \5930 );
buf \U$5196 ( \5932 , \5848 );
nand \U$5197 ( \5933 , \5931 , \5932 );
buf \U$5198 ( \5934 , \5933 );
buf \U$5199 ( \5935 , \5934 );
not \U$5200 ( \5936 , \5935 );
buf \U$5201 ( \5937 , \5843 );
not \U$5202 ( \5938 , \5937 );
and \U$5203 ( \5939 , \5936 , \5938 );
buf \U$5204 ( \5940 , \5851 );
buf \U$5205 ( \5941 , \5843 );
and \U$5206 ( \5942 , \5940 , \5941 );
nor \U$5207 ( \5943 , \5939 , \5942 );
buf \U$5208 ( \5944 , \5943 );
buf \U$5209 ( \5945 , \5944 );
not \U$5210 ( \5946 , \5945 );
buf \U$5211 ( \5947 , \5890 );
not \U$5212 ( \5948 , \5947 );
and \U$5213 ( \5949 , \5946 , \5948 );
buf \U$5214 ( \5950 , \5890 );
buf \U$5215 ( \5951 , \5944 );
and \U$5216 ( \5952 , \5950 , \5951 );
nor \U$5217 ( \5953 , \5949 , \5952 );
buf \U$5218 ( \5954 , \5953 );
buf \U$5219 ( \5955 , \5954 );
not \U$5220 ( \5956 , \5955 );
xor \U$5221 ( \5957 , \5235 , \5275 );
xor \U$5222 ( \5958 , \5957 , \5413 );
buf \U$5223 ( \5959 , \5958 );
buf \U$5224 ( \5960 , \5959 );
not \U$5225 ( \5961 , \5960 );
xor \U$5226 ( \5962 , \5859 , \5872 );
xor \U$5227 ( \5963 , \5962 , \5886 );
buf \U$5228 ( \5964 , \5963 );
buf \U$5229 ( \5965 , \5964 );
not \U$5230 ( \5966 , \5965 );
or \U$5231 ( \5967 , \5961 , \5966 );
buf \U$5232 ( \5968 , \5964 );
buf \U$5233 ( \5969 , \5959 );
or \U$5234 ( \5970 , \5968 , \5969 );
xor \U$5235 ( \5971 , \5014 , \5042 );
xor \U$5236 ( \5972 , \5971 , \5086 );
buf \U$5237 ( \5973 , \5972 );
buf \U$5238 ( \5974 , \5973 );
nand \U$5239 ( \5975 , \5970 , \5974 );
buf \U$5240 ( \5976 , \5975 );
buf \U$5241 ( \5977 , \5976 );
nand \U$5242 ( \5978 , \5967 , \5977 );
buf \U$5243 ( \5979 , \5978 );
buf \U$5244 ( \5980 , \5979 );
not \U$5245 ( \5981 , \5980 );
buf \U$5246 ( \5982 , \5981 );
buf \U$5247 ( \5983 , \5982 );
not \U$5248 ( \5984 , \5983 );
or \U$5249 ( \5985 , \5956 , \5984 );
and \U$5250 ( \5986 , \5090 , \4984 );
not \U$5251 ( \5987 , \5090 );
and \U$5252 ( \5988 , \5987 , \4978 );
nor \U$5253 ( \5989 , \5986 , \5988 );
buf \U$5256 ( \5990 , \4971 );
xor \U$5257 ( \5991 , \5989 , \5990 );
buf \U$5258 ( \5992 , \5991 );
nand \U$5259 ( \5993 , \5985 , \5992 );
buf \U$5260 ( \5994 , \5993 );
buf \U$5261 ( \5995 , \5994 );
buf \U$5262 ( \5996 , \5954 );
not \U$5263 ( \5997 , \5996 );
buf \U$5264 ( \5998 , \5979 );
nand \U$5265 ( \5999 , \5997 , \5998 );
buf \U$5266 ( \6000 , \5999 );
buf \U$5267 ( \6001 , \6000 );
and \U$5268 ( \6002 , \5995 , \6001 );
buf \U$5269 ( \6003 , \6002 );
buf \U$5270 ( \6004 , \6003 );
xor \U$5271 ( \6005 , \5929 , \6004 );
buf \U$5272 ( \6006 , \5092 );
buf \U$5273 ( \6007 , \5196 );
xor \U$5274 ( \6008 , \6006 , \6007 );
buf \U$5275 ( \6009 , \5779 );
xnor \U$5276 ( \6010 , \6008 , \6009 );
buf \U$5277 ( \6011 , \6010 );
buf \U$5278 ( \6012 , \6011 );
and \U$5279 ( \6013 , \6005 , \6012 );
and \U$5280 ( \6014 , \5929 , \6004 );
or \U$5281 ( \6015 , \6013 , \6014 );
buf \U$5282 ( \6016 , \6015 );
buf \U$5283 ( \6017 , \6016 );
or \U$5284 ( \6018 , \5922 , \6017 );
buf \U$5285 ( \6019 , \6018 );
buf \U$5286 ( \6020 , \6019 );
nand \U$5287 ( \6021 , \4958 , \6020 );
buf \U$5288 ( \6022 , \6021 );
buf \U$5289 ( \6023 , \6022 );
buf \U$5290 ( \6024 , \5921 );
buf \U$5291 ( \6025 , \6016 );
nand \U$5292 ( \6026 , \6024 , \6025 );
buf \U$5293 ( \6027 , \6026 );
buf \U$5294 ( \6028 , \6027 );
xor \U$5295 ( \6029 , \5929 , \6004 );
xor \U$5296 ( \6030 , \6029 , \6012 );
buf \U$5297 ( \6031 , \6030 );
buf \U$5298 ( \6032 , \6031 );
buf \U$5299 ( \6033 , \5954 );
buf \U$5300 ( \6034 , \5979 );
xor \U$5301 ( \6035 , \6033 , \6034 );
buf \U$5302 ( \6036 , \5991 );
xnor \U$5303 ( \6037 , \6035 , \6036 );
buf \U$5304 ( \6038 , \6037 );
buf \U$5305 ( \6039 , \6038 );
xor \U$5306 ( \6040 , \5417 , \5208 );
xor \U$5307 ( \6041 , \6040 , \5773 );
buf \U$5308 ( \6042 , \6041 );
not \U$5309 ( \6043 , \6042 );
buf \U$5310 ( \6044 , \6043 );
buf \U$5311 ( \6045 , \6044 );
or \U$5312 ( \6046 , \6039 , \6045 );
not \U$5313 ( \6047 , RI9154a98_642);
nor \U$5314 ( \6048 , \6047 , \976 );
not \U$5315 ( \6049 , RI9155218_658);
nor \U$5316 ( \6050 , \6049 , \983 );
nor \U$5317 ( \6051 , \6048 , \6050 );
not \U$5318 ( \6052 , \1205 );
and \U$5319 ( \6053 , \6052 , RI9155998_674);
and \U$5320 ( \6054 , \5430 , RI9156118_690);
nor \U$5321 ( \6055 , \6053 , \6054 );
and \U$5322 ( \6056 , \4003 , RI9156898_706);
and \U$5323 ( \6057 , \2052 , RI9157018_722);
nor \U$5324 ( \6058 , \6056 , \6057 );
and \U$5325 ( \6059 , \1014 , RI9157798_738);
and \U$5326 ( \6060 , \5439 , RI9157f18_754);
nor \U$5327 ( \6061 , \6059 , \6060 );
and \U$5328 ( \6062 , \6051 , \6055 , \6058 , \6061 );
not \U$5329 ( \6063 , RI9152c98_578);
nor \U$5330 ( \6064 , \6063 , \1282 );
not \U$5331 ( \6065 , RI9153418_594);
nor \U$5332 ( \6066 , \6065 , \957 );
nor \U$5333 ( \6067 , \6064 , \6066 );
not \U$5334 ( \6068 , RI9153b98_610);
not \U$5335 ( \6069 , \1226 );
nor \U$5336 ( \6070 , \6068 , \6069 );
and \U$5337 ( \6071 , RI9154318_626, \5453 );
nor \U$5338 ( \6072 , \6070 , \6071 );
nand \U$5339 ( \6073 , \6067 , \6072 );
not \U$5340 ( \6074 , RI9151d98_546);
nor \U$5341 ( \6075 , \6074 , \922 );
not \U$5342 ( \6076 , RI9152518_562);
nor \U$5343 ( \6077 , \6076 , \929 );
nor \U$5344 ( \6078 , \6075 , \6077 );
and \U$5345 ( \6079 , \963 , RI9151618_530);
not \U$5346 ( \6080 , RI9150e98_514);
nor \U$5347 ( \6081 , \6080 , \5464 );
nor \U$5348 ( \6082 , \6079 , \6081 );
nand \U$5349 ( \6083 , \6078 , \6082 );
nor \U$5350 ( \6084 , \6073 , \6083 );
nand \U$5351 ( \6085 , \6062 , \6084 );
buf \U$5352 ( \6086 , \6085 );
not \U$5353 ( \6087 , \6086 );
buf \U$5354 ( \6088 , \1882 );
buf \U$5355 ( \6089 , \5321 );
nand \U$5356 ( \6090 , \6088 , \6089 );
buf \U$5357 ( \6091 , \6090 );
buf \U$5358 ( \6092 , \6091 );
nand \U$5359 ( \6093 , \6087 , \6092 );
buf \U$5360 ( \6094 , \6093 );
buf \U$5361 ( \6095 , \6094 );
not \U$5362 ( \6096 , \6095 );
not \U$5363 ( \6097 , \4794 );
buf \U$5364 ( \6098 , \6097 );
not \U$5365 ( \6099 , \6098 );
buf \U$5366 ( \6100 , \1328 );
not \U$5367 ( \6101 , \6100 );
or \U$5368 ( \6102 , \6099 , \6101 );
buf \U$5369 ( \6103 , \4794 );
buf \U$5370 ( \6104 , \1331 );
nand \U$5371 ( \6105 , \6103 , \6104 );
buf \U$5372 ( \6106 , \6105 );
buf \U$5373 ( \6107 , \6106 );
nand \U$5374 ( \6108 , \6102 , \6107 );
buf \U$5375 ( \6109 , \6108 );
buf \U$5376 ( \6110 , \6109 );
not \U$5377 ( \6111 , \6110 );
buf \U$5378 ( \6112 , \5506 );
not \U$5379 ( \6113 , \6112 );
or \U$5380 ( \6114 , \6111 , \6113 );
buf \U$5381 ( \6115 , \5520 );
buf \U$5382 ( \6116 , \5398 );
nand \U$5383 ( \6117 , \6115 , \6116 );
buf \U$5384 ( \6118 , \6117 );
buf \U$5385 ( \6119 , \6118 );
nand \U$5386 ( \6120 , \6114 , \6119 );
buf \U$5387 ( \6121 , \6120 );
buf \U$5388 ( \6122 , \6121 );
not \U$5389 ( \6123 , \6122 );
or \U$5390 ( \6124 , \6096 , \6123 );
buf \U$5391 ( \6125 , \6091 );
not \U$5392 ( \6126 , \6125 );
buf \U$5393 ( \6127 , \6085 );
nand \U$5394 ( \6128 , \6126 , \6127 );
buf \U$5395 ( \6129 , \6128 );
buf \U$5396 ( \6130 , \6129 );
nand \U$5397 ( \6131 , \6124 , \6130 );
buf \U$5398 ( \6132 , \6131 );
buf \U$5399 ( \6133 , \6132 );
not \U$5400 ( \6134 , \6133 );
buf \U$5401 ( \6135 , \6134 );
buf \U$5402 ( \6136 , \6135 );
not \U$5403 ( \6137 , \6136 );
and \U$5404 ( \6138 , \1669 , \2479 );
not \U$5405 ( \6139 , \1669 );
and \U$5406 ( \6140 , \6139 , \4070 );
or \U$5407 ( \6141 , \6138 , \6140 );
buf \U$5408 ( \6142 , \6141 );
not \U$5409 ( \6143 , \6142 );
buf \U$5410 ( \6144 , \3288 );
not \U$5411 ( \6145 , \6144 );
or \U$5412 ( \6146 , \6143 , \6145 );
buf \U$5413 ( \6147 , \5544 );
buf \U$5414 ( \6148 , \2473 );
nand \U$5415 ( \6149 , \6147 , \6148 );
buf \U$5416 ( \6150 , \6149 );
buf \U$5417 ( \6151 , \6150 );
nand \U$5418 ( \6152 , \6146 , \6151 );
buf \U$5419 ( \6153 , \6152 );
buf \U$5420 ( \6154 , \6153 );
buf \U$5421 ( \6155 , \5017 );
not \U$5422 ( \6156 , \6155 );
buf \U$5423 ( \6157 , \4516 );
not \U$5424 ( \6158 , \6157 );
or \U$5425 ( \6159 , \6156 , \6158 );
buf \U$5426 ( \6160 , \3134 );
buf \U$5427 ( \6161 , \1865 );
nand \U$5428 ( \6162 , \6160 , \6161 );
buf \U$5429 ( \6163 , \6162 );
buf \U$5430 ( \6164 , \6163 );
nand \U$5431 ( \6165 , \6159 , \6164 );
buf \U$5432 ( \6166 , \6165 );
buf \U$5433 ( \6167 , \6166 );
not \U$5434 ( \6168 , \6167 );
buf \U$5435 ( \6169 , \5615 );
not \U$5436 ( \6170 , \6169 );
or \U$5437 ( \6171 , \6168 , \6170 );
buf \U$5438 ( \6172 , \3095 );
buf \U$5439 ( \6173 , \5610 );
nand \U$5440 ( \6174 , \6172 , \6173 );
buf \U$5441 ( \6175 , \6174 );
buf \U$5442 ( \6176 , \6175 );
nand \U$5443 ( \6177 , \6171 , \6176 );
buf \U$5444 ( \6178 , \6177 );
buf \U$5445 ( \6179 , \6178 );
or \U$5446 ( \6180 , \6154 , \6179 );
buf \U$5447 ( \6181 , \6180 );
buf \U$5448 ( \6182 , \6181 );
buf \U$5449 ( \6183 , \1178 );
not \U$5450 ( \6184 , \6183 );
buf \U$5451 ( \6185 , \4848 );
not \U$5452 ( \6186 , \6185 );
or \U$5453 ( \6187 , \6184 , \6186 );
buf \U$5454 ( \6188 , \4991 );
buf \U$5455 ( \6189 , \3329 );
nand \U$5456 ( \6190 , \6188 , \6189 );
buf \U$5457 ( \6191 , \6190 );
buf \U$5458 ( \6192 , \6191 );
nand \U$5459 ( \6193 , \6187 , \6192 );
buf \U$5460 ( \6194 , \6193 );
buf \U$5461 ( \6195 , \6194 );
not \U$5462 ( \6196 , \6195 );
buf \U$5463 ( \6197 , \1187 );
not \U$5464 ( \6198 , \6197 );
or \U$5465 ( \6199 , \6196 , \6198 );
buf \U$5466 ( \6200 , \5658 );
buf \U$5467 ( \6201 , \1194 );
nand \U$5468 ( \6202 , \6200 , \6201 );
buf \U$5469 ( \6203 , \6202 );
buf \U$5470 ( \6204 , \6203 );
nand \U$5471 ( \6205 , \6199 , \6204 );
buf \U$5472 ( \6206 , \6205 );
buf \U$5473 ( \6207 , \6206 );
and \U$5474 ( \6208 , \6182 , \6207 );
buf \U$5475 ( \6209 , \6178 );
buf \U$5476 ( \6210 , \6153 );
and \U$5477 ( \6211 , \6209 , \6210 );
buf \U$5478 ( \6212 , \6211 );
buf \U$5479 ( \6213 , \6212 );
nor \U$5480 ( \6214 , \6208 , \6213 );
buf \U$5481 ( \6215 , \6214 );
buf \U$5482 ( \6216 , \6215 );
not \U$5483 ( \6217 , \6216 );
or \U$5484 ( \6218 , \6137 , \6217 );
buf \U$5485 ( \6219 , \5319 );
not \U$5486 ( \6220 , \6219 );
buf \U$5487 ( \6221 , \1165 );
nand \U$5488 ( \6222 , \6220 , \6221 );
buf \U$5489 ( \6223 , \6222 );
buf \U$5490 ( \6224 , \6223 );
buf \U$5491 ( \6225 , \1107 );
and \U$5492 ( \6226 , \6224 , \6225 );
buf \U$5493 ( \6227 , \5319 );
not \U$5494 ( \6228 , \6227 );
buf \U$5495 ( \6229 , \1162 );
not \U$5496 ( \6230 , \6229 );
or \U$5497 ( \6231 , \6228 , \6230 );
buf \U$5498 ( \6232 , \909 );
nand \U$5499 ( \6233 , \6231 , \6232 );
buf \U$5500 ( \6234 , \6233 );
buf \U$5501 ( \6235 , \6234 );
nor \U$5502 ( \6236 , \6226 , \6235 );
buf \U$5503 ( \6237 , \6236 );
buf \U$5504 ( \6238 , \6237 );
buf \U$5505 ( \6239 , \1014 );
and \U$5506 ( \6240 , \6239 , RI9157810_739);
and \U$5507 ( \6241 , \4011 , RI9157f90_755);
nor \U$5508 ( \6242 , \6240 , \6241 );
not \U$5509 ( \6243 , \6242 );
not \U$5510 ( \6244 , RI9156910_707);
nor \U$5511 ( \6245 , \6244 , \1524 );
not \U$5512 ( \6246 , RI9157090_723);
nor \U$5513 ( \6247 , \6246 , \1847 );
not \U$5514 ( \6248 , RI9155a10_675);
nor \U$5515 ( \6249 , \6248 , \989 );
not \U$5516 ( \6250 , RI9156190_691);
nor \U$5517 ( \6251 , \6250 , \994 );
nor \U$5518 ( \6252 , \6249 , \6251 );
not \U$5519 ( \6253 , RI9154b10_643);
nor \U$5520 ( \6254 , \6253 , \976 );
not \U$5521 ( \6255 , RI9155290_659);
nor \U$5522 ( \6256 , \6255 , \983 );
nor \U$5523 ( \6257 , \6254 , \6256 );
nand \U$5524 ( \6258 , \6252 , \6257 );
nor \U$5525 ( \6259 , \6243 , \6245 , \6247 , \6258 );
not \U$5526 ( \6260 , RI9152d10_579);
nor \U$5527 ( \6261 , \6260 , \952 );
not \U$5528 ( \6262 , RI9153490_595);
nor \U$5529 ( \6263 , \6262 , \1285 );
nor \U$5530 ( \6264 , \6261 , \6263 );
and \U$5531 ( \6265 , \5453 , RI9154390_627);
not \U$5532 ( \6266 , RI9153c10_611);
nor \U$5533 ( \6267 , \6266 , \6069 );
nor \U$5534 ( \6268 , \6265 , \6267 );
nand \U$5535 ( \6269 , \6264 , \6268 );
not \U$5536 ( \6270 , RI9152590_563);
nor \U$5537 ( \6271 , \6270 , \929 );
not \U$5538 ( \6272 , \6271 );
not \U$5539 ( \6273 , \1302 );
not \U$5540 ( \6274 , \6273 );
nand \U$5541 ( \6275 , \6274 , RI9151e10_547);
and \U$5542 ( \6276 , \963 , RI9151690_531);
and \U$5543 ( \6277 , \968 , RI9150f10_515);
nor \U$5544 ( \6278 , \6276 , \6277 );
nand \U$5545 ( \6279 , \6272 , \6275 , \6278 );
nor \U$5546 ( \6280 , \6269 , \6279 );
nand \U$5547 ( \6281 , \6259 , \6280 );
buf \U$5548 ( \6282 , \6281 );
and \U$5549 ( \6283 , \6238 , \6282 );
buf \U$5550 ( \6284 , \6283 );
buf \U$5551 ( \6285 , \6284 );
not \U$5552 ( \6286 , \6285 );
buf \U$5553 ( \6287 , \3223 );
not \U$5554 ( \6288 , \6287 );
buf \U$5555 ( \6289 , \2071 );
not \U$5556 ( \6290 , \6289 );
or \U$5557 ( \6291 , \6288 , \6290 );
buf \U$5558 ( \6292 , \2068 );
buf \U$5559 ( \6293 , \3459 );
nand \U$5560 ( \6294 , \6292 , \6293 );
buf \U$5561 ( \6295 , \6294 );
buf \U$5562 ( \6296 , \6295 );
nand \U$5563 ( \6297 , \6291 , \6296 );
buf \U$5564 ( \6298 , \6297 );
buf \U$5565 ( \6299 , \6298 );
not \U$5566 ( \6300 , \6299 );
buf \U$5567 ( \6301 , \2503 );
not \U$5568 ( \6302 , \6301 );
or \U$5569 ( \6303 , \6300 , \6302 );
buf \U$5570 ( \6304 , \2897 );
buf \U$5571 ( \6305 , \5690 );
nand \U$5572 ( \6306 , \6304 , \6305 );
buf \U$5573 ( \6307 , \6306 );
buf \U$5574 ( \6308 , \6307 );
nand \U$5575 ( \6309 , \6303 , \6308 );
buf \U$5576 ( \6310 , \6309 );
buf \U$5577 ( \6311 , \6310 );
not \U$5578 ( \6312 , \6311 );
or \U$5579 ( \6313 , \6286 , \6312 );
buf \U$5580 ( \6314 , \6310 );
buf \U$5581 ( \6315 , \6284 );
or \U$5582 ( \6316 , \6314 , \6315 );
buf \U$5583 ( \6317 , \1027 );
not \U$5584 ( \6318 , \6317 );
buf \U$5585 ( \6319 , \4281 );
not \U$5586 ( \6320 , \6319 );
or \U$5587 ( \6321 , \6318 , \6320 );
buf \U$5588 ( \6322 , \4278 );
buf \U$5589 ( \6323 , \1024 );
nand \U$5590 ( \6324 , \6322 , \6323 );
buf \U$5591 ( \6325 , \6324 );
buf \U$5592 ( \6326 , \6325 );
nand \U$5593 ( \6327 , \6321 , \6326 );
buf \U$5594 ( \6328 , \6327 );
buf \U$5595 ( \6329 , \6328 );
not \U$5596 ( \6330 , \6329 );
buf \U$5597 ( \6331 , \4543 );
not \U$5598 ( \6332 , \6331 );
or \U$5599 ( \6333 , \6330 , \6332 );
buf \U$5600 ( \6334 , \4581 );
buf \U$5601 ( \6335 , \5754 );
nand \U$5602 ( \6336 , \6334 , \6335 );
buf \U$5603 ( \6337 , \6336 );
buf \U$5604 ( \6338 , \6337 );
nand \U$5605 ( \6339 , \6333 , \6338 );
buf \U$5606 ( \6340 , \6339 );
buf \U$5607 ( \6341 , \6340 );
nand \U$5608 ( \6342 , \6316 , \6341 );
buf \U$5609 ( \6343 , \6342 );
buf \U$5610 ( \6344 , \6343 );
nand \U$5611 ( \6345 , \6313 , \6344 );
buf \U$5612 ( \6346 , \6345 );
buf \U$5613 ( \6347 , \6346 );
nand \U$5614 ( \6348 , \6218 , \6347 );
buf \U$5615 ( \6349 , \6348 );
buf \U$5616 ( \6350 , \6349 );
buf \U$5617 ( \6351 , \6215 );
not \U$5618 ( \6352 , \6351 );
buf \U$5619 ( \6353 , \6352 );
buf \U$5620 ( \6354 , \6353 );
buf \U$5621 ( \6355 , \6132 );
nand \U$5622 ( \6356 , \6354 , \6355 );
buf \U$5623 ( \6357 , \6356 );
buf \U$5624 ( \6358 , \6357 );
nand \U$5625 ( \6359 , \6350 , \6358 );
buf \U$5626 ( \6360 , \6359 );
buf \U$5627 ( \6361 , \6360 );
not \U$5628 ( \6362 , \6361 );
xor \U$5629 ( \6363 , \5568 , \5677 );
xor \U$5630 ( \6364 , \6363 , \5769 );
buf \U$5631 ( \6365 , \6364 );
buf \U$5632 ( \6366 , \6365 );
not \U$5633 ( \6367 , \6366 );
or \U$5634 ( \6368 , \6362 , \6367 );
buf \U$5635 ( \6369 , \6360 );
buf \U$5636 ( \6370 , \6365 );
or \U$5637 ( \6371 , \6369 , \6370 );
buf \U$5638 ( \6372 , \5530 );
buf \U$5639 ( \6373 , \5502 );
xor \U$5640 ( \6374 , \6372 , \6373 );
buf \U$5641 ( \6375 , \6374 );
buf \U$5644 ( \6376 , \5556 );
xnor \U$5645 ( \6377 , \6375 , \6376 );
buf \U$5646 ( \6378 , \6377 );
not \U$5647 ( \6379 , \6378 );
buf \U$5648 ( \6380 , \6379 );
buf \U$5649 ( \6381 , \6380 );
not \U$5650 ( \6382 , \6381 );
and \U$5651 ( \6383 , \5766 , \5740 );
not \U$5652 ( \6384 , \5766 );
and \U$5653 ( \6385 , \6384 , \5706 );
or \U$5654 ( \6386 , \6383 , \6385 );
buf \U$5655 ( \6387 , \6386 );
buf \U$5658 ( \6388 , \5731 );
buf \U$5659 ( \6389 , \6388 );
and \U$5660 ( \6390 , \6387 , \6389 );
not \U$5661 ( \6391 , \6387 );
buf \U$5662 ( \6392 , \6388 );
not \U$5663 ( \6393 , \6392 );
buf \U$5664 ( \6394 , \6393 );
buf \U$5665 ( \6395 , \6394 );
and \U$5666 ( \6396 , \6391 , \6395 );
nor \U$5667 ( \6397 , \6390 , \6396 );
buf \U$5668 ( \6398 , \6397 );
buf \U$5669 ( \6399 , \6398 );
not \U$5670 ( \6400 , \6399 );
or \U$5671 ( \6401 , \6382 , \6400 );
buf \U$5672 ( \6402 , \6380 );
buf \U$5673 ( \6403 , \6398 );
or \U$5674 ( \6404 , \6402 , \6403 );
buf \U$5675 ( \6405 , \5640 );
buf \U$5676 ( \6406 , \5595 );
xor \U$5677 ( \6407 , \6405 , \6406 );
buf \U$5678 ( \6408 , \6407 );
buf \U$5679 ( \6409 , \6408 );
buf \U$5680 ( \6410 , \5670 );
xor \U$5681 ( \6411 , \6409 , \6410 );
buf \U$5682 ( \6412 , \6411 );
buf \U$5683 ( \6413 , \6412 );
nand \U$5684 ( \6414 , \6404 , \6413 );
buf \U$5685 ( \6415 , \6414 );
buf \U$5686 ( \6416 , \6415 );
nand \U$5687 ( \6417 , \6401 , \6416 );
buf \U$5688 ( \6418 , \6417 );
buf \U$5689 ( \6419 , \6418 );
nand \U$5690 ( \6420 , \6371 , \6419 );
buf \U$5691 ( \6421 , \6420 );
buf \U$5692 ( \6422 , \6421 );
nand \U$5693 ( \6423 , \6368 , \6422 );
buf \U$5694 ( \6424 , \6423 );
buf \U$5695 ( \6425 , \6424 );
nand \U$5696 ( \6426 , \6046 , \6425 );
buf \U$5697 ( \6427 , \6426 );
buf \U$5698 ( \6428 , \6427 );
buf \U$5699 ( \6429 , \6038 );
buf \U$5700 ( \6430 , \6044 );
nand \U$5701 ( \6431 , \6429 , \6430 );
buf \U$5702 ( \6432 , \6431 );
buf \U$5703 ( \6433 , \6432 );
and \U$5704 ( \6434 , \6428 , \6433 );
buf \U$5705 ( \6435 , \6434 );
buf \U$5706 ( \6436 , \6435 );
nor \U$5707 ( \6437 , \6032 , \6436 );
buf \U$5708 ( \6438 , \6437 );
buf \U$5709 ( \6439 , \6438 );
and \U$5710 ( \6440 , \6028 , \6439 );
buf \U$5711 ( \6441 , \6440 );
buf \U$5712 ( \6442 , \6441 );
nor \U$5713 ( \6443 , \6023 , \6442 );
buf \U$5714 ( \6444 , \6443 );
buf \U$5715 ( \6445 , \6444 );
buf \U$5716 ( \6446 , \5959 );
not \U$5717 ( \6447 , \6446 );
buf \U$5718 ( \6448 , \6447 );
buf \U$5719 ( \6449 , \6448 );
not \U$5720 ( \6450 , \6449 );
xor \U$5721 ( \6451 , \5964 , \5973 );
buf \U$5722 ( \6452 , \6451 );
not \U$5723 ( \6453 , \6452 );
or \U$5724 ( \6454 , \6450 , \6453 );
buf \U$5725 ( \6455 , \6451 );
buf \U$5726 ( \6456 , \6448 );
or \U$5727 ( \6457 , \6455 , \6456 );
nand \U$5728 ( \6458 , \6454 , \6457 );
buf \U$5729 ( \6459 , \6458 );
buf \U$5730 ( \6460 , \6459 );
buf \U$5731 ( \6461 , \6091 );
not \U$5732 ( \6462 , \6461 );
buf \U$5733 ( \6463 , \6085 );
not \U$5734 ( \6464 , \6463 );
and \U$5735 ( \6465 , \6462 , \6464 );
buf \U$5736 ( \6466 , \6091 );
buf \U$5737 ( \6467 , \6085 );
and \U$5738 ( \6468 , \6466 , \6467 );
nor \U$5739 ( \6469 , \6465 , \6468 );
buf \U$5740 ( \6470 , \6469 );
xor \U$5741 ( \6471 , \6121 , \6470 );
buf \U$5742 ( \6472 , \6471 );
buf \U$5743 ( \6473 , \4768 );
not \U$5744 ( \6474 , \6473 );
buf \U$5745 ( \6475 , \2273 );
not \U$5746 ( \6476 , \6475 );
or \U$5747 ( \6477 , \6474 , \6476 );
buf \U$5748 ( \6478 , \2276 );
buf \U$5749 ( \6479 , \4029 );
nand \U$5750 ( \6480 , \6478 , \6479 );
buf \U$5751 ( \6481 , \6480 );
buf \U$5752 ( \6482 , \6481 );
nand \U$5753 ( \6483 , \6477 , \6482 );
buf \U$5754 ( \6484 , \6483 );
buf \U$5755 ( \6485 , \6484 );
not \U$5756 ( \6486 , \6485 );
buf \U$5757 ( \6487 , \1478 );
not \U$5758 ( \6488 , \6487 );
or \U$5759 ( \6489 , \6486 , \6488 );
buf \U$5760 ( \6490 , \1904 );
buf \U$5761 ( \6491 , \5719 );
nand \U$5762 ( \6492 , \6490 , \6491 );
buf \U$5763 ( \6493 , \6492 );
buf \U$5764 ( \6494 , \6493 );
nand \U$5765 ( \6495 , \6489 , \6494 );
buf \U$5766 ( \6496 , \6495 );
buf \U$5767 ( \6497 , \6496 );
not \U$5768 ( \6498 , \6497 );
buf \U$5769 ( \6499 , \6498 );
buf \U$5770 ( \6500 , \6499 );
nand \U$5771 ( \6501 , \6472 , \6500 );
buf \U$5772 ( \6502 , \6501 );
buf \U$5773 ( \6503 , \6502 );
not \U$5774 ( \6504 , \6503 );
buf \U$5775 ( \6505 , \4516 );
not \U$5776 ( \6506 , \6505 );
buf \U$5777 ( \6507 , \1795 );
not \U$5778 ( \6508 , \6507 );
or \U$5779 ( \6509 , \6506 , \6508 );
buf \U$5780 ( \6510 , \5603 );
buf \U$5781 ( \6511 , \1931 );
nand \U$5782 ( \6512 , \6510 , \6511 );
buf \U$5783 ( \6513 , \6512 );
buf \U$5784 ( \6514 , \6513 );
nand \U$5785 ( \6515 , \6509 , \6514 );
buf \U$5786 ( \6516 , \6515 );
buf \U$5787 ( \6517 , \6516 );
not \U$5788 ( \6518 , \6517 );
buf \U$5789 ( \6519 , \5143 );
not \U$5790 ( \6520 , \6519 );
or \U$5791 ( \6521 , \6518 , \6520 );
buf \U$5792 ( \6522 , \6166 );
buf \U$5793 ( \6523 , \3095 );
nand \U$5794 ( \6524 , \6522 , \6523 );
buf \U$5795 ( \6525 , \6524 );
buf \U$5796 ( \6526 , \6525 );
nand \U$5797 ( \6527 , \6521 , \6526 );
buf \U$5798 ( \6528 , \6527 );
buf \U$5799 ( \6529 , \6528 );
not \U$5800 ( \6530 , \6529 );
buf \U$5801 ( \6531 , \6530 );
buf \U$5802 ( \6532 , \6531 );
not \U$5803 ( \6533 , \6532 );
buf \U$5804 ( \6534 , \3288 );
not \U$5805 ( \6535 , \6534 );
buf \U$5806 ( \6536 , \2758 );
not \U$5807 ( \6537 , \6536 );
buf \U$5808 ( \6538 , \2627 );
not \U$5809 ( \6539 , \6538 );
or \U$5810 ( \6540 , \6537 , \6539 );
buf \U$5811 ( \6541 , \3276 );
buf \U$5812 ( \6542 , \2853 );
nand \U$5813 ( \6543 , \6541 , \6542 );
buf \U$5814 ( \6544 , \6543 );
buf \U$5815 ( \6545 , \6544 );
nand \U$5816 ( \6546 , \6540 , \6545 );
buf \U$5817 ( \6547 , \6546 );
buf \U$5818 ( \6548 , \6547 );
not \U$5819 ( \6549 , \6548 );
or \U$5820 ( \6550 , \6535 , \6549 );
buf \U$5821 ( \6551 , \6141 );
buf \U$5822 ( \6552 , \2473 );
nand \U$5823 ( \6553 , \6551 , \6552 );
buf \U$5824 ( \6554 , \6553 );
buf \U$5825 ( \6555 , \6554 );
nand \U$5826 ( \6556 , \6550 , \6555 );
buf \U$5827 ( \6557 , \6556 );
buf \U$5828 ( \6558 , \6557 );
not \U$5829 ( \6559 , \6558 );
buf \U$5830 ( \6560 , \6559 );
buf \U$5831 ( \6561 , \6560 );
not \U$5832 ( \6562 , \6561 );
or \U$5833 ( \6563 , \6533 , \6562 );
buf \U$5834 ( \6564 , \2521 );
not \U$5835 ( \6565 , \6564 );
buf \U$5836 ( \6566 , \4550 );
not \U$5837 ( \6567 , \6566 );
or \U$5838 ( \6568 , \6565 , \6567 );
buf \U$5839 ( \6569 , \4278 );
buf \U$5840 ( \6570 , \1999 );
nand \U$5841 ( \6571 , \6569 , \6570 );
buf \U$5842 ( \6572 , \6571 );
buf \U$5843 ( \6573 , \6572 );
nand \U$5844 ( \6574 , \6568 , \6573 );
buf \U$5845 ( \6575 , \6574 );
buf \U$5846 ( \6576 , \6575 );
not \U$5847 ( \6577 , \6576 );
buf \U$5850 ( \6578 , \4543 );
buf \U$5851 ( \6579 , \6578 );
not \U$5852 ( \6580 , \6579 );
or \U$5853 ( \6581 , \6577 , \6580 );
buf \U$5856 ( \6582 , \4581 );
buf \U$5857 ( \6583 , \6582 );
buf \U$5858 ( \6584 , \6328 );
nand \U$5859 ( \6585 , \6583 , \6584 );
buf \U$5860 ( \6586 , \6585 );
buf \U$5861 ( \6587 , \6586 );
nand \U$5862 ( \6588 , \6581 , \6587 );
buf \U$5863 ( \6589 , \6588 );
buf \U$5864 ( \6590 , \6589 );
nand \U$5865 ( \6591 , \6563 , \6590 );
buf \U$5866 ( \6592 , \6591 );
buf \U$5867 ( \6593 , \6592 );
buf \U$5868 ( \6594 , \6557 );
buf \U$5869 ( \6595 , \6528 );
nand \U$5870 ( \6596 , \6594 , \6595 );
buf \U$5871 ( \6597 , \6596 );
buf \U$5872 ( \6598 , \6597 );
nand \U$5873 ( \6599 , \6593 , \6598 );
buf \U$5874 ( \6600 , \6599 );
buf \U$5875 ( \6601 , \6600 );
not \U$5876 ( \6602 , \6601 );
or \U$5877 ( \6603 , \6504 , \6602 );
buf \U$5878 ( \6604 , \6471 );
not \U$5879 ( \6605 , \6604 );
buf \U$5880 ( \6606 , \6496 );
nand \U$5881 ( \6607 , \6605 , \6606 );
buf \U$5882 ( \6608 , \6607 );
buf \U$5883 ( \6609 , \6608 );
nand \U$5884 ( \6610 , \6603 , \6609 );
buf \U$5885 ( \6611 , \6610 );
buf \U$5886 ( \6612 , \6611 );
not \U$5887 ( \6613 , \6612 );
buf \U$5888 ( \6614 , \6132 );
buf \U$5889 ( \6615 , \6346 );
xor \U$5890 ( \6616 , \6614 , \6615 );
buf \U$5891 ( \6617 , \6353 );
xnor \U$5892 ( \6618 , \6616 , \6617 );
buf \U$5893 ( \6619 , \6618 );
buf \U$5894 ( \6620 , \6619 );
not \U$5895 ( \6621 , \6620 );
buf \U$5896 ( \6622 , \6621 );
buf \U$5897 ( \6623 , \6622 );
not \U$5898 ( \6624 , \6623 );
or \U$5899 ( \6625 , \6613 , \6624 );
buf \U$5900 ( \6626 , \6611 );
not \U$5901 ( \6627 , \6626 );
buf \U$5902 ( \6628 , \6627 );
buf \U$5903 ( \6629 , \6628 );
not \U$5904 ( \6630 , \6629 );
buf \U$5905 ( \6631 , \6619 );
not \U$5906 ( \6632 , \6631 );
or \U$5907 ( \6633 , \6630 , \6632 );
buf \U$5908 ( \6634 , \6284 );
buf \U$5909 ( \6635 , \6340 );
xor \U$5910 ( \6636 , \6634 , \6635 );
buf \U$5911 ( \6637 , \6310 );
xnor \U$5912 ( \6638 , \6636 , \6637 );
buf \U$5913 ( \6639 , \6638 );
buf \U$5914 ( \6640 , \6639 );
not \U$5915 ( \6641 , \6640 );
buf \U$5916 ( \6642 , \6641 );
not \U$5917 ( \6643 , \6642 );
buf \U$5918 ( \6644 , \5506 );
not \U$5919 ( \6645 , \6644 );
and \U$5920 ( \6646 , \1255 , \5330 );
not \U$5921 ( \6647 , \1255 );
and \U$5922 ( \6648 , \6647 , \4794 );
or \U$5923 ( \6649 , \6646 , \6648 );
buf \U$5924 ( \6650 , \6649 );
not \U$5925 ( \6651 , \6650 );
or \U$5926 ( \6652 , \6645 , \6651 );
buf \U$5927 ( \6653 , \6109 );
buf \U$5928 ( \6654 , \5398 );
nand \U$5929 ( \6655 , \6653 , \6654 );
buf \U$5930 ( \6656 , \6655 );
buf \U$5931 ( \6657 , \6656 );
nand \U$5932 ( \6658 , \6652 , \6657 );
buf \U$5933 ( \6659 , \6658 );
buf \U$5936 ( \6660 , \6659 );
buf \U$5937 ( \6661 , \6660 );
not \U$5938 ( \6662 , \6661 );
buf \U$5939 ( \6663 , \6223 );
buf \U$5940 ( \6664 , \1107 );
and \U$5941 ( \6665 , \6663 , \6664 );
buf \U$5942 ( \6666 , \6234 );
nor \U$5943 ( \6667 , \6665 , \6666 );
buf \U$5944 ( \6668 , \6667 );
buf \U$5945 ( \6669 , \6668 );
not \U$5946 ( \6670 , \6669 );
buf \U$5947 ( \6671 , \6281 );
not \U$5948 ( \6672 , \6671 );
buf \U$5949 ( \6673 , \6672 );
buf \U$5950 ( \6674 , \6673 );
not \U$5951 ( \6675 , \6674 );
and \U$5952 ( \6676 , \6670 , \6675 );
buf \U$5953 ( \6677 , \6673 );
buf \U$5954 ( \6678 , \6237 );
and \U$5955 ( \6679 , \6677 , \6678 );
nor \U$5956 ( \6680 , \6676 , \6679 );
buf \U$5957 ( \6681 , \6680 );
buf \U$5958 ( \6682 , \6681 );
not \U$5959 ( \6683 , \6682 );
buf \U$5960 ( \6684 , \6683 );
buf \U$5961 ( \6685 , \6684 );
not \U$5962 ( \6686 , \6685 );
or \U$5963 ( \6687 , \6662 , \6686 );
buf \U$5964 ( \6688 , \6660 );
buf \U$5965 ( \6689 , \6684 );
or \U$5966 ( \6690 , \6688 , \6689 );
buf \U$5967 ( \6691 , \3329 );
buf \U$5968 ( \6692 , \5321 );
and \U$5969 ( \6693 , \6691 , \6692 );
not \U$5970 ( \6694 , \6691 );
buf \U$5971 ( \6695 , \5573 );
and \U$5972 ( \6696 , \6694 , \6695 );
nor \U$5973 ( \6697 , \6693 , \6696 );
buf \U$5974 ( \6698 , \6697 );
buf \U$5975 ( \6699 , \6698 );
not \U$5976 ( \6700 , \6699 );
buf \U$5977 ( \6701 , \1186 );
not \U$5978 ( \6702 , \6701 );
or \U$5979 ( \6703 , \6700 , \6702 );
buf \U$5980 ( \6704 , \6194 );
buf \U$5981 ( \6705 , \1193 );
nand \U$5982 ( \6706 , \6704 , \6705 );
buf \U$5983 ( \6707 , \6706 );
buf \U$5984 ( \6708 , \6707 );
nand \U$5985 ( \6709 , \6703 , \6708 );
buf \U$5986 ( \6710 , \6709 );
buf \U$5987 ( \6711 , \6710 );
nand \U$5988 ( \6712 , \6690 , \6711 );
buf \U$5989 ( \6713 , \6712 );
buf \U$5990 ( \6714 , \6713 );
nand \U$5991 ( \6715 , \6687 , \6714 );
buf \U$5992 ( \6716 , \6715 );
not \U$5993 ( \6717 , \6716 );
or \U$5994 ( \6718 , \6643 , \6717 );
buf \U$5995 ( \6719 , \6716 );
not \U$5996 ( \6720 , \6719 );
buf \U$5997 ( \6721 , \6720 );
not \U$5998 ( \6722 , \6721 );
not \U$5999 ( \6723 , \6639 );
or \U$6000 ( \6724 , \6722 , \6723 );
xor \U$6001 ( \6725 , \6209 , \6210 );
buf \U$6002 ( \6726 , \6725 );
xor \U$6003 ( \6727 , \6206 , \6726 );
nand \U$6004 ( \6728 , \6724 , \6727 );
nand \U$6005 ( \6729 , \6718 , \6728 );
buf \U$6006 ( \6730 , \6729 );
nand \U$6007 ( \6731 , \6633 , \6730 );
buf \U$6008 ( \6732 , \6731 );
buf \U$6009 ( \6733 , \6732 );
nand \U$6010 ( \6734 , \6625 , \6733 );
buf \U$6011 ( \6735 , \6734 );
buf \U$6012 ( \6736 , \6735 );
xor \U$6013 ( \6737 , \6460 , \6736 );
buf \U$6014 ( \6738 , \6360 );
buf \U$6015 ( \6739 , \6365 );
and \U$6016 ( \6740 , \6738 , \6739 );
not \U$6017 ( \6741 , \6738 );
buf \U$6018 ( \6742 , \6365 );
not \U$6019 ( \6743 , \6742 );
buf \U$6020 ( \6744 , \6743 );
buf \U$6021 ( \6745 , \6744 );
and \U$6022 ( \6746 , \6741 , \6745 );
nor \U$6023 ( \6747 , \6740 , \6746 );
buf \U$6024 ( \6748 , \6747 );
buf \U$6025 ( \6749 , \6748 );
buf \U$6026 ( \6750 , \6418 );
and \U$6027 ( \6751 , \6749 , \6750 );
not \U$6028 ( \6752 , \6749 );
buf \U$6029 ( \6753 , \6418 );
not \U$6030 ( \6754 , \6753 );
buf \U$6031 ( \6755 , \6754 );
buf \U$6032 ( \6756 , \6755 );
and \U$6033 ( \6757 , \6752 , \6756 );
nor \U$6034 ( \6758 , \6751 , \6757 );
buf \U$6035 ( \6759 , \6758 );
buf \U$6036 ( \6760 , \6759 );
xor \U$6037 ( \6761 , \6737 , \6760 );
buf \U$6038 ( \6762 , \6761 );
buf \U$6039 ( \6763 , \6762 );
buf \U$6040 ( \6764 , \4691 );
not \U$6041 ( \6765 , \6764 );
buf \U$6042 ( \6766 , \6765 );
buf \U$6043 ( \6767 , \6766 );
not \U$6044 ( \6768 , \6767 );
buf \U$6045 ( \6769 , \4675 );
not \U$6046 ( \6770 , \6769 );
or \U$6047 ( \6771 , \6768 , \6770 );
buf \U$6048 ( \6772 , \4855 );
buf \U$6049 ( \6773 , \4691 );
nand \U$6050 ( \6774 , \6772 , \6773 );
buf \U$6051 ( \6775 , \6774 );
buf \U$6052 ( \6776 , \6775 );
nand \U$6053 ( \6777 , \6771 , \6776 );
buf \U$6054 ( \6778 , \6777 );
buf \U$6055 ( \6779 , \6778 );
not \U$6056 ( \6780 , \6779 );
buf \U$6057 ( \6781 , \1472 );
not \U$6058 ( \6782 , \6781 );
or \U$6059 ( \6783 , \6780 , \6782 );
buf \U$6060 ( \6784 , \6484 );
buf \U$6061 ( \6785 , \1485 );
nand \U$6062 ( \6786 , \6784 , \6785 );
buf \U$6063 ( \6787 , \6786 );
buf \U$6064 ( \6788 , \6787 );
nand \U$6065 ( \6789 , \6783 , \6788 );
buf \U$6066 ( \6790 , \6789 );
buf \U$6067 ( \6791 , \6790 );
not \U$6068 ( \6792 , \6791 );
buf \U$6069 ( \6793 , \3444 );
not \U$6070 ( \6794 , \6793 );
buf \U$6071 ( \6795 , \2488 );
not \U$6072 ( \6796 , \6795 );
or \U$6073 ( \6797 , \6794 , \6796 );
buf \U$6074 ( \6798 , \2068 );
buf \U$6075 ( \6799 , \4381 );
nand \U$6076 ( \6800 , \6798 , \6799 );
buf \U$6077 ( \6801 , \6800 );
buf \U$6078 ( \6802 , \6801 );
nand \U$6079 ( \6803 , \6797 , \6802 );
buf \U$6080 ( \6804 , \6803 );
buf \U$6081 ( \6805 , \6804 );
not \U$6082 ( \6806 , \6805 );
buf \U$6083 ( \6807 , \2503 );
not \U$6084 ( \6808 , \6807 );
or \U$6085 ( \6809 , \6806 , \6808 );
buf \U$6086 ( \6810 , \2214 );
buf \U$6087 ( \6811 , \6298 );
nand \U$6088 ( \6812 , \6810 , \6811 );
buf \U$6089 ( \6813 , \6812 );
buf \U$6090 ( \6814 , \6813 );
nand \U$6091 ( \6815 , \6809 , \6814 );
buf \U$6092 ( \6816 , \6815 );
buf \U$6093 ( \6817 , \6816 );
not \U$6094 ( \6818 , \6817 );
buf \U$6095 ( \6819 , \6818 );
buf \U$6096 ( \6820 , \6819 );
nand \U$6097 ( \6821 , \6792 , \6820 );
buf \U$6098 ( \6822 , \6821 );
buf \U$6099 ( \6823 , \6822 );
not \U$6100 ( \6824 , \6823 );
buf \U$6101 ( \6825 , \1547 );
not \U$6102 ( \6826 , \6825 );
buf \U$6103 ( \6827 , \4848 );
not \U$6104 ( \6828 , \6827 );
or \U$6105 ( \6829 , \6826 , \6828 );
buf \U$6106 ( \6830 , \4991 );
buf \U$6107 ( \6831 , \6766 );
nand \U$6108 ( \6832 , \6830 , \6831 );
buf \U$6109 ( \6833 , \6832 );
buf \U$6110 ( \6834 , \6833 );
nand \U$6111 ( \6835 , \6829 , \6834 );
buf \U$6112 ( \6836 , \6835 );
buf \U$6113 ( \6837 , \6836 );
not \U$6114 ( \6838 , \6837 );
buf \U$6115 ( \6839 , \1472 );
not \U$6116 ( \6840 , \6839 );
or \U$6117 ( \6841 , \6838 , \6840 );
buf \U$6118 ( \6842 , \1482 );
not \U$6119 ( \6843 , \6842 );
buf \U$6120 ( \6844 , \6778 );
nand \U$6121 ( \6845 , \6843 , \6844 );
buf \U$6122 ( \6846 , \6845 );
buf \U$6123 ( \6847 , \6846 );
nand \U$6124 ( \6848 , \6841 , \6847 );
buf \U$6125 ( \6849 , \6848 );
buf \U$6128 ( \6850 , \6849 );
buf \U$6129 ( \6851 , \6850 );
not \U$6130 ( \6852 , \6851 );
buf \U$6131 ( \6853 , \4032 );
not \U$6132 ( \6854 , \6853 );
buf \U$6133 ( \6855 , \2878 );
not \U$6134 ( \6856 , \6855 );
or \U$6135 ( \6857 , \6854 , \6856 );
buf \U$6136 ( \6858 , \2068 );
buf \U$6137 ( \6859 , \4029 );
nand \U$6138 ( \6860 , \6858 , \6859 );
buf \U$6139 ( \6861 , \6860 );
buf \U$6140 ( \6862 , \6861 );
nand \U$6141 ( \6863 , \6857 , \6862 );
buf \U$6142 ( \6864 , \6863 );
buf \U$6143 ( \6865 , \6864 );
not \U$6144 ( \6866 , \6865 );
buf \U$6145 ( \6867 , \2200 );
not \U$6146 ( \6868 , \6867 );
or \U$6147 ( \6869 , \6866 , \6868 );
buf \U$6148 ( \6870 , \2214 );
buf \U$6149 ( \6871 , \6804 );
nand \U$6150 ( \6872 , \6870 , \6871 );
buf \U$6151 ( \6873 , \6872 );
buf \U$6152 ( \6874 , \6873 );
nand \U$6153 ( \6875 , \6869 , \6874 );
buf \U$6154 ( \6876 , \6875 );
buf \U$6155 ( \6877 , \6876 );
not \U$6156 ( \6878 , \6877 );
or \U$6157 ( \6879 , \6852 , \6878 );
buf \U$6158 ( \6880 , \6850 );
buf \U$6159 ( \6881 , \6876 );
or \U$6160 ( \6882 , \6880 , \6881 );
buf \U$6161 ( \6883 , \1868 );
not \U$6162 ( \6884 , \6883 );
buf \U$6163 ( \6885 , \4282 );
not \U$6164 ( \6886 , \6885 );
or \U$6165 ( \6887 , \6884 , \6886 );
buf \U$6166 ( \6888 , \4278 );
buf \U$6167 ( \6889 , \2670 );
nand \U$6168 ( \6890 , \6888 , \6889 );
buf \U$6169 ( \6891 , \6890 );
buf \U$6170 ( \6892 , \6891 );
nand \U$6171 ( \6893 , \6887 , \6892 );
buf \U$6172 ( \6894 , \6893 );
buf \U$6173 ( \6895 , \6894 );
not \U$6174 ( \6896 , \6895 );
buf \U$6175 ( \6897 , \6578 );
not \U$6176 ( \6898 , \6897 );
or \U$6177 ( \6899 , \6896 , \6898 );
buf \U$6178 ( \6900 , \4581 );
buf \U$6179 ( \6901 , \6575 );
nand \U$6180 ( \6902 , \6900 , \6901 );
buf \U$6181 ( \6903 , \6902 );
buf \U$6182 ( \6904 , \6903 );
nand \U$6183 ( \6905 , \6899 , \6904 );
buf \U$6184 ( \6906 , \6905 );
buf \U$6185 ( \6907 , \6906 );
nand \U$6186 ( \6908 , \6882 , \6907 );
buf \U$6187 ( \6909 , \6908 );
buf \U$6188 ( \6910 , \6909 );
nand \U$6189 ( \6911 , \6879 , \6910 );
buf \U$6190 ( \6912 , \6911 );
buf \U$6191 ( \6913 , \6912 );
not \U$6192 ( \6914 , \6913 );
or \U$6193 ( \6915 , \6824 , \6914 );
buf \U$6194 ( \6916 , \6816 );
buf \U$6195 ( \6917 , \6790 );
nand \U$6196 ( \6918 , \6916 , \6917 );
buf \U$6197 ( \6919 , \6918 );
buf \U$6198 ( \6920 , \6919 );
nand \U$6199 ( \6921 , \6915 , \6920 );
buf \U$6200 ( \6922 , \6921 );
buf \U$6201 ( \6923 , \6922 );
not \U$6202 ( \6924 , \6923 );
buf \U$6203 ( \6925 , \6924 );
buf \U$6204 ( \6926 , \6925 );
not \U$6205 ( \6927 , \6926 );
xor \U$6206 ( \6928 , \6121 , \6470 );
xnor \U$6207 ( \6929 , \6928 , \6499 );
buf \U$6208 ( \6930 , \6929 );
not \U$6209 ( \6931 , \6930 );
buf \U$6210 ( \6932 , \6600 );
not \U$6211 ( \6933 , \6932 );
and \U$6212 ( \6934 , \6931 , \6933 );
buf \U$6213 ( \6935 , \6600 );
buf \U$6214 ( \6936 , \6929 );
and \U$6215 ( \6937 , \6935 , \6936 );
nor \U$6216 ( \6938 , \6934 , \6937 );
buf \U$6217 ( \6939 , \6938 );
buf \U$6218 ( \6940 , \6939 );
not \U$6219 ( \6941 , \6940 );
or \U$6220 ( \6942 , \6927 , \6941 );
and \U$6221 ( \6943 , \1669 , \4516 );
not \U$6222 ( \6944 , \1669 );
and \U$6223 ( \6945 , \6944 , \5603 );
or \U$6224 ( \6946 , \6943 , \6945 );
buf \U$6225 ( \6947 , \6946 );
not \U$6226 ( \6948 , \6947 );
buf \U$6227 ( \6949 , \5143 );
not \U$6228 ( \6950 , \6949 );
or \U$6229 ( \6951 , \6948 , \6950 );
buf \U$6230 ( \6952 , \3095 );
buf \U$6231 ( \6953 , \6516 );
nand \U$6232 ( \6954 , \6952 , \6953 );
buf \U$6233 ( \6955 , \6954 );
buf \U$6234 ( \6956 , \6955 );
nand \U$6235 ( \6957 , \6951 , \6956 );
buf \U$6236 ( \6958 , \6957 );
buf \U$6237 ( \6959 , \6958 );
not \U$6238 ( \6960 , \6959 );
not \U$6239 ( \6961 , \1400 );
nand \U$6240 ( \6962 , \6961 , \5573 );
buf \U$6241 ( \6963 , \6962 );
buf \U$6242 ( \6964 , \2067 );
and \U$6243 ( \6965 , \6963 , \6964 );
buf \U$6244 ( \6966 , \1400 );
not \U$6245 ( \6967 , \6966 );
buf \U$6246 ( \6968 , \5321 );
not \U$6247 ( \6969 , \6968 );
or \U$6248 ( \6970 , \6967 , \6969 );
buf \U$6249 ( \6971 , \1107 );
nand \U$6250 ( \6972 , \6970 , \6971 );
buf \U$6251 ( \6973 , \6972 );
buf \U$6252 ( \6974 , \6973 );
nor \U$6253 ( \6975 , \6965 , \6974 );
buf \U$6254 ( \6976 , \6975 );
buf \U$6255 ( \6977 , \6976 );
and \U$6256 ( \6978 , \6052 , RI9155b00_677);
and \U$6257 ( \6979 , \5430 , RI9156280_693);
nor \U$6258 ( \6980 , \6978 , \6979 );
and \U$6259 ( \6981 , \4644 , RI9154c00_645);
and \U$6260 ( \6982 , \1765 , RI9155380_661);
nor \U$6261 ( \6983 , \6981 , \6982 );
nand \U$6262 ( \6984 , \6980 , \6983 );
and \U$6263 ( \6985 , \5434 , RI9156a00_709);
not \U$6264 ( \6986 , RI9157180_725);
nor \U$6265 ( \6987 , \6986 , \1199 );
nor \U$6266 ( \6988 , \6985 , \6987 );
and \U$6267 ( \6989 , \1014 , RI9157900_741);
and \U$6268 ( \6990 , \5439 , RI9158080_757);
nor \U$6269 ( \6991 , \6989 , \6990 );
nand \U$6270 ( \6992 , \6988 , \6991 );
nor \U$6271 ( \6993 , \6984 , \6992 );
nand \U$6272 ( \6994 , \5463 , RI9151000_517);
nand \U$6273 ( \6995 , \5453 , RI9154480_629);
nand \U$6274 ( \6996 , \5451 , RI9153d00_613);
nand \U$6275 ( \6997 , \963 , RI9151780_533);
nand \U$6276 ( \6998 , \6994 , \6995 , \6996 , \6997 );
not \U$6277 ( \6999 , RI9152e00_581);
nor \U$6278 ( \7000 , \6999 , \1282 );
not \U$6279 ( \7001 , RI9153580_597);
nor \U$6280 ( \7002 , \7001 , \1285 );
nor \U$6281 ( \7003 , \7000 , \7002 );
and \U$6282 ( \7004 , \1302 , RI9151f00_549);
and \U$6283 ( \7005 , \928 , RI9152680_565);
nor \U$6284 ( \7006 , \7004 , \7005 );
nand \U$6285 ( \7007 , \7003 , \7006 );
nor \U$6286 ( \7008 , \6998 , \7007 );
nand \U$6287 ( \7009 , \6993 , \7008 );
buf \U$6288 ( \7010 , \7009 );
nand \U$6289 ( \7011 , \6977 , \7010 );
buf \U$6290 ( \7012 , \7011 );
buf \U$6291 ( \7013 , \7012 );
nand \U$6292 ( \7014 , \6960 , \7013 );
buf \U$6293 ( \7015 , \7014 );
buf \U$6294 ( \7016 , \7015 );
buf \U$6295 ( \7017 , \3223 );
not \U$6296 ( \7018 , \7017 );
buf \U$6297 ( \7019 , \2479 );
not \U$6298 ( \7020 , \7019 );
or \U$6299 ( \7021 , \7018 , \7020 );
buf \U$6300 ( \7022 , \3459 );
buf \U$6301 ( \7023 , \3276 );
nand \U$6302 ( \7024 , \7022 , \7023 );
buf \U$6303 ( \7025 , \7024 );
buf \U$6304 ( \7026 , \7025 );
nand \U$6305 ( \7027 , \7021 , \7026 );
buf \U$6306 ( \7028 , \7027 );
buf \U$6307 ( \7029 , \7028 );
not \U$6308 ( \7030 , \7029 );
buf \U$6309 ( \7031 , \2645 );
not \U$6310 ( \7032 , \7031 );
or \U$6311 ( \7033 , \7030 , \7032 );
buf \U$6312 ( \7034 , \2473 );
buf \U$6313 ( \7035 , \6547 );
nand \U$6314 ( \7036 , \7034 , \7035 );
buf \U$6315 ( \7037 , \7036 );
buf \U$6316 ( \7038 , \7037 );
nand \U$6317 ( \7039 , \7033 , \7038 );
buf \U$6318 ( \7040 , \7039 );
buf \U$6319 ( \7041 , \7040 );
and \U$6320 ( \7042 , \7016 , \7041 );
buf \U$6321 ( \7043 , \6958 );
not \U$6322 ( \7044 , \7043 );
buf \U$6323 ( \7045 , \7012 );
nor \U$6324 ( \7046 , \7044 , \7045 );
buf \U$6325 ( \7047 , \7046 );
buf \U$6326 ( \7048 , \7047 );
nor \U$6327 ( \7049 , \7042 , \7048 );
buf \U$6328 ( \7050 , \7049 );
buf \U$6329 ( \7051 , \7050 );
not \U$6330 ( \7052 , \7051 );
buf \U$6331 ( \7053 , \6684 );
not \U$6332 ( \7054 , \7053 );
buf \U$6333 ( \7055 , \6659 );
not \U$6334 ( \7056 , \7055 );
buf \U$6335 ( \7057 , \7056 );
buf \U$6336 ( \7058 , \7057 );
not \U$6337 ( \7059 , \7058 );
or \U$6338 ( \7060 , \7054 , \7059 );
buf \U$6339 ( \7061 , \6681 );
buf \U$6340 ( \7062 , \6659 );
nand \U$6341 ( \7063 , \7061 , \7062 );
buf \U$6342 ( \7064 , \7063 );
buf \U$6343 ( \7065 , \7064 );
nand \U$6344 ( \7066 , \7060 , \7065 );
buf \U$6345 ( \7067 , \7066 );
buf \U$6346 ( \7068 , \7067 );
buf \U$6347 ( \7069 , \6710 );
not \U$6348 ( \7070 , \7069 );
buf \U$6349 ( \7071 , \7070 );
buf \U$6350 ( \7072 , \7071 );
and \U$6351 ( \7073 , \7068 , \7072 );
not \U$6352 ( \7074 , \7068 );
buf \U$6353 ( \7075 , \6710 );
and \U$6354 ( \7076 , \7074 , \7075 );
nor \U$6355 ( \7077 , \7073 , \7076 );
buf \U$6356 ( \7078 , \7077 );
buf \U$6357 ( \7079 , \7078 );
and \U$6358 ( \7080 , \4644 , RI9154b88_644);
and \U$6359 ( \7081 , \984 , RI9155308_660);
nor \U$6360 ( \7082 , \7080 , \7081 );
and \U$6361 ( \7083 , \5428 , RI9155a88_676);
and \U$6362 ( \7084 , \5430 , RI9156208_692);
nor \U$6363 ( \7085 , \7083 , \7084 );
and \U$6364 ( \7086 , \5434 , RI9156988_708);
and \U$6365 ( \7087 , \2052 , RI9157108_724);
nor \U$6366 ( \7088 , \7086 , \7087 );
and \U$6367 ( \7089 , \1014 , RI9157888_740);
and \U$6368 ( \7090 , \5439 , RI9158008_756);
nor \U$6369 ( \7091 , \7089 , \7090 );
and \U$6370 ( \7092 , \7082 , \7085 , \7088 , \7091 );
and \U$6371 ( \7093 , RI9153508_596, \1218 );
not \U$6372 ( \7094 , \952 );
and \U$6373 ( \7095 , RI9152d88_580, \7094 );
not \U$6374 ( \7096 , RI9154408_628);
not \U$6375 ( \7097 , \5453 );
or \U$6376 ( \7098 , \7096 , \7097 );
not \U$6377 ( \7099 , \6069 );
nand \U$6378 ( \7100 , \7099 , RI9153c88_612);
nand \U$6379 ( \7101 , \7098 , \7100 );
nor \U$6380 ( \7102 , \7093 , \7095 , \7101 );
and \U$6381 ( \7103 , \5463 , RI9150f88_516);
and \U$6382 ( \7104 , \963 , RI9151708_532);
nor \U$6383 ( \7105 , \7103 , \7104 );
not \U$6384 ( \7106 , \922 );
and \U$6385 ( \7107 , \7106 , RI9151e88_548);
and \U$6386 ( \7108 , \1623 , RI9152608_564);
nor \U$6387 ( \7109 , \7107 , \7108 );
and \U$6388 ( \7110 , \7102 , \7105 , \7109 );
nand \U$6389 ( \7111 , \7092 , \7110 );
buf \U$6390 ( \7112 , \7111 );
buf \U$6391 ( \7113 , \1193 );
buf \U$6392 ( \7114 , \5321 );
and \U$6393 ( \7115 , \7113 , \7114 );
buf \U$6394 ( \7116 , \7115 );
buf \U$6395 ( \7117 , \7116 );
xor \U$6396 ( \7118 , \7112 , \7117 );
buf \U$6397 ( \7119 , \5388 );
not \U$6398 ( \7120 , \7119 );
buf \U$6399 ( \7121 , \7120 );
buf \U$6400 ( \7122 , \7121 );
not \U$6401 ( \7123 , \7122 );
buf \U$6402 ( \7124 , \6097 );
not \U$6403 ( \7125 , \7124 );
buf \U$6404 ( \7126 , \5621 );
not \U$6405 ( \7127 , \7126 );
or \U$6406 ( \7128 , \7125 , \7127 );
buf \U$6407 ( \7129 , \5334 );
buf \U$6408 ( \7130 , \1024 );
nand \U$6409 ( \7131 , \7129 , \7130 );
buf \U$6410 ( \7132 , \7131 );
buf \U$6411 ( \7133 , \7132 );
nand \U$6412 ( \7134 , \7128 , \7133 );
buf \U$6413 ( \7135 , \7134 );
buf \U$6414 ( \7136 , \7135 );
not \U$6415 ( \7137 , \7136 );
or \U$6416 ( \7138 , \7123 , \7137 );
buf \U$6417 ( \7139 , \6649 );
buf \U$6418 ( \7140 , \5398 );
nand \U$6419 ( \7141 , \7139 , \7140 );
buf \U$6420 ( \7142 , \7141 );
buf \U$6421 ( \7143 , \7142 );
nand \U$6422 ( \7144 , \7138 , \7143 );
buf \U$6423 ( \7145 , \7144 );
buf \U$6424 ( \7146 , \7145 );
and \U$6425 ( \7147 , \7118 , \7146 );
and \U$6426 ( \7148 , \7112 , \7117 );
or \U$6427 ( \7149 , \7147 , \7148 );
buf \U$6428 ( \7150 , \7149 );
buf \U$6429 ( \7151 , \7150 );
not \U$6430 ( \7152 , \7151 );
buf \U$6431 ( \7153 , \7152 );
buf \U$6432 ( \7154 , \7153 );
nand \U$6433 ( \7155 , \7079 , \7154 );
buf \U$6434 ( \7156 , \7155 );
buf \U$6435 ( \7157 , \7156 );
nand \U$6436 ( \7158 , \7052 , \7157 );
buf \U$6437 ( \7159 , \7158 );
buf \U$6438 ( \7160 , \7159 );
buf \U$6439 ( \7161 , \7078 );
not \U$6440 ( \7162 , \7161 );
buf \U$6441 ( \7163 , \7162 );
buf \U$6442 ( \7164 , \7163 );
buf \U$6443 ( \7165 , \7150 );
nand \U$6444 ( \7166 , \7164 , \7165 );
buf \U$6445 ( \7167 , \7166 );
buf \U$6446 ( \7168 , \7167 );
nand \U$6447 ( \7169 , \7160 , \7168 );
buf \U$6448 ( \7170 , \7169 );
buf \U$6452 ( \7171 , \7170 );
nand \U$6453 ( \7172 , \6942 , \7171 );
buf \U$6454 ( \7173 , \7172 );
buf \U$6455 ( \7174 , \7173 );
buf \U$6456 ( \7175 , \6925 );
not \U$6457 ( \7176 , \7175 );
buf \U$6458 ( \7177 , \6939 );
not \U$6459 ( \7178 , \7177 );
buf \U$6460 ( \7179 , \7178 );
buf \U$6461 ( \7180 , \7179 );
nand \U$6462 ( \7181 , \7176 , \7180 );
buf \U$6463 ( \7182 , \7181 );
buf \U$6464 ( \7183 , \7182 );
nand \U$6465 ( \7184 , \7174 , \7183 );
buf \U$6466 ( \7185 , \7184 );
buf \U$6467 ( \7186 , \7185 );
not \U$6468 ( \7187 , \7186 );
buf \U$6469 ( \7188 , \7187 );
buf \U$6470 ( \7189 , \7188 );
buf \U$6471 ( \7190 , \6380 );
not \U$6472 ( \7191 , \7190 );
buf \U$6473 ( \7192 , \6398 );
not \U$6474 ( \7193 , \7192 );
buf \U$6475 ( \7194 , \7193 );
buf \U$6476 ( \7195 , \7194 );
not \U$6477 ( \7196 , \7195 );
or \U$6478 ( \7197 , \7191 , \7196 );
buf \U$6479 ( \7198 , \6398 );
buf \U$6480 ( \7199 , \6377 );
nand \U$6481 ( \7200 , \7198 , \7199 );
buf \U$6482 ( \7201 , \7200 );
buf \U$6483 ( \7202 , \7201 );
nand \U$6484 ( \7203 , \7197 , \7202 );
buf \U$6485 ( \7204 , \7203 );
buf \U$6486 ( \7205 , \7204 );
buf \U$6487 ( \7206 , \6412 );
not \U$6488 ( \7207 , \7206 );
buf \U$6489 ( \7208 , \7207 );
buf \U$6490 ( \7209 , \7208 );
and \U$6491 ( \7210 , \7205 , \7209 );
not \U$6492 ( \7211 , \7205 );
buf \U$6493 ( \7212 , \6412 );
and \U$6494 ( \7213 , \7211 , \7212 );
nor \U$6495 ( \7214 , \7210 , \7213 );
buf \U$6496 ( \7215 , \7214 );
buf \U$6497 ( \7216 , \7215 );
nand \U$6498 ( \7217 , \7189 , \7216 );
buf \U$6499 ( \7218 , \7217 );
buf \U$6500 ( \7219 , \7218 );
not \U$6501 ( \7220 , \7219 );
buf \U$6502 ( \7221 , \6611 );
not \U$6503 ( \7222 , \7221 );
buf \U$6504 ( \7223 , \6729 );
not \U$6505 ( \7224 , \7223 );
buf \U$6506 ( \7225 , \7224 );
buf \U$6507 ( \7226 , \7225 );
not \U$6508 ( \7227 , \7226 );
or \U$6509 ( \7228 , \7222 , \7227 );
buf \U$6510 ( \7229 , \7225 );
buf \U$6511 ( \7230 , \6611 );
or \U$6512 ( \7231 , \7229 , \7230 );
nand \U$6513 ( \7232 , \7228 , \7231 );
buf \U$6514 ( \7233 , \7232 );
buf \U$6515 ( \7234 , \7233 );
buf \U$6516 ( \7235 , \6622 );
and \U$6517 ( \7236 , \7234 , \7235 );
not \U$6518 ( \7237 , \7234 );
buf \U$6519 ( \7238 , \6619 );
and \U$6520 ( \7239 , \7237 , \7238 );
nor \U$6521 ( \7240 , \7236 , \7239 );
buf \U$6522 ( \7241 , \7240 );
buf \U$6523 ( \7242 , \7241 );
not \U$6524 ( \7243 , \7242 );
or \U$6525 ( \7244 , \7220 , \7243 );
buf \U$6526 ( \7245 , \7188 );
not \U$6527 ( \7246 , \7245 );
buf \U$6528 ( \7247 , \7215 );
not \U$6529 ( \7248 , \7247 );
buf \U$6530 ( \7249 , \7248 );
buf \U$6531 ( \7250 , \7249 );
nand \U$6532 ( \7251 , \7246 , \7250 );
buf \U$6533 ( \7252 , \7251 );
buf \U$6534 ( \7253 , \7252 );
nand \U$6535 ( \7254 , \7244 , \7253 );
buf \U$6536 ( \7255 , \7254 );
buf \U$6537 ( \7256 , \7255 );
nand \U$6538 ( \7257 , \6763 , \7256 );
buf \U$6539 ( \7258 , \7257 );
buf \U$6540 ( \7259 , \7258 );
buf \U$6541 ( \7260 , \6041 );
buf \U$6542 ( \7261 , \6424 );
xor \U$6543 ( \7262 , \7260 , \7261 );
buf \U$6544 ( \7263 , \6038 );
xnor \U$6545 ( \7264 , \7262 , \7263 );
buf \U$6546 ( \7265 , \7264 );
buf \U$6547 ( \7266 , \7265 );
xor \U$6548 ( \7267 , \6460 , \6736 );
and \U$6549 ( \7268 , \7267 , \6760 );
and \U$6550 ( \7269 , \6460 , \6736 );
or \U$6551 ( \7270 , \7268 , \7269 );
buf \U$6552 ( \7271 , \7270 );
buf \U$6553 ( \7272 , \7271 );
nand \U$6554 ( \7273 , \7266 , \7272 );
buf \U$6555 ( \7274 , \7273 );
buf \U$6556 ( \7275 , \7274 );
nand \U$6557 ( \7276 , \7259 , \7275 );
buf \U$6558 ( \7277 , \7276 );
buf \U$6559 ( \7278 , \7277 );
buf \U$6560 ( \7279 , \6031 );
buf \U$6561 ( \7280 , \6435 );
nand \U$6562 ( \7281 , \7279 , \7280 );
buf \U$6563 ( \7282 , \7281 );
buf \U$6564 ( \7283 , \7282 );
buf \U$6565 ( \7284 , \6027 );
buf \U$6566 ( \7285 , \7271 );
not \U$6567 ( \7286 , \7285 );
buf \U$6568 ( \7287 , \7265 );
not \U$6569 ( \7288 , \7287 );
buf \U$6570 ( \7289 , \7288 );
buf \U$6571 ( \7290 , \7289 );
nand \U$6572 ( \7291 , \7286 , \7290 );
buf \U$6573 ( \7292 , \7291 );
buf \U$6574 ( \7293 , \7292 );
nand \U$6575 ( \7294 , \7278 , \7283 , \7284 , \7293 );
buf \U$6576 ( \7295 , \7294 );
buf \U$6577 ( \7296 , \7295 );
buf \U$6578 ( \7297 , \4505 );
buf \U$6579 ( \7298 , \4944 );
xor \U$6580 ( \7299 , \7297 , \7298 );
buf \U$6581 ( \7300 , \4340 );
xnor \U$6582 ( \7301 , \7299 , \7300 );
buf \U$6583 ( \7302 , \7301 );
buf \U$6584 ( \7303 , \7302 );
buf \U$6585 ( \7304 , \4934 );
not \U$6586 ( \7305 , \7304 );
buf \U$6587 ( \7306 , \4741 );
not \U$6588 ( \7307 , \7306 );
buf \U$6589 ( \7308 , \4751 );
not \U$6590 ( \7309 , \7308 );
or \U$6591 ( \7310 , \7307 , \7309 );
buf \U$6592 ( \7311 , \4741 );
buf \U$6593 ( \7312 , \4751 );
or \U$6594 ( \7313 , \7311 , \7312 );
nand \U$6595 ( \7314 , \7310 , \7313 );
buf \U$6596 ( \7315 , \7314 );
buf \U$6597 ( \7316 , \7315 );
not \U$6598 ( \7317 , \7316 );
buf \U$6599 ( \7318 , \7317 );
buf \U$6600 ( \7319 , \7318 );
not \U$6601 ( \7320 , \7319 );
or \U$6602 ( \7321 , \7305 , \7320 );
nand \U$6603 ( \7322 , \4922 , \4931 , \7315 );
buf \U$6604 ( \7323 , \7322 );
nand \U$6605 ( \7324 , \7321 , \7323 );
buf \U$6606 ( \7325 , \7324 );
buf \U$6607 ( \7326 , \7325 );
xor \U$6608 ( \7327 , \4368 , \4375 );
xor \U$6609 ( \7328 , \7327 , \4501 );
buf \U$6610 ( \7329 , \7328 );
buf \U$6611 ( \7330 , \7329 );
or \U$6612 ( \7331 , \7326 , \7330 );
buf \U$6613 ( \7332 , \7331 );
buf \U$6614 ( \7333 , \7332 );
buf \U$6615 ( \7334 , \5796 );
not \U$6616 ( \7335 , \7334 );
not \U$6617 ( \7336 , \5804 );
buf \U$6618 ( \7337 , \7336 );
not \U$6619 ( \7338 , \7337 );
or \U$6620 ( \7339 , \7335 , \7338 );
buf \U$6621 ( \7340 , \5907 );
buf \U$6622 ( \7341 , \5804 );
buf \U$6623 ( \7342 , \5793 );
nand \U$6624 ( \7343 , \7341 , \7342 );
buf \U$6625 ( \7344 , \7343 );
buf \U$6626 ( \7345 , \7344 );
nand \U$6627 ( \7346 , \7340 , \7345 );
buf \U$6628 ( \7347 , \7346 );
buf \U$6629 ( \7348 , \7347 );
nand \U$6630 ( \7349 , \7339 , \7348 );
buf \U$6631 ( \7350 , \7349 );
buf \U$6632 ( \7351 , \7350 );
not \U$6633 ( \7352 , \7351 );
buf \U$6634 ( \7353 , \7352 );
buf \U$6635 ( \7354 , \7353 );
not \U$6636 ( \7355 , \7354 );
buf \U$6637 ( \7356 , \7355 );
buf \U$6638 ( \7357 , \7356 );
and \U$6639 ( \7358 , \7333 , \7357 );
buf \U$6640 ( \7359 , \7329 );
buf \U$6641 ( \7360 , \7325 );
and \U$6642 ( \7361 , \7359 , \7360 );
buf \U$6643 ( \7362 , \7361 );
buf \U$6644 ( \7363 , \7362 );
nor \U$6645 ( \7364 , \7358 , \7363 );
buf \U$6646 ( \7365 , \7364 );
buf \U$6647 ( \7366 , \7365 );
nand \U$6648 ( \7367 , \7303 , \7366 );
buf \U$6649 ( \7368 , \7367 );
buf \U$6650 ( \7369 , \7368 );
not \U$6651 ( \7370 , \7369 );
buf \U$6652 ( \7371 , \7353 );
not \U$6653 ( \7372 , \7371 );
xor \U$6654 ( \7373 , \7359 , \7360 );
buf \U$6655 ( \7374 , \7373 );
buf \U$6656 ( \7375 , \7374 );
not \U$6657 ( \7376 , \7375 );
or \U$6658 ( \7377 , \7372 , \7376 );
buf \U$6659 ( \7378 , \7374 );
buf \U$6660 ( \7379 , \7353 );
or \U$6661 ( \7380 , \7378 , \7379 );
nand \U$6662 ( \7381 , \7377 , \7380 );
buf \U$6663 ( \7382 , \7381 );
buf \U$6664 ( \7383 , \7382 );
not \U$6665 ( \7384 , \5918 );
buf \U$6666 ( \7385 , \4964 );
not \U$6667 ( \7386 , \7385 );
or \U$6668 ( \7387 , \7384 , \7386 );
not \U$6669 ( \7388 , \7385 );
not \U$6670 ( \7389 , \7388 );
not \U$6671 ( \7390 , \5917 );
or \U$6672 ( \7391 , \7389 , \7390 );
buf \U$6675 ( \7392 , \5785 );
nand \U$6676 ( \7393 , \7391 , \7392 );
nand \U$6677 ( \7394 , \7387 , \7393 );
buf \U$6678 ( \7395 , \7394 );
and \U$6679 ( \7396 , \7383 , \7395 );
buf \U$6680 ( \7397 , \7396 );
buf \U$6681 ( \7398 , \7397 );
not \U$6682 ( \7399 , \7398 );
or \U$6683 ( \7400 , \7370 , \7399 );
buf \U$6684 ( \7401 , \7302 );
not \U$6685 ( \7402 , \7401 );
buf \U$6686 ( \7403 , \7402 );
buf \U$6687 ( \7404 , \7403 );
buf \U$6688 ( \7405 , \7365 );
not \U$6689 ( \7406 , \7405 );
buf \U$6690 ( \7407 , \7406 );
buf \U$6691 ( \7408 , \7407 );
nand \U$6692 ( \7409 , \7404 , \7408 );
buf \U$6693 ( \7410 , \7409 );
buf \U$6694 ( \7411 , \7410 );
nand \U$6695 ( \7412 , \7400 , \7411 );
buf \U$6696 ( \7413 , \7412 );
buf \U$6697 ( \7414 , \7413 );
not \U$6698 ( \7415 , \7414 );
buf \U$6699 ( \7416 , \7415 );
buf \U$6700 ( \7417 , \7416 );
nand \U$6701 ( \7418 , \6445 , \7296 , \7417 );
buf \U$6702 ( \7419 , \7418 );
buf \U$6703 ( \7420 , \7419 );
not \U$6704 ( \7421 , \7420 );
buf \U$6705 ( \7422 , \7416 );
buf \U$6706 ( \7423 , \7382 );
not \U$6707 ( \7424 , \7423 );
buf \U$6708 ( \7425 , \7424 );
buf \U$6709 ( \7426 , \7425 );
buf \U$6710 ( \7427 , \7394 );
not \U$6711 ( \7428 , \7427 );
buf \U$6712 ( \7429 , \7428 );
buf \U$6713 ( \7430 , \7429 );
nand \U$6714 ( \7431 , \7426 , \7430 );
buf \U$6715 ( \7432 , \7431 );
and \U$6716 ( \7433 , \7432 , \7368 );
not \U$6717 ( \7434 , \7433 );
buf \U$6718 ( \7435 , \7434 );
buf \U$6719 ( \7436 , \4957 );
and \U$6720 ( \7437 , \7422 , \7435 , \7436 );
buf \U$6722 ( \7438 , \3924 );
buf \U$6723 ( \7439 , \4312 );
nor \U$6724 ( \7440 , \7438 , \7439 );
buf \U$6725 ( \7441 , \7440 );
buf \U$6726 ( \7442 , \7441 );
not \U$6727 ( \7443 , \7442 );
or \U$6728 ( \7444 , 1'b0 , \7443 );
buf \U$6729 ( \7445 , \4954 );
buf \U$6730 ( \7446 , \4319 );
not \U$6731 ( \7447 , \7446 );
buf \U$6732 ( \7448 , \7447 );
buf \U$6733 ( \7449 , \7448 );
not \U$6734 ( \7450 , \4948 );
buf \U$6735 ( \7451 , \7450 );
nand \U$6736 ( \7452 , \7449 , \7451 );
buf \U$6737 ( \7453 , \7452 );
buf \U$6738 ( \7454 , \7453 );
or \U$6739 ( \7455 , \7445 , \7454 );
nand \U$6740 ( \7456 , \7444 , \7455 );
buf \U$6741 ( \7457 , \7456 );
buf \U$6742 ( \7458 , \7457 );
nor \U$6743 ( \7459 , \7437 , \7458 );
buf \U$6744 ( \7460 , \7459 );
buf \U$6745 ( \7461 , \7460 );
not \U$6746 ( \7462 , \7461 );
or \U$6747 ( \7463 , \7421 , \7462 );
buf \U$6748 ( \7464 , \7433 );
and \U$6749 ( \7465 , \7448 , \7450 );
nor \U$6750 ( \7466 , \7465 , \7441 );
buf \U$6751 ( \7467 , \7466 );
and \U$6752 ( \7468 , \7464 , \7467 );
buf \U$6753 ( \7469 , \7468 );
buf \U$6754 ( \7470 , \7469 );
not \U$6755 ( \7471 , \6762 );
buf \U$6756 ( \7472 , \7471 );
buf \U$6757 ( \7473 , \7255 );
not \U$6758 ( \7474 , \7473 );
buf \U$6759 ( \7475 , \7474 );
buf \U$6760 ( \7476 , \7475 );
nand \U$6761 ( \7477 , \7472 , \7476 );
buf \U$6762 ( \7478 , \7477 );
and \U$6763 ( \7479 , \7292 , \7478 , \6027 , \7282 );
buf \U$6764 ( \7480 , \7479 );
xor \U$6765 ( \7481 , \7112 , \7117 );
xor \U$6766 ( \7482 , \7481 , \7146 );
buf \U$6767 ( \7483 , \7482 );
buf \U$6768 ( \7484 , \7483 );
buf \U$6769 ( \7485 , \7121 );
not \U$6770 ( \7486 , \7485 );
buf \U$6771 ( \7487 , \2521 );
not \U$6772 ( \7488 , \7487 );
buf \U$6773 ( \7489 , \5330 );
not \U$6774 ( \7490 , \7489 );
or \U$6775 ( \7491 , \7488 , \7490 );
buf \U$6776 ( \7492 , \4794 );
buf \U$6777 ( \7493 , \1999 );
nand \U$6778 ( \7494 , \7492 , \7493 );
buf \U$6779 ( \7495 , \7494 );
buf \U$6780 ( \7496 , \7495 );
nand \U$6781 ( \7497 , \7491 , \7496 );
buf \U$6782 ( \7498 , \7497 );
buf \U$6783 ( \7499 , \7498 );
not \U$6784 ( \7500 , \7499 );
or \U$6785 ( \7501 , \7486 , \7500 );
buf \U$6786 ( \7502 , \7135 );
buf \U$6787 ( \7503 , \5398 );
nand \U$6788 ( \7504 , \7502 , \7503 );
buf \U$6789 ( \7505 , \7504 );
buf \U$6790 ( \7506 , \7505 );
nand \U$6791 ( \7507 , \7501 , \7506 );
buf \U$6792 ( \7508 , \7507 );
buf \U$6793 ( \7509 , \7508 );
not \U$6794 ( \7510 , \7509 );
buf \U$6795 ( \7511 , \7510 );
buf \U$6796 ( \7512 , \7511 );
not \U$6797 ( \7513 , \7512 );
buf \U$6798 ( \7514 , \6976 );
not \U$6799 ( \7515 , \7514 );
buf \U$6800 ( \7516 , \7009 );
not \U$6801 ( \7517 , \7516 );
buf \U$6802 ( \7518 , \7517 );
buf \U$6803 ( \7519 , \7518 );
not \U$6804 ( \7520 , \7519 );
and \U$6805 ( \7521 , \7515 , \7520 );
buf \U$6806 ( \7522 , \6976 );
buf \U$6807 ( \7523 , \7518 );
and \U$6808 ( \7524 , \7522 , \7523 );
nor \U$6809 ( \7525 , \7521 , \7524 );
buf \U$6810 ( \7526 , \7525 );
buf \U$6811 ( \7527 , \7526 );
not \U$6812 ( \7528 , \7527 );
or \U$6813 ( \7529 , \7513 , \7528 );
buf \U$6814 ( \7530 , \2758 );
not \U$6815 ( \7531 , \7530 );
buf \U$6816 ( \7532 , \4516 );
not \U$6817 ( \7533 , \7532 );
or \U$6818 ( \7534 , \7531 , \7533 );
buf \U$6819 ( \7535 , \5603 );
buf \U$6820 ( \7536 , \2853 );
nand \U$6821 ( \7537 , \7535 , \7536 );
buf \U$6822 ( \7538 , \7537 );
buf \U$6823 ( \7539 , \7538 );
nand \U$6824 ( \7540 , \7534 , \7539 );
buf \U$6825 ( \7541 , \7540 );
buf \U$6826 ( \7542 , \7541 );
not \U$6827 ( \7543 , \7542 );
buf \U$6828 ( \7544 , \5615 );
not \U$6829 ( \7545 , \7544 );
or \U$6830 ( \7546 , \7543 , \7545 );
buf \U$6831 ( \7547 , \3095 );
buf \U$6832 ( \7548 , \6946 );
nand \U$6833 ( \7549 , \7547 , \7548 );
buf \U$6834 ( \7550 , \7549 );
buf \U$6835 ( \7551 , \7550 );
nand \U$6836 ( \7552 , \7546 , \7551 );
buf \U$6837 ( \7553 , \7552 );
buf \U$6838 ( \7554 , \7553 );
nand \U$6839 ( \7555 , \7529 , \7554 );
buf \U$6840 ( \7556 , \7555 );
buf \U$6841 ( \7557 , \7556 );
buf \U$6842 ( \7558 , \7526 );
buf \U$6843 ( \7559 , \7511 );
or \U$6844 ( \7560 , \7558 , \7559 );
buf \U$6845 ( \7561 , \7560 );
buf \U$6846 ( \7562 , \7561 );
nand \U$6847 ( \7563 , \7557 , \7562 );
buf \U$6848 ( \7564 , \7563 );
buf \U$6849 ( \7565 , \7564 );
xor \U$6850 ( \7566 , \7484 , \7565 );
buf \U$6851 ( \7567 , \4070 );
not \U$6852 ( \7568 , \7567 );
buf \U$6853 ( \7569 , \4381 );
not \U$6854 ( \7570 , \7569 );
or \U$6855 ( \7571 , \7568 , \7570 );
buf \U$6856 ( \7572 , \2479 );
buf \U$6857 ( \7573 , \3444 );
nand \U$6858 ( \7574 , \7572 , \7573 );
buf \U$6859 ( \7575 , \7574 );
buf \U$6860 ( \7576 , \7575 );
nand \U$6861 ( \7577 , \7571 , \7576 );
buf \U$6862 ( \7578 , \7577 );
buf \U$6863 ( \7579 , \7578 );
not \U$6864 ( \7580 , \7579 );
buf \U$6865 ( \7581 , \3288 );
not \U$6866 ( \7582 , \7581 );
or \U$6867 ( \7583 , \7580 , \7582 );
buf \U$6868 ( \7584 , \7028 );
buf \U$6869 ( \7585 , \2473 );
nand \U$6870 ( \7586 , \7584 , \7585 );
buf \U$6871 ( \7587 , \7586 );
buf \U$6872 ( \7588 , \7587 );
nand \U$6873 ( \7589 , \7583 , \7588 );
buf \U$6874 ( \7590 , \7589 );
buf \U$6875 ( \7591 , \7590 );
buf \U$6876 ( \7592 , \4678 );
not \U$6877 ( \7593 , \7592 );
buf \U$6878 ( \7594 , \2071 );
not \U$6879 ( \7595 , \7594 );
or \U$6880 ( \7596 , \7593 , \7595 );
buf \U$6881 ( \7597 , \2068 );
buf \U$6882 ( \7598 , \4863 );
nand \U$6883 ( \7599 , \7597 , \7598 );
buf \U$6884 ( \7600 , \7599 );
buf \U$6885 ( \7601 , \7600 );
nand \U$6886 ( \7602 , \7596 , \7601 );
buf \U$6887 ( \7603 , \7602 );
buf \U$6888 ( \7604 , \7603 );
not \U$6889 ( \7605 , \7604 );
buf \U$6890 ( \7606 , \2503 );
not \U$6891 ( \7607 , \7606 );
or \U$6892 ( \7608 , \7605 , \7607 );
buf \U$6893 ( \7609 , \2897 );
buf \U$6894 ( \7610 , \6864 );
nand \U$6895 ( \7611 , \7609 , \7610 );
buf \U$6896 ( \7612 , \7611 );
buf \U$6897 ( \7613 , \7612 );
nand \U$6898 ( \7614 , \7608 , \7613 );
buf \U$6899 ( \7615 , \7614 );
buf \U$6900 ( \7616 , \7615 );
xor \U$6901 ( \7617 , \7591 , \7616 );
buf \U$6902 ( \7618 , \1934 );
not \U$6903 ( \7619 , \7618 );
buf \U$6904 ( \7620 , \4282 );
not \U$6905 ( \7621 , \7620 );
or \U$6906 ( \7622 , \7619 , \7621 );
buf \U$6907 ( \7623 , \4278 );
buf \U$6908 ( \7624 , \1931 );
nand \U$6909 ( \7625 , \7623 , \7624 );
buf \U$6910 ( \7626 , \7625 );
buf \U$6911 ( \7627 , \7626 );
nand \U$6912 ( \7628 , \7622 , \7627 );
buf \U$6913 ( \7629 , \7628 );
buf \U$6914 ( \7630 , \7629 );
not \U$6915 ( \7631 , \7630 );
buf \U$6916 ( \7632 , \6578 );
not \U$6917 ( \7633 , \7632 );
or \U$6918 ( \7634 , \7631 , \7633 );
buf \U$6919 ( \7635 , \4581 );
buf \U$6920 ( \7636 , \6894 );
nand \U$6921 ( \7637 , \7635 , \7636 );
buf \U$6922 ( \7638 , \7637 );
buf \U$6923 ( \7639 , \7638 );
nand \U$6924 ( \7640 , \7634 , \7639 );
buf \U$6925 ( \7641 , \7640 );
buf \U$6926 ( \7642 , \7641 );
and \U$6927 ( \7643 , \7617 , \7642 );
and \U$6928 ( \7644 , \7591 , \7616 );
or \U$6929 ( \7645 , \7643 , \7644 );
buf \U$6930 ( \7646 , \7645 );
buf \U$6931 ( \7647 , \7646 );
xor \U$6932 ( \7648 , \7566 , \7647 );
buf \U$6933 ( \7649 , \7648 );
buf \U$6934 ( \7650 , \7649 );
and \U$6935 ( \7651 , \1669 , \4281 );
not \U$6936 ( \7652 , \1669 );
and \U$6937 ( \7653 , \7652 , \4278 );
or \U$6938 ( \7654 , \7651 , \7653 );
buf \U$6939 ( \7655 , \7654 );
not \U$6940 ( \7656 , \7655 );
buf \U$6941 ( \7657 , \5046 );
not \U$6942 ( \7658 , \7657 );
buf \U$6943 ( \7659 , \7658 );
buf \U$6944 ( \7660 , \7659 );
not \U$6945 ( \7661 , \7660 );
or \U$6946 ( \7662 , \7656 , \7661 );
buf \U$6947 ( \7663 , \7629 );
buf \U$6948 ( \7664 , \6582 );
nand \U$6949 ( \7665 , \7663 , \7664 );
buf \U$6950 ( \7666 , \7665 );
buf \U$6951 ( \7667 , \7666 );
nand \U$6952 ( \7668 , \7662 , \7667 );
buf \U$6953 ( \7669 , \7668 );
buf \U$6954 ( \7670 , \7669 );
not \U$6955 ( \7671 , \7670 );
buf \U$6956 ( \7672 , \4848 );
not \U$6957 ( \7673 , \7672 );
buf \U$6958 ( \7674 , \2071 );
not \U$6959 ( \7675 , \7674 );
or \U$6960 ( \7676 , \7673 , \7675 );
buf \U$6961 ( \7677 , \2884 );
buf \U$6962 ( \7678 , \4991 );
nand \U$6963 ( \7679 , \7677 , \7678 );
buf \U$6964 ( \7680 , \7679 );
buf \U$6965 ( \7681 , \7680 );
nand \U$6966 ( \7682 , \7676 , \7681 );
buf \U$6967 ( \7683 , \7682 );
buf \U$6968 ( \7684 , \7683 );
not \U$6969 ( \7685 , \7684 );
buf \U$6970 ( \7686 , \2201 );
not \U$6971 ( \7687 , \7686 );
or \U$6972 ( \7688 , \7685 , \7687 );
buf \U$6973 ( \7689 , \2214 );
buf \U$6974 ( \7690 , \7603 );
nand \U$6975 ( \7691 , \7689 , \7690 );
buf \U$6976 ( \7692 , \7691 );
buf \U$6977 ( \7693 , \7692 );
nand \U$6978 ( \7694 , \7688 , \7693 );
buf \U$6979 ( \7695 , \7694 );
buf \U$6980 ( \7696 , \7695 );
not \U$6981 ( \7697 , \7696 );
buf \U$6982 ( \7698 , \7697 );
buf \U$6983 ( \7699 , \7698 );
nand \U$6984 ( \7700 , \7671 , \7699 );
buf \U$6985 ( \7701 , \7700 );
buf \U$6986 ( \7702 , \7701 );
not \U$6987 ( \7703 , \7702 );
buf \U$6988 ( \7704 , \1795 );
not \U$6989 ( \7705 , \7704 );
buf \U$6990 ( \7706 , \5330 );
not \U$6991 ( \7707 , \7706 );
or \U$6992 ( \7708 , \7705 , \7707 );
buf \U$6993 ( \7709 , \4794 );
buf \U$6994 ( \7710 , \1792 );
nand \U$6995 ( \7711 , \7709 , \7710 );
buf \U$6996 ( \7712 , \7711 );
buf \U$6997 ( \7713 , \7712 );
nand \U$6998 ( \7714 , \7708 , \7713 );
buf \U$6999 ( \7715 , \7714 );
buf \U$7000 ( \7716 , \7715 );
not \U$7001 ( \7717 , \7716 );
buf \U$7002 ( \7718 , \7121 );
not \U$7003 ( \7719 , \7718 );
or \U$7004 ( \7720 , \7717 , \7719 );
buf \U$7005 ( \7721 , \1862 );
not \U$7006 ( \7722 , \7721 );
buf \U$7007 ( \7723 , \5330 );
not \U$7008 ( \7724 , \7723 );
or \U$7009 ( \7725 , \7722 , \7724 );
buf \U$7010 ( \7726 , \5334 );
buf \U$7011 ( \7727 , \2670 );
nand \U$7012 ( \7728 , \7726 , \7727 );
buf \U$7013 ( \7729 , \7728 );
buf \U$7014 ( \7730 , \7729 );
nand \U$7015 ( \7731 , \7725 , \7730 );
buf \U$7016 ( \7732 , \7731 );
buf \U$7017 ( \7733 , \7732 );
buf \U$7018 ( \7734 , \5398 );
nand \U$7019 ( \7735 , \7733 , \7734 );
buf \U$7020 ( \7736 , \7735 );
buf \U$7021 ( \7737 , \7736 );
nand \U$7022 ( \7738 , \7720 , \7737 );
buf \U$7023 ( \7739 , \7738 );
buf \U$7026 ( \7740 , \7739 );
buf \U$7027 ( \7741 , \7740 );
not \U$7028 ( \7742 , \7741 );
buf \U$7029 ( \7743 , \7742 );
buf \U$7030 ( \7744 , \7743 );
not \U$7031 ( \7745 , \7744 );
and \U$7032 ( \7746 , \4644 , RI9154cf0_647);
and \U$7033 ( \7747 , \1765 , RI9155470_663);
nor \U$7034 ( \7748 , \7746 , \7747 );
and \U$7035 ( \7749 , \6052 , RI9155bf0_679);
and \U$7036 ( \7750 , \5430 , RI9156370_695);
nor \U$7037 ( \7751 , \7749 , \7750 );
and \U$7038 ( \7752 , \4003 , RI9156af0_711);
and \U$7039 ( \7753 , \2052 , RI9157270_727);
nor \U$7040 ( \7754 , \7752 , \7753 );
and \U$7041 ( \7755 , \6239 , RI91579f0_743);
and \U$7042 ( \7756 , \4011 , RI9158170_759);
nor \U$7043 ( \7757 , \7755 , \7756 );
and \U$7044 ( \7758 , \7748 , \7751 , \7754 , \7757 );
and \U$7045 ( \7759 , \5463 , RI91510f0_519);
and \U$7046 ( \7760 , \963 , RI9151870_535);
nor \U$7047 ( \7761 , \7759 , \7760 );
not \U$7048 ( \7762 , \929 );
and \U$7049 ( \7763 , \7762 , RI9152770_567);
not \U$7050 ( \7764 , RI9151ff0_551);
nor \U$7051 ( \7765 , \7764 , \6273 );
nor \U$7052 ( \7766 , \7763 , \7765 );
and \U$7053 ( \7767 , \7094 , RI9152ef0_583);
and \U$7054 ( \7768 , \1500 , RI9153670_599);
nor \U$7055 ( \7769 , \7767 , \7768 );
and \U$7056 ( \7770 , \5451 , RI9153df0_615);
and \U$7057 ( \7771 , \5453 , RI9154570_631);
nor \U$7058 ( \7772 , \7770 , \7771 );
and \U$7059 ( \7773 , \7761 , \7766 , \7769 , \7772 );
nand \U$7060 ( \7774 , \7758 , \7773 );
buf \U$7061 ( \7775 , \7774 );
not \U$7062 ( \7776 , \7775 );
buf \U$7063 ( \7777 , \7776 );
buf \U$7064 ( \7778 , \7777 );
not \U$7065 ( \7779 , \7778 );
buf \U$7066 ( \7780 , \2187 );
not \U$7067 ( \7781 , \7780 );
buf \U$7068 ( \7782 , \7781 );
buf \U$7069 ( \7783 , \7782 );
not \U$7070 ( \7784 , \7783 );
buf \U$7071 ( \7785 , \5472 );
not \U$7072 ( \7786 , \7785 );
or \U$7073 ( \7787 , \7784 , \7786 );
buf \U$7074 ( \7788 , \2067 );
nand \U$7075 ( \7789 , \7787 , \7788 );
buf \U$7076 ( \7790 , \7789 );
buf \U$7077 ( \7791 , \7790 );
not \U$7078 ( \7792 , \7791 );
buf \U$7079 ( \7793 , \7782 );
not \U$7080 ( \7794 , \7793 );
buf \U$7081 ( \7795 , \7794 );
buf \U$7082 ( \7796 , \7795 );
not \U$7083 ( \7797 , \7796 );
buf \U$7084 ( \7798 , \5321 );
not \U$7085 ( \7799 , \7798 );
buf \U$7086 ( \7800 , \7799 );
buf \U$7087 ( \7801 , \7800 );
not \U$7088 ( \7802 , \7801 );
or \U$7089 ( \7803 , \7797 , \7802 );
buf \U$7090 ( \7804 , \3276 );
nand \U$7091 ( \7805 , \7803 , \7804 );
buf \U$7092 ( \7806 , \7805 );
buf \U$7093 ( \7807 , \7806 );
nand \U$7094 ( \7808 , \7792 , \7807 );
buf \U$7095 ( \7809 , \7808 );
buf \U$7096 ( \7810 , \7809 );
not \U$7097 ( \7811 , \7810 );
buf \U$7098 ( \7812 , \7811 );
buf \U$7099 ( \7813 , \7812 );
not \U$7100 ( \7814 , \7813 );
or \U$7101 ( \7815 , \7779 , \7814 );
buf \U$7102 ( \7816 , \7809 );
buf \U$7103 ( \7817 , \7774 );
nand \U$7104 ( \7818 , \7816 , \7817 );
buf \U$7105 ( \7819 , \7818 );
buf \U$7106 ( \7820 , \7819 );
nand \U$7107 ( \7821 , \7815 , \7820 );
buf \U$7108 ( \7822 , \7821 );
buf \U$7109 ( \7823 , \7822 );
not \U$7110 ( \7824 , \7823 );
buf \U$7111 ( \7825 , \7824 );
buf \U$7112 ( \7826 , \7825 );
not \U$7113 ( \7827 , \7826 );
or \U$7114 ( \7828 , \7745 , \7827 );
buf \U$7115 ( \7829 , \3444 );
not \U$7116 ( \7830 , \7829 );
buf \U$7117 ( \7831 , \3134 );
not \U$7118 ( \7832 , \7831 );
buf \U$7119 ( \7833 , \7832 );
buf \U$7120 ( \7834 , \7833 );
not \U$7121 ( \7835 , \7834 );
or \U$7122 ( \7836 , \7830 , \7835 );
buf \U$7123 ( \7837 , \4516 );
not \U$7124 ( \7838 , \7837 );
buf \U$7125 ( \7839 , \7838 );
buf \U$7126 ( \7840 , \7839 );
buf \U$7127 ( \7841 , \4381 );
nand \U$7128 ( \7842 , \7840 , \7841 );
buf \U$7129 ( \7843 , \7842 );
buf \U$7130 ( \7844 , \7843 );
nand \U$7131 ( \7845 , \7836 , \7844 );
buf \U$7132 ( \7846 , \7845 );
buf \U$7133 ( \7847 , \7846 );
not \U$7134 ( \7848 , \7847 );
buf \U$7135 ( \7849 , \5615 );
not \U$7136 ( \7850 , \7849 );
or \U$7137 ( \7851 , \7848 , \7850 );
buf \U$7138 ( \7852 , \3095 );
buf \U$7139 ( \7853 , \3223 );
not \U$7140 ( \7854 , \7853 );
buf \U$7141 ( \7855 , \4516 );
not \U$7142 ( \7856 , \7855 );
or \U$7143 ( \7857 , \7854 , \7856 );
buf \U$7144 ( \7858 , \5603 );
buf \U$7145 ( \7859 , \3459 );
nand \U$7146 ( \7860 , \7858 , \7859 );
buf \U$7147 ( \7861 , \7860 );
buf \U$7148 ( \7862 , \7861 );
nand \U$7149 ( \7863 , \7857 , \7862 );
buf \U$7150 ( \7864 , \7863 );
buf \U$7151 ( \7865 , \7864 );
nand \U$7152 ( \7866 , \7852 , \7865 );
buf \U$7153 ( \7867 , \7866 );
buf \U$7154 ( \7868 , \7867 );
nand \U$7155 ( \7869 , \7851 , \7868 );
buf \U$7156 ( \7870 , \7869 );
buf \U$7157 ( \7871 , \7870 );
nand \U$7158 ( \7872 , \7828 , \7871 );
buf \U$7159 ( \7873 , \7872 );
buf \U$7160 ( \7874 , \7873 );
buf \U$7161 ( \7875 , \7825 );
not \U$7162 ( \7876 , \7875 );
buf \U$7163 ( \7877 , \7740 );
nand \U$7164 ( \7878 , \7876 , \7877 );
buf \U$7165 ( \7879 , \7878 );
buf \U$7166 ( \7880 , \7879 );
nand \U$7167 ( \7881 , \7874 , \7880 );
buf \U$7168 ( \7882 , \7881 );
buf \U$7169 ( \7883 , \7882 );
not \U$7170 ( \7884 , \7883 );
or \U$7171 ( \7885 , \7703 , \7884 );
buf \U$7172 ( \7886 , \7695 );
buf \U$7173 ( \7887 , \7669 );
nand \U$7174 ( \7888 , \7886 , \7887 );
buf \U$7175 ( \7889 , \7888 );
buf \U$7176 ( \7890 , \7889 );
nand \U$7177 ( \7891 , \7885 , \7890 );
buf \U$7178 ( \7892 , \7891 );
not \U$7179 ( \7893 , \7892 );
xor \U$7180 ( \7894 , \7591 , \7616 );
xor \U$7181 ( \7895 , \7894 , \7642 );
buf \U$7182 ( \7896 , \7895 );
buf \U$7183 ( \7897 , \7896 );
not \U$7184 ( \7898 , \7897 );
buf \U$7185 ( \7899 , \7508 );
not \U$7186 ( \7900 , \7899 );
buf \U$7187 ( \7901 , \7526 );
not \U$7188 ( \7902 , \7901 );
or \U$7189 ( \7903 , \7900 , \7902 );
buf \U$7190 ( \7904 , \7526 );
buf \U$7191 ( \7905 , \7508 );
or \U$7192 ( \7906 , \7904 , \7905 );
nand \U$7193 ( \7907 , \7903 , \7906 );
buf \U$7194 ( \7908 , \7907 );
buf \U$7195 ( \7909 , \7908 );
not \U$7196 ( \7910 , \7909 );
buf \U$7197 ( \7911 , \7553 );
not \U$7198 ( \7912 , \7911 );
buf \U$7199 ( \7913 , \7912 );
buf \U$7200 ( \7914 , \7913 );
not \U$7201 ( \7915 , \7914 );
and \U$7202 ( \7916 , \7910 , \7915 );
buf \U$7203 ( \7917 , \7908 );
buf \U$7204 ( \7918 , \7913 );
and \U$7205 ( \7919 , \7917 , \7918 );
nor \U$7206 ( \7920 , \7916 , \7919 );
buf \U$7207 ( \7921 , \7920 );
buf \U$7208 ( \7922 , \7921 );
nand \U$7209 ( \7923 , \7898 , \7922 );
buf \U$7210 ( \7924 , \7923 );
not \U$7211 ( \7925 , \7924 );
or \U$7212 ( \7926 , \7893 , \7925 );
not \U$7213 ( \7927 , \7921 );
nand \U$7214 ( \7928 , \7927 , \7896 );
nand \U$7215 ( \7929 , \7926 , \7928 );
buf \U$7216 ( \7930 , \7929 );
xor \U$7217 ( \7931 , \7650 , \7930 );
buf \U$7218 ( \7932 , \6849 );
buf \U$7219 ( \7933 , \6876 );
xor \U$7220 ( \7934 , \7932 , \7933 );
buf \U$7221 ( \7935 , \6906 );
xnor \U$7222 ( \7936 , \7934 , \7935 );
buf \U$7223 ( \7937 , \7936 );
buf \U$7224 ( \7938 , \7937 );
not \U$7225 ( \7939 , \7938 );
buf \U$7226 ( \7940 , \7012 );
buf \U$7227 ( \7941 , \6958 );
xor \U$7228 ( \7942 , \7940 , \7941 );
buf \U$7229 ( \7943 , \7040 );
xor \U$7230 ( \7944 , \7942 , \7943 );
buf \U$7231 ( \7945 , \7944 );
buf \U$7232 ( \7946 , \7945 );
not \U$7233 ( \7947 , \7946 );
buf \U$7234 ( \7948 , \7947 );
buf \U$7235 ( \7949 , \7948 );
not \U$7236 ( \7950 , \7949 );
or \U$7237 ( \7951 , \7939 , \7950 );
buf \U$7238 ( \7952 , \7937 );
not \U$7239 ( \7953 , \7952 );
buf \U$7240 ( \7954 , \7953 );
buf \U$7241 ( \7955 , \7954 );
buf \U$7242 ( \7956 , \7945 );
nand \U$7243 ( \7957 , \7955 , \7956 );
buf \U$7244 ( \7958 , \7957 );
buf \U$7245 ( \7959 , \7958 );
nand \U$7246 ( \7960 , \7951 , \7959 );
buf \U$7247 ( \7961 , \7960 );
buf \U$7248 ( \7962 , \7961 );
buf \U$7249 ( \7963 , \5321 );
not \U$7250 ( \7964 , \7963 );
buf \U$7251 ( \7965 , \2273 );
not \U$7252 ( \7966 , \7965 );
or \U$7253 ( \7967 , \7964 , \7966 );
buf \U$7254 ( \7968 , \7800 );
buf \U$7255 ( \7969 , \1337 );
nand \U$7256 ( \7970 , \7968 , \7969 );
buf \U$7257 ( \7971 , \7970 );
buf \U$7258 ( \7972 , \7971 );
nand \U$7259 ( \7973 , \7967 , \7972 );
buf \U$7260 ( \7974 , \7973 );
buf \U$7261 ( \7975 , \7974 );
not \U$7262 ( \7976 , \7975 );
buf \U$7263 ( \7977 , \1478 );
not \U$7264 ( \7978 , \7977 );
or \U$7265 ( \7979 , \7976 , \7978 );
buf \U$7266 ( \7980 , \1485 );
buf \U$7267 ( \7981 , \6836 );
nand \U$7268 ( \7982 , \7980 , \7981 );
buf \U$7269 ( \7983 , \7982 );
buf \U$7270 ( \7984 , \7983 );
nand \U$7271 ( \7985 , \7979 , \7984 );
buf \U$7272 ( \7986 , \7985 );
buf \U$7273 ( \7987 , \7986 );
not \U$7274 ( \7988 , \7987 );
buf \U$7275 ( \7989 , \7988 );
buf \U$7276 ( \7990 , \7989 );
not \U$7277 ( \7991 , \7990 );
and \U$7278 ( \7992 , \4644 , RI9154c78_646);
and \U$7279 ( \7993 , \984 , RI91553f8_662);
nor \U$7280 ( \7994 , \7992 , \7993 );
and \U$7281 ( \7995 , \6052 , RI9155b78_678);
and \U$7282 ( \7996 , \5430 , RI91562f8_694);
nor \U$7283 ( \7997 , \7995 , \7996 );
and \U$7284 ( \7998 , \4003 , RI9156a78_710);
and \U$7285 ( \7999 , \1200 , RI91571f8_726);
nor \U$7286 ( \8000 , \7998 , \7999 );
and \U$7287 ( \8001 , \1014 , RI9157978_742);
and \U$7288 ( \8002 , \5439 , RI91580f8_758);
nor \U$7289 ( \8003 , \8001 , \8002 );
and \U$7290 ( \8004 , \7994 , \7997 , \8000 , \8003 );
not \U$7291 ( \8005 , \1285 );
and \U$7292 ( \8006 , RI91535f8_598, \8005 );
and \U$7293 ( \8007 , \7094 , RI9152e78_582);
not \U$7294 ( \8008 , RI91544f8_630);
not \U$7295 ( \8009 , \5453 );
or \U$7296 ( \8010 , \8008 , \8009 );
nand \U$7297 ( \8011 , \7099 , RI9153d78_614);
nand \U$7298 ( \8012 , \8010 , \8011 );
nor \U$7299 ( \8013 , \8006 , \8007 , \8012 );
and \U$7300 ( \8014 , \5463 , RI9151078_518);
and \U$7301 ( \8015 , \963 , RI91517f8_534);
nor \U$7302 ( \8016 , \8014 , \8015 );
and \U$7303 ( \8017 , \7106 , RI9151f78_550);
and \U$7304 ( \8018 , \1623 , RI91526f8_566);
nor \U$7305 ( \8019 , \8017 , \8018 );
and \U$7306 ( \8020 , \8013 , \8016 , \8019 );
nand \U$7307 ( \8021 , \8004 , \8020 );
buf \U$7308 ( \8022 , \8021 );
buf \U$7309 ( \8023 , \5321 );
not \U$7310 ( \8024 , \8023 );
buf \U$7311 ( \8025 , \1482 );
nor \U$7312 ( \8026 , \8024 , \8025 );
buf \U$7313 ( \8027 , \8026 );
buf \U$7314 ( \8028 , \8027 );
xor \U$7315 ( \8029 , \8022 , \8028 );
buf \U$7316 ( \8030 , \7121 );
not \U$7317 ( \8031 , \8030 );
buf \U$7318 ( \8032 , \7732 );
not \U$7319 ( \8033 , \8032 );
or \U$7320 ( \8034 , \8031 , \8033 );
buf \U$7321 ( \8035 , \7498 );
buf \U$7322 ( \8036 , \5398 );
nand \U$7323 ( \8037 , \8035 , \8036 );
buf \U$7324 ( \8038 , \8037 );
buf \U$7325 ( \8039 , \8038 );
nand \U$7326 ( \8040 , \8034 , \8039 );
buf \U$7327 ( \8041 , \8040 );
buf \U$7328 ( \8042 , \8041 );
and \U$7329 ( \8043 , \8029 , \8042 );
and \U$7330 ( \8044 , \8022 , \8028 );
or \U$7331 ( \8045 , \8043 , \8044 );
buf \U$7332 ( \8046 , \8045 );
buf \U$7333 ( \8047 , \8046 );
not \U$7334 ( \8048 , \8047 );
buf \U$7335 ( \8049 , \8048 );
buf \U$7336 ( \8050 , \8049 );
not \U$7337 ( \8051 , \8050 );
or \U$7338 ( \8052 , \7991 , \8051 );
buf \U$7339 ( \8053 , \7864 );
not \U$7340 ( \8054 , \8053 );
buf \U$7341 ( \8055 , \5143 );
not \U$7342 ( \8056 , \8055 );
or \U$7343 ( \8057 , \8054 , \8056 );
buf \U$7344 ( \8058 , \7541 );
buf \U$7345 ( \8059 , \3095 );
nand \U$7346 ( \8060 , \8058 , \8059 );
buf \U$7347 ( \8061 , \8060 );
buf \U$7348 ( \8062 , \8061 );
nand \U$7349 ( \8063 , \8057 , \8062 );
buf \U$7350 ( \8064 , \8063 );
not \U$7351 ( \8065 , \8064 );
buf \U$7352 ( \8066 , \7812 );
buf \U$7353 ( \8067 , \7774 );
nand \U$7354 ( \8068 , \8066 , \8067 );
buf \U$7355 ( \8069 , \8068 );
buf \U$7356 ( \8070 , \8069 );
not \U$7357 ( \8071 , \8070 );
buf \U$7358 ( \8072 , \8071 );
not \U$7359 ( \8073 , \8072 );
or \U$7360 ( \8074 , \8065 , \8073 );
not \U$7361 ( \8075 , \8069 );
buf \U$7362 ( \8076 , \8064 );
not \U$7363 ( \8077 , \8076 );
buf \U$7364 ( \8078 , \8077 );
not \U$7365 ( \8079 , \8078 );
or \U$7366 ( \8080 , \8075 , \8079 );
buf \U$7367 ( \8081 , \4032 );
not \U$7368 ( \8082 , \8081 );
buf \U$7369 ( \8083 , \2479 );
not \U$7370 ( \8084 , \8083 );
or \U$7371 ( \8085 , \8082 , \8084 );
buf \U$7372 ( \8086 , \2627 );
not \U$7373 ( \8087 , \8086 );
buf \U$7374 ( \8088 , \8087 );
buf \U$7375 ( \8089 , \8088 );
buf \U$7376 ( \8090 , \4029 );
nand \U$7377 ( \8091 , \8089 , \8090 );
buf \U$7378 ( \8092 , \8091 );
buf \U$7379 ( \8093 , \8092 );
nand \U$7380 ( \8094 , \8085 , \8093 );
buf \U$7381 ( \8095 , \8094 );
buf \U$7382 ( \8096 , \8095 );
not \U$7383 ( \8097 , \8096 );
buf \U$7384 ( \8098 , \2983 );
not \U$7385 ( \8099 , \8098 );
or \U$7386 ( \8100 , \8097 , \8099 );
buf \U$7387 ( \8101 , \2473 );
buf \U$7388 ( \8102 , \7578 );
nand \U$7389 ( \8103 , \8101 , \8102 );
buf \U$7390 ( \8104 , \8103 );
buf \U$7391 ( \8105 , \8104 );
nand \U$7392 ( \8106 , \8100 , \8105 );
buf \U$7393 ( \8107 , \8106 );
nand \U$7394 ( \8108 , \8080 , \8107 );
nand \U$7395 ( \8109 , \8074 , \8108 );
buf \U$7396 ( \8110 , \8109 );
nand \U$7397 ( \8111 , \8052 , \8110 );
buf \U$7398 ( \8112 , \8111 );
buf \U$7399 ( \8113 , \8112 );
buf \U$7400 ( \8114 , \8046 );
buf \U$7401 ( \8115 , \7986 );
nand \U$7402 ( \8116 , \8114 , \8115 );
buf \U$7403 ( \8117 , \8116 );
buf \U$7404 ( \8118 , \8117 );
nand \U$7405 ( \8119 , \8113 , \8118 );
buf \U$7406 ( \8120 , \8119 );
buf \U$7409 ( \8121 , \8120 );
buf \U$7410 ( \8122 , \8121 );
and \U$7411 ( \8123 , \7962 , \8122 );
not \U$7412 ( \8124 , \7962 );
buf \U$7413 ( \8125 , \8121 );
not \U$7414 ( \8126 , \8125 );
buf \U$7415 ( \8127 , \8126 );
buf \U$7416 ( \8128 , \8127 );
and \U$7417 ( \8129 , \8124 , \8128 );
nor \U$7418 ( \8130 , \8123 , \8129 );
buf \U$7419 ( \8131 , \8130 );
buf \U$7420 ( \8132 , \8131 );
xor \U$7421 ( \8133 , \7931 , \8132 );
buf \U$7422 ( \8134 , \8133 );
buf \U$7423 ( \8135 , \8134 );
xor \U$7424 ( \8136 , \7989 , \8046 );
xor \U$7425 ( \8137 , \8136 , \8109 );
buf \U$7426 ( \8138 , \8137 );
not \U$7427 ( \8139 , \8138 );
buf \U$7428 ( \8140 , \8139 );
buf \U$7429 ( \8141 , \8140 );
not \U$7430 ( \8142 , \8141 );
buf \U$7431 ( \8143 , \7896 );
not \U$7432 ( \8144 , \8143 );
buf \U$7433 ( \8145 , \7921 );
not \U$7434 ( \8146 , \8145 );
or \U$7435 ( \8147 , \8144 , \8146 );
buf \U$7436 ( \8148 , \7896 );
buf \U$7437 ( \8149 , \7921 );
or \U$7438 ( \8150 , \8148 , \8149 );
nand \U$7439 ( \8151 , \8147 , \8150 );
buf \U$7440 ( \8152 , \8151 );
buf \U$7441 ( \8153 , \8152 );
buf \U$7442 ( \8154 , \7892 );
not \U$7443 ( \8155 , \8154 );
buf \U$7444 ( \8156 , \8155 );
buf \U$7445 ( \8157 , \8156 );
and \U$7446 ( \8158 , \8153 , \8157 );
not \U$7447 ( \8159 , \8153 );
buf \U$7448 ( \8160 , \7892 );
and \U$7449 ( \8161 , \8159 , \8160 );
nor \U$7450 ( \8162 , \8158 , \8161 );
buf \U$7451 ( \8163 , \8162 );
buf \U$7452 ( \8164 , \8163 );
not \U$7453 ( \8165 , \8164 );
buf \U$7454 ( \8166 , \8165 );
buf \U$7455 ( \8167 , \8166 );
not \U$7456 ( \8168 , \8167 );
or \U$7457 ( \8169 , \8142 , \8168 );
buf \U$7458 ( \8170 , \8137 );
not \U$7459 ( \8171 , \8170 );
buf \U$7460 ( \8172 , \8163 );
not \U$7461 ( \8173 , \8172 );
or \U$7462 ( \8174 , \8171 , \8173 );
xor \U$7463 ( \8175 , \8022 , \8028 );
xor \U$7464 ( \8176 , \8175 , \8042 );
buf \U$7465 ( \8177 , \8176 );
buf \U$7466 ( \8178 , \8177 );
not \U$7467 ( \8179 , \8178 );
buf \U$7468 ( \8180 , \8072 );
not \U$7469 ( \8181 , \8180 );
buf \U$7470 ( \8182 , \8078 );
not \U$7471 ( \8183 , \8182 );
or \U$7472 ( \8184 , \8181 , \8183 );
buf \U$7473 ( \8185 , \8064 );
buf \U$7474 ( \8186 , \8069 );
nand \U$7475 ( \8187 , \8185 , \8186 );
buf \U$7476 ( \8188 , \8187 );
buf \U$7477 ( \8189 , \8188 );
nand \U$7478 ( \8190 , \8184 , \8189 );
buf \U$7479 ( \8191 , \8190 );
buf \U$7480 ( \8192 , \8191 );
buf \U$7481 ( \8193 , \8107 );
not \U$7482 ( \8194 , \8193 );
buf \U$7483 ( \8195 , \8194 );
buf \U$7484 ( \8196 , \8195 );
and \U$7485 ( \8197 , \8192 , \8196 );
not \U$7486 ( \8198 , \8192 );
buf \U$7487 ( \8199 , \8107 );
and \U$7488 ( \8200 , \8198 , \8199 );
nor \U$7489 ( \8201 , \8197 , \8200 );
buf \U$7490 ( \8202 , \8201 );
buf \U$7491 ( \8203 , \8202 );
not \U$7492 ( \8204 , \8203 );
buf \U$7493 ( \8205 , \8204 );
buf \U$7494 ( \8206 , \8205 );
not \U$7495 ( \8207 , \8206 );
or \U$7496 ( \8208 , \8179 , \8207 );
buf \U$7497 ( \8209 , \8202 );
buf \U$7498 ( \8210 , \8177 );
not \U$7499 ( \8211 , \8210 );
buf \U$7500 ( \8212 , \8211 );
buf \U$7501 ( \8213 , \8212 );
nand \U$7502 ( \8214 , \8209 , \8213 );
buf \U$7503 ( \8215 , \8214 );
buf \U$7504 ( \8216 , \8215 );
buf \U$7505 ( \8217 , \8095 );
not \U$7506 ( \8218 , \8217 );
buf \U$7507 ( \8219 , \8218 );
buf \U$7508 ( \8220 , \8219 );
buf \U$7509 ( \8221 , \2476 );
or \U$7510 ( \8222 , \8220 , \8221 );
buf \U$7511 ( \8223 , \2425 );
buf \U$7512 ( \8224 , \2476 );
buf \U$7513 ( \8225 , \4855 );
not \U$7514 ( \8226 , \8225 );
buf \U$7515 ( \8227 , \2627 );
not \U$7516 ( \8228 , \8227 );
or \U$7517 ( \8229 , \8226 , \8228 );
buf \U$7518 ( \8230 , \3276 );
buf \U$7519 ( \8231 , \4863 );
nand \U$7520 ( \8232 , \8230 , \8231 );
buf \U$7521 ( \8233 , \8232 );
buf \U$7522 ( \8234 , \8233 );
nand \U$7523 ( \8235 , \8229 , \8234 );
buf \U$7524 ( \8236 , \8235 );
buf \U$7525 ( \8237 , \8236 );
nand \U$7526 ( \8238 , \8223 , \8224 , \8237 );
buf \U$7527 ( \8239 , \8238 );
buf \U$7528 ( \8240 , \8239 );
nand \U$7529 ( \8241 , \8222 , \8240 );
buf \U$7530 ( \8242 , \8241 );
buf \U$7531 ( \8243 , \8242 );
not \U$7532 ( \8244 , \8243 );
buf \U$7533 ( \8245 , \2068 );
buf \U$7534 ( \8246 , \7800 );
nand \U$7535 ( \8247 , \8245 , \8246 );
buf \U$7536 ( \8248 , \8247 );
buf \U$7537 ( \8249 , \8248 );
buf \U$7538 ( \8250 , \2884 );
not \U$7539 ( \8251 , \8250 );
buf \U$7540 ( \8252 , \5321 );
nand \U$7541 ( \8253 , \8251 , \8252 );
buf \U$7542 ( \8254 , \8253 );
buf \U$7543 ( \8255 , \8254 );
and \U$7544 ( \8256 , \8249 , \8255 );
buf \U$7545 ( \8257 , \4127 );
nor \U$7546 ( \8258 , \8256 , \8257 );
buf \U$7547 ( \8259 , \8258 );
buf \U$7548 ( \8260 , \8259 );
not \U$7549 ( \8261 , \8260 );
buf \U$7550 ( \8262 , \4814 );
not \U$7551 ( \8263 , \8262 );
or \U$7552 ( \8264 , \8261 , \8263 );
buf \U$7553 ( \8265 , \2897 );
buf \U$7554 ( \8266 , \7683 );
nand \U$7555 ( \8267 , \8265 , \8266 );
buf \U$7556 ( \8268 , \8267 );
buf \U$7557 ( \8269 , \8268 );
nand \U$7558 ( \8270 , \8264 , \8269 );
buf \U$7559 ( \8271 , \8270 );
buf \U$7560 ( \8272 , \8271 );
not \U$7561 ( \8273 , \8272 );
or \U$7562 ( \8274 , \8244 , \8273 );
buf \U$7563 ( \8275 , \8242 );
not \U$7564 ( \8276 , \8275 );
buf \U$7565 ( \8277 , \8276 );
buf \U$7566 ( \8278 , \8277 );
not \U$7567 ( \8279 , \8278 );
buf \U$7568 ( \8280 , \8271 );
not \U$7569 ( \8281 , \8280 );
buf \U$7570 ( \8282 , \8281 );
buf \U$7571 ( \8283 , \8282 );
not \U$7572 ( \8284 , \8283 );
or \U$7573 ( \8285 , \8279 , \8284 );
buf \U$7574 ( \8286 , \2758 );
not \U$7575 ( \8287 , \8286 );
buf \U$7576 ( \8288 , \4550 );
not \U$7577 ( \8289 , \8288 );
or \U$7578 ( \8290 , \8287 , \8289 );
buf \U$7579 ( \8291 , \2853 );
buf \U$7580 ( \8292 , \4278 );
nand \U$7581 ( \8293 , \8291 , \8292 );
buf \U$7582 ( \8294 , \8293 );
buf \U$7583 ( \8295 , \8294 );
nand \U$7584 ( \8296 , \8290 , \8295 );
buf \U$7585 ( \8297 , \8296 );
buf \U$7586 ( \8298 , \8297 );
not \U$7587 ( \8299 , \8298 );
buf \U$7588 ( \8300 , \4543 );
not \U$7589 ( \8301 , \8300 );
or \U$7590 ( \8302 , \8299 , \8301 );
buf \U$7591 ( \8303 , \7654 );
buf \U$7592 ( \8304 , \4581 );
nand \U$7593 ( \8305 , \8303 , \8304 );
buf \U$7594 ( \8306 , \8305 );
buf \U$7595 ( \8307 , \8306 );
nand \U$7596 ( \8308 , \8302 , \8307 );
buf \U$7597 ( \8309 , \8308 );
buf \U$7598 ( \8310 , \8309 );
nand \U$7599 ( \8311 , \8285 , \8310 );
buf \U$7600 ( \8312 , \8311 );
buf \U$7601 ( \8313 , \8312 );
nand \U$7602 ( \8314 , \8274 , \8313 );
buf \U$7603 ( \8315 , \8314 );
buf \U$7604 ( \8316 , \8315 );
nand \U$7605 ( \8317 , \8216 , \8316 );
buf \U$7606 ( \8318 , \8317 );
buf \U$7607 ( \8319 , \8318 );
nand \U$7608 ( \8320 , \8208 , \8319 );
buf \U$7609 ( \8321 , \8320 );
buf \U$7610 ( \8322 , \8321 );
nand \U$7611 ( \8323 , \8174 , \8322 );
buf \U$7612 ( \8324 , \8323 );
buf \U$7613 ( \8325 , \8324 );
nand \U$7614 ( \8326 , \8169 , \8325 );
buf \U$7615 ( \8327 , \8326 );
buf \U$7616 ( \8328 , \8327 );
nor \U$7617 ( \8329 , \8135 , \8328 );
buf \U$7618 ( \8330 , \8329 );
buf \U$7619 ( \8331 , \8330 );
buf \U$7620 ( \8332 , \7954 );
not \U$7621 ( \8333 , \8332 );
buf \U$7622 ( \8334 , \7948 );
not \U$7623 ( \8335 , \8334 );
or \U$7624 ( \8336 , \8333 , \8335 );
buf \U$7625 ( \8337 , \7945 );
not \U$7626 ( \8338 , \8337 );
buf \U$7627 ( \8339 , \7937 );
not \U$7628 ( \8340 , \8339 );
or \U$7629 ( \8341 , \8338 , \8340 );
buf \U$7630 ( \8342 , \8120 );
nand \U$7631 ( \8343 , \8341 , \8342 );
buf \U$7632 ( \8344 , \8343 );
buf \U$7633 ( \8345 , \8344 );
nand \U$7634 ( \8346 , \8336 , \8345 );
buf \U$7635 ( \8347 , \8346 );
buf \U$7636 ( \8348 , \8347 );
not \U$7637 ( \8349 , \8348 );
buf \U$7638 ( \8350 , \7150 );
buf \U$7639 ( \8351 , \7078 );
xor \U$7640 ( \8352 , \8350 , \8351 );
buf \U$7641 ( \8353 , \7050 );
xnor \U$7642 ( \8354 , \8352 , \8353 );
buf \U$7643 ( \8355 , \8354 );
buf \U$7644 ( \8356 , \8355 );
not \U$7645 ( \8357 , \8356 );
and \U$7646 ( \8358 , \8349 , \8357 );
buf \U$7649 ( \8359 , \8355 );
buf \U$7650 ( \8360 , \8359 );
buf \U$7651 ( \8361 , \8347 );
and \U$7652 ( \8362 , \8360 , \8361 );
nor \U$7653 ( \8363 , \8358 , \8362 );
buf \U$7654 ( \8364 , \8363 );
buf \U$7655 ( \8365 , \8364 );
not \U$7656 ( \8366 , \8365 );
not \U$7657 ( \8367 , \6528 );
not \U$7658 ( \8368 , \6560 );
or \U$7659 ( \8369 , \8367 , \8368 );
buf \U$7660 ( \8370 , \6531 );
buf \U$7661 ( \8371 , \6557 );
nand \U$7662 ( \8372 , \8370 , \8371 );
buf \U$7663 ( \8373 , \8372 );
nand \U$7664 ( \8374 , \8369 , \8373 );
xor \U$7665 ( \8375 , \8374 , \6589 );
buf \U$7666 ( \8376 , \8375 );
buf \U$7667 ( \8377 , \6819 );
buf \U$7668 ( \8378 , \6790 );
xor \U$7669 ( \8379 , \8377 , \8378 );
buf \U$7670 ( \8380 , \8379 );
buf \U$7671 ( \8381 , \8380 );
not \U$7672 ( \8382 , \8381 );
buf \U$7673 ( \8383 , \6912 );
not \U$7674 ( \8384 , \8383 );
or \U$7675 ( \8385 , \8382 , \8384 );
buf \U$7676 ( \8386 , \8380 );
buf \U$7677 ( \8387 , \6912 );
or \U$7678 ( \8388 , \8386 , \8387 );
nand \U$7679 ( \8389 , \8385 , \8388 );
buf \U$7680 ( \8390 , \8389 );
buf \U$7681 ( \8391 , \8390 );
xor \U$7682 ( \8392 , \8376 , \8391 );
xor \U$7683 ( \8393 , \7484 , \7565 );
and \U$7684 ( \8394 , \8393 , \7647 );
and \U$7685 ( \8395 , \7484 , \7565 );
or \U$7686 ( \8396 , \8394 , \8395 );
buf \U$7687 ( \8397 , \8396 );
buf \U$7688 ( \8398 , \8397 );
xor \U$7689 ( \8399 , \8392 , \8398 );
buf \U$7690 ( \8400 , \8399 );
buf \U$7691 ( \8401 , \8400 );
not \U$7692 ( \8402 , \8401 );
or \U$7693 ( \8403 , \8366 , \8402 );
buf \U$7694 ( \8404 , \8400 );
buf \U$7695 ( \8405 , \8364 );
or \U$7696 ( \8406 , \8404 , \8405 );
nand \U$7697 ( \8407 , \8403 , \8406 );
buf \U$7698 ( \8408 , \8407 );
buf \U$7699 ( \8409 , \8408 );
xor \U$7700 ( \8410 , \7650 , \7930 );
and \U$7701 ( \8411 , \8410 , \8132 );
and \U$7702 ( \8412 , \7650 , \7930 );
or \U$7703 ( \8413 , \8411 , \8412 );
buf \U$7704 ( \8414 , \8413 );
buf \U$7705 ( \8415 , \8414 );
nor \U$7706 ( \8416 , \8409 , \8415 );
buf \U$7707 ( \8417 , \8416 );
buf \U$7708 ( \8418 , \8417 );
nor \U$7709 ( \8419 , \8331 , \8418 );
buf \U$7710 ( \8420 , \8419 );
buf \U$7711 ( \8421 , \8420 );
buf \U$7712 ( \8422 , \7249 );
not \U$7713 ( \8423 , \8422 );
buf \U$7714 ( \8424 , \7188 );
not \U$7715 ( \8425 , \8424 );
or \U$7716 ( \8426 , \8423 , \8425 );
buf \U$7717 ( \8427 , \7185 );
buf \U$7718 ( \8428 , \7215 );
nand \U$7719 ( \8429 , \8427 , \8428 );
buf \U$7720 ( \8430 , \8429 );
buf \U$7721 ( \8431 , \8430 );
nand \U$7722 ( \8432 , \8426 , \8431 );
buf \U$7723 ( \8433 , \8432 );
buf \U$7724 ( \8434 , \8433 );
buf \U$7725 ( \8435 , \7241 );
not \U$7726 ( \8436 , \8435 );
buf \U$7727 ( \8437 , \8436 );
buf \U$7728 ( \8438 , \8437 );
and \U$7729 ( \8439 , \8434 , \8438 );
not \U$7730 ( \8440 , \8434 );
buf \U$7731 ( \8441 , \7241 );
and \U$7732 ( \8442 , \8440 , \8441 );
nor \U$7733 ( \8443 , \8439 , \8442 );
buf \U$7734 ( \8444 , \8443 );
buf \U$7735 ( \8445 , \8444 );
buf \U$7736 ( \8446 , \7170 );
buf \U$7737 ( \8447 , \6922 );
and \U$7738 ( \8448 , \8446 , \8447 );
not \U$7739 ( \8449 , \8446 );
buf \U$7740 ( \8450 , \6925 );
and \U$7741 ( \8451 , \8449 , \8450 );
nor \U$7742 ( \8452 , \8448 , \8451 );
buf \U$7743 ( \8453 , \8452 );
buf \U$7744 ( \8454 , \8453 );
buf \U$7745 ( \8455 , \6939 );
and \U$7746 ( \8456 , \8454 , \8455 );
not \U$7747 ( \8457 , \8454 );
buf \U$7748 ( \8458 , \7179 );
and \U$7749 ( \8459 , \8457 , \8458 );
nor \U$7750 ( \8460 , \8456 , \8459 );
buf \U$7751 ( \8461 , \8460 );
buf \U$7752 ( \8462 , \8461 );
not \U$7753 ( \8463 , \8462 );
buf \U$7754 ( \8464 , \8463 );
not \U$7755 ( \8465 , \8464 );
buf \U$7756 ( \8466 , \6716 );
buf \U$7757 ( \8467 , \6642 );
xor \U$7758 ( \8468 , \8466 , \8467 );
buf \U$7759 ( \8469 , \6727 );
xnor \U$7760 ( \8470 , \8468 , \8469 );
buf \U$7761 ( \8471 , \8470 );
buf \U$7762 ( \8472 , \8471 );
not \U$7763 ( \8473 , \8472 );
buf \U$7764 ( \8474 , \8473 );
not \U$7765 ( \8475 , \8474 );
or \U$7766 ( \8476 , \8465 , \8475 );
not \U$7767 ( \8477 , \8471 );
not \U$7768 ( \8478 , \8461 );
or \U$7769 ( \8479 , \8477 , \8478 );
xor \U$7770 ( \8480 , \8376 , \8391 );
and \U$7771 ( \8481 , \8480 , \8398 );
and \U$7772 ( \8482 , \8376 , \8391 );
or \U$7773 ( \8483 , \8481 , \8482 );
buf \U$7774 ( \8484 , \8483 );
nand \U$7775 ( \8485 , \8479 , \8484 );
nand \U$7776 ( \8486 , \8476 , \8485 );
buf \U$7777 ( \8487 , \8486 );
not \U$7778 ( \8488 , \8487 );
buf \U$7779 ( \8489 , \8488 );
buf \U$7780 ( \8490 , \8489 );
nand \U$7781 ( \8491 , \8445 , \8490 );
buf \U$7782 ( \8492 , \8491 );
buf \U$7783 ( \8493 , \8492 );
buf \U$7784 ( \8494 , \8474 );
not \U$7785 ( \8495 , \8494 );
buf \U$7786 ( \8496 , \8484 );
not \U$7787 ( \8497 , \8496 );
buf \U$7788 ( \8498 , \8497 );
buf \U$7789 ( \8499 , \8498 );
not \U$7790 ( \8500 , \8499 );
or \U$7791 ( \8501 , \8495 , \8500 );
buf \U$7792 ( \8502 , \8484 );
buf \U$7793 ( \8503 , \8471 );
nand \U$7794 ( \8504 , \8502 , \8503 );
buf \U$7795 ( \8505 , \8504 );
buf \U$7796 ( \8506 , \8505 );
nand \U$7797 ( \8507 , \8501 , \8506 );
buf \U$7798 ( \8508 , \8507 );
buf \U$7799 ( \8509 , \8508 );
buf \U$7800 ( \8510 , \8461 );
and \U$7801 ( \8511 , \8509 , \8510 );
not \U$7802 ( \8512 , \8509 );
buf \U$7803 ( \8513 , \8464 );
and \U$7804 ( \8514 , \8512 , \8513 );
nor \U$7805 ( \8515 , \8511 , \8514 );
buf \U$7806 ( \8516 , \8515 );
buf \U$7807 ( \8517 , \8516 );
buf \U$7808 ( \8518 , \8400 );
not \U$7809 ( \8519 , \8518 );
buf \U$7810 ( \8520 , \8347 );
not \U$7811 ( \8521 , \8520 );
buf \U$7812 ( \8522 , \8359 );
nand \U$7813 ( \8523 , \8521 , \8522 );
buf \U$7814 ( \8524 , \8523 );
buf \U$7815 ( \8525 , \8524 );
not \U$7816 ( \8526 , \8525 );
or \U$7817 ( \8527 , \8519 , \8526 );
buf \U$7818 ( \8528 , \8359 );
not \U$7819 ( \8529 , \8528 );
buf \U$7820 ( \8530 , \8347 );
nand \U$7821 ( \8531 , \8529 , \8530 );
buf \U$7822 ( \8532 , \8531 );
buf \U$7823 ( \8533 , \8532 );
nand \U$7824 ( \8534 , \8527 , \8533 );
buf \U$7825 ( \8535 , \8534 );
buf \U$7826 ( \8536 , \8535 );
not \U$7827 ( \8537 , \8536 );
buf \U$7828 ( \8538 , \8537 );
buf \U$7829 ( \8539 , \8538 );
nand \U$7830 ( \8540 , \8517 , \8539 );
buf \U$7831 ( \8541 , \8540 );
buf \U$7832 ( \8542 , \8541 );
nand \U$7833 ( \8543 , \8421 , \8493 , \8542 );
buf \U$7834 ( \8544 , \8543 );
buf \U$7835 ( \8545 , \8544 );
not \U$7836 ( \8546 , \8545 );
buf \U$7837 ( \8547 , \8546 );
buf \U$7838 ( \8548 , \8547 );
not \U$7839 ( \8549 , \8548 );
buf \U$7840 ( \8550 , \8321 );
not \U$7841 ( \8551 , \8550 );
buf \U$7842 ( \8552 , \8137 );
not \U$7843 ( \8553 , \8552 );
and \U$7844 ( \8554 , \8551 , \8553 );
buf \U$7845 ( \8555 , \8321 );
buf \U$7846 ( \8556 , \8137 );
and \U$7847 ( \8557 , \8555 , \8556 );
nor \U$7848 ( \8558 , \8554 , \8557 );
buf \U$7849 ( \8559 , \8558 );
buf \U$7850 ( \8560 , \8559 );
buf \U$7851 ( \8561 , \8166 );
and \U$7852 ( \8562 , \8560 , \8561 );
not \U$7853 ( \8563 , \8560 );
buf \U$7854 ( \8564 , \8163 );
and \U$7855 ( \8565 , \8563 , \8564 );
nor \U$7856 ( \8566 , \8562 , \8565 );
buf \U$7857 ( \8567 , \8566 );
buf \U$7858 ( \8568 , \8567 );
xor \U$7859 ( \8569 , \7698 , \7669 );
xor \U$7860 ( \8570 , \8569 , \7882 );
buf \U$7861 ( \8571 , \8570 );
and \U$7862 ( \8572 , \4644 , RI9154d68_648);
not \U$7863 ( \8573 , \983 );
and \U$7864 ( \8574 , \8573 , RI91554e8_664);
nor \U$7865 ( \8575 , \8572 , \8574 );
and \U$7866 ( \8576 , \5434 , RI9156b68_712);
and \U$7867 ( \8577 , \1200 , RI91572e8_728);
nor \U$7868 ( \8578 , \8576 , \8577 );
and \U$7869 ( \8579 , \8575 , \8578 );
and \U$7870 ( \8580 , \7094 , RI9152f68_584);
and \U$7871 ( \8581 , \1500 , RI91536e8_600);
nor \U$7872 ( \8582 , \8580 , \8581 );
and \U$7873 ( \8583 , \5451 , RI9153e68_616);
and \U$7874 ( \8584 , \5453 , RI91545e8_632);
nor \U$7875 ( \8585 , \8583 , \8584 );
and \U$7876 ( \8586 , \8582 , \8585 );
and \U$7877 ( \8587 , \5463 , RI9151168_520);
and \U$7878 ( \8588 , \963 , RI91518e8_536);
nor \U$7879 ( \8589 , \8587 , \8588 );
and \U$7880 ( \8590 , \7106 , RI9152068_552);
and \U$7881 ( \8591 , \1623 , RI91527e8_568);
nor \U$7882 ( \8592 , \8590 , \8591 );
and \U$7883 ( \8593 , \8589 , \8592 );
and \U$7884 ( \8594 , \5428 , RI9155c68_680);
and \U$7885 ( \8595 , \5430 , RI91563e8_696);
nor \U$7886 ( \8596 , \8594 , \8595 );
and \U$7887 ( \8597 , \1014 , RI9157a68_744);
and \U$7888 ( \8598 , \4011 , RI91581e8_760);
nor \U$7889 ( \8599 , \8597 , \8598 );
and \U$7890 ( \8600 , \8596 , \8599 );
nand \U$7891 ( \8601 , \8579 , \8586 , \8593 , \8600 );
buf \U$7892 ( \8602 , \8601 );
buf \U$7893 ( \8603 , \2211 );
buf \U$7894 ( \8604 , \7800 );
nor \U$7895 ( \8605 , \8603 , \8604 );
buf \U$7896 ( \8606 , \8605 );
buf \U$7897 ( \8607 , \8606 );
xor \U$7898 ( \8608 , \8602 , \8607 );
buf \U$7899 ( \8609 , \5391 );
not \U$7900 ( \8610 , \8609 );
and \U$7901 ( \8611 , \1669 , \4795 );
not \U$7902 ( \8612 , \1669 );
and \U$7903 ( \8613 , \8612 , \4794 );
or \U$7904 ( \8614 , \8611 , \8613 );
buf \U$7905 ( \8615 , \8614 );
not \U$7906 ( \8616 , \8615 );
or \U$7907 ( \8617 , \8610 , \8616 );
buf \U$7908 ( \8618 , \7715 );
buf \U$7909 ( \8619 , \5398 );
nand \U$7910 ( \8620 , \8618 , \8619 );
buf \U$7911 ( \8621 , \8620 );
buf \U$7912 ( \8622 , \8621 );
nand \U$7913 ( \8623 , \8617 , \8622 );
buf \U$7914 ( \8624 , \8623 );
buf \U$7915 ( \8625 , \8624 );
and \U$7916 ( \8626 , \8608 , \8625 );
and \U$7917 ( \8627 , \8602 , \8607 );
or \U$7918 ( \8628 , \8626 , \8627 );
buf \U$7919 ( \8629 , \8628 );
buf \U$7920 ( \8630 , \8629 );
not \U$7921 ( \8631 , \8630 );
buf \U$7922 ( \8632 , \7739 );
buf \U$7923 ( \8633 , \7822 );
xor \U$7924 ( \8634 , \8632 , \8633 );
buf \U$7925 ( \8635 , \7870 );
xnor \U$7926 ( \8636 , \8634 , \8635 );
buf \U$7927 ( \8637 , \8636 );
buf \U$7928 ( \8638 , \8637 );
nand \U$7929 ( \8639 , \8631 , \8638 );
buf \U$7930 ( \8640 , \8639 );
buf \U$7931 ( \8641 , \8640 );
and \U$7932 ( \8642 , RI9152fe0_585, \7094 );
and \U$7933 ( \8643 , \8005 , RI9153760_601);
not \U$7934 ( \8644 , RI9154660_633);
not \U$7935 ( \8645 , \5453 );
or \U$7936 ( \8646 , \8644 , \8645 );
nand \U$7937 ( \8647 , \7099 , RI9153ee0_617);
nand \U$7938 ( \8648 , \8646 , \8647 );
nor \U$7939 ( \8649 , \8642 , \8643 , \8648 );
and \U$7940 ( \8650 , \5463 , RI91511e0_521);
and \U$7941 ( \8651 , \963 , RI9151960_537);
nor \U$7942 ( \8652 , \8650 , \8651 );
and \U$7943 ( \8653 , \7106 , RI91520e0_553);
and \U$7944 ( \8654 , \1623 , RI9152860_569);
nor \U$7945 ( \8655 , \8653 , \8654 );
and \U$7946 ( \8656 , \4644 , RI9154de0_649);
and \U$7947 ( \8657 , \984 , RI9155560_665);
nor \U$7948 ( \8658 , \8656 , \8657 );
and \U$7949 ( \8659 , \6052 , RI9155ce0_681);
and \U$7950 ( \8660 , \5430 , RI9156460_697);
nor \U$7951 ( \8661 , \8659 , \8660 );
and \U$7952 ( \8662 , \4003 , RI9156be0_713);
and \U$7953 ( \8663 , \2052 , RI9157360_729);
nor \U$7954 ( \8664 , \8662 , \8663 );
and \U$7955 ( \8665 , \1014 , RI9157ae0_745);
and \U$7956 ( \8666 , \5439 , RI9158260_761);
nor \U$7957 ( \8667 , \8665 , \8666 );
and \U$7958 ( \8668 , \8658 , \8661 , \8664 , \8667 );
nand \U$7959 ( \8669 , \8649 , \8652 , \8655 , \8668 );
not \U$7960 ( \8670 , \8669 );
buf \U$7961 ( \8671 , \2407 );
not \U$7962 ( \8672 , \8671 );
buf \U$7963 ( \8673 , \8672 );
buf \U$7964 ( \8674 , \8673 );
not \U$7965 ( \8675 , \8674 );
buf \U$7966 ( \8676 , \8675 );
buf \U$7967 ( \8677 , \8676 );
not \U$7968 ( \8678 , \8677 );
buf \U$7969 ( \8679 , \5573 );
not \U$7970 ( \8680 , \8679 );
or \U$7971 ( \8681 , \8678 , \8680 );
buf \U$7972 ( \8682 , \4100 );
nand \U$7973 ( \8683 , \8681 , \8682 );
buf \U$7974 ( \8684 , \8683 );
buf \U$7975 ( \8685 , \8684 );
buf \U$7976 ( \8686 , \5472 );
buf \U$7977 ( \8687 , \8673 );
nand \U$7978 ( \8688 , \8686 , \8687 );
buf \U$7979 ( \8689 , \8688 );
buf \U$7980 ( \8690 , \8689 );
buf \U$7981 ( \8691 , \2633 );
and \U$7982 ( \8692 , \8690 , \8691 );
buf \U$7983 ( \8693 , \8692 );
buf \U$7984 ( \8694 , \8693 );
nand \U$7985 ( \8695 , \8685 , \8694 );
buf \U$7986 ( \8696 , \8695 );
nor \U$7987 ( \8697 , \8670 , \8696 );
buf \U$7988 ( \8698 , \8697 );
not \U$7989 ( \8699 , \8698 );
buf \U$7990 ( \8700 , \4032 );
not \U$7991 ( \8701 , \8700 );
buf \U$7992 ( \8702 , \7833 );
not \U$7993 ( \8703 , \8702 );
or \U$7994 ( \8704 , \8701 , \8703 );
buf \U$7995 ( \8705 , \7839 );
buf \U$7996 ( \8706 , \5243 );
nand \U$7997 ( \8707 , \8705 , \8706 );
buf \U$7998 ( \8708 , \8707 );
buf \U$7999 ( \8709 , \8708 );
nand \U$8000 ( \8710 , \8704 , \8709 );
buf \U$8001 ( \8711 , \8710 );
buf \U$8002 ( \8712 , \8711 );
not \U$8003 ( \8713 , \8712 );
buf \U$8004 ( \8714 , \5615 );
not \U$8005 ( \8715 , \8714 );
or \U$8006 ( \8716 , \8713 , \8715 );
buf \U$8007 ( \8717 , \3095 );
buf \U$8008 ( \8718 , \7846 );
nand \U$8009 ( \8719 , \8717 , \8718 );
buf \U$8010 ( \8720 , \8719 );
buf \U$8011 ( \8721 , \8720 );
nand \U$8012 ( \8722 , \8716 , \8721 );
buf \U$8013 ( \8723 , \8722 );
buf \U$8014 ( \8724 , \8723 );
not \U$8015 ( \8725 , \8724 );
or \U$8016 ( \8726 , \8699 , \8725 );
buf \U$8017 ( \8727 , \8723 );
buf \U$8018 ( \8728 , \8697 );
or \U$8019 ( \8729 , \8727 , \8728 );
buf \U$8020 ( \8730 , \4848 );
not \U$8021 ( \8731 , \8730 );
buf \U$8022 ( \8732 , \2479 );
not \U$8023 ( \8733 , \8732 );
or \U$8024 ( \8734 , \8731 , \8733 );
buf \U$8025 ( \8735 , \4070 );
buf \U$8026 ( \8736 , \4991 );
nand \U$8027 ( \8737 , \8735 , \8736 );
buf \U$8028 ( \8738 , \8737 );
buf \U$8029 ( \8739 , \8738 );
nand \U$8030 ( \8740 , \8734 , \8739 );
buf \U$8031 ( \8741 , \8740 );
buf \U$8032 ( \8742 , \8741 );
not \U$8033 ( \8743 , \8742 );
buf \U$8034 ( \8744 , \2645 );
not \U$8035 ( \8745 , \8744 );
or \U$8036 ( \8746 , \8743 , \8745 );
buf \U$8037 ( \8747 , \2473 );
buf \U$8038 ( \8748 , \8236 );
nand \U$8039 ( \8749 , \8747 , \8748 );
buf \U$8040 ( \8750 , \8749 );
buf \U$8041 ( \8751 , \8750 );
nand \U$8042 ( \8752 , \8746 , \8751 );
buf \U$8043 ( \8753 , \8752 );
buf \U$8044 ( \8754 , \8753 );
nand \U$8045 ( \8755 , \8729 , \8754 );
buf \U$8046 ( \8756 , \8755 );
buf \U$8047 ( \8757 , \8756 );
nand \U$8048 ( \8758 , \8726 , \8757 );
buf \U$8049 ( \8759 , \8758 );
buf \U$8050 ( \8760 , \8759 );
and \U$8051 ( \8761 , \8641 , \8760 );
buf \U$8052 ( \8762 , \8629 );
not \U$8053 ( \8763 , \8762 );
buf \U$8054 ( \8764 , \8637 );
nor \U$8055 ( \8765 , \8763 , \8764 );
buf \U$8056 ( \8766 , \8765 );
buf \U$8057 ( \8767 , \8766 );
nor \U$8058 ( \8768 , \8761 , \8767 );
buf \U$8059 ( \8769 , \8768 );
buf \U$8060 ( \8770 , \8769 );
xor \U$8061 ( \8771 , \8571 , \8770 );
buf \U$8062 ( \8772 , \8315 );
buf \U$8063 ( \8773 , \8177 );
and \U$8064 ( \8774 , \8772 , \8773 );
not \U$8065 ( \8775 , \8772 );
buf \U$8066 ( \8776 , \8212 );
and \U$8067 ( \8777 , \8775 , \8776 );
nor \U$8068 ( \8778 , \8774 , \8777 );
buf \U$8069 ( \8779 , \8778 );
buf \U$8070 ( \8780 , \8779 );
buf \U$8071 ( \8781 , \8205 );
not \U$8072 ( \8782 , \8781 );
buf \U$8073 ( \8783 , \8782 );
buf \U$8074 ( \8784 , \8783 );
and \U$8075 ( \8785 , \8780 , \8784 );
not \U$8076 ( \8786 , \8780 );
buf \U$8077 ( \8787 , \8205 );
and \U$8078 ( \8788 , \8786 , \8787 );
nor \U$8079 ( \8789 , \8785 , \8788 );
buf \U$8080 ( \8790 , \8789 );
buf \U$8081 ( \8791 , \8790 );
and \U$8082 ( \8792 , \8771 , \8791 );
and \U$8083 ( \8793 , \8571 , \8770 );
or \U$8084 ( \8794 , \8792 , \8793 );
buf \U$8085 ( \8795 , \8794 );
buf \U$8086 ( \8796 , \8795 );
nand \U$8087 ( \8797 , \8568 , \8796 );
buf \U$8088 ( \8798 , \8797 );
buf \U$8089 ( \8799 , \8798 );
xor \U$8090 ( \8800 , \8571 , \8770 );
xor \U$8091 ( \8801 , \8800 , \8791 );
buf \U$8092 ( \8802 , \8801 );
buf \U$8093 ( \8803 , \8802 );
xor \U$8094 ( \8804 , \8629 , \8759 );
xor \U$8095 ( \8805 , \8804 , \8637 );
buf \U$8096 ( \8806 , \8309 );
buf \U$8097 ( \8807 , \8271 );
and \U$8098 ( \8808 , \8806 , \8807 );
not \U$8099 ( \8809 , \8806 );
buf \U$8100 ( \8810 , \8282 );
and \U$8101 ( \8811 , \8809 , \8810 );
nor \U$8102 ( \8812 , \8808 , \8811 );
buf \U$8103 ( \8813 , \8812 );
buf \U$8104 ( \8814 , \8813 );
buf \U$8108 ( \8815 , \8242 );
xnor \U$8109 ( \8816 , \8814 , \8815 );
buf \U$8110 ( \8817 , \8816 );
buf \U$8113 ( \8818 , \8817 );
nand \U$8114 ( \8819 , \8805 , \8818 );
buf \U$8115 ( \8820 , \8819 );
buf \U$8116 ( \8821 , \3223 );
not \U$8117 ( \8822 , \8821 );
buf \U$8118 ( \8823 , \4282 );
not \U$8119 ( \8824 , \8823 );
or \U$8120 ( \8825 , \8822 , \8824 );
buf \U$8121 ( \8826 , \4278 );
buf \U$8122 ( \8827 , \3459 );
nand \U$8123 ( \8828 , \8826 , \8827 );
buf \U$8124 ( \8829 , \8828 );
buf \U$8125 ( \8830 , \8829 );
nand \U$8126 ( \8831 , \8825 , \8830 );
buf \U$8127 ( \8832 , \8831 );
buf \U$8128 ( \8833 , \8832 );
not \U$8129 ( \8834 , \8833 );
buf \U$8130 ( \8835 , \7659 );
not \U$8131 ( \8836 , \8835 );
or \U$8132 ( \8837 , \8834 , \8836 );
buf \U$8133 ( \8838 , \6582 );
buf \U$8134 ( \8839 , \8297 );
nand \U$8135 ( \8840 , \8838 , \8839 );
buf \U$8136 ( \8841 , \8840 );
buf \U$8137 ( \8842 , \8841 );
nand \U$8138 ( \8843 , \8837 , \8842 );
buf \U$8139 ( \8844 , \8843 );
buf \U$8140 ( \8845 , \8844 );
not \U$8141 ( \8846 , \8845 );
buf \U$8142 ( \8847 , \8846 );
buf \U$8143 ( \8848 , \8847 );
not \U$8144 ( \8849 , \8848 );
buf \U$8145 ( \8850 , \8696 );
not \U$8146 ( \8851 , \8850 );
buf \U$8147 ( \8852 , \8669 );
not \U$8148 ( \8853 , \8852 );
and \U$8149 ( \8854 , \8851 , \8853 );
buf \U$8150 ( \8855 , \8696 );
buf \U$8151 ( \8856 , \8669 );
and \U$8152 ( \8857 , \8855 , \8856 );
nor \U$8153 ( \8858 , \8854 , \8857 );
buf \U$8154 ( \8859 , \8858 );
buf \U$8155 ( \8860 , \8859 );
buf \U$8156 ( \8861 , \2853 );
buf \U$8157 ( \8862 , \4794 );
and \U$8158 ( \8863 , \8861 , \8862 );
not \U$8159 ( \8864 , \8861 );
buf \U$8160 ( \8865 , \4795 );
and \U$8161 ( \8866 , \8864 , \8865 );
nor \U$8162 ( \8867 , \8863 , \8866 );
buf \U$8163 ( \8868 , \8867 );
buf \U$8164 ( \8869 , \8868 );
not \U$8165 ( \8870 , \8869 );
buf \U$8166 ( \8871 , \5388 );
not \U$8167 ( \8872 , \8871 );
and \U$8168 ( \8873 , \8870 , \8872 );
buf \U$8169 ( \8874 , \8614 );
buf \U$8170 ( \8875 , \5398 );
and \U$8171 ( \8876 , \8874 , \8875 );
nor \U$8172 ( \8877 , \8873 , \8876 );
buf \U$8173 ( \8878 , \8877 );
buf \U$8174 ( \8879 , \8878 );
nand \U$8175 ( \8880 , \8860 , \8879 );
buf \U$8176 ( \8881 , \8880 );
buf \U$8177 ( \8882 , \8881 );
buf \U$8178 ( \8883 , \4863 );
buf \U$8179 ( \8884 , \3134 );
or \U$8180 ( \8885 , \8883 , \8884 );
buf \U$8181 ( \8886 , \7833 );
buf \U$8182 ( \8887 , \4855 );
or \U$8183 ( \8888 , \8886 , \8887 );
nand \U$8184 ( \8889 , \8885 , \8888 );
buf \U$8185 ( \8890 , \8889 );
buf \U$8186 ( \8891 , \8890 );
not \U$8187 ( \8892 , \8891 );
buf \U$8188 ( \8893 , \5615 );
not \U$8189 ( \8894 , \8893 );
or \U$8190 ( \8895 , \8892 , \8894 );
buf \U$8191 ( \8896 , \8711 );
buf \U$8192 ( \8897 , \3095 );
nand \U$8193 ( \8898 , \8896 , \8897 );
buf \U$8194 ( \8899 , \8898 );
buf \U$8195 ( \8900 , \8899 );
nand \U$8196 ( \8901 , \8895 , \8900 );
buf \U$8197 ( \8902 , \8901 );
buf \U$8198 ( \8903 , \8902 );
and \U$8199 ( \8904 , \8882 , \8903 );
buf \U$8200 ( \8905 , \8859 );
buf \U$8201 ( \8906 , \8878 );
nor \U$8202 ( \8907 , \8905 , \8906 );
buf \U$8203 ( \8908 , \8907 );
buf \U$8204 ( \8909 , \8908 );
nor \U$8205 ( \8910 , \8904 , \8909 );
buf \U$8206 ( \8911 , \8910 );
buf \U$8207 ( \8912 , \8911 );
not \U$8208 ( \8913 , \8912 );
or \U$8209 ( \8914 , \8849 , \8913 );
xor \U$8210 ( \8915 , \8602 , \8607 );
xor \U$8211 ( \8916 , \8915 , \8625 );
buf \U$8212 ( \8917 , \8916 );
buf \U$8213 ( \8918 , \8917 );
nand \U$8214 ( \8919 , \8914 , \8918 );
buf \U$8215 ( \8920 , \8919 );
buf \U$8216 ( \8921 , \8920 );
or \U$8217 ( \8922 , \8911 , \8847 );
buf \U$8218 ( \8923 , \8922 );
nand \U$8219 ( \8924 , \8921 , \8923 );
buf \U$8220 ( \8925 , \8924 );
buf \U$8224 ( \8926 , \8925 );
and \U$8225 ( \8927 , \8820 , \8926 );
buf \U$8226 ( \8928 , \8629 );
buf \U$8227 ( \8929 , \8759 );
xor \U$8228 ( \8930 , \8928 , \8929 );
buf \U$8229 ( \8931 , \8637 );
xnor \U$8230 ( \8932 , \8930 , \8931 );
buf \U$8231 ( \8933 , \8932 );
buf \U$8232 ( \8934 , \8933 );
not \U$8233 ( \8935 , \8934 );
buf \U$8234 ( \8936 , \8935 );
buf \U$8235 ( \8937 , \8936 );
buf \U$8236 ( \8938 , \8818 );
nor \U$8237 ( \8939 , \8937 , \8938 );
buf \U$8238 ( \8940 , \8939 );
buf \U$8239 ( \8941 , \8940 );
nor \U$8240 ( \8942 , \8927 , \8941 );
buf \U$8241 ( \8943 , \8942 );
buf \U$8242 ( \8944 , \8943 );
nand \U$8243 ( \8945 , \8803 , \8944 );
buf \U$8244 ( \8946 , \8945 );
buf \U$8245 ( \8947 , \8946 );
nand \U$8246 ( \8948 , \8799 , \8947 );
buf \U$8247 ( \8949 , \8948 );
buf \U$8248 ( \8950 , \8949 );
not \U$8249 ( \8951 , \8950 );
buf \U$8250 ( \8952 , \8951 );
buf \U$8251 ( \8953 , \8952 );
buf \U$8252 ( \8954 , \8925 );
not \U$8253 ( \8955 , \8954 );
buf \U$8254 ( \8956 , \8817 );
not \U$8255 ( \8957 , \8956 );
and \U$8256 ( \8958 , \8955 , \8957 );
buf \U$8257 ( \8959 , \8925 );
buf \U$8258 ( \8960 , \8817 );
and \U$8259 ( \8961 , \8959 , \8960 );
nor \U$8260 ( \8962 , \8958 , \8961 );
buf \U$8261 ( \8963 , \8962 );
buf \U$8262 ( \8964 , \8963 );
not \U$8263 ( \8965 , \8964 );
buf \U$8264 ( \8966 , \8933 );
not \U$8265 ( \8967 , \8966 );
or \U$8266 ( \8968 , \8965 , \8967 );
buf \U$8267 ( \8969 , \8933 );
buf \U$8268 ( \8970 , \8963 );
or \U$8269 ( \8971 , \8969 , \8970 );
nand \U$8270 ( \8972 , \8968 , \8971 );
buf \U$8271 ( \8973 , \8972 );
buf \U$8272 ( \8974 , \8973 );
buf \U$8273 ( \8975 , \5321 );
not \U$8274 ( \8976 , \8975 );
buf \U$8275 ( \8977 , \2479 );
not \U$8276 ( \8978 , \8977 );
or \U$8277 ( \8979 , \8976 , \8978 );
buf \U$8278 ( \8980 , \7800 );
buf \U$8279 ( \8981 , \3276 );
nand \U$8280 ( \8982 , \8980 , \8981 );
buf \U$8281 ( \8983 , \8982 );
buf \U$8282 ( \8984 , \8983 );
nand \U$8283 ( \8985 , \8979 , \8984 );
buf \U$8284 ( \8986 , \8985 );
buf \U$8285 ( \8987 , \8986 );
not \U$8286 ( \8988 , \8987 );
buf \U$8287 ( \8989 , \2645 );
not \U$8288 ( \8990 , \8989 );
or \U$8289 ( \8991 , \8988 , \8990 );
buf \U$8290 ( \8992 , \2473 );
buf \U$8291 ( \8993 , \8741 );
nand \U$8292 ( \8994 , \8992 , \8993 );
buf \U$8293 ( \8995 , \8994 );
buf \U$8294 ( \8996 , \8995 );
nand \U$8295 ( \8997 , \8991 , \8996 );
buf \U$8296 ( \8998 , \8997 );
buf \U$8297 ( \8999 , \8998 );
not \U$8298 ( \9000 , \8999 );
buf \U$8299 ( \9001 , \3444 );
not \U$8300 ( \9002 , \9001 );
buf \U$8301 ( \9003 , \4282 );
not \U$8302 ( \9004 , \9003 );
or \U$8303 ( \9005 , \9002 , \9004 );
buf \U$8304 ( \9006 , \4381 );
buf \U$8305 ( \9007 , \4278 );
nand \U$8306 ( \9008 , \9006 , \9007 );
buf \U$8307 ( \9009 , \9008 );
buf \U$8308 ( \9010 , \9009 );
nand \U$8309 ( \9011 , \9005 , \9010 );
buf \U$8310 ( \9012 , \9011 );
buf \U$8311 ( \9013 , \9012 );
not \U$8312 ( \9014 , \9013 );
buf \U$8313 ( \9015 , \7659 );
not \U$8314 ( \9016 , \9015 );
or \U$8315 ( \9017 , \9014 , \9016 );
buf \U$8316 ( \9018 , \6582 );
buf \U$8317 ( \9019 , \8832 );
nand \U$8318 ( \9020 , \9018 , \9019 );
buf \U$8319 ( \9021 , \9020 );
buf \U$8320 ( \9022 , \9021 );
nand \U$8321 ( \9023 , \9017 , \9022 );
buf \U$8322 ( \9024 , \9023 );
buf \U$8323 ( \9025 , \9024 );
not \U$8324 ( \9026 , \9025 );
or \U$8325 ( \9027 , \9000 , \9026 );
buf \U$8326 ( \9028 , \8998 );
not \U$8327 ( \9029 , \9028 );
buf \U$8328 ( \9030 , \9024 );
not \U$8329 ( \9031 , \9030 );
buf \U$8330 ( \9032 , \9031 );
buf \U$8331 ( \9033 , \9032 );
nand \U$8332 ( \9034 , \9029 , \9033 );
buf \U$8333 ( \9035 , \9034 );
buf \U$8334 ( \9036 , \9035 );
buf \U$8335 ( \9037 , \2473 );
buf \U$8336 ( \9038 , \5321 );
nand \U$8337 ( \9039 , \9037 , \9038 );
buf \U$8338 ( \9040 , \9039 );
buf \U$8339 ( \9041 , \9040 );
and \U$8340 ( \9042 , \5463 , RI9151258_522);
and \U$8341 ( \9043 , \963 , RI91519d8_538);
nor \U$8342 ( \9044 , \9042 , \9043 );
not \U$8343 ( \9045 , \6273 );
and \U$8344 ( \9046 , \9045 , RI9152158_554);
and \U$8345 ( \9047 , \7762 , RI91528d8_570);
nor \U$8346 ( \9048 , \9046 , \9047 );
and \U$8347 ( \9049 , \7094 , RI9153058_586);
and \U$8348 ( \9050 , \1635 , RI91537d8_602);
nor \U$8349 ( \9051 , \9049 , \9050 );
and \U$8350 ( \9052 , \5451 , RI9153f58_618);
and \U$8351 ( \9053 , \5453 , RI91546d8_634);
nor \U$8352 ( \9054 , \9052 , \9053 );
nand \U$8353 ( \9055 , \9044 , \9048 , \9051 , \9054 );
and \U$8354 ( \9056 , \4644 , RI9154e58_650);
and \U$8355 ( \9057 , \8573 , RI91555d8_666);
nor \U$8356 ( \9058 , \9056 , \9057 );
and \U$8357 ( \9059 , \5428 , RI9155d58_682);
and \U$8358 ( \9060 , \5430 , RI91564d8_698);
nor \U$8359 ( \9061 , \9059 , \9060 );
and \U$8360 ( \9062 , \5434 , RI9156c58_714);
and \U$8361 ( \9063 , \1200 , RI91573d8_730);
nor \U$8362 ( \9064 , \9062 , \9063 );
and \U$8363 ( \9065 , \1014 , RI9157b58_746);
and \U$8364 ( \9066 , \4011 , RI91582d8_762);
nor \U$8365 ( \9067 , \9065 , \9066 );
nand \U$8366 ( \9068 , \9058 , \9061 , \9064 , \9067 );
or \U$8367 ( \9069 , \9055 , \9068 );
buf \U$8368 ( \9070 , \9069 );
not \U$8369 ( \9071 , \9070 );
buf \U$8370 ( \9072 , \9071 );
buf \U$8371 ( \9073 , \9072 );
nand \U$8372 ( \9074 , \9041 , \9073 );
buf \U$8373 ( \9075 , \9074 );
buf \U$8374 ( \9076 , \9075 );
not \U$8375 ( \9077 , \9076 );
buf \U$8376 ( \9078 , \4848 );
not \U$8377 ( \9079 , \9078 );
buf \U$8378 ( \9080 , \7833 );
not \U$8379 ( \9081 , \9080 );
or \U$8380 ( \9082 , \9079 , \9081 );
buf \U$8381 ( \9083 , \4991 );
buf \U$8382 ( \9084 , \3134 );
nand \U$8383 ( \9085 , \9083 , \9084 );
buf \U$8384 ( \9086 , \9085 );
buf \U$8385 ( \9087 , \9086 );
nand \U$8386 ( \9088 , \9082 , \9087 );
buf \U$8387 ( \9089 , \9088 );
buf \U$8388 ( \9090 , \9089 );
not \U$8389 ( \9091 , \9090 );
buf \U$8390 ( \9092 , \5615 );
not \U$8391 ( \9093 , \9092 );
or \U$8392 ( \9094 , \9091 , \9093 );
buf \U$8393 ( \9095 , \3095 );
buf \U$8394 ( \9096 , \8890 );
nand \U$8395 ( \9097 , \9095 , \9096 );
buf \U$8396 ( \9098 , \9097 );
buf \U$8397 ( \9099 , \9098 );
nand \U$8398 ( \9100 , \9094 , \9099 );
buf \U$8399 ( \9101 , \9100 );
buf \U$8400 ( \9102 , \9101 );
not \U$8401 ( \9103 , \9102 );
or \U$8402 ( \9104 , \9077 , \9103 );
buf \U$8403 ( \9105 , \9040 );
not \U$8404 ( \9106 , \9105 );
buf \U$8405 ( \9107 , \9106 );
buf \U$8406 ( \9108 , \9107 );
buf \U$8407 ( \9109 , \9069 );
nand \U$8408 ( \9110 , \9108 , \9109 );
buf \U$8409 ( \9111 , \9110 );
buf \U$8410 ( \9112 , \9111 );
nand \U$8411 ( \9113 , \9104 , \9112 );
buf \U$8412 ( \9114 , \9113 );
buf \U$8413 ( \9115 , \9114 );
nand \U$8414 ( \9116 , \9036 , \9115 );
buf \U$8415 ( \9117 , \9116 );
buf \U$8416 ( \9118 , \9117 );
nand \U$8417 ( \9119 , \9027 , \9118 );
buf \U$8418 ( \9120 , \9119 );
buf \U$8419 ( \9121 , \9120 );
xor \U$8420 ( \9122 , \8697 , \8723 );
xor \U$8421 ( \9123 , \9122 , \8753 );
buf \U$8422 ( \9124 , \9123 );
xor \U$8423 ( \9125 , \9121 , \9124 );
buf \U$8424 ( \9126 , \8844 );
buf \U$8425 ( \9127 , \8917 );
xor \U$8426 ( \9128 , \9126 , \9127 );
buf \U$8427 ( \9129 , \8911 );
xnor \U$8428 ( \9130 , \9128 , \9129 );
buf \U$8429 ( \9131 , \9130 );
buf \U$8430 ( \9132 , \9131 );
and \U$8431 ( \9133 , \9125 , \9132 );
and \U$8432 ( \9134 , \9121 , \9124 );
or \U$8433 ( \9135 , \9133 , \9134 );
buf \U$8434 ( \9136 , \9135 );
buf \U$8435 ( \9137 , \9136 );
nand \U$8436 ( \9138 , \8974 , \9137 );
buf \U$8437 ( \9139 , \9138 );
not \U$8438 ( \9140 , \9139 );
xor \U$8439 ( \9141 , \9121 , \9124 );
xor \U$8440 ( \9142 , \9141 , \9132 );
buf \U$8441 ( \9143 , \9142 );
buf \U$8442 ( \9144 , \9143 );
buf \U$8443 ( \9145 , \5391 );
not \U$8444 ( \9146 , \9145 );
buf \U$8445 ( \9147 , \3223 );
not \U$8446 ( \9148 , \9147 );
buf \U$8447 ( \9149 , \4795 );
not \U$8448 ( \9150 , \9149 );
or \U$8449 ( \9151 , \9148 , \9150 );
buf \U$8450 ( \9152 , \3459 );
not \U$8451 ( \9153 , \4794 );
not \U$8452 ( \9154 , \9153 );
buf \U$8453 ( \9155 , \9154 );
nand \U$8454 ( \9156 , \9152 , \9155 );
buf \U$8455 ( \9157 , \9156 );
buf \U$8456 ( \9158 , \9157 );
nand \U$8457 ( \9159 , \9151 , \9158 );
buf \U$8458 ( \9160 , \9159 );
buf \U$8459 ( \9161 , \9160 );
not \U$8460 ( \9162 , \9161 );
or \U$8461 ( \9163 , \9146 , \9162 );
buf \U$8462 ( \9164 , \8868 );
not \U$8463 ( \9165 , \9164 );
buf \U$8464 ( \9166 , \5398 );
nand \U$8465 ( \9167 , \9165 , \9166 );
buf \U$8466 ( \9168 , \9167 );
buf \U$8467 ( \9169 , \9168 );
nand \U$8468 ( \9170 , \9163 , \9169 );
buf \U$8469 ( \9171 , \9170 );
buf \U$8470 ( \9172 , \9171 );
and \U$8471 ( \9173 , \4644 , RI9154ed0_651);
and \U$8472 ( \9174 , \8573 , RI9155650_667);
nor \U$8473 ( \9175 , \9173 , \9174 );
and \U$8474 ( \9176 , \5428 , RI9155dd0_683);
and \U$8475 ( \9177 , \5430 , RI9156550_699);
nor \U$8476 ( \9178 , \9176 , \9177 );
and \U$8477 ( \9179 , \9175 , \9178 );
and \U$8478 ( \9180 , \7094 , RI91530d0_587);
and \U$8479 ( \9181 , \1635 , RI9153850_603);
nor \U$8480 ( \9182 , \9180 , \9181 );
and \U$8481 ( \9183 , \5451 , RI9153fd0_619);
and \U$8482 ( \9184 , \5453 , RI9154750_635);
nor \U$8483 ( \9185 , \9183 , \9184 );
and \U$8484 ( \9186 , \9182 , \9185 );
and \U$8485 ( \9187 , \5463 , RI91512d0_523);
and \U$8486 ( \9188 , \963 , RI9151a50_539);
nor \U$8487 ( \9189 , \9187 , \9188 );
and \U$8488 ( \9190 , \7106 , RI91521d0_555);
and \U$8489 ( \9191 , \1623 , RI9152950_571);
nor \U$8490 ( \9192 , \9190 , \9191 );
and \U$8491 ( \9193 , \9189 , \9192 );
and \U$8492 ( \9194 , \5434 , RI9156cd0_715);
and \U$8493 ( \9195 , \1200 , RI9157450_731);
nor \U$8494 ( \9196 , \9194 , \9195 );
and \U$8495 ( \9197 , \1014 , RI9157bd0_747);
and \U$8496 ( \9198 , \4011 , RI9158350_763);
nor \U$8497 ( \9199 , \9197 , \9198 );
and \U$8498 ( \9200 , \9196 , \9199 );
nand \U$8499 ( \9201 , \9179 , \9186 , \9193 , \9200 );
buf \U$8500 ( \9202 , \9201 );
buf \U$8501 ( \9203 , \3115 );
not \U$8502 ( \9204 , \9203 );
buf \U$8503 ( \9205 , \7800 );
not \U$8504 ( \9206 , \9205 );
or \U$8505 ( \9207 , \9204 , \9206 );
buf \U$8506 ( \9208 , \4278 );
nand \U$8507 ( \9209 , \9207 , \9208 );
buf \U$8508 ( \9210 , \9209 );
buf \U$8509 ( \9211 , \9210 );
buf \U$8510 ( \9212 , \3115 );
not \U$8511 ( \9213 , \9212 );
buf \U$8512 ( \9214 , \5321 );
nand \U$8513 ( \9215 , \9213 , \9214 );
buf \U$8514 ( \9216 , \9215 );
buf \U$8515 ( \9217 , \9216 );
buf \U$8516 ( \9218 , \7839 );
and \U$8517 ( \9219 , \9211 , \9217 , \9218 );
buf \U$8518 ( \9220 , \9219 );
buf \U$8519 ( \9221 , \9220 );
and \U$8520 ( \9222 , \9202 , \9221 );
buf \U$8521 ( \9223 , \9222 );
buf \U$8522 ( \9224 , \9223 );
xor \U$8523 ( \9225 , \9172 , \9224 );
buf \U$8524 ( \9226 , \4032 );
not \U$8525 ( \9227 , \9226 );
buf \U$8526 ( \9228 , \4282 );
not \U$8527 ( \9229 , \9228 );
or \U$8528 ( \9230 , \9227 , \9229 );
buf \U$8529 ( \9231 , \4029 );
buf \U$8530 ( \9232 , \4278 );
nand \U$8531 ( \9233 , \9231 , \9232 );
buf \U$8532 ( \9234 , \9233 );
buf \U$8533 ( \9235 , \9234 );
nand \U$8534 ( \9236 , \9230 , \9235 );
buf \U$8535 ( \9237 , \9236 );
buf \U$8536 ( \9238 , \9237 );
not \U$8537 ( \9239 , \9238 );
buf \U$8538 ( \9240 , \6578 );
not \U$8539 ( \9241 , \9240 );
or \U$8540 ( \9242 , \9239 , \9241 );
buf \U$8541 ( \9243 , \9012 );
buf \U$8542 ( \9244 , \4581 );
nand \U$8543 ( \9245 , \9243 , \9244 );
buf \U$8544 ( \9246 , \9245 );
buf \U$8545 ( \9247 , \9246 );
nand \U$8546 ( \9248 , \9242 , \9247 );
buf \U$8547 ( \9249 , \9248 );
buf \U$8548 ( \9250 , \9249 );
and \U$8549 ( \9251 , \9225 , \9250 );
and \U$8550 ( \9252 , \9172 , \9224 );
or \U$8551 ( \9253 , \9251 , \9252 );
buf \U$8552 ( \9254 , \9253 );
buf \U$8553 ( \9255 , \9254 );
xor \U$8554 ( \9256 , \8878 , \8859 );
xor \U$8555 ( \9257 , \8902 , \9256 );
buf \U$8556 ( \9258 , \9257 );
xor \U$8557 ( \9259 , \9255 , \9258 );
xor \U$8558 ( \9260 , \8998 , \9032 );
xnor \U$8559 ( \9261 , \9260 , \9114 );
buf \U$8560 ( \9262 , \9261 );
and \U$8561 ( \9263 , \9259 , \9262 );
and \U$8562 ( \9264 , \9255 , \9258 );
or \U$8563 ( \9265 , \9263 , \9264 );
buf \U$8564 ( \9266 , \9265 );
buf \U$8565 ( \9267 , \9266 );
nand \U$8566 ( \9268 , \9144 , \9267 );
buf \U$8567 ( \9269 , \9268 );
not \U$8568 ( \9270 , \9269 );
or \U$8569 ( \9271 , \9140 , \9270 );
buf \U$8570 ( \9272 , \8973 );
not \U$8571 ( \9273 , \9272 );
buf \U$8572 ( \9274 , \9273 );
buf \U$8573 ( \9275 , \9274 );
buf \U$8574 ( \9276 , \9136 );
not \U$8575 ( \9277 , \9276 );
buf \U$8576 ( \9278 , \9277 );
buf \U$8577 ( \9279 , \9278 );
nand \U$8578 ( \9280 , \9275 , \9279 );
buf \U$8579 ( \9281 , \9280 );
nand \U$8580 ( \9282 , \9271 , \9281 );
buf \U$8581 ( \9283 , \9282 );
buf \U$8582 ( \9284 , \8802 );
not \U$8583 ( \9285 , \9284 );
buf \U$8584 ( \9286 , \9285 );
buf \U$8585 ( \9287 , \9286 );
buf \U$8586 ( \9288 , \8943 );
not \U$8587 ( \9289 , \9288 );
buf \U$8588 ( \9290 , \9289 );
buf \U$8589 ( \9291 , \9290 );
nand \U$8590 ( \9292 , \9287 , \9291 );
buf \U$8591 ( \9293 , \9292 );
buf \U$8592 ( \9294 , \9293 );
nand \U$8593 ( \9295 , \9283 , \9294 );
buf \U$8594 ( \9296 , \9295 );
buf \U$8595 ( \9297 , \9296 );
and \U$8596 ( \9298 , \8953 , \9297 );
buf \U$8600 ( \9299 , \8567 );
buf \U$8601 ( \9300 , \8795 );
nor \U$8602 ( \9301 , \9299 , \9300 );
buf \U$8603 ( \9302 , \9301 );
buf \U$8604 ( \9303 , \9302 );
nor \U$8605 ( \9304 , \9298 , \9303 );
buf \U$8606 ( \9305 , \9304 );
buf \U$8607 ( \9306 , \9305 );
buf \U$8608 ( \9307 , \8952 );
buf \U$8609 ( \9308 , \9281 );
buf \U$8610 ( \9309 , \9143 );
not \U$8611 ( \9310 , \9309 );
buf \U$8612 ( \9311 , \9310 );
buf \U$8613 ( \9312 , \9311 );
buf \U$8614 ( \9313 , \9266 );
not \U$8615 ( \9314 , \9313 );
buf \U$8616 ( \9315 , \9314 );
buf \U$8617 ( \9316 , \9315 );
nand \U$8618 ( \9317 , \9312 , \9316 );
buf \U$8619 ( \9318 , \9317 );
buf \U$8620 ( \9319 , \9318 );
and \U$8621 ( \9320 , \9308 , \9319 );
buf \U$8622 ( \9321 , \9320 );
buf \U$8623 ( \9322 , \9321 );
xor \U$8624 ( \9323 , \9172 , \9224 );
xor \U$8625 ( \9324 , \9323 , \9250 );
buf \U$8626 ( \9325 , \9324 );
buf \U$8629 ( \9326 , \9325 );
buf \U$8630 ( \9327 , \9326 );
buf \U$8631 ( \9328 , \9072 );
not \U$8632 ( \9329 , \9328 );
buf \U$8633 ( \9330 , \9107 );
not \U$8634 ( \9331 , \9330 );
or \U$8635 ( \9332 , \9329 , \9331 );
buf \U$8636 ( \9333 , \9040 );
buf \U$8637 ( \9334 , \9069 );
nand \U$8638 ( \9335 , \9333 , \9334 );
buf \U$8639 ( \9336 , \9335 );
buf \U$8640 ( \9337 , \9336 );
nand \U$8641 ( \9338 , \9332 , \9337 );
buf \U$8642 ( \9339 , \9338 );
buf \U$8643 ( \9340 , \9339 );
buf \U$8644 ( \9341 , \9101 );
xor \U$8645 ( \9342 , \9340 , \9341 );
buf \U$8646 ( \9343 , \9342 );
buf \U$8647 ( \9344 , \9343 );
or \U$8648 ( \9345 , \9327 , \9344 );
buf \U$8649 ( \9346 , \5506 );
not \U$8650 ( \9347 , \9346 );
buf \U$8651 ( \9348 , \3444 );
not \U$8652 ( \9349 , \9348 );
buf \U$8653 ( \9350 , \5330 );
not \U$8654 ( \9351 , \9350 );
or \U$8655 ( \9352 , \9349 , \9351 );
buf \U$8656 ( \9353 , \9154 );
buf \U$8657 ( \9354 , \4381 );
nand \U$8658 ( \9355 , \9353 , \9354 );
buf \U$8659 ( \9356 , \9355 );
buf \U$8660 ( \9357 , \9356 );
nand \U$8661 ( \9358 , \9352 , \9357 );
buf \U$8662 ( \9359 , \9358 );
buf \U$8663 ( \9360 , \9359 );
not \U$8664 ( \9361 , \9360 );
or \U$8665 ( \9362 , \9347 , \9361 );
buf \U$8666 ( \9363 , \9160 );
buf \U$8667 ( \9364 , \5398 );
nand \U$8668 ( \9365 , \9363 , \9364 );
buf \U$8669 ( \9366 , \9365 );
buf \U$8670 ( \9367 , \9366 );
nand \U$8671 ( \9368 , \9362 , \9367 );
buf \U$8672 ( \9369 , \9368 );
buf \U$8673 ( \9370 , \9369 );
xor \U$8674 ( \9371 , \9202 , \9221 );
buf \U$8675 ( \9372 , \9371 );
buf \U$8676 ( \9373 , \9372 );
xor \U$8677 ( \9374 , \9370 , \9373 );
buf \U$8678 ( \9375 , \5321 );
not \U$8679 ( \9376 , \9375 );
buf \U$8680 ( \9377 , \7833 );
not \U$8681 ( \9378 , \9377 );
or \U$8682 ( \9379 , \9376 , \9378 );
buf \U$8683 ( \9380 , \7800 );
buf \U$8684 ( \9381 , \3134 );
nand \U$8685 ( \9382 , \9380 , \9381 );
buf \U$8686 ( \9383 , \9382 );
buf \U$8687 ( \9384 , \9383 );
nand \U$8688 ( \9385 , \9379 , \9384 );
buf \U$8689 ( \9386 , \9385 );
buf \U$8690 ( \9387 , \9386 );
not \U$8691 ( \9388 , \9387 );
buf \U$8692 ( \9389 , \5615 );
not \U$8693 ( \9390 , \9389 );
or \U$8694 ( \9391 , \9388 , \9390 );
buf \U$8695 ( \9392 , \3095 );
buf \U$8696 ( \9393 , \9089 );
nand \U$8697 ( \9394 , \9392 , \9393 );
buf \U$8698 ( \9395 , \9394 );
buf \U$8699 ( \9396 , \9395 );
nand \U$8700 ( \9397 , \9391 , \9396 );
buf \U$8701 ( \9398 , \9397 );
buf \U$8702 ( \9399 , \9398 );
and \U$8703 ( \9400 , \9374 , \9399 );
and \U$8704 ( \9401 , \9370 , \9373 );
or \U$8705 ( \9402 , \9400 , \9401 );
buf \U$8706 ( \9403 , \9402 );
buf \U$8707 ( \9404 , \9403 );
nand \U$8708 ( \9405 , \9345 , \9404 );
buf \U$8709 ( \9406 , \9405 );
buf \U$8710 ( \9407 , \9406 );
buf \U$8711 ( \9408 , \9326 );
buf \U$8712 ( \9409 , \9343 );
nand \U$8713 ( \9410 , \9408 , \9409 );
buf \U$8714 ( \9411 , \9410 );
buf \U$8715 ( \9412 , \9411 );
nand \U$8716 ( \9413 , \9407 , \9412 );
buf \U$8717 ( \9414 , \9413 );
buf \U$8718 ( \9415 , \9414 );
xor \U$8719 ( \9416 , \9255 , \9258 );
xor \U$8720 ( \9417 , \9416 , \9262 );
buf \U$8721 ( \9418 , \9417 );
buf \U$8722 ( \9419 , \9418 );
xor \U$8723 ( \9420 , \9415 , \9419 );
buf \U$8724 ( \9421 , \9403 );
not \U$8725 ( \9422 , \9421 );
buf \U$8726 ( \9423 , \9422 );
buf \U$8727 ( \9424 , \9423 );
not \U$8728 ( \9425 , \9424 );
buf \U$8729 ( \9426 , \9325 );
not \U$8730 ( \9427 , \9426 );
or \U$8731 ( \9428 , \9425 , \9427 );
buf \U$8732 ( \9429 , \9423 );
buf \U$8733 ( \9430 , \9325 );
or \U$8734 ( \9431 , \9429 , \9430 );
nand \U$8735 ( \9432 , \9428 , \9431 );
buf \U$8736 ( \9433 , \9432 );
buf \U$8737 ( \9434 , \9433 );
buf \U$8738 ( \9435 , \9343 );
not \U$8739 ( \9436 , \9435 );
buf \U$8740 ( \9437 , \9436 );
buf \U$8741 ( \9438 , \9437 );
and \U$8742 ( \9439 , \9434 , \9438 );
not \U$8743 ( \9440 , \9434 );
buf \U$8744 ( \9441 , \9343 );
and \U$8745 ( \9442 , \9440 , \9441 );
nor \U$8746 ( \9443 , \9439 , \9442 );
buf \U$8747 ( \9444 , \9443 );
buf \U$8748 ( \9445 , \9444 );
xor \U$8749 ( \9446 , \9370 , \9373 );
xor \U$8750 ( \9447 , \9446 , \9399 );
buf \U$8751 ( \9448 , \9447 );
buf \U$8752 ( \9449 , \9448 );
buf \U$8753 ( \9450 , \4863 );
not \U$8754 ( \9451 , \9450 );
buf \U$8755 ( \9452 , \4278 );
not \U$8756 ( \9453 , \9452 );
or \U$8757 ( \9454 , \9451 , \9453 );
buf \U$8758 ( \9455 , \4281 );
buf \U$8759 ( \9456 , \4678 );
nand \U$8760 ( \9457 , \9455 , \9456 );
buf \U$8761 ( \9458 , \9457 );
buf \U$8762 ( \9459 , \9458 );
nand \U$8763 ( \9460 , \9454 , \9459 );
buf \U$8764 ( \9461 , \9460 );
buf \U$8765 ( \9462 , \9461 );
not \U$8766 ( \9463 , \9462 );
buf \U$8767 ( \9464 , \7659 );
not \U$8768 ( \9465 , \9464 );
or \U$8769 ( \9466 , \9463 , \9465 );
buf \U$8770 ( \9467 , \9237 );
buf \U$8771 ( \9468 , \6582 );
nand \U$8772 ( \9469 , \9467 , \9468 );
buf \U$8773 ( \9470 , \9469 );
buf \U$8774 ( \9471 , \9470 );
nand \U$8775 ( \9472 , \9466 , \9471 );
buf \U$8776 ( \9473 , \9472 );
buf \U$8777 ( \9474 , \9473 );
or \U$8778 ( \9475 , \9449 , \9474 );
buf \U$8779 ( \9476 , \9475 );
buf \U$8780 ( \9477 , \9476 );
buf \U$8781 ( \9478 , \4260 );
not \U$8782 ( \9479 , \9478 );
buf \U$8783 ( \9480 , \5475 );
nand \U$8784 ( \9481 , \9479 , \9480 );
buf \U$8785 ( \9482 , \9481 );
buf \U$8786 ( \9483 , \9482 );
buf \U$8787 ( \9484 , \4794 );
and \U$8788 ( \9485 , \9483 , \9484 );
buf \U$8789 ( \9486 , \5321 );
not \U$8790 ( \9487 , \9486 );
buf \U$8791 ( \9488 , \4260 );
not \U$8792 ( \9489 , \9488 );
or \U$8793 ( \9490 , \9487 , \9489 );
buf \U$8794 ( \9491 , \4278 );
nand \U$8795 ( \9492 , \9490 , \9491 );
buf \U$8796 ( \9493 , \9492 );
buf \U$8797 ( \9494 , \9493 );
nor \U$8798 ( \9495 , \9485 , \9494 );
buf \U$8799 ( \9496 , \9495 );
buf \U$8800 ( \9497 , \9496 );
and \U$8801 ( \9498 , \4003 , RI9156dc0_717);
and \U$8802 ( \9499 , \1200 , RI9157540_733);
nor \U$8803 ( \9500 , \9498 , \9499 );
and \U$8804 ( \9501 , \5428 , RI9155ec0_685);
and \U$8805 ( \9502 , \5430 , RI9156640_701);
nor \U$8806 ( \9503 , \9501 , \9502 );
nand \U$8807 ( \9504 , \9500 , \9503 );
and \U$8808 ( \9505 , \4644 , RI9154fc0_653);
and \U$8809 ( \9506 , \8573 , RI9155740_669);
nor \U$8810 ( \9507 , \9505 , \9506 );
and \U$8811 ( \9508 , \1014 , RI9157cc0_749);
and \U$8812 ( \9509 , \4011 , RI9158440_765);
nor \U$8813 ( \9510 , \9508 , \9509 );
nand \U$8814 ( \9511 , \9507 , \9510 );
nor \U$8815 ( \9512 , \9504 , \9511 );
and \U$8816 ( \9513 , \5463 , RI91513c0_525);
and \U$8817 ( \9514 , \963 , RI9151b40_541);
nor \U$8818 ( \9515 , \9513 , \9514 );
not \U$8819 ( \9516 , RI91522c0_557);
nor \U$8820 ( \9517 , \9516 , \922 );
not \U$8821 ( \9518 , RI9152a40_573);
nor \U$8822 ( \9519 , \9518 , \929 );
nor \U$8823 ( \9520 , \9517 , \9519 );
nand \U$8824 ( \9521 , \9515 , \9520 );
not \U$8825 ( \9522 , RI91531c0_589);
nor \U$8826 ( \9523 , \9522 , \1282 );
not \U$8827 ( \9524 , RI9153940_605);
nor \U$8828 ( \9525 , \9524 , \957 );
nor \U$8829 ( \9526 , \9523 , \9525 );
and \U$8830 ( \9527 , \5451 , RI91540c0_621);
and \U$8831 ( \9528 , \5453 , RI9154840_637);
nor \U$8832 ( \9529 , \9527 , \9528 );
nand \U$8833 ( \9530 , \9526 , \9529 );
nor \U$8834 ( \9531 , \9521 , \9530 );
nand \U$8835 ( \9532 , \9512 , \9531 );
buf \U$8836 ( \9533 , \9532 );
nand \U$8837 ( \9534 , \9497 , \9533 );
buf \U$8838 ( \9535 , \9534 );
buf \U$8839 ( \9536 , \9535 );
not \U$8840 ( \9537 , \9536 );
buf \U$8841 ( \9538 , \9537 );
buf \U$8842 ( \9539 , \9538 );
and \U$8843 ( \9540 , \7094 , RI9153148_588);
and \U$8844 ( \9541 , \1500 , RI91538c8_604);
nor \U$8845 ( \9542 , \9540 , \9541 );
and \U$8846 ( \9543 , \9045 , RI9152248_556);
and \U$8847 ( \9544 , \7762 , RI91529c8_572);
nor \U$8848 ( \9545 , \9543 , \9544 );
and \U$8849 ( \9546 , \9542 , \9545 );
and \U$8850 ( \9547 , \4644 , RI9154f48_652);
and \U$8851 ( \9548 , \8573 , RI91556c8_668);
nor \U$8852 ( \9549 , \9547 , \9548 );
and \U$8853 ( \9550 , \5434 , RI9156d48_716);
and \U$8854 ( \9551 , \1200 , RI91574c8_732);
nor \U$8855 ( \9552 , \9550 , \9551 );
and \U$8856 ( \9553 , \9549 , \9552 );
and \U$8857 ( \9554 , \5428 , RI9155e48_684);
and \U$8858 ( \9555 , \5430 , RI91565c8_700);
nor \U$8859 ( \9556 , \9554 , \9555 );
and \U$8860 ( \9557 , \1014 , RI9157c48_748);
and \U$8861 ( \9558 , \4011 , RI91583c8_764);
nor \U$8862 ( \9559 , \9557 , \9558 );
and \U$8863 ( \9560 , \9556 , \9559 );
and \U$8864 ( \9561 , \5463 , RI9151348_524);
and \U$8865 ( \9562 , \963 , RI9151ac8_540);
nor \U$8866 ( \9563 , \9561 , \9562 );
and \U$8867 ( \9564 , \5451 , RI9154048_620);
and \U$8868 ( \9565 , \5453 , RI91547c8_636);
nor \U$8869 ( \9566 , \9564 , \9565 );
and \U$8870 ( \9567 , \9563 , \9566 );
nand \U$8871 ( \9568 , \9546 , \9553 , \9560 , \9567 );
buf \U$8872 ( \9569 , \9568 );
buf \U$8873 ( \9570 , \3094 );
buf \U$8874 ( \9571 , \5321 );
and \U$8875 ( \9572 , \9570 , \9571 );
buf \U$8876 ( \9573 , \9572 );
buf \U$8877 ( \9574 , \9573 );
or \U$8878 ( \9575 , \9569 , \9574 );
buf \U$8879 ( \9576 , \9575 );
buf \U$8880 ( \9577 , \9576 );
and \U$8881 ( \9578 , \9539 , \9577 );
buf \U$8882 ( \9579 , \9568 );
buf \U$8883 ( \9580 , \9573 );
and \U$8884 ( \9581 , \9579 , \9580 );
buf \U$8885 ( \9582 , \9581 );
buf \U$8886 ( \9583 , \9582 );
nor \U$8887 ( \9584 , \9578 , \9583 );
buf \U$8888 ( \9585 , \9584 );
buf \U$8889 ( \9586 , \9585 );
not \U$8890 ( \9587 , \9586 );
buf \U$8891 ( \9588 , \9587 );
buf \U$8892 ( \9589 , \9588 );
and \U$8893 ( \9590 , \9477 , \9589 );
buf \U$8894 ( \9591 , \9448 );
buf \U$8895 ( \9592 , \9473 );
and \U$8896 ( \9593 , \9591 , \9592 );
buf \U$8897 ( \9594 , \9593 );
buf \U$8898 ( \9595 , \9594 );
nor \U$8899 ( \9596 , \9590 , \9595 );
buf \U$8900 ( \9597 , \9596 );
buf \U$8901 ( \9598 , \9597 );
nand \U$8902 ( \9599 , \9445 , \9598 );
buf \U$8903 ( \9600 , \9599 );
buf \U$8904 ( \9601 , \9600 );
not \U$8905 ( \9602 , \9601 );
buf \U$8906 ( \9603 , \4848 );
not \U$8907 ( \9604 , \9603 );
buf \U$8908 ( \9605 , \4281 );
not \U$8909 ( \9606 , \9605 );
or \U$8910 ( \9607 , \9604 , \9606 );
buf \U$8911 ( \9608 , \4278 );
buf \U$8912 ( \9609 , \4991 );
nand \U$8913 ( \9610 , \9608 , \9609 );
buf \U$8914 ( \9611 , \9610 );
buf \U$8915 ( \9612 , \9611 );
nand \U$8916 ( \9613 , \9607 , \9612 );
buf \U$8917 ( \9614 , \9613 );
buf \U$8918 ( \9615 , \9614 );
not \U$8919 ( \9616 , \9615 );
buf \U$8920 ( \9617 , \4248 );
buf \U$8921 ( \9618 , \4270 );
nand \U$8922 ( \9619 , \9617 , \9618 );
buf \U$8923 ( \9620 , \9619 );
buf \U$8924 ( \9621 , \9620 );
not \U$8925 ( \9622 , \9621 );
buf \U$8926 ( \9623 , \9622 );
buf \U$8927 ( \9624 , \9623 );
not \U$8928 ( \9625 , \9624 );
or \U$8929 ( \9626 , \9616 , \9625 );
buf \U$8930 ( \9627 , \9461 );
buf \U$8931 ( \9628 , \4581 );
nand \U$8932 ( \9629 , \9627 , \9628 );
buf \U$8933 ( \9630 , \9629 );
buf \U$8934 ( \9631 , \9630 );
nand \U$8935 ( \9632 , \9626 , \9631 );
buf \U$8936 ( \9633 , \9632 );
buf \U$8937 ( \9634 , \9633 );
not \U$8938 ( \9635 , \9634 );
buf \U$8939 ( \9636 , \5398 );
not \U$8940 ( \9637 , \9636 );
buf \U$8941 ( \9638 , \9359 );
not \U$8942 ( \9639 , \9638 );
or \U$8943 ( \9640 , \9637 , \9639 );
buf \U$8944 ( \9641 , \5506 );
and \U$8945 ( \9642 , \4026 , \4795 );
not \U$8946 ( \9643 , \4026 );
and \U$8947 ( \9644 , \9643 , \4794 );
or \U$8948 ( \9645 , \9642 , \9644 );
buf \U$8949 ( \9646 , \9645 );
nand \U$8950 ( \9647 , \9641 , \9646 );
buf \U$8951 ( \9648 , \9647 );
buf \U$8952 ( \9649 , \9648 );
nand \U$8953 ( \9650 , \9640 , \9649 );
buf \U$8954 ( \9651 , \9650 );
buf \U$8955 ( \9652 , \9651 );
not \U$8956 ( \9653 , \9652 );
buf \U$8957 ( \9654 , \9653 );
buf \U$8958 ( \9655 , \9654 );
not \U$8959 ( \9656 , \9655 );
and \U$8960 ( \9657 , \9635 , \9656 );
buf \U$8961 ( \9658 , \9654 );
buf \U$8962 ( \9659 , \9633 );
and \U$8963 ( \9660 , \9658 , \9659 );
nor \U$8964 ( \9661 , \9657 , \9660 );
buf \U$8965 ( \9662 , \9661 );
buf \U$8966 ( \9663 , \9662 );
not \U$8967 ( \9664 , \9663 );
buf \U$8968 ( \9665 , \9538 );
not \U$8969 ( \9666 , \9665 );
xor \U$8970 ( \9667 , \9579 , \9580 );
buf \U$8971 ( \9668 , \9667 );
buf \U$8972 ( \9669 , \9668 );
not \U$8973 ( \9670 , \9669 );
buf \U$8974 ( \9671 , \9670 );
buf \U$8975 ( \9672 , \9671 );
not \U$8976 ( \9673 , \9672 );
or \U$8977 ( \9674 , \9666 , \9673 );
buf \U$8978 ( \9675 , \9668 );
buf \U$8979 ( \9676 , \9535 );
nand \U$8980 ( \9677 , \9675 , \9676 );
buf \U$8981 ( \9678 , \9677 );
buf \U$8982 ( \9679 , \9678 );
nand \U$8983 ( \9680 , \9674 , \9679 );
buf \U$8984 ( \9681 , \9680 );
buf \U$8985 ( \9682 , \9681 );
not \U$8986 ( \9683 , \9682 );
and \U$8987 ( \9684 , \9664 , \9683 );
buf \U$8988 ( \9685 , \9662 );
buf \U$8989 ( \9686 , \9681 );
and \U$8990 ( \9687 , \9685 , \9686 );
nor \U$8991 ( \9688 , \9684 , \9687 );
buf \U$8992 ( \9689 , \9688 );
buf \U$8993 ( \9690 , \9689 );
buf \U$8994 ( \9691 , \5398 );
not \U$8995 ( \9692 , \9691 );
buf \U$8996 ( \9693 , \9645 );
not \U$8997 ( \9694 , \9693 );
or \U$8998 ( \9695 , \9692 , \9694 );
buf \U$8999 ( \9696 , \4855 );
not \U$9000 ( \9697 , \9696 );
buf \U$9001 ( \9698 , \9153 );
not \U$9002 ( \9699 , \9698 );
or \U$9003 ( \9700 , \9697 , \9699 );
buf \U$9004 ( \9701 , \4794 );
buf \U$9005 ( \9702 , \4675 );
nand \U$9006 ( \9703 , \9701 , \9702 );
buf \U$9007 ( \9704 , \9703 );
buf \U$9008 ( \9705 , \9704 );
nand \U$9009 ( \9706 , \9700 , \9705 );
buf \U$9010 ( \9707 , \9706 );
buf \U$9011 ( \9708 , \9707 );
buf \U$9012 ( \9709 , \5506 );
nand \U$9013 ( \9710 , \9708 , \9709 );
buf \U$9014 ( \9711 , \9710 );
buf \U$9015 ( \9712 , \9711 );
nand \U$9016 ( \9713 , \9695 , \9712 );
buf \U$9017 ( \9714 , \9713 );
buf \U$9018 ( \9715 , \9714 );
not \U$9019 ( \9716 , \9715 );
buf \U$9020 ( \9717 , \9716 );
buf \U$9021 ( \9718 , \9717 );
buf \U$9022 ( \9719 , \9496 );
not \U$9023 ( \9720 , \9719 );
buf \U$9024 ( \9721 , \9532 );
not \U$9025 ( \9722 , \9721 );
buf \U$9026 ( \9723 , \9722 );
buf \U$9027 ( \9724 , \9723 );
not \U$9028 ( \9725 , \9724 );
and \U$9029 ( \9726 , \9720 , \9725 );
buf \U$9030 ( \9727 , \9496 );
buf \U$9031 ( \9728 , \9723 );
and \U$9032 ( \9729 , \9727 , \9728 );
nor \U$9033 ( \9730 , \9726 , \9729 );
buf \U$9034 ( \9731 , \9730 );
buf \U$9035 ( \9732 , \9731 );
xor \U$9036 ( \9733 , \9718 , \9732 );
not \U$9037 ( \9734 , \9620 );
buf \U$9038 ( \9735 , \4278 );
buf \U$9039 ( \9736 , \7800 );
and \U$9040 ( \9737 , \9735 , \9736 );
not \U$9041 ( \9738 , \9735 );
buf \U$9042 ( \9739 , \5321 );
and \U$9043 ( \9740 , \9738 , \9739 );
nor \U$9044 ( \9741 , \9737 , \9740 );
buf \U$9045 ( \9742 , \9741 );
not \U$9046 ( \9743 , \9742 );
and \U$9047 ( \9744 , \9734 , \9743 );
buf \U$9048 ( \9745 , \9614 );
not \U$9049 ( \9746 , \9745 );
buf \U$9050 ( \9747 , \5065 );
nor \U$9051 ( \9748 , \9746 , \9747 );
buf \U$9052 ( \9749 , \9748 );
nor \U$9053 ( \9750 , \9744 , \9749 );
buf \U$9054 ( \9751 , \9750 );
and \U$9055 ( \9752 , \9733 , \9751 );
and \U$9056 ( \9753 , \9718 , \9732 );
or \U$9057 ( \9754 , \9752 , \9753 );
buf \U$9058 ( \9755 , \9754 );
buf \U$9059 ( \9756 , \9755 );
nand \U$9060 ( \9757 , \9690 , \9756 );
buf \U$9061 ( \9758 , \9757 );
buf \U$9062 ( \9759 , \9758 );
not \U$9063 ( \9760 , \9759 );
xor \U$9064 ( \9761 , \9718 , \9732 );
xor \U$9065 ( \9762 , \9761 , \9751 );
buf \U$9066 ( \9763 , \9762 );
buf \U$9067 ( \9764 , \9763 );
and \U$9068 ( \9765 , \5434 , RI9156e38_718);
and \U$9069 ( \9766 , \2052 , RI91575b8_734);
nor \U$9070 ( \9767 , \9765 , \9766 );
and \U$9071 ( \9768 , \5428 , RI9155f38_686);
and \U$9072 ( \9769 , \5430 , RI91566b8_702);
nor \U$9073 ( \9770 , \9768 , \9769 );
nand \U$9074 ( \9771 , \9767 , \9770 );
and \U$9075 ( \9772 , \4644 , RI9155038_654);
and \U$9076 ( \9773 , \1765 , RI91557b8_670);
nor \U$9077 ( \9774 , \9772 , \9773 );
and \U$9078 ( \9775 , \6239 , RI9157d38_750);
and \U$9079 ( \9776 , \4011 , RI91584b8_766);
nor \U$9080 ( \9777 , \9775 , \9776 );
nand \U$9081 ( \9778 , \9774 , \9777 );
nor \U$9082 ( \9779 , \9771 , \9778 );
not \U$9083 ( \9780 , \957 );
not \U$9084 ( \9781 , RI91539b8_606);
not \U$9085 ( \9782 , \9781 );
and \U$9086 ( \9783 , \9780 , \9782 );
not \U$9087 ( \9784 , RI9153238_590);
nor \U$9088 ( \9785 , \9784 , \952 );
nor \U$9089 ( \9786 , \9783 , \9785 );
and \U$9090 ( \9787 , \9045 , RI9152338_558);
and \U$9091 ( \9788 , \1623 , RI9152ab8_574);
nor \U$9092 ( \9789 , \9787 , \9788 );
nand \U$9093 ( \9790 , \9786 , \9789 );
and \U$9094 ( \9791 , \5463 , RI9151438_526);
and \U$9095 ( \9792 , \963 , RI9151bb8_542);
nor \U$9096 ( \9793 , \9791 , \9792 );
and \U$9097 ( \9794 , \5451 , RI9154138_622);
and \U$9098 ( \9795 , \5453 , RI91548b8_638);
nor \U$9099 ( \9796 , \9794 , \9795 );
nand \U$9100 ( \9797 , \9793 , \9796 );
nor \U$9101 ( \9798 , \9790 , \9797 );
and \U$9102 ( \9799 , \9779 , \9798 );
buf \U$9103 ( \9800 , \9799 );
buf \U$9104 ( \9801 , \4581 );
buf \U$9105 ( \9802 , \5321 );
nand \U$9106 ( \9803 , \9801 , \9802 );
buf \U$9107 ( \9804 , \9803 );
buf \U$9108 ( \9805 , \9804 );
xor \U$9109 ( \9806 , \9800 , \9805 );
buf \U$9110 ( \9807 , \5397 );
buf \U$9111 ( \9808 , \5321 );
nand \U$9112 ( \9809 , \9807 , \9808 );
buf \U$9113 ( \9810 , \9809 );
buf \U$9114 ( \9811 , \9810 );
not \U$9115 ( \9812 , \4795 );
buf \U$9116 ( \9813 , \9812 );
and \U$9117 ( \9814 , \9811 , \9813 );
buf \U$9118 ( \9815 , \9814 );
buf \U$9119 ( \9816 , \9815 );
and \U$9120 ( \9817 , \4644 , RI91550b0_655);
and \U$9121 ( \9818 , \8573 , RI9155830_671);
nor \U$9122 ( \9819 , \9817 , \9818 );
and \U$9123 ( \9820 , \6052 , RI9155fb0_687);
and \U$9124 ( \9821 , \5430 , RI9156730_703);
nor \U$9125 ( \9822 , \9820 , \9821 );
and \U$9126 ( \9823 , \5434 , RI9156eb0_719);
and \U$9127 ( \9824 , \2052 , RI9157630_735);
nor \U$9128 ( \9825 , \9823 , \9824 );
and \U$9129 ( \9826 , \1014 , RI9157db0_751);
and \U$9130 ( \9827 , \5439 , RI9158530_767);
nor \U$9131 ( \9828 , \9826 , \9827 );
and \U$9132 ( \9829 , \9819 , \9822 , \9825 , \9828 );
and \U$9133 ( \9830 , \5463 , RI91514b0_527);
and \U$9134 ( \9831 , \963 , RI9151c30_543);
nor \U$9135 ( \9832 , \9830 , \9831 );
and \U$9136 ( \9833 , \7762 , RI9152b30_575);
not \U$9137 ( \9834 , RI91523b0_559);
nor \U$9138 ( \9835 , \9834 , \6273 );
nor \U$9139 ( \9836 , \9833 , \9835 );
not \U$9140 ( \9837 , \957 );
not \U$9141 ( \9838 , RI9153a30_607);
not \U$9142 ( \9839 , \9838 );
and \U$9143 ( \9840 , \9837 , \9839 );
not \U$9144 ( \9841 , RI91532b0_591);
nor \U$9145 ( \9842 , \9841 , \1282 );
nor \U$9146 ( \9843 , \9840 , \9842 );
and \U$9147 ( \9844 , \5451 , RI91541b0_623);
and \U$9148 ( \9845 , \5453 , RI9154930_639);
nor \U$9149 ( \9846 , \9844 , \9845 );
and \U$9150 ( \9847 , \9832 , \9836 , \9843 , \9846 );
nand \U$9151 ( \9848 , \9829 , \9847 );
buf \U$9152 ( \9849 , \9848 );
nand \U$9153 ( \9850 , \9816 , \9849 );
buf \U$9154 ( \9851 , \9850 );
buf \U$9155 ( \9852 , \9851 );
and \U$9156 ( \9853 , \9806 , \9852 );
and \U$9157 ( \9854 , \9800 , \9805 );
or \U$9158 ( \9855 , \9853 , \9854 );
buf \U$9159 ( \9856 , \9855 );
buf \U$9160 ( \9857 , \9856 );
nand \U$9161 ( \9858 , \9764 , \9857 );
buf \U$9162 ( \9859 , \9858 );
not \U$9163 ( \9860 , \9859 );
and \U$9164 ( \9861 , \1206 , RI9156028_688);
and \U$9165 ( \9862 , \5430 , RI91567a8_704);
nor \U$9166 ( \9863 , \9861 , \9862 );
and \U$9167 ( \9864 , \4644 , RI9155128_656);
and \U$9168 ( \9865 , \984 , RI91558a8_672);
nor \U$9169 ( \9866 , \9864 , \9865 );
nand \U$9170 ( \9867 , \9863 , \9866 );
and \U$9171 ( \9868 , \4003 , RI9156f28_720);
and \U$9172 ( \9869 , \2052 , RI91576a8_736);
nor \U$9173 ( \9870 , \9868 , \9869 );
and \U$9174 ( \9871 , \6239 , RI9157e28_752);
and \U$9175 ( \9872 , \4011 , RI91585a8_768);
nor \U$9176 ( \9873 , \9871 , \9872 );
nand \U$9177 ( \9874 , \9870 , \9873 );
nor \U$9178 ( \9875 , \9867 , \9874 );
nand \U$9179 ( \9876 , \5463 , RI9151528_528);
nand \U$9180 ( \9877 , \1623 , RI9152ba8_576);
nand \U$9181 ( \9878 , \7106 , RI9152428_560);
nand \U$9182 ( \9879 , RI9151ca8_544, \963 );
nand \U$9183 ( \9880 , \9876 , \9877 , \9878 , \9879 );
nand \U$9184 ( \9881 , \7094 , RI9153328_592);
nand \U$9185 ( \9882 , \5453 , RI91549a8_640);
nand \U$9186 ( \9883 , \8005 , RI9153aa8_608);
nand \U$9187 ( \9884 , \7099 , RI9154228_624);
nand \U$9188 ( \9885 , \9881 , \9882 , \9883 , \9884 );
nor \U$9189 ( \9886 , \9880 , \9885 );
and \U$9190 ( \9887 , \9875 , \9886 );
nor \U$9191 ( \9888 , \9887 , \9810 );
buf \U$9192 ( \9889 , \9888 );
buf \U$9193 ( \9890 , \5398 );
not \U$9194 ( \9891 , \9890 );
buf \U$9195 ( \9892 , \4848 );
not \U$9196 ( \9893 , \9892 );
buf \U$9197 ( \9894 , \5330 );
not \U$9198 ( \9895 , \9894 );
or \U$9199 ( \9896 , \9893 , \9895 );
buf \U$9200 ( \9897 , \9812 );
buf \U$9201 ( \9898 , \4991 );
nand \U$9202 ( \9899 , \9897 , \9898 );
buf \U$9203 ( \9900 , \9899 );
buf \U$9204 ( \9901 , \9900 );
nand \U$9205 ( \9902 , \9896 , \9901 );
buf \U$9206 ( \9903 , \9902 );
buf \U$9207 ( \9904 , \9903 );
not \U$9208 ( \9905 , \9904 );
or \U$9209 ( \9906 , \9891 , \9905 );
buf \U$9210 ( \9907 , \7121 );
buf \U$9211 ( \9908 , \5573 );
nand \U$9212 ( \9909 , \9907 , \9908 );
buf \U$9213 ( \9910 , \9909 );
buf \U$9214 ( \9911 , \9910 );
nand \U$9215 ( \9912 , \9906 , \9911 );
buf \U$9216 ( \9913 , \9912 );
buf \U$9217 ( \9914 , \9913 );
xor \U$9218 ( \9915 , \9889 , \9914 );
xor \U$9219 ( \9916 , \9848 , \9815 );
buf \U$9220 ( \9917 , \9916 );
and \U$9221 ( \9918 , \9915 , \9917 );
and \U$9222 ( \9919 , \9889 , \9914 );
or \U$9223 ( \9920 , \9918 , \9919 );
buf \U$9224 ( \9921 , \9920 );
not \U$9225 ( \9922 , \9921 );
xor \U$9226 ( \9923 , \9800 , \9805 );
xor \U$9227 ( \9924 , \9923 , \9852 );
buf \U$9228 ( \9925 , \9924 );
buf \U$9229 ( \9926 , \9925 );
buf \U$9230 ( \9927 , \5391 );
buf \U$9231 ( \9928 , \9903 );
and \U$9232 ( \9929 , \9927 , \9928 );
buf \U$9233 ( \9930 , \9707 );
buf \U$9234 ( \9931 , \5398 );
and \U$9235 ( \9932 , \9930 , \9931 );
nor \U$9236 ( \9933 , \9929 , \9932 );
buf \U$9237 ( \9934 , \9933 );
buf \U$9238 ( \9935 , \9934 );
nand \U$9239 ( \9936 , \9926 , \9935 );
buf \U$9240 ( \9937 , \9936 );
not \U$9241 ( \9938 , \9937 );
or \U$9242 ( \9939 , \9922 , \9938 );
buf \U$9243 ( \9940 , \9925 );
not \U$9244 ( \9941 , \9940 );
buf \U$9245 ( \9942 , \9941 );
buf \U$9246 ( \9943 , \9942 );
buf \U$9247 ( \9944 , \9934 );
not \U$9248 ( \9945 , \9944 );
buf \U$9249 ( \9946 , \9945 );
buf \U$9250 ( \9947 , \9946 );
nand \U$9251 ( \9948 , \9943 , \9947 );
buf \U$9252 ( \9949 , \9948 );
nand \U$9253 ( \9950 , \9939 , \9949 );
not \U$9254 ( \9951 , \9950 );
or \U$9255 ( \9952 , \9860 , \9951 );
buf \U$9256 ( \9953 , \9763 );
not \U$9257 ( \9954 , \9953 );
buf \U$9258 ( \9955 , \9954 );
buf \U$9259 ( \9956 , \9955 );
buf \U$9260 ( \9957 , \9856 );
not \U$9261 ( \9958 , \9957 );
buf \U$9262 ( \9959 , \9958 );
buf \U$9263 ( \9960 , \9959 );
nand \U$9264 ( \9961 , \9956 , \9960 );
buf \U$9265 ( \9962 , \9961 );
nand \U$9266 ( \9963 , \9952 , \9962 );
buf \U$9267 ( \9964 , \9963 );
not \U$9268 ( \9965 , \9964 );
or \U$9269 ( \9966 , \9760 , \9965 );
buf \U$9270 ( \9967 , \9689 );
not \U$9271 ( \9968 , \9967 );
buf \U$9272 ( \9969 , \9968 );
buf \U$9273 ( \9970 , \9969 );
buf \U$9274 ( \9971 , \9755 );
not \U$9275 ( \9972 , \9971 );
buf \U$9276 ( \9973 , \9972 );
buf \U$9277 ( \9974 , \9973 );
nand \U$9278 ( \9975 , \9970 , \9974 );
buf \U$9279 ( \9976 , \9975 );
buf \U$9280 ( \9977 , \9976 );
nand \U$9281 ( \9978 , \9966 , \9977 );
buf \U$9282 ( \9979 , \9978 );
buf \U$9283 ( \9980 , \9979 );
not \U$9284 ( \9981 , \9980 );
buf \U$9285 ( \9982 , \9448 );
not \U$9286 ( \9983 , \9982 );
buf \U$9287 ( \9984 , \9585 );
not \U$9288 ( \9985 , \9984 );
buf \U$9289 ( \9986 , \9473 );
not \U$9290 ( \9987 , \9986 );
and \U$9291 ( \9988 , \9985 , \9987 );
buf \U$9292 ( \9989 , \9585 );
buf \U$9293 ( \9990 , \9473 );
and \U$9294 ( \9991 , \9989 , \9990 );
nor \U$9295 ( \9992 , \9988 , \9991 );
buf \U$9296 ( \9993 , \9992 );
buf \U$9297 ( \9994 , \9993 );
not \U$9298 ( \9995 , \9994 );
and \U$9299 ( \9996 , \9983 , \9995 );
buf \U$9300 ( \9997 , \9448 );
buf \U$9301 ( \9998 , \9993 );
and \U$9302 ( \9999 , \9997 , \9998 );
nor \U$9303 ( \10000 , \9996 , \9999 );
buf \U$9304 ( \10001 , \10000 );
buf \U$9305 ( \10002 , \10001 );
buf \U$9306 ( \10003 , \9681 );
buf \U$9307 ( \10004 , \9633 );
buf \U$9308 ( \10005 , \9651 );
or \U$9309 ( \10006 , \10004 , \10005 );
buf \U$9310 ( \10007 , \10006 );
buf \U$9311 ( \10008 , \10007 );
and \U$9312 ( \10009 , \10003 , \10008 );
buf \U$9313 ( \10010 , \9633 );
buf \U$9314 ( \10011 , \9651 );
and \U$9315 ( \10012 , \10010 , \10011 );
buf \U$9316 ( \10013 , \10012 );
buf \U$9317 ( \10014 , \10013 );
nor \U$9318 ( \10015 , \10009 , \10014 );
buf \U$9319 ( \10016 , \10015 );
buf \U$9320 ( \10017 , \10016 );
nand \U$9321 ( \10018 , \10002 , \10017 );
buf \U$9322 ( \10019 , \10018 );
buf \U$9323 ( \10020 , \10019 );
not \U$9324 ( \10021 , \10020 );
or \U$9325 ( \10022 , \9981 , \10021 );
buf \U$9326 ( \10023 , \10001 );
not \U$9327 ( \10024 , \10023 );
buf \U$9328 ( \10025 , \10024 );
buf \U$9329 ( \10026 , \10025 );
buf \U$9330 ( \10027 , \10016 );
not \U$9331 ( \10028 , \10027 );
buf \U$9332 ( \10029 , \10028 );
buf \U$9333 ( \10030 , \10029 );
nand \U$9334 ( \10031 , \10026 , \10030 );
buf \U$9335 ( \10032 , \10031 );
buf \U$9336 ( \10033 , \10032 );
nand \U$9337 ( \10034 , \10022 , \10033 );
buf \U$9338 ( \10035 , \10034 );
buf \U$9339 ( \10036 , \10035 );
not \U$9340 ( \10037 , \10036 );
or \U$9341 ( \10038 , \9602 , \10037 );
buf \U$9342 ( \10039 , \9444 );
not \U$9343 ( \10040 , \10039 );
buf \U$9344 ( \10041 , \10040 );
buf \U$9345 ( \10042 , \10041 );
buf \U$9346 ( \10043 , \9597 );
not \U$9347 ( \10044 , \10043 );
buf \U$9348 ( \10045 , \10044 );
buf \U$9349 ( \10046 , \10045 );
nand \U$9350 ( \10047 , \10042 , \10046 );
buf \U$9351 ( \10048 , \10047 );
buf \U$9352 ( \10049 , \10048 );
nand \U$9353 ( \10050 , \10038 , \10049 );
buf \U$9354 ( \10051 , \10050 );
buf \U$9355 ( \10052 , \10051 );
and \U$9356 ( \10053 , \9420 , \10052 );
and \U$9357 ( \10054 , \9415 , \9419 );
or \U$9358 ( \10055 , \10053 , \10054 );
buf \U$9359 ( \10056 , \10055 );
buf \U$9360 ( \10057 , \10056 );
nand \U$9361 ( \10058 , \9307 , \9322 , \10057 );
buf \U$9362 ( \10059 , \10058 );
buf \U$9363 ( \10060 , \10059 );
nand \U$9364 ( \10061 , \9306 , \10060 );
buf \U$9365 ( \10062 , \10061 );
buf \U$9366 ( \10063 , \10062 );
not \U$9367 ( \10064 , \10063 );
or \U$9368 ( \10065 , \8549 , \10064 );
buf \U$9370 ( \10066 , \8492 );
not \U$9371 ( \10067 , \10066 );
buf \U$9372 ( \10068 , \10067 );
buf \U$9373 ( \10069 , \10068 );
not \U$9374 ( \10070 , \10069 );
or \U$9375 ( \10071 , 1'b0 , \10070 );
buf \U$9376 ( \10072 , \8541 );
buf \U$9377 ( \10073 , \8408 );
buf \U$9378 ( \10074 , \8414 );
nand \U$9379 ( \10075 , \10073 , \10074 );
buf \U$9380 ( \10076 , \10075 );
buf \U$9381 ( \10077 , \10076 );
buf \U$9382 ( \10078 , \8134 );
buf \U$9383 ( \10079 , \8327 );
nand \U$9384 ( \10080 , \10078 , \10079 );
buf \U$9385 ( \10081 , \10080 );
buf \U$9386 ( \10082 , \10081 );
nand \U$9387 ( \10083 , \10077 , \10082 );
buf \U$9388 ( \10084 , \10083 );
buf \U$9389 ( \10085 , \10084 );
buf \U$9390 ( \10086 , \8417 );
not \U$9391 ( \10087 , \10086 );
buf \U$9392 ( \10088 , \10087 );
buf \U$9393 ( \10089 , \10088 );
nand \U$9394 ( \10090 , \10072 , \10085 , \10089 );
buf \U$9395 ( \10091 , \10090 );
buf \U$9396 ( \10092 , \10091 );
buf \U$9397 ( \10093 , \8444 );
not \U$9398 ( \10094 , \10093 );
buf \U$9399 ( \10095 , \10094 );
buf \U$9400 ( \10096 , \10095 );
buf \U$9401 ( \10097 , \8486 );
nand \U$9402 ( \10098 , \10096 , \10097 );
buf \U$9403 ( \10099 , \10098 );
buf \U$9404 ( \10100 , \10099 );
buf \U$9405 ( \10101 , \8516 );
not \U$9406 ( \10102 , \10101 );
buf \U$9407 ( \10103 , \10102 );
buf \U$9408 ( \10104 , \10103 );
buf \U$9409 ( \10105 , \8535 );
nand \U$9410 ( \10106 , \10104 , \10105 );
buf \U$9411 ( \10107 , \10106 );
buf \U$9412 ( \10108 , \10107 );
nand \U$9413 ( \10109 , \10092 , \10100 , \10108 );
buf \U$9414 ( \10110 , \10109 );
buf \U$9415 ( \10111 , \10110 );
nand \U$9416 ( \10112 , \10071 , \10111 );
buf \U$9417 ( \10113 , \10112 );
buf \U$9418 ( \10114 , \10113 );
nand \U$9419 ( \10115 , \10065 , \10114 );
buf \U$9420 ( \10116 , \10115 );
buf \U$9421 ( \10117 , \10116 );
nand \U$9422 ( \10118 , \7470 , \7480 , \10117 );
buf \U$9423 ( \10119 , \10118 );
buf \U$9424 ( \10120 , \10119 );
nand \U$9425 ( \10121 , \7463 , \10120 );
buf \U$9426 ( \10122 , \10121 );
buf \U$9427 ( \10123 , \10122 );
not \U$9428 ( \10124 , \10123 );
or \U$9429 ( \10125 , \3918 , \10124 );
buf \U$9430 ( \10126 , \3752 );
buf \U$9431 ( \10127 , \3816 );
buf \U$9432 ( \10128 , \3877 );
and \U$9433 ( \10129 , \10126 , \10127 , \10128 );
buf \U$9434 ( \10130 , \10129 );
buf \U$9435 ( \10131 , \10130 );
not \U$9436 ( \10132 , \10131 );
buf \U$9437 ( \10133 , \3645 );
not \U$9438 ( \10134 , \10133 );
buf \U$9439 ( \10135 , \10134 );
buf \U$9440 ( \10136 , \10135 );
not \U$9441 ( \10137 , \10136 );
buf \U$9445 ( \10138 , \3531 );
buf \U$9446 ( \10139 , \2818 );
nor \U$9447 ( \10140 , \10138 , \10139 );
buf \U$9448 ( \10141 , \10140 );
not \U$9449 ( \10142 , \10141 );
not \U$9450 ( \10143 , \2814 );
or \U$9451 ( \10144 , \10142 , \10143 );
buf \U$9452 ( \10145 , \2561 );
buf \U$9453 ( \10146 , \2811 );
or \U$9454 ( \10147 , \10145 , \10146 );
buf \U$9455 ( \10148 , \10147 );
nand \U$9456 ( \10149 , \10144 , \10148 );
buf \U$9457 ( \10150 , \10149 );
not \U$9458 ( \10151 , \10150 );
or \U$9459 ( \10152 , \10137 , \10151 );
buf \U$9460 ( \10153 , \3548 );
buf \U$9461 ( \10154 , \3642 );
nand \U$9462 ( \10155 , \10153 , \10154 );
buf \U$9463 ( \10156 , \10155 );
buf \U$9464 ( \10157 , \10156 );
nand \U$9465 ( \10158 , \10152 , \10157 );
buf \U$9466 ( \10159 , \10158 );
buf \U$9467 ( \10160 , \10159 );
not \U$9468 ( \10161 , \10160 );
or \U$9469 ( \10162 , \10132 , \10161 );
buf \U$9470 ( \10163 , \3749 );
buf \U$9471 ( \10164 , \3743 );
nand \U$9472 ( \10165 , \10163 , \10164 );
buf \U$9473 ( \10166 , \10165 );
buf \U$9474 ( \10167 , \10166 );
buf \U$9475 ( \10168 , \3813 );
or \U$9476 ( \10169 , \10167 , \10168 );
buf \U$9477 ( \10170 , \3810 );
buf \U$9478 ( \10171 , \3804 );
nand \U$9479 ( \10172 , \10170 , \10171 );
buf \U$9480 ( \10173 , \10172 );
buf \U$9481 ( \10174 , \10173 );
nand \U$9482 ( \10175 , \10169 , \10174 );
buf \U$9483 ( \10176 , \10175 );
buf \U$9484 ( \10177 , \10176 );
buf \U$9485 ( \10178 , \3877 );
and \U$9486 ( \10179 , \10177 , \10178 );
buf \U$9487 ( \10180 , \3874 );
buf \U$9488 ( \10181 , \3868 );
and \U$9489 ( \10182 , \10180 , \10181 );
buf \U$9490 ( \10183 , \10182 );
buf \U$9491 ( \10184 , \10183 );
nor \U$9492 ( \10185 , \10179 , \10184 );
buf \U$9493 ( \10186 , \10185 );
buf \U$9494 ( \10187 , \10186 );
nand \U$9495 ( \10188 , \10162 , \10187 );
buf \U$9496 ( \10189 , \10188 );
buf \U$9497 ( \10190 , \10189 );
buf \U$9498 ( \10191 , \3913 );
not \U$9499 ( \10192 , \10191 );
buf \U$9500 ( \10193 , \10192 );
buf \U$9501 ( \10194 , \10193 );
and \U$9502 ( \10195 , \10190 , \10194 );
buf \U$9503 ( \10196 , \3886 );
buf \U$9504 ( \10197 , \3910 );
and \U$9505 ( \10198 , \10196 , \10197 );
buf \U$9506 ( \10199 , \10198 );
buf \U$9507 ( \10200 , \10199 );
nor \U$9508 ( \10201 , \10195 , \10200 );
buf \U$9509 ( \10202 , \10201 );
buf \U$9510 ( \10203 , \10202 );
nand \U$9511 ( \10204 , \10125 , \10203 );
buf \U$9512 ( \10205 , \10204 );
buf \U$9513 ( \10206 , \10205 );
buf \U$9514 ( \10207 , \3900 );
not \U$9515 ( \10208 , \10207 );
buf \U$9516 ( \10209 , \1619 );
buf \U$9517 ( \10210 , \2063 );
nand \U$9518 ( \10211 , \10209 , \10210 );
buf \U$9519 ( \10212 , \10211 );
buf \U$9520 ( \10213 , \10212 );
not \U$9521 ( \10214 , \10213 );
buf \U$9522 ( \10215 , \2296 );
buf \U$9523 ( \10216 , \1950 );
or \U$9524 ( \10217 , \10215 , \10216 );
buf \U$9525 ( \10218 , \1619 );
nand \U$9526 ( \10219 , \10217 , \10218 );
buf \U$9527 ( \10220 , \10219 );
buf \U$9528 ( \10221 , \10220 );
not \U$9529 ( \10222 , \10221 );
or \U$9530 ( \10223 , \10214 , \10222 );
buf \U$9531 ( \10224 , \10220 );
buf \U$9532 ( \10225 , \10212 );
or \U$9533 ( \10226 , \10224 , \10225 );
nand \U$9534 ( \10227 , \10223 , \10226 );
buf \U$9535 ( \10228 , \10227 );
buf \U$9536 ( \10229 , \10228 );
not \U$9537 ( \10230 , \10229 );
or \U$9538 ( \10231 , \10208 , \10230 );
buf \U$9539 ( \10232 , \10228 );
buf \U$9540 ( \10233 , \3900 );
or \U$9541 ( \10234 , \10232 , \10233 );
nand \U$9542 ( \10235 , \10231 , \10234 );
buf \U$9543 ( \10236 , \10235 );
buf \U$9544 ( \10237 , \10236 );
not \U$9545 ( \10238 , \10237 );
xor \U$9546 ( \10239 , \3896 , \3901 );
and \U$9547 ( \10240 , \10239 , \3908 );
and \U$9548 ( \10241 , \3896 , \3901 );
or \U$9549 ( \10242 , \10240 , \10241 );
buf \U$9550 ( \10243 , \10242 );
buf \U$9551 ( \10244 , \10243 );
not \U$9552 ( \10245 , \10244 );
or \U$9553 ( \10246 , \10238 , \10245 );
buf \U$9554 ( \10247 , \10243 );
buf \U$9555 ( \10248 , \10236 );
or \U$9556 ( \10249 , \10247 , \10248 );
nand \U$9557 ( \10250 , \10246 , \10249 );
buf \U$9558 ( \10251 , \10250 );
buf \U$9559 ( \10252 , \10251 );
not \U$9560 ( \10253 , \10252 );
buf \U$9561 ( \10254 , \10253 );
buf \U$9562 ( \10255 , \10254 );
and \U$9563 ( \10256 , \10206 , \10255 );
not \U$9564 ( \10257 , \10206 );
buf \U$9565 ( \10258 , \10251 );
and \U$9566 ( \10259 , \10257 , \10258 );
nor \U$9567 ( \10260 , \10256 , \10259 );
buf \U$9568 ( \10261 , \10260 );
buf \U$9569 ( \10262 , \10261 );
buf \U$9570 ( \10263 , \3880 );
not \U$9571 ( \10264 , \10263 );
buf \U$9572 ( \10265 , \10264 );
buf \U$9573 ( \10266 , \10265 );
not \U$9574 ( \10267 , \10266 );
buf \U$9575 ( \10268 , \10122 );
not \U$9576 ( \10269 , \10268 );
or \U$9577 ( \10270 , \10267 , \10269 );
buf \U$9578 ( \10271 , \10189 );
not \U$9579 ( \10272 , \10271 );
buf \U$9580 ( \10273 , \10272 );
buf \U$9581 ( \10274 , \10273 );
nand \U$9582 ( \10275 , \10270 , \10274 );
buf \U$9583 ( \10276 , \10275 );
buf \U$9584 ( \10277 , \10276 );
buf \U$9585 ( \10278 , \3913 );
buf \U$9586 ( \10279 , \10199 );
nor \U$9587 ( \10280 , \10278 , \10279 );
buf \U$9588 ( \10281 , \10280 );
buf \U$9589 ( \10282 , \10281 );
and \U$9590 ( \10283 , \10277 , \10282 );
not \U$9591 ( \10284 , \10277 );
buf \U$9592 ( \10285 , \10281 );
not \U$9593 ( \10286 , \10285 );
buf \U$9594 ( \10287 , \10286 );
buf \U$9595 ( \10288 , \10287 );
and \U$9596 ( \10289 , \10284 , \10288 );
nor \U$9597 ( \10290 , \10283 , \10289 );
buf \U$9598 ( \10291 , \10290 );
buf \U$9599 ( \10292 , \10291 );
buf \U$9600 ( \10293 , \3819 );
not \U$9601 ( \10294 , \10293 );
buf \U$9602 ( \10295 , \10122 );
not \U$9603 ( \10296 , \10295 );
or \U$9604 ( \10297 , \10294 , \10296 );
buf \U$9605 ( \10298 , \3752 );
not \U$9606 ( \10299 , \10298 );
buf \U$9607 ( \10300 , \10159 );
not \U$9608 ( \10301 , \10300 );
or \U$9609 ( \10302 , \10299 , \10301 );
buf \U$9610 ( \10303 , \10166 );
nand \U$9611 ( \10304 , \10302 , \10303 );
buf \U$9612 ( \10305 , \10304 );
buf \U$9613 ( \10306 , \10305 );
buf \U$9614 ( \10307 , \3816 );
and \U$9615 ( \10308 , \10306 , \10307 );
buf \U$9616 ( \10309 , \10173 );
not \U$9617 ( \10310 , \10309 );
buf \U$9618 ( \10311 , \10310 );
buf \U$9619 ( \10312 , \10311 );
nor \U$9620 ( \10313 , \10308 , \10312 );
buf \U$9621 ( \10314 , \10313 );
buf \U$9622 ( \10315 , \10314 );
nand \U$9623 ( \10316 , \10297 , \10315 );
buf \U$9624 ( \10317 , \10316 );
buf \U$9625 ( \10318 , \10317 );
buf \U$9626 ( \10319 , \10183 );
not \U$9627 ( \10320 , \10319 );
buf \U$9628 ( \10321 , \3877 );
nand \U$9629 ( \10322 , \10320 , \10321 );
buf \U$9630 ( \10323 , \10322 );
buf \U$9631 ( \10324 , \10323 );
not \U$9632 ( \10325 , \10324 );
buf \U$9633 ( \10326 , \10325 );
buf \U$9634 ( \10327 , \10326 );
and \U$9635 ( \10328 , \10318 , \10327 );
not \U$9636 ( \10329 , \10318 );
buf \U$9637 ( \10330 , \10323 );
and \U$9638 ( \10331 , \10329 , \10330 );
nor \U$9639 ( \10332 , \10328 , \10331 );
buf \U$9640 ( \10333 , \10332 );
buf \U$9641 ( \10334 , \10333 );
buf \U$9642 ( \10335 , \3755 );
not \U$9643 ( \10336 , \10335 );
buf \U$9644 ( \10337 , \10122 );
not \U$9645 ( \10338 , \10337 );
or \U$9646 ( \10339 , \10336 , \10338 );
buf \U$9647 ( \10340 , \10305 );
not \U$9648 ( \10341 , \10340 );
buf \U$9649 ( \10342 , \10341 );
buf \U$9650 ( \10343 , \10342 );
nand \U$9651 ( \10344 , \10339 , \10343 );
buf \U$9652 ( \10345 , \10344 );
buf \U$9653 ( \10346 , \10345 );
buf \U$9654 ( \10347 , \10173 );
buf \U$9655 ( \10348 , \3816 );
nand \U$9656 ( \10349 , \10347 , \10348 );
buf \U$9657 ( \10350 , \10349 );
buf \U$9658 ( \10351 , \10350 );
not \U$9659 ( \10352 , \10351 );
buf \U$9660 ( \10353 , \10352 );
buf \U$9661 ( \10354 , \10353 );
and \U$9662 ( \10355 , \10346 , \10354 );
not \U$9663 ( \10356 , \10346 );
buf \U$9664 ( \10357 , \10350 );
and \U$9665 ( \10358 , \10356 , \10357 );
nor \U$9666 ( \10359 , \10355 , \10358 );
buf \U$9667 ( \10360 , \10359 );
buf \U$9668 ( \10361 , \10360 );
buf \U$9669 ( \10362 , \3648 );
not \U$9670 ( \10363 , \10362 );
buf \U$9671 ( \10364 , \10122 );
not \U$9672 ( \10365 , \10364 );
or \U$9673 ( \10366 , \10363 , \10365 );
buf \U$9674 ( \10367 , \10159 );
not \U$9675 ( \10368 , \10367 );
buf \U$9676 ( \10369 , \10368 );
buf \U$9677 ( \10370 , \10369 );
nand \U$9678 ( \10371 , \10366 , \10370 );
buf \U$9679 ( \10372 , \10371 );
buf \U$9680 ( \10373 , \10372 );
buf \U$9681 ( \10374 , \3752 );
buf \U$9682 ( \10375 , \10166 );
nand \U$9683 ( \10376 , \10374 , \10375 );
buf \U$9684 ( \10377 , \10376 );
buf \U$9685 ( \10378 , \10377 );
not \U$9686 ( \10379 , \10378 );
buf \U$9687 ( \10380 , \10379 );
buf \U$9688 ( \10381 , \10380 );
and \U$9689 ( \10382 , \10373 , \10381 );
not \U$9690 ( \10383 , \10373 );
buf \U$9691 ( \10384 , \10377 );
and \U$9692 ( \10385 , \10383 , \10384 );
nor \U$9693 ( \10386 , \10382 , \10385 );
buf \U$9694 ( \10387 , \10386 );
buf \U$9695 ( \10388 , \10387 );
buf \U$9696 ( \10389 , \7479 );
not \U$9697 ( \10390 , \10389 );
buf \U$9698 ( \10391 , \10116 );
not \U$9699 ( \10392 , \10391 );
or \U$9700 ( \10393 , \10390 , \10392 );
buf \U$9701 ( \10394 , \7295 );
buf \U$9702 ( \10395 , \6441 );
not \U$9703 ( \10396 , \10395 );
buf \U$9704 ( \10397 , \10396 );
buf \U$9705 ( \10398 , \10397 );
buf \U$9706 ( \10399 , \6019 );
and \U$9707 ( \10400 , \10394 , \10398 , \10399 );
buf \U$9708 ( \10401 , \10400 );
buf \U$9709 ( \10402 , \10401 );
nand \U$9710 ( \10403 , \10393 , \10402 );
buf \U$9711 ( \10404 , \10403 );
buf \U$9712 ( \10405 , \10404 );
not \U$9713 ( \10406 , \7469 );
buf \U$9714 ( \10407 , \10406 );
buf \U$9715 ( \10408 , \3537 );
nor \U$9716 ( \10409 , \10407 , \10408 );
buf \U$9717 ( \10410 , \10409 );
buf \U$9718 ( \10411 , \10410 );
nand \U$9719 ( \10412 , \10405 , \10411 );
buf \U$9720 ( \10413 , \10412 );
buf \U$9721 ( \10414 , \10413 );
buf \U$9722 ( \10415 , \7416 );
not \U$9723 ( \10416 , \10415 );
buf \U$9724 ( \10417 , \10416 );
buf \U$9725 ( \10418 , \10417 );
buf \U$9728 ( \10419 , \7453 );
buf \U$9729 ( \10420 , \10419 );
and \U$9730 ( \10421 , \10418 , \10420 );
buf \U$9733 ( \10422 , \4951 );
buf \U$9734 ( \10423 , \10422 );
not \U$9735 ( \10424 , \10423 );
buf \U$9736 ( \10425 , \10424 );
buf \U$9737 ( \10426 , \10425 );
nor \U$9738 ( \10427 , \10421 , \10426 );
buf \U$9739 ( \10428 , \10427 );
buf \U$9740 ( \10429 , \10428 );
buf \U$9743 ( \10430 , \7441 );
buf \U$9744 ( \10431 , \10430 );
or \U$9745 ( \10432 , \10429 , \10431 );
buf \U$9748 ( \10433 , \4315 );
buf \U$9749 ( \10434 , \10433 );
nand \U$9750 ( \10435 , \10432 , \10434 );
buf \U$9751 ( \10436 , \10435 );
buf \U$9752 ( \10437 , \10436 );
buf \U$9753 ( \10438 , \3537 );
not \U$9754 ( \10439 , \10438 );
buf \U$9755 ( \10440 , \10439 );
buf \U$9756 ( \10441 , \10440 );
nand \U$9757 ( \10442 , \10437 , \10441 );
buf \U$9758 ( \10443 , \10442 );
buf \U$9759 ( \10444 , \10443 );
buf \U$9760 ( \10445 , \10149 );
not \U$9761 ( \10446 , \10445 );
buf \U$9762 ( \10447 , \10446 );
buf \U$9763 ( \10448 , \10447 );
nand \U$9764 ( \10449 , \10414 , \10444 , \10448 );
buf \U$9765 ( \10450 , \10449 );
buf \U$9766 ( \10451 , \10450 );
buf \U$9767 ( \10452 , \10135 );
buf \U$9768 ( \10453 , \10156 );
nand \U$9769 ( \10454 , \10452 , \10453 );
buf \U$9770 ( \10455 , \10454 );
buf \U$9771 ( \10456 , \10455 );
not \U$9772 ( \10457 , \10456 );
buf \U$9773 ( \10458 , \10457 );
buf \U$9774 ( \10459 , \10458 );
and \U$9775 ( \10460 , \10451 , \10459 );
not \U$9776 ( \10461 , \10451 );
buf \U$9777 ( \10462 , \10455 );
and \U$9778 ( \10463 , \10461 , \10462 );
nor \U$9779 ( \10464 , \10460 , \10463 );
buf \U$9780 ( \10465 , \10464 );
buf \U$9781 ( \10466 , \10465 );
buf \U$9782 ( \10467 , \10404 );
buf \U$9785 ( \10468 , \3534 );
buf \U$9786 ( \10469 , \10468 );
not \U$9787 ( \10470 , \10469 );
buf \U$9788 ( \10471 , \10406 );
nor \U$9789 ( \10472 , \10470 , \10471 );
buf \U$9790 ( \10473 , \10472 );
buf \U$9791 ( \10474 , \10473 );
nand \U$9792 ( \10475 , \10467 , \10474 );
buf \U$9793 ( \10476 , \10475 );
buf \U$9794 ( \10477 , \10476 );
buf \U$9795 ( \10478 , \10436 );
buf \U$9796 ( \10479 , \10468 );
nand \U$9797 ( \10480 , \10478 , \10479 );
buf \U$9798 ( \10481 , \10480 );
buf \U$9799 ( \10482 , \10481 );
buf \U$9800 ( \10483 , \10141 );
not \U$9801 ( \10484 , \10483 );
buf \U$9802 ( \10485 , \10484 );
buf \U$9803 ( \10486 , \10485 );
nand \U$9804 ( \10487 , \10477 , \10482 , \10486 );
buf \U$9805 ( \10488 , \10487 );
buf \U$9806 ( \10489 , \10488 );
buf \U$9807 ( \10490 , \2814 );
buf \U$9808 ( \10491 , \10148 );
nand \U$9809 ( \10492 , \10490 , \10491 );
buf \U$9810 ( \10493 , \10492 );
buf \U$9811 ( \10494 , \10493 );
not \U$9812 ( \10495 , \10494 );
buf \U$9813 ( \10496 , \10495 );
buf \U$9814 ( \10497 , \10496 );
and \U$9815 ( \10498 , \10489 , \10497 );
not \U$9816 ( \10499 , \10489 );
buf \U$9817 ( \10500 , \10493 );
and \U$9818 ( \10501 , \10499 , \10500 );
nor \U$9819 ( \10502 , \10498 , \10501 );
buf \U$9820 ( \10503 , \10502 );
buf \U$9821 ( \10504 , \10503 );
buf \U$9822 ( \10505 , \10468 );
buf \U$9823 ( \10506 , \10485 );
nand \U$9824 ( \10507 , \10505 , \10506 );
buf \U$9825 ( \10508 , \10507 );
buf \U$9826 ( \10509 , \10508 );
not \U$9827 ( \10510 , \10509 );
buf \U$9828 ( \10511 , \10122 );
buf \U$9829 ( \10512 , \10511 );
not \U$9830 ( \10513 , \10512 );
or \U$9831 ( \10514 , \10510 , \10513 );
buf \U$9832 ( \10515 , \10508 );
buf \U$9833 ( \10516 , \10511 );
or \U$9834 ( \10517 , \10515 , \10516 );
nand \U$9835 ( \10518 , \10514 , \10517 );
buf \U$9836 ( \10519 , \10518 );
buf \U$9837 ( \10520 , \10519 );
buf \U$9838 ( \10521 , \10419 );
not \U$9839 ( \10522 , \10521 );
buf \U$9840 ( \10523 , \7434 );
buf \U$9841 ( \10524 , \10523 );
nor \U$9842 ( \10525 , \10522 , \10524 );
buf \U$9843 ( \10526 , \10525 );
buf \U$9844 ( \10527 , \10526 );
not \U$9845 ( \10528 , \10527 );
buf \U$9846 ( \10529 , \10404 );
not \U$9847 ( \10530 , \10529 );
or \U$9848 ( \10531 , \10528 , \10530 );
buf \U$9850 ( \10532 , \10428 );
nand \U$9851 ( \10533 , \10531 , \10532 );
buf \U$9852 ( \10534 , \10533 );
buf \U$9853 ( \10535 , \10534 );
buf \U$9854 ( \10536 , \10430 );
not \U$9855 ( \10537 , \10536 );
buf \U$9856 ( \10538 , \10433 );
nand \U$9857 ( \10539 , \10537 , \10538 );
buf \U$9858 ( \10540 , \10539 );
buf \U$9859 ( \10541 , \10540 );
not \U$9860 ( \10542 , \10541 );
buf \U$9861 ( \10543 , \10542 );
buf \U$9862 ( \10544 , \10543 );
and \U$9863 ( \10545 , \10535 , \10544 );
not \U$9864 ( \10546 , \10535 );
buf \U$9865 ( \10547 , \10540 );
and \U$9866 ( \10548 , \10546 , \10547 );
nor \U$9867 ( \10549 , \10545 , \10548 );
buf \U$9868 ( \10550 , \10549 );
buf \U$9869 ( \10551 , \10550 );
not \U$9870 ( \10552 , \10523 );
buf \U$9871 ( \10553 , \10552 );
not \U$9872 ( \10554 , \10553 );
buf \U$9873 ( \10555 , \10404 );
not \U$9874 ( \10556 , \10555 );
or \U$9875 ( \10557 , \10554 , \10556 );
buf \U$9876 ( \10558 , \10417 );
not \U$9877 ( \10559 , \10558 );
buf \U$9878 ( \10560 , \10559 );
buf \U$9879 ( \10561 , \10560 );
nand \U$9880 ( \10562 , \10557 , \10561 );
buf \U$9881 ( \10563 , \10562 );
buf \U$9882 ( \10564 , \10563 );
buf \U$9883 ( \10565 , \10422 );
buf \U$9884 ( \10566 , \10419 );
nand \U$9885 ( \10567 , \10565 , \10566 );
buf \U$9886 ( \10568 , \10567 );
buf \U$9887 ( \10569 , \10568 );
not \U$9888 ( \10570 , \10569 );
buf \U$9889 ( \10571 , \10570 );
buf \U$9890 ( \10572 , \10571 );
and \U$9891 ( \10573 , \10564 , \10572 );
not \U$9892 ( \10574 , \10564 );
buf \U$9893 ( \10575 , \10568 );
and \U$9894 ( \10576 , \10574 , \10575 );
nor \U$9895 ( \10577 , \10573 , \10576 );
buf \U$9896 ( \10578 , \10577 );
buf \U$9897 ( \10579 , \10578 );
buf \U$9898 ( \10580 , \7432 );
not \U$9899 ( \10581 , \10580 );
buf \U$9900 ( \10582 , \10404 );
not \U$9901 ( \10583 , \10582 );
or \U$9902 ( \10584 , \10581 , \10583 );
buf \U$9903 ( \10585 , \7397 );
not \U$9904 ( \10586 , \10585 );
buf \U$9905 ( \10587 , \10586 );
buf \U$9906 ( \10588 , \10587 );
nand \U$9907 ( \10589 , \10584 , \10588 );
buf \U$9908 ( \10590 , \10589 );
buf \U$9909 ( \10591 , \10590 );
buf \U$9910 ( \10592 , \7368 );
buf \U$9911 ( \10593 , \7410 );
nand \U$9912 ( \10594 , \10592 , \10593 );
buf \U$9913 ( \10595 , \10594 );
buf \U$9914 ( \10596 , \10595 );
not \U$9915 ( \10597 , \10596 );
buf \U$9916 ( \10598 , \10597 );
buf \U$9917 ( \10599 , \10598 );
and \U$9918 ( \10600 , \10591 , \10599 );
not \U$9919 ( \10601 , \10591 );
buf \U$9920 ( \10602 , \10595 );
and \U$9921 ( \10603 , \10601 , \10602 );
nor \U$9922 ( \10604 , \10600 , \10603 );
buf \U$9923 ( \10605 , \10604 );
buf \U$9924 ( \10606 , \10605 );
buf \U$9925 ( \10607 , \10587 );
buf \U$9926 ( \10608 , \7432 );
nand \U$9927 ( \10609 , \10607 , \10608 );
buf \U$9928 ( \10610 , \10609 );
buf \U$9929 ( \10611 , \10610 );
not \U$9930 ( \10612 , \10611 );
buf \U$9931 ( \10613 , \10404 );
buf \U$9932 ( \10614 , \10613 );
not \U$9933 ( \10615 , \10614 );
or \U$9934 ( \10616 , \10612 , \10615 );
buf \U$9935 ( \10617 , \10610 );
buf \U$9936 ( \10618 , \10613 );
or \U$9937 ( \10619 , \10617 , \10618 );
nand \U$9938 ( \10620 , \10616 , \10619 );
buf \U$9939 ( \10621 , \10620 );
buf \U$9940 ( \10622 , \10621 );
buf \U$9941 ( \10623 , \7292 );
buf \U$9942 ( \10624 , \7478 );
and \U$9943 ( \10625 , \10623 , \10624 );
buf \U$9944 ( \10626 , \10625 );
buf \U$9945 ( \10627 , \10626 );
not \U$9946 ( \10628 , \10627 );
buf \U$9947 ( \10629 , \10116 );
not \U$9948 ( \10630 , \10629 );
or \U$9949 ( \10631 , \10628 , \10630 );
buf \U$9950 ( \10632 , \7277 );
buf \U$9953 ( \10633 , \7292 );
buf \U$9954 ( \10634 , \10633 );
nand \U$9955 ( \10635 , \10632 , \10634 );
buf \U$9956 ( \10636 , \10635 );
buf \U$9957 ( \10637 , \10636 );
nand \U$9958 ( \10638 , \10631 , \10637 );
buf \U$9959 ( \10639 , \10638 );
buf \U$9960 ( \10640 , \10639 );
buf \U$9963 ( \10641 , \7282 );
buf \U$9964 ( \10642 , \10641 );
and \U$9965 ( \10643 , \10640 , \10642 );
buf \U$9968 ( \10644 , \6438 );
buf \U$9969 ( \10645 , \10644 );
nor \U$9970 ( \10646 , \10643 , \10645 );
buf \U$9971 ( \10647 , \10646 );
buf \U$9972 ( \10648 , \10647 );
buf \U$9973 ( \10649 , \6027 );
buf \U$9974 ( \10650 , \6019 );
nand \U$9975 ( \10651 , \10649 , \10650 );
buf \U$9976 ( \10652 , \10651 );
buf \U$9977 ( \10653 , \10652 );
and \U$9978 ( \10654 , \10648 , \10653 );
not \U$9979 ( \10655 , \10648 );
buf \U$9980 ( \10656 , \10652 );
not \U$9981 ( \10657 , \10656 );
buf \U$9982 ( \10658 , \10657 );
buf \U$9983 ( \10659 , \10658 );
and \U$9984 ( \10660 , \10655 , \10659 );
nor \U$9985 ( \10661 , \10654 , \10660 );
buf \U$9986 ( \10662 , \10661 );
buf \U$9987 ( \10663 , \10662 );
buf \U$9988 ( \10664 , \10639 );
buf \U$9989 ( \10665 , \10644 );
not \U$9990 ( \10666 , \10665 );
buf \U$9991 ( \10667 , \10641 );
nand \U$9992 ( \10668 , \10666 , \10667 );
buf \U$9993 ( \10669 , \10668 );
buf \U$9994 ( \10670 , \10669 );
not \U$9995 ( \10671 , \10670 );
buf \U$9996 ( \10672 , \10671 );
buf \U$9997 ( \10673 , \10672 );
and \U$9998 ( \10674 , \10664 , \10673 );
not \U$9999 ( \10675 , \10664 );
buf \U$10000 ( \10676 , \10669 );
and \U$10001 ( \10677 , \10675 , \10676 );
nor \U$10002 ( \10678 , \10674 , \10677 );
buf \U$10003 ( \10679 , \10678 );
buf \U$10004 ( \10680 , \10679 );
buf \U$10007 ( \10681 , \7478 );
buf \U$10008 ( \10682 , \10681 );
not \U$10009 ( \10683 , \10682 );
buf \U$10010 ( \10684 , \10116 );
buf \U$10011 ( \10685 , \10684 );
not \U$10012 ( \10686 , \10685 );
or \U$10013 ( \10687 , \10683 , \10686 );
buf \U$10014 ( \10688 , \7258 );
nand \U$10015 ( \10689 , \10687 , \10688 );
buf \U$10016 ( \10690 , \10689 );
buf \U$10017 ( \10691 , \10690 );
buf \U$10018 ( \10692 , \7274 );
buf \U$10019 ( \10693 , \10633 );
nand \U$10020 ( \10694 , \10692 , \10693 );
buf \U$10021 ( \10695 , \10694 );
buf \U$10022 ( \10696 , \10695 );
not \U$10023 ( \10697 , \10696 );
buf \U$10024 ( \10698 , \10697 );
buf \U$10025 ( \10699 , \10698 );
and \U$10026 ( \10700 , \10691 , \10699 );
not \U$10027 ( \10701 , \10691 );
buf \U$10028 ( \10702 , \10695 );
and \U$10029 ( \10703 , \10701 , \10702 );
nor \U$10030 ( \10704 , \10700 , \10703 );
buf \U$10031 ( \10705 , \10704 );
buf \U$10032 ( \10706 , \10705 );
buf \U$10033 ( \10707 , \7258 );
buf \U$10034 ( \10708 , \10681 );
nand \U$10035 ( \10709 , \10707 , \10708 );
buf \U$10036 ( \10710 , \10709 );
not \U$10037 ( \10711 , \10684 );
xor \U$10038 ( \10712 , \10710 , \10711 );
buf \U$10039 ( \10713 , \10712 );
buf \U$10042 ( \10714 , \8541 );
buf \U$10043 ( \10715 , \10714 );
not \U$10044 ( \10716 , \10715 );
buf \U$10045 ( \10717 , \8420 );
not \U$10046 ( \10718 , \10717 );
buf \U$10047 ( \10719 , \10062 );
not \U$10048 ( \10720 , \10719 );
or \U$10049 ( \10721 , \10718 , \10720 );
buf \U$10052 ( \10722 , \10088 );
buf \U$10053 ( \10723 , \10722 );
buf \U$10054 ( \10724 , \10084 );
nand \U$10055 ( \10725 , \10723 , \10724 );
buf \U$10056 ( \10726 , \10725 );
buf \U$10057 ( \10727 , \10726 );
nand \U$10058 ( \10728 , \10721 , \10727 );
buf \U$10059 ( \10729 , \10728 );
buf \U$10060 ( \10730 , \10729 );
not \U$10061 ( \10731 , \10730 );
or \U$10062 ( \10732 , \10716 , \10731 );
buf \U$10063 ( \10733 , \10107 );
nand \U$10064 ( \10734 , \10732 , \10733 );
buf \U$10065 ( \10735 , \10734 );
buf \U$10066 ( \10736 , \10735 );
buf \U$10067 ( \10737 , \10068 );
not \U$10068 ( \10738 , \10737 );
buf \U$10069 ( \10739 , \10099 );
nand \U$10070 ( \10740 , \10738 , \10739 );
buf \U$10071 ( \10741 , \10740 );
buf \U$10072 ( \10742 , \10741 );
not \U$10073 ( \10743 , \10742 );
buf \U$10074 ( \10744 , \10743 );
buf \U$10075 ( \10745 , \10744 );
and \U$10076 ( \10746 , \10736 , \10745 );
not \U$10077 ( \10747 , \10736 );
buf \U$10078 ( \10748 , \10741 );
and \U$10079 ( \10749 , \10747 , \10748 );
nor \U$10080 ( \10750 , \10746 , \10749 );
buf \U$10081 ( \10751 , \10750 );
buf \U$10082 ( \10752 , \10751 );
buf \U$10083 ( \10753 , \10714 );
buf \U$10084 ( \10754 , \10107 );
nand \U$10085 ( \10755 , \10753 , \10754 );
buf \U$10086 ( \10756 , \10755 );
buf \U$10087 ( \10757 , \10756 );
buf \U$10088 ( \10758 , \10729 );
not \U$10089 ( \10759 , \10758 );
buf \U$10090 ( \10760 , \10759 );
buf \U$10091 ( \10761 , \10760 );
and \U$10092 ( \10762 , \10757 , \10761 );
not \U$10093 ( \10763 , \10757 );
buf \U$10094 ( \10764 , \10729 );
and \U$10095 ( \10765 , \10763 , \10764 );
nor \U$10096 ( \10766 , \10762 , \10765 );
buf \U$10097 ( \10767 , \10766 );
buf \U$10098 ( \10768 , \10767 );
buf \U$10099 ( \10769 , \8330 );
not \U$10100 ( \10770 , \10769 );
buf \U$10101 ( \10771 , \10770 );
buf \U$10102 ( \10772 , \10771 );
not \U$10103 ( \10773 , \10772 );
buf \U$10104 ( \10774 , \10062 );
not \U$10105 ( \10775 , \10774 );
or \U$10106 ( \10776 , \10773 , \10775 );
buf \U$10107 ( \10777 , \10081 );
nand \U$10108 ( \10778 , \10776 , \10777 );
buf \U$10109 ( \10779 , \10778 );
buf \U$10110 ( \10780 , \10779 );
buf \U$10111 ( \10781 , \10722 );
buf \U$10112 ( \10782 , \10076 );
nand \U$10113 ( \10783 , \10781 , \10782 );
buf \U$10114 ( \10784 , \10783 );
buf \U$10115 ( \10785 , \10784 );
not \U$10116 ( \10786 , \10785 );
buf \U$10117 ( \10787 , \10786 );
buf \U$10118 ( \10788 , \10787 );
and \U$10119 ( \10789 , \10780 , \10788 );
not \U$10120 ( \10790 , \10780 );
buf \U$10121 ( \10791 , \10784 );
and \U$10122 ( \10792 , \10790 , \10791 );
nor \U$10123 ( \10793 , \10789 , \10792 );
buf \U$10124 ( \10794 , \10793 );
buf \U$10125 ( \10795 , \10794 );
buf \U$10126 ( \10796 , \10062 );
buf \U$10127 ( \10797 , \10771 );
buf \U$10128 ( \10798 , \10081 );
nand \U$10129 ( \10799 , \10797 , \10798 );
buf \U$10130 ( \10800 , \10799 );
buf \U$10131 ( \10801 , \10800 );
not \U$10132 ( \10802 , \10801 );
buf \U$10133 ( \10803 , \10802 );
buf \U$10134 ( \10804 , \10803 );
and \U$10135 ( \10805 , \10796 , \10804 );
not \U$10136 ( \10806 , \10796 );
buf \U$10137 ( \10807 , \10800 );
and \U$10138 ( \10808 , \10806 , \10807 );
nor \U$10139 ( \10809 , \10805 , \10808 );
buf \U$10140 ( \10810 , \10809 );
buf \U$10141 ( \10811 , \10810 );
buf \U$10142 ( \10812 , \10056 );
buf \U$10143 ( \10813 , \9321 );
nand \U$10144 ( \10814 , \10812 , \10813 );
buf \U$10145 ( \10815 , \10814 );
buf \U$10146 ( \10816 , \10815 );
buf \U$10147 ( \10817 , \9282 );
buf \U$10150 ( \10818 , \10817 );
nand \U$10151 ( \10819 , \10816 , \10818 );
buf \U$10152 ( \10820 , \10819 );
buf \U$10153 ( \10821 , \10820 );
buf \U$10156 ( \10822 , \8946 );
buf \U$10157 ( \10823 , \10822 );
and \U$10158 ( \10824 , \10821 , \10823 );
buf \U$10159 ( \10825 , \9293 );
not \U$10160 ( \10826 , \10825 );
buf \U$10161 ( \10827 , \10826 );
buf \U$10162 ( \10828 , \10827 );
nor \U$10163 ( \10829 , \10824 , \10828 );
buf \U$10164 ( \10830 , \10829 );
buf \U$10165 ( \10831 , \10830 );
buf \U$10166 ( \10832 , \9302 );
not \U$10167 ( \10833 , \10832 );
buf \U$10168 ( \10834 , \8798 );
nand \U$10169 ( \10835 , \10833 , \10834 );
buf \U$10170 ( \10836 , \10835 );
buf \U$10171 ( \10837 , \10836 );
and \U$10172 ( \10838 , \10831 , \10837 );
not \U$10173 ( \10839 , \10831 );
buf \U$10174 ( \10840 , \10836 );
not \U$10175 ( \10841 , \10840 );
buf \U$10176 ( \10842 , \10841 );
buf \U$10177 ( \10843 , \10842 );
and \U$10178 ( \10844 , \10839 , \10843 );
nor \U$10179 ( \10845 , \10838 , \10844 );
buf \U$10180 ( \10846 , \10845 );
buf \U$10181 ( \10847 , \10846 );
buf \U$10182 ( \10848 , \9293 );
buf \U$10183 ( \10849 , \10822 );
and \U$10184 ( \10850 , \10848 , \10849 );
buf \U$10185 ( \10851 , \10850 );
buf \U$10186 ( \10852 , \10851 );
buf \U$10187 ( \10853 , \10820 );
and \U$10188 ( \10854 , \10852 , \10853 );
not \U$10189 ( \10855 , \10852 );
buf \U$10190 ( \10856 , \10820 );
not \U$10191 ( \10857 , \10856 );
buf \U$10192 ( \10858 , \10857 );
buf \U$10193 ( \10859 , \10858 );
and \U$10194 ( \10860 , \10855 , \10859 );
nor \U$10195 ( \10861 , \10854 , \10860 );
buf \U$10196 ( \10862 , \10861 );
buf \U$10197 ( \10863 , \10862 );
buf \U$10198 ( \10864 , \10056 );
not \U$10199 ( \10865 , \10864 );
buf \U$10200 ( \10866 , \10865 );
buf \U$10201 ( \10867 , \10866 );
not \U$10202 ( \10868 , \10867 );
buf \U$10203 ( \10869 , \10868 );
buf \U$10204 ( \10870 , \10869 );
buf \U$10207 ( \10871 , \9318 );
buf \U$10208 ( \10872 , \10871 );
and \U$10209 ( \10873 , \10870 , \10872 );
buf \U$10210 ( \10874 , \9269 );
not \U$10211 ( \10875 , \10874 );
buf \U$10212 ( \10876 , \10875 );
buf \U$10213 ( \10877 , \10876 );
nor \U$10214 ( \10878 , \10873 , \10877 );
buf \U$10215 ( \10879 , \10878 );
buf \U$10216 ( \10880 , \10879 );
buf \U$10217 ( \10881 , \9139 );
buf \U$10218 ( \10882 , \9281 );
nand \U$10219 ( \10883 , \10881 , \10882 );
buf \U$10220 ( \10884 , \10883 );
buf \U$10221 ( \10885 , \10884 );
and \U$10222 ( \10886 , \10880 , \10885 );
not \U$10223 ( \10887 , \10880 );
buf \U$10224 ( \10888 , \10884 );
not \U$10225 ( \10889 , \10888 );
buf \U$10226 ( \10890 , \10889 );
buf \U$10227 ( \10891 , \10890 );
and \U$10228 ( \10892 , \10887 , \10891 );
nor \U$10229 ( \10893 , \10886 , \10892 );
buf \U$10230 ( \10894 , \10893 );
buf \U$10231 ( \10895 , \10894 );
buf \U$10232 ( \10896 , \10866 );
buf \U$10233 ( \10897 , \10871 );
buf \U$10234 ( \10898 , \9269 );
nand \U$10235 ( \10899 , \10897 , \10898 );
buf \U$10236 ( \10900 , \10899 );
buf \U$10237 ( \10901 , \10900 );
and \U$10238 ( \10902 , \10896 , \10901 );
not \U$10239 ( \10903 , \10896 );
buf \U$10240 ( \10904 , \10900 );
not \U$10241 ( \10905 , \10904 );
buf \U$10242 ( \10906 , \10905 );
buf \U$10243 ( \10907 , \10906 );
and \U$10244 ( \10908 , \10903 , \10907 );
nor \U$10245 ( \10909 , \10902 , \10908 );
buf \U$10246 ( \10910 , \10909 );
buf \U$10247 ( \10911 , \10910 );
xor \U$10248 ( \10912 , \9415 , \9419 );
xor \U$10249 ( \10913 , \10912 , \10052 );
buf \U$10250 ( \10914 , \10913 );
buf \U$10251 ( \10915 , \10914 );
buf \U$10252 ( \10916 , \10048 );
buf \U$10253 ( \10917 , \9600 );
nand \U$10254 ( \10918 , \10916 , \10917 );
buf \U$10255 ( \10919 , \10918 );
buf \U$10256 ( \10920 , \10919 );
buf \U$10257 ( \10921 , \10035 );
not \U$10258 ( \10922 , \10921 );
buf \U$10259 ( \10923 , \10922 );
buf \U$10260 ( \10924 , \10923 );
and \U$10261 ( \10925 , \10920 , \10924 );
not \U$10262 ( \10926 , \10920 );
buf \U$10263 ( \10927 , \10035 );
and \U$10264 ( \10928 , \10926 , \10927 );
nor \U$10265 ( \10929 , \10925 , \10928 );
buf \U$10266 ( \10930 , \10929 );
buf \U$10267 ( \10931 , \10930 );
buf \U$10268 ( \10932 , \9979 );
buf \U$10269 ( \10933 , \10032 );
buf \U$10270 ( \10934 , \10019 );
nand \U$10271 ( \10935 , \10933 , \10934 );
buf \U$10272 ( \10936 , \10935 );
buf \U$10273 ( \10937 , \10936 );
xnor \U$10274 ( \10938 , \10932 , \10937 );
buf \U$10275 ( \10939 , \10938 );
buf \U$10276 ( \10940 , \10939 );
endmodule

