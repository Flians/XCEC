//
// Conformal-LEC Version 20.10-d211 (31-Aug-2020)
//
module top(RI8929640_33,RI8929dc0_49,RI8929730_35,RI8929eb0_51,RI8929fa0_53,RI8929820_37,RI8929910_39,RI892a090_55,RI8929a00_41,
        RI892a180_57,RI8929a78_42,RI892a1f8_58,RI8929af0_43,RI892a270_59,RI892a2e8_60,RI8929b68_44,RI8929d48_48,RI892a4c8_64,RI8929cd0_47,
        RI892a450_63,RI8929c58_46,RI892a3d8_62,RI8929be0_45,RI892a360_61,RI8929988_40,RI892a108_56,RI8929898_38,RI892a018_54,RI89297a8_36,
        RI8929f28_52,RI89296b8_34,RI8929e38_50,RI8928b00_9,RI89293e8_28,RI8929460_29,RI8928e48_16,RI8928ce0_13,RI8929550_31,RI89295c8_32,
        RI8928c68_12,RI8928dd0_15,RI89294d8_30,RI8928d58_14,RI8928bf0_11,RI8929370_27,RI8928b78_10,RI89292f8_26,RI8929190_23,RI8929208_24,
        RI8929280_25,RI8928a88_8,RI8928a10_7,RI8928998_6,RI8929118_22,RI8928920_5,RI89290a0_21,RI89288a8_4,RI8929028_20,RI8928fb0_19,
        RI8928830_3,RI8928f38_18,RI8928ec0_17,RI8928740_1,RI89287b8_2,R_41_7a88898,R_42_7a83a80,R_43_7a83bd0,R_44_7a87788,R_45_7a88be0,
        R_46_7a81ef0,R_47_7a889e8,R_48_7a84a40,R_49_7a882b0,R_4a_7a82c10,R_4b_7a82d60,R_4c_7a87b78,R_4d_7a84b90,R_4e_7a86f00,R_4f_7a84ce0,
        R_50_7a87440,R_51_7a88160,R_52_7a83d20,R_53_7a88c88,R_54_7a82040,R_55_7a84e30,R_56_7a876e0,R_57_7a87f68,R_58_7a82eb0,R_59_7a88dd8,
        R_5a_7a86e58,R_5b_7a83e70);
input RI8929640_33,RI8929dc0_49,RI8929730_35,RI8929eb0_51,RI8929fa0_53,RI8929820_37,RI8929910_39,RI892a090_55,RI8929a00_41,
        RI892a180_57,RI8929a78_42,RI892a1f8_58,RI8929af0_43,RI892a270_59,RI892a2e8_60,RI8929b68_44,RI8929d48_48,RI892a4c8_64,RI8929cd0_47,
        RI892a450_63,RI8929c58_46,RI892a3d8_62,RI8929be0_45,RI892a360_61,RI8929988_40,RI892a108_56,RI8929898_38,RI892a018_54,RI89297a8_36,
        RI8929f28_52,RI89296b8_34,RI8929e38_50,RI8928b00_9,RI89293e8_28,RI8929460_29,RI8928e48_16,RI8928ce0_13,RI8929550_31,RI89295c8_32,
        RI8928c68_12,RI8928dd0_15,RI89294d8_30,RI8928d58_14,RI8928bf0_11,RI8929370_27,RI8928b78_10,RI89292f8_26,RI8929190_23,RI8929208_24,
        RI8929280_25,RI8928a88_8,RI8928a10_7,RI8928998_6,RI8929118_22,RI8928920_5,RI89290a0_21,RI89288a8_4,RI8929028_20,RI8928fb0_19,
        RI8928830_3,RI8928f38_18,RI8928ec0_17,RI8928740_1,RI89287b8_2;
output R_41_7a88898,R_42_7a83a80,R_43_7a83bd0,R_44_7a87788,R_45_7a88be0,R_46_7a81ef0,R_47_7a889e8,R_48_7a84a40,R_49_7a882b0,
        R_4a_7a82c10,R_4b_7a82d60,R_4c_7a87b78,R_4d_7a84b90,R_4e_7a86f00,R_4f_7a84ce0,R_50_7a87440,R_51_7a88160,R_52_7a83d20,R_53_7a88c88,
        R_54_7a82040,R_55_7a84e30,R_56_7a876e0,R_57_7a87f68,R_58_7a82eb0,R_59_7a88dd8,R_5a_7a86e58,R_5b_7a83e70;

wire \92_ZERO , \93_ONE , \94 , \95 , \96 , \97 , \98 , \99 , \100 ,
         \101 , \102 , \103 , \104 , \105 , \106 , \107 , \108 , \109 , \110 ,
         \111 , \112 , \113 , \114 , \115 , \116 , \117 , \118 , \119 , \120 ,
         \121 , \122 , \123 , \124 , \125 , \126 , \127 , \128 , \129 , \130 ,
         \131 , \132 , \133 , \134 , \135 , \136 , \137 , \138 , \139 , \140 ,
         \141 , \142 , \143 , \144 , \145 , \146 , \147 , \148 , \149 , \150 ,
         \151 , \152 , \153 , \154 , \155 , \156 , \157 , \158 , \159 , \160 ,
         \161 , \162 , \163 , \164 , \165 , \166 , \167 , \168 , \169 , \170 ,
         \171 , \172 , \173 , \174 , \175 , \176 , \177 , \178 , \179 , \180 ,
         \181 , \182 , \183 , \184 , \185 , \186 , \187 , \188 , \189 , \190 ,
         \191 , \192 , \193 , \194 , \195 , \196 , \197 , \198 , \199 , \200 ,
         \201 , \202 , \203 , \204 , \205 , \206 , \207 , \208 , \209 , \210 ,
         \211 , \212 , \213 , \214 , \215 , \216 , \217 , \218 , \219 , \220 ,
         \221 , \222 , \223 , \224 , \225 , \226 , \227 , \228 , \229 , \230 ,
         \231 , \232 , \233 , \234 , \235 , \236 , \237 , \238 , \239 , \240 ,
         \241 , \242 , \243 , \244 , \245 , \246 , \247 , \248 , \249 , \250 ,
         \251 , \252 , \253 , \254 , \255 , \256 , \257 , \258 , \259 , \260 ,
         \261 , \262 , \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 ,
         \271 , \272 , \273 , \274 , \275 , \276 , \277 , \278 , \279 , \280 ,
         \281 , \282 , \283 , \284 , \285 , \286 , \287 , \288 , \289 , \290 ,
         \291 , \292 , \293 , \294 , \295 , \296 , \297 , \298 , \299 , \300 ,
         \301 , \302 , \303 , \304 , \305 , \306 , \307 , \308 , \309 , \310 ,
         \311 , \312 , \313 , \314 , \315 , \316 , \317 , \318 , \319 , \320 ,
         \321 , \322 , \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 ,
         \331 , \332 , \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 ,
         \341 , \342 , \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 ,
         \351 , \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 ,
         \361 , \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 ,
         \371 , \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 ,
         \381 , \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 ,
         \391 , \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 ,
         \401 , \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 ,
         \411 , \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 ,
         \421 , \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 ,
         \431 , \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 ,
         \441 , \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 ,
         \451 , \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 ,
         \461 , \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 ,
         \471 , \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 ,
         \481 , \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 ,
         \491 , \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 ,
         \501 , \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 ,
         \511 , \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 ,
         \521 , \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 ,
         \531 , \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 ,
         \541 , \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 ,
         \551 , \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 ,
         \561 , \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 ,
         \571 , \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 ,
         \581 , \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 ,
         \591 , \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 ,
         \601 , \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 ,
         \611 , \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 ,
         \621 , \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 ,
         \631 , \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 ,
         \641 , \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 ,
         \651 , \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 ,
         \661 , \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 ,
         \671 , \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 ,
         \681 , \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 ,
         \691 , \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 ,
         \701 , \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 ,
         \711 , \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 ,
         \721 , \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 ,
         \731 , \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 ,
         \741 , \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 ,
         \751 , \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 ,
         \761 , \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 ,
         \771 , \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 ,
         \781 , \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 ,
         \791 , \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 ,
         \801 , \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 ,
         \811 , \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 ,
         \821 , \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 ,
         \831 , \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 ,
         \841 , \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 ,
         \851 , \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 ,
         \861 , \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 ,
         \871 , \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 ,
         \881 , \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 ,
         \891 , \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 ,
         \901 , \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 ,
         \911 , \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 ,
         \921 , \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 ,
         \931 , \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 ,
         \941 , \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 ,
         \951 , \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 ,
         \961 , \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 ,
         \971 , \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 ,
         \981 , \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 ,
         \991 , \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 ,
         \1001 , \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 ,
         \1011 , \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 ,
         \1021 , \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 ,
         \1031 , \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 ,
         \1041 , \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 ,
         \1051 , \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 ,
         \1061 , \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 ,
         \1071 , \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 ,
         \1081 , \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 ,
         \1091 , \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 ,
         \1101 , \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 ,
         \1111 , \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 ,
         \1121 , \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 ,
         \1131 , \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 ,
         \1141 , \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 ,
         \1151 , \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 ,
         \1161 , \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 ,
         \1171 , \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 ,
         \1181 , \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 ,
         \1191 , \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 ,
         \1201 , \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 ,
         \1211 , \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 ,
         \1221 , \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 ,
         \1231 , \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 ,
         \1241 , \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 ,
         \1251 , \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 ,
         \1261 , \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 ,
         \1271 , \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 ,
         \1281 , \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 ,
         \1291 , \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 ,
         \1301 , \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 ,
         \1311 , \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 ,
         \1321 , \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 ,
         \1331 , \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 ,
         \1341 , \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 ,
         \1351 , \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 ,
         \1361 , \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 ,
         \1371 , \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 ,
         \1381 , \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 ,
         \1391 , \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 ,
         \1401 , \1402 , \1403 , \1404 , \1405 , \1406 , \1407 , \1408 , \1409 , \1410 ,
         \1411 , \1412 , \1413 , \1414 , \1415 , \1416 , \1417 , \1418 , \1419 , \1420 ,
         \1421 , \1422 , \1423 , \1424 , \1425 , \1426 , \1427 , \1428 , \1429 , \1430 ,
         \1431 , \1432 , \1433 , \1434 , \1435 , \1436 , \1437 , \1438 , \1439 , \1440 ,
         \1441 , \1442 , \1443 , \1444 , \1445 , \1446 , \1447 , \1448 , \1449 , \1450 ,
         \1451 , \1452 , \1453 , \1454 , \1455 , \1456 , \1457 , \1458 , \1459 , \1460 ,
         \1461 , \1462 , \1463 , \1464 , \1465 , \1466 , \1467 , \1468 , \1469 , \1470 ,
         \1471 , \1472 , \1473 , \1474 , \1475 , \1476 , \1477 , \1478 , \1479 , \1480 ,
         \1481 , \1482 , \1483 , \1484 , \1485 , \1486 , \1487 , \1488 , \1489 , \1490 ,
         \1491 , \1492 , \1493 , \1494 , \1495 , \1496 , \1497 , \1498 , \1499 , \1500 ,
         \1501 , \1502 , \1503 , \1504 , \1505 , \1506 , \1507 , \1508 , \1509 , \1510 ,
         \1511 , \1512 , \1513 , \1514 , \1515 , \1516 , \1517 , \1518 , \1519 , \1520 ,
         \1521 , \1522 , \1523 , \1524 , \1525 , \1526 , \1527 , \1528 , \1529 , \1530 ,
         \1531 , \1532 , \1533 , \1534 , \1535 , \1536 , \1537 , \1538 , \1539 , \1540 ,
         \1541 , \1542 , \1543 , \1544 , \1545 , \1546 , \1547 , \1548 , \1549 , \1550 ,
         \1551 , \1552 , \1553 , \1554 , \1555 , \1556 , \1557 , \1558 , \1559 , \1560 ,
         \1561 , \1562 , \1563 , \1564 , \1565 , \1566 , \1567 , \1568 , \1569 , \1570 ,
         \1571 , \1572 , \1573 , \1574 , \1575 , \1576 , \1577 , \1578 , \1579 , \1580 ,
         \1581 , \1582 , \1583 , \1584 , \1585 , \1586 , \1587 , \1588 , \1589 , \1590 ,
         \1591 , \1592 , \1593 , \1594 , \1595 , \1596 , \1597 , \1598 , \1599 , \1600 ,
         \1601 , \1602 , \1603 , \1604 , \1605 , \1606 , \1607 , \1608 , \1609 , \1610 ,
         \1611 , \1612 , \1613 , \1614 , \1615 , \1616 , \1617 , \1618 , \1619 , \1620 ,
         \1621 , \1622 , \1623 , \1624 , \1625 , \1626 , \1627 , \1628 , \1629 , \1630 ,
         \1631 , \1632 , \1633 , \1634 , \1635 , \1636 , \1637 , \1638 , \1639 , \1640 ,
         \1641 , \1642 , \1643 , \1644 , \1645 , \1646 , \1647 , \1648 , \1649 , \1650 ,
         \1651 , \1652 , \1653 , \1654 , \1655 , \1656 , \1657 , \1658 , \1659 , \1660 ,
         \1661 , \1662 , \1663 , \1664 , \1665 , \1666 , \1667 , \1668 , \1669 , \1670 ,
         \1671 , \1672 , \1673 , \1674 , \1675 , \1676 , \1677 , \1678 , \1679 , \1680 ,
         \1681 , \1682 , \1683 , \1684 , \1685 , \1686 , \1687 , \1688 , \1689 , \1690 ,
         \1691 , \1692 , \1693 , \1694 , \1695 , \1696 , \1697 , \1698 , \1699 , \1700 ,
         \1701 , \1702 , \1703 , \1704 , \1705 , \1706 , \1707 , \1708 , \1709 , \1710 ,
         \1711 , \1712 , \1713 , \1714 , \1715 , \1716 , \1717 , \1718 , \1719 , \1720 ,
         \1721 , \1722 , \1723 , \1724 , \1725 , \1726 , \1727 , \1728 , \1729 , \1730 ,
         \1731 , \1732 , \1733 , \1734 , \1735 , \1736 , \1737 , \1738 , \1739 , \1740 ,
         \1741 , \1742 , \1743 , \1744 , \1745 , \1746 , \1747 , \1748 , \1749 , \1750 ,
         \1751 , \1752 , \1753 , \1754 , \1755 , \1756 , \1757 , \1758 , \1759 , \1760 ,
         \1761 , \1762 , \1763 , \1764 , \1765 , \1766 , \1767 , \1768 , \1769 , \1770 ,
         \1771 , \1772 , \1773 , \1774 , \1775 , \1776 , \1777 , \1778 , \1779 , \1780 ,
         \1781 , \1782 , \1783 , \1784 , \1785 , \1786 , \1787 , \1788 , \1789 , \1790 ,
         \1791 , \1792 , \1793 , \1794 , \1795 , \1796 , \1797 , \1798 , \1799 , \1800 ,
         \1801 , \1802 , \1803 , \1804 , \1805 , \1806 , \1807 , \1808 , \1809 , \1810 ,
         \1811 , \1812 , \1813 , \1814 , \1815 , \1816 , \1817 , \1818 , \1819 , \1820 ,
         \1821 , \1822 , \1823 , \1824 , \1825 , \1826 , \1827 , \1828 , \1829 , \1830 ,
         \1831 , \1832 , \1833 , \1834 , \1835 , \1836 , \1837 , \1838 , \1839 , \1840 ,
         \1841 , \1842 , \1843 , \1844 , \1845 , \1846 , \1847 , \1848 , \1849 , \1850 ,
         \1851 , \1852 , \1853 , \1854 , \1855 , \1856 , \1857 , \1858 , \1859 , \1860 ,
         \1861 , \1862 , \1863 , \1864 , \1865 , \1866 , \1867 , \1868 , \1869 , \1870 ,
         \1871 , \1872 , \1873 , \1874 , \1875 , \1876 , \1877 , \1878 , \1879 , \1880 ,
         \1881 , \1882 , \1883 , \1884 , \1885 , \1886 , \1887 , \1888 , \1889 , \1890 ,
         \1891 , \1892 , \1893 , \1894 , \1895 , \1896 , \1897 , \1898 , \1899 , \1900 ,
         \1901 , \1902 , \1903 , \1904 , \1905 , \1906 , \1907 , \1908 , \1909 , \1910 ,
         \1911 , \1912 , \1913 , \1914 , \1915 , \1916 , \1917 , \1918 , \1919 , \1920 ,
         \1921 , \1922 , \1923 , \1924 , \1925 , \1926 , \1927 , \1928 , \1929 , \1930 ,
         \1931 , \1932 , \1933 , \1934 , \1935 , \1936 , \1937 , \1938 , \1939 , \1940 ,
         \1941 , \1942 , \1943 , \1944 , \1945 , \1946 , \1947 , \1948 , \1949 , \1950 ,
         \1951 , \1952 , \1953 , \1954 , \1955 , \1956 , \1957 , \1958 , \1959 , \1960 ,
         \1961 , \1962 , \1963 , \1964 , \1965 , \1966 , \1967 , \1968 , \1969 , \1970 ,
         \1971 , \1972 , \1973 , \1974 , \1975 , \1976 , \1977 , \1978 , \1979 , \1980 ,
         \1981 , \1982 , \1983 , \1984 , \1985 , \1986 , \1987 , \1988 , \1989 , \1990 ,
         \1991 , \1992 , \1993 , \1994 , \1995 , \1996 , \1997 , \1998 , \1999 , \2000 ,
         \2001 , \2002 , \2003 , \2004 , \2005 , \2006 , \2007 , \2008 , \2009 , \2010 ,
         \2011 , \2012 , \2013 , \2014 , \2015 , \2016 , \2017 , \2018 , \2019 , \2020 ,
         \2021 , \2022 , \2023 , \2024 , \2025 , \2026 , \2027 , \2028 , \2029 , \2030 ,
         \2031 , \2032 , \2033 , \2034 , \2035 , \2036 , \2037 , \2038 , \2039 , \2040 ,
         \2041 , \2042 , \2043 , \2044 , \2045 , \2046 , \2047 , \2048 , \2049 , \2050 ,
         \2051 , \2052 , \2053 , \2054 , \2055 , \2056 , \2057 , \2058 , \2059 , \2060 ,
         \2061 , \2062 , \2063 , \2064 , \2065 , \2066 , \2067 , \2068 , \2069 , \2070 ,
         \2071 , \2072 , \2073 , \2074 , \2075 , \2076 , \2077 , \2078 , \2079 , \2080 ,
         \2081 , \2082 , \2083 , \2084 , \2085 , \2086 , \2087 , \2088 , \2089 , \2090 ,
         \2091 , \2092 , \2093 , \2094 , \2095 , \2096 , \2097 , \2098 , \2099 , \2100 ,
         \2101 , \2102 , \2103 , \2104 , \2105 , \2106 , \2107 , \2108 , \2109 , \2110 ,
         \2111 , \2112 , \2113 , \2114 , \2115 , \2116 , \2117 , \2118 , \2119 , \2120 ,
         \2121 , \2122 , \2123 , \2124 , \2125 , \2126 , \2127 , \2128 , \2129 , \2130 ,
         \2131 , \2132 , \2133 , \2134 , \2135 , \2136 , \2137 , \2138 , \2139 , \2140 ,
         \2141 , \2142 , \2143 , \2144 , \2145 , \2146 , \2147 , \2148 , \2149 , \2150 ,
         \2151 , \2152 , \2153 , \2154 , \2155 , \2156 , \2157 , \2158 , \2159 , \2160 ,
         \2161 , \2162 , \2163 , \2164 , \2165 , \2166 , \2167 , \2168 , \2169 , \2170 ,
         \2171 , \2172 , \2173 , \2174 , \2175 , \2176 , \2177 , \2178 , \2179 , \2180 ,
         \2181 , \2182 , \2183 , \2184 , \2185 , \2186 , \2187 , \2188 , \2189 , \2190 ,
         \2191 , \2192 , \2193 , \2194 , \2195 , \2196 , \2197 , \2198 , \2199 , \2200 ,
         \2201 , \2202 , \2203 , \2204 , \2205 , \2206 , \2207 , \2208 , \2209 , \2210 ,
         \2211 , \2212 , \2213 , \2214 , \2215 , \2216 , \2217 , \2218 , \2219 , \2220 ,
         \2221 , \2222 , \2223 , \2224 , \2225 , \2226 , \2227 , \2228 , \2229 , \2230 ,
         \2231 , \2232 , \2233 , \2234 , \2235 , \2236 , \2237 , \2238 , \2239 , \2240 ,
         \2241 , \2242 , \2243 , \2244 , \2245 , \2246 , \2247 , \2248 , \2249 , \2250 ,
         \2251 , \2252 , \2253 , \2254 , \2255 , \2256 , \2257 , \2258 , \2259 , \2260 ,
         \2261 , \2262 , \2263 , \2264 , \2265 , \2266 , \2267 , \2268 , \2269 , \2270 ,
         \2271 , \2272 , \2273 , \2274 , \2275 , \2276 , \2277 , \2278 , \2279 , \2280 ,
         \2281 , \2282 , \2283 , \2284 , \2285 , \2286 , \2287 , \2288 , \2289 , \2290 ,
         \2291 , \2292 , \2293 , \2294 , \2295 , \2296 , \2297 , \2298 , \2299 , \2300 ,
         \2301 , \2302 , \2303 , \2304 , \2305 , \2306 , \2307 , \2308 , \2309 , \2310 ,
         \2311 , \2312 , \2313 , \2314 , \2315 , \2316 , \2317 , \2318 , \2319 , \2320 ,
         \2321 , \2322 , \2323 , \2324 , \2325 , \2326 , \2327 , \2328 , \2329 , \2330 ,
         \2331 , \2332 , \2333 , \2334 , \2335 , \2336 , \2337 , \2338 , \2339 , \2340 ,
         \2341 , \2342 , \2343 , \2344 , \2345 , \2346 , \2347 , \2348 , \2349 , \2350 ,
         \2351 , \2352 , \2353 , \2354 , \2355 , \2356 , \2357 , \2358 , \2359 , \2360 ,
         \2361 , \2362 , \2363 , \2364 , \2365 , \2366 , \2367 , \2368 , \2369 , \2370 ,
         \2371 , \2372 , \2373 , \2374 , \2375 , \2376 , \2377 , \2378 , \2379 , \2380 ,
         \2381 , \2382 , \2383 , \2384 , \2385 , \2386 , \2387 , \2388 , \2389 , \2390 ,
         \2391 , \2392 , \2393 , \2394 , \2395 , \2396 , \2397 , \2398 , \2399 , \2400 ,
         \2401 , \2402 , \2403 , \2404 , \2405 , \2406 , \2407 , \2408 , \2409 , \2410 ,
         \2411 , \2412 , \2413 , \2414 , \2415 , \2416 , \2417 , \2418 , \2419 , \2420 ,
         \2421 , \2422 , \2423 , \2424 , \2425 , \2426 , \2427 , \2428 , \2429 , \2430 ,
         \2431 , \2432 , \2433 , \2434 , \2435 , \2436 , \2437 , \2438 , \2439 , \2440 ,
         \2441 , \2442 , \2443 , \2444 , \2445 , \2446 , \2447 , \2448 , \2449 , \2450 ,
         \2451 , \2452 , \2453 , \2454 , \2455 , \2456 , \2457 , \2458 , \2459 , \2460 ,
         \2461 , \2462 , \2463 , \2464 , \2465 , \2466 , \2467 , \2468 , \2469 , \2470 ,
         \2471 , \2472 , \2473 , \2474 , \2475 , \2476 , \2477 , \2478 , \2479 , \2480 ,
         \2481 , \2482 , \2483 , \2484 , \2485 , \2486 , \2487 , \2488 , \2489 , \2490 ,
         \2491 , \2492 , \2493 , \2494 , \2495 , \2496 , \2497 , \2498 , \2499 , \2500 ,
         \2501 , \2502 , \2503 , \2504 , \2505 , \2506 , \2507 , \2508 , \2509 , \2510 ,
         \2511 , \2512 , \2513 , \2514 , \2515 , \2516 , \2517 , \2518 , \2519 , \2520 ,
         \2521 , \2522 , \2523 , \2524 , \2525 , \2526 , \2527 , \2528 , \2529 , \2530 ,
         \2531 , \2532 , \2533 , \2534 , \2535 , \2536 , \2537 , \2538 , \2539 , \2540 ,
         \2541 , \2542 , \2543 , \2544 , \2545 , \2546 , \2547 , \2548 , \2549 , \2550 ,
         \2551 , \2552 , \2553 , \2554 , \2555 , \2556 , \2557 , \2558 , \2559 , \2560 ,
         \2561 , \2562 , \2563 , \2564 , \2565 , \2566 , \2567 , \2568 , \2569 , \2570 ,
         \2571 , \2572 , \2573 , \2574 , \2575 , \2576 , \2577 , \2578 , \2579 , \2580 ,
         \2581 , \2582 , \2583 , \2584 , \2585 , \2586 , \2587 , \2588 , \2589 , \2590 ,
         \2591 , \2592 , \2593 , \2594 , \2595 , \2596 , \2597 , \2598 , \2599 , \2600 ,
         \2601 , \2602 , \2603 , \2604 , \2605 , \2606 , \2607 , \2608 , \2609 , \2610 ,
         \2611 , \2612 , \2613 , \2614 , \2615 , \2616 , \2617 , \2618 , \2619 , \2620 ,
         \2621 , \2622 , \2623 , \2624 , \2625 , \2626 , \2627 , \2628 , \2629 , \2630 ,
         \2631 , \2632 , \2633 , \2634 , \2635 , \2636 , \2637 , \2638 , \2639 , \2640 ,
         \2641 , \2642 , \2643 , \2644 , \2645 , \2646 , \2647 , \2648 , \2649 , \2650 ,
         \2651 , \2652 , \2653 , \2654 , \2655 , \2656 , \2657 , \2658 , \2659 , \2660 ,
         \2661 , \2662 , \2663 , \2664 , \2665 , \2666 , \2667 , \2668 , \2669 , \2670 ,
         \2671 , \2672 , \2673 , \2674 , \2675 , \2676 , \2677 , \2678 , \2679 , \2680 ,
         \2681 , \2682 , \2683 , \2684 , \2685 , \2686 , \2687 , \2688 , \2689 , \2690 ,
         \2691 , \2692 , \2693 , \2694 , \2695 , \2696 , \2697 , \2698 , \2699 , \2700 ,
         \2701 , \2702 , \2703 , \2704 , \2705 , \2706 , \2707 , \2708 , \2709 , \2710 ,
         \2711 , \2712 , \2713 , \2714 , \2715 , \2716 , \2717 , \2718 , \2719 , \2720 ,
         \2721 , \2722 , \2723 , \2724 , \2725 , \2726 , \2727 , \2728 , \2729 , \2730 ,
         \2731 , \2732 , \2733 , \2734 , \2735 , \2736 , \2737 , \2738 , \2739 , \2740 ,
         \2741 , \2742 , \2743 , \2744 , \2745 , \2746 , \2747 , \2748 , \2749 , \2750 ,
         \2751 , \2752 , \2753 , \2754 , \2755 , \2756 , \2757 , \2758 , \2759 , \2760 ,
         \2761 , \2762 , \2763 , \2764 , \2765 , \2766 , \2767 , \2768 , \2769 , \2770 ,
         \2771 , \2772 , \2773 , \2774 , \2775 , \2776 , \2777 , \2778 , \2779 , \2780 ,
         \2781 , \2782 , \2783 , \2784 , \2785 , \2786 , \2787 , \2788 , \2789 , \2790 ,
         \2791 , \2792 , \2793 , \2794 , \2795 , \2796 , \2797 , \2798 , \2799 , \2800 ,
         \2801 , \2802 , \2803 , \2804 , \2805 , \2806 , \2807 , \2808 , \2809 , \2810 ,
         \2811 , \2812 , \2813 , \2814 , \2815 , \2816 , \2817 , \2818 , \2819 , \2820 ,
         \2821 , \2822 , \2823 , \2824 , \2825 , \2826 , \2827 , \2828 , \2829 , \2830 ,
         \2831 , \2832 , \2833 , \2834 , \2835 , \2836 , \2837 , \2838 , \2839 , \2840 ,
         \2841 , \2842 , \2843 , \2844 , \2845 , \2846 , \2847 , \2848 , \2849 , \2850 ,
         \2851 , \2852 , \2853 , \2854 , \2855 , \2856 , \2857 , \2858 , \2859 , \2860 ,
         \2861 , \2862 , \2863 , \2864 , \2865 , \2866 , \2867 , \2868 , \2869 , \2870 ,
         \2871 , \2872 , \2873 , \2874 , \2875 , \2876 , \2877 , \2878 , \2879 , \2880 ,
         \2881 , \2882 , \2883 , \2884 , \2885 , \2886 , \2887 , \2888 , \2889 , \2890 ,
         \2891 , \2892 , \2893 , \2894 , \2895 , \2896 , \2897 , \2898 , \2899 , \2900 ,
         \2901 , \2902 , \2903 , \2904 , \2905 , \2906 , \2907 , \2908 , \2909 , \2910 ,
         \2911 , \2912 , \2913 , \2914 , \2915 , \2916 , \2917 , \2918 , \2919 , \2920 ,
         \2921 , \2922 , \2923 , \2924 , \2925 , \2926 , \2927 , \2928 , \2929 , \2930 ,
         \2931 , \2932 , \2933 , \2934 , \2935 , \2936 , \2937 , \2938 , \2939 , \2940 ,
         \2941 , \2942 , \2943 , \2944 , \2945 , \2946 , \2947 , \2948 , \2949 , \2950 ,
         \2951 , \2952 , \2953 , \2954 , \2955 , \2956 , \2957 , \2958 , \2959 , \2960 ,
         \2961 , \2962 , \2963 , \2964 , \2965 , \2966 , \2967 , \2968 , \2969 , \2970 ,
         \2971 , \2972 , \2973 , \2974 , \2975 , \2976 , \2977 , \2978 , \2979 , \2980 ,
         \2981 , \2982 , \2983 , \2984 , \2985 , \2986 , \2987 , \2988 , \2989 , \2990 ,
         \2991 , \2992 , \2993 , \2994 , \2995 , \2996 , \2997 , \2998 , \2999 , \3000 ,
         \3001 , \3002 , \3003 , \3004 , \3005 , \3006 , \3007 , \3008 , \3009 , \3010 ,
         \3011 , \3012 , \3013 , \3014 , \3015 , \3016 , \3017 , \3018 , \3019 , \3020 ,
         \3021 , \3022 , \3023 , \3024 , \3025 , \3026 , \3027 , \3028 , \3029 , \3030 ,
         \3031 , \3032 , \3033 , \3034 , \3035 , \3036 , \3037 , \3038 , \3039 , \3040 ,
         \3041 , \3042 , \3043 , \3044 , \3045 , \3046 , \3047 , \3048 , \3049 , \3050 ,
         \3051 , \3052 , \3053 , \3054 , \3055 , \3056 , \3057 , \3058 , \3059 , \3060 ,
         \3061 , \3062 , \3063 , \3064 , \3065 , \3066 , \3067 , \3068 , \3069 , \3070 ,
         \3071 , \3072 , \3073 , \3074 , \3075 , \3076 , \3077 , \3078 , \3079 , \3080 ,
         \3081 , \3082 , \3083 , \3084 , \3085 , \3086 , \3087 , \3088 , \3089 , \3090 ,
         \3091 , \3092 , \3093 , \3094 , \3095 , \3096 , \3097 , \3098 , \3099 , \3100 ,
         \3101 , \3102 , \3103 , \3104 , \3105 , \3106 , \3107 , \3108 , \3109 , \3110 ,
         \3111 , \3112 , \3113 , \3114 , \3115 , \3116 , \3117 , \3118 , \3119 , \3120 ,
         \3121 , \3122 , \3123 , \3124 , \3125 , \3126 , \3127 , \3128 , \3129 , \3130 ,
         \3131 , \3132 , \3133 , \3134 , \3135 , \3136 , \3137 , \3138 , \3139 , \3140 ,
         \3141 , \3142 , \3143 , \3144 , \3145 , \3146 , \3147 , \3148 , \3149 , \3150 ,
         \3151 , \3152 , \3153 , \3154 , \3155 , \3156 , \3157 , \3158 , \3159 , \3160 ,
         \3161 , \3162 , \3163 , \3164 , \3165 , \3166 , \3167 , \3168 , \3169 , \3170 ,
         \3171 , \3172 , \3173 , \3174 , \3175 , \3176 , \3177 , \3178 , \3179 , \3180 ,
         \3181 , \3182 , \3183 , \3184 , \3185 , \3186 , \3187 , \3188 , \3189 , \3190 ,
         \3191 , \3192 , \3193 , \3194 , \3195 , \3196 , \3197 , \3198 , \3199 , \3200 ,
         \3201 , \3202 , \3203 , \3204 , \3205 , \3206 , \3207 , \3208 , \3209 , \3210 ,
         \3211 , \3212 , \3213 , \3214 , \3215 , \3216 , \3217 , \3218 , \3219 , \3220 ,
         \3221 , \3222 , \3223 , \3224 , \3225 , \3226 , \3227 , \3228 , \3229 , \3230 ,
         \3231 , \3232 , \3233 , \3234 , \3235 , \3236 , \3237 , \3238 , \3239 , \3240 ,
         \3241 , \3242 , \3243 , \3244 , \3245 , \3246 , \3247 , \3248 , \3249 , \3250 ,
         \3251 , \3252 , \3253 , \3254 , \3255 , \3256 , \3257 , \3258 , \3259 , \3260 ,
         \3261 , \3262 , \3263 , \3264 , \3265 , \3266 , \3267 , \3268 , \3269 , \3270 ,
         \3271 , \3272 , \3273 , \3274 , \3275 , \3276 , \3277 , \3278 , \3279 , \3280 ,
         \3281 , \3282 , \3283 , \3284 , \3285 , \3286 , \3287 , \3288 , \3289 , \3290 ,
         \3291 , \3292 , \3293 , \3294 , \3295 , \3296 , \3297 , \3298 , \3299 , \3300 ,
         \3301 , \3302 , \3303 , \3304 , \3305 , \3306 , \3307 , \3308 , \3309 , \3310 ,
         \3311 , \3312 , \3313 , \3314 , \3315 , \3316 , \3317 , \3318 , \3319 , \3320 ,
         \3321 , \3322 , \3323 , \3324 , \3325 , \3326 , \3327 , \3328 , \3329 , \3330 ,
         \3331 , \3332 , \3333 , \3334 , \3335 , \3336 , \3337 , \3338 , \3339 , \3340 ,
         \3341 , \3342 , \3343 , \3344 , \3345 , \3346 , \3347 , \3348 , \3349 , \3350 ,
         \3351 , \3352 , \3353 , \3354 , \3355 , \3356 , \3357 , \3358 , \3359 , \3360 ,
         \3361 , \3362 , \3363 , \3364 , \3365 , \3366 , \3367 , \3368 , \3369 , \3370 ,
         \3371 , \3372 , \3373 , \3374 , \3375 , \3376 , \3377 , \3378 , \3379 , \3380 ,
         \3381 , \3382 , \3383 , \3384 , \3385 , \3386 , \3387 , \3388 , \3389 , \3390 ,
         \3391 , \3392 , \3393 , \3394 , \3395 , \3396 , \3397 , \3398 , \3399 , \3400 ,
         \3401 , \3402 , \3403 , \3404 , \3405 , \3406 , \3407 , \3408 , \3409 , \3410 ,
         \3411 , \3412 , \3413 , \3414 , \3415 , \3416 , \3417 , \3418 , \3419 , \3420 ,
         \3421 , \3422 , \3423 , \3424 , \3425 , \3426 , \3427 , \3428 , \3429 , \3430 ,
         \3431 , \3432 , \3433 , \3434 , \3435 , \3436 , \3437 , \3438 , \3439 , \3440 ,
         \3441 , \3442 , \3443 , \3444 , \3445 , \3446 , \3447 , \3448 , \3449 , \3450 ,
         \3451 , \3452 , \3453 , \3454 , \3455 , \3456 , \3457 , \3458 , \3459 , \3460 ,
         \3461 , \3462 , \3463 , \3464 , \3465 , \3466 , \3467 , \3468 , \3469 , \3470 ,
         \3471 , \3472 , \3473 , \3474 , \3475 , \3476 , \3477 , \3478 , \3479 , \3480 ,
         \3481 , \3482 , \3483 , \3484 , \3485 , \3486 , \3487 , \3488 , \3489 , \3490 ,
         \3491 , \3492 , \3493 , \3494 , \3495 , \3496 , \3497 , \3498 , \3499 , \3500 ,
         \3501 , \3502 , \3503 , \3504 , \3505 , \3506 , \3507 , \3508 , \3509 , \3510 ,
         \3511 , \3512 , \3513 , \3514 , \3515 , \3516 , \3517 , \3518 , \3519 , \3520 ,
         \3521 , \3522 , \3523 , \3524 , \3525 , \3526 , \3527 , \3528 , \3529 , \3530 ,
         \3531 , \3532 , \3533 , \3534 , \3535 , \3536 , \3537 , \3538 , \3539 , \3540 ,
         \3541 , \3542 , \3543 , \3544 , \3545 , \3546 , \3547 , \3548 , \3549 , \3550 ,
         \3551 , \3552 , \3553 , \3554 , \3555 , \3556 , \3557 , \3558 , \3559 , \3560 ,
         \3561 , \3562 , \3563 , \3564 , \3565 , \3566 , \3567 , \3568 , \3569 , \3570 ,
         \3571 , \3572 , \3573 , \3574 , \3575 , \3576 , \3577 , \3578 , \3579 , \3580 ,
         \3581 , \3582 , \3583 , \3584 , \3585 , \3586 , \3587 , \3588 , \3589 , \3590 ,
         \3591 , \3592 , \3593 , \3594 , \3595 , \3596 , \3597 , \3598 , \3599 , \3600 ,
         \3601 , \3602 , \3603 , \3604 , \3605 , \3606 , \3607 , \3608 , \3609 , \3610 ,
         \3611 , \3612 , \3613 , \3614 , \3615 , \3616 , \3617 , \3618 , \3619 , \3620 ,
         \3621 , \3622 , \3623 , \3624 , \3625 , \3626 , \3627 , \3628 , \3629 , \3630 ,
         \3631 , \3632 , \3633 , \3634 , \3635 , \3636 , \3637 , \3638 , \3639 , \3640 ,
         \3641 , \3642 , \3643 , \3644 , \3645 , \3646 , \3647 , \3648 , \3649 , \3650 ,
         \3651 , \3652 , \3653 , \3654 , \3655 , \3656 , \3657 , \3658 , \3659 , \3660 ,
         \3661 , \3662 , \3663 , \3664 , \3665 , \3666 , \3667 , \3668 , \3669 , \3670 ,
         \3671 , \3672 , \3673 , \3674 , \3675 , \3676 , \3677 , \3678 , \3679 , \3680 ,
         \3681 , \3682 , \3683 , \3684 , \3685 , \3686 , \3687 , \3688 , \3689 , \3690 ,
         \3691 , \3692 , \3693 , \3694 , \3695 , \3696 , \3697 , \3698 , \3699 , \3700 ,
         \3701 , \3702 , \3703 , \3704 , \3705 , \3706 , \3707 , \3708 , \3709 , \3710 ,
         \3711 , \3712 , \3713 , \3714 , \3715 , \3716 , \3717 , \3718 , \3719 , \3720 ,
         \3721 , \3722 , \3723 , \3724 , \3725 , \3726 , \3727 , \3728 , \3729 , \3730 ,
         \3731 , \3732 , \3733 , \3734 , \3735 , \3736 , \3737 , \3738 , \3739 , \3740 ,
         \3741 , \3742 , \3743 , \3744 , \3745 , \3746 , \3747 , \3748 , \3749 , \3750 ,
         \3751 , \3752 , \3753 , \3754 , \3755 , \3756 , \3757 , \3758 , \3759 , \3760 ,
         \3761 , \3762 , \3763 , \3764 , \3765 , \3766 , \3767 , \3768 , \3769 , \3770 ,
         \3771 , \3772 , \3773 , \3774 , \3775 , \3776 , \3777 , \3778 , \3779 , \3780 ,
         \3781 , \3782 , \3783 , \3784 , \3785 , \3786 , \3787 , \3788 , \3789 , \3790 ,
         \3791 , \3792 , \3793 , \3794 , \3795 , \3796 , \3797 , \3798 , \3799 , \3800 ,
         \3801 , \3802 , \3803 , \3804 , \3805 , \3806 , \3807 , \3808 , \3809 , \3810 ,
         \3811 , \3812 , \3813 , \3814 , \3815 , \3816 , \3817 , \3818 , \3819 , \3820 ,
         \3821 , \3822 , \3823 , \3824 , \3825 , \3826 , \3827 , \3828 , \3829 , \3830 ,
         \3831 , \3832 , \3833 , \3834 , \3835 , \3836 , \3837 , \3838 , \3839 , \3840 ,
         \3841 , \3842 , \3843 , \3844 , \3845 , \3846 , \3847 , \3848 , \3849 , \3850 ,
         \3851 , \3852 , \3853 , \3854 , \3855 , \3856 , \3857 , \3858 , \3859 , \3860 ,
         \3861 , \3862 , \3863 , \3864 , \3865 , \3866 , \3867 , \3868 , \3869 , \3870 ,
         \3871 , \3872 , \3873 , \3874 , \3875 , \3876 , \3877 , \3878 , \3879 , \3880 ,
         \3881 , \3882 , \3883 , \3884 , \3885 , \3886 , \3887 , \3888 , \3889 , \3890 ,
         \3891 , \3892 , \3893 , \3894 , \3895 , \3896 , \3897 , \3898 , \3899 , \3900 ,
         \3901 , \3902 , \3903 , \3904 , \3905 , \3906 , \3907 , \3908 , \3909 , \3910 ,
         \3911 , \3912 , \3913 , \3914 , \3915 , \3916 , \3917 , \3918 , \3919 , \3920 ,
         \3921 , \3922 , \3923 , \3924 , \3925 , \3926 , \3927 , \3928 , \3929 , \3930 ,
         \3931 , \3932 , \3933 , \3934 , \3935 , \3936 , \3937 , \3938 , \3939 , \3940 ,
         \3941 , \3942 , \3943 , \3944 , \3945 , \3946 , \3947 , \3948 , \3949 , \3950 ,
         \3951 , \3952 , \3953 , \3954 , \3955 , \3956 , \3957 , \3958 , \3959 , \3960 ,
         \3961 , \3962 , \3963 , \3964 , \3965 , \3966 , \3967 , \3968 , \3969 , \3970 ,
         \3971 , \3972 , \3973 , \3974 , \3975 , \3976 , \3977 , \3978 , \3979 , \3980 ,
         \3981 , \3982 , \3983 , \3984 , \3985 , \3986 , \3987 , \3988 , \3989 , \3990 ,
         \3991 , \3992 , \3993 , \3994 , \3995 , \3996 , \3997 , \3998 , \3999 , \4000 ,
         \4001 , \4002 , \4003 , \4004 , \4005 , \4006 , \4007 , \4008 , \4009 , \4010 ,
         \4011 , \4012 , \4013 , \4014 , \4015 , \4016 , \4017 , \4018 , \4019 , \4020 ,
         \4021 , \4022 , \4023 , \4024 , \4025 , \4026 , \4027 , \4028 , \4029 , \4030 ,
         \4031 , \4032 , \4033 , \4034 , \4035 , \4036 , \4037 , \4038 , \4039 , \4040 ,
         \4041 , \4042 , \4043 , \4044 , \4045 , \4046 , \4047 , \4048 , \4049 , \4050 ,
         \4051 , \4052 , \4053 , \4054 , \4055 , \4056 , \4057 , \4058 , \4059 , \4060 ,
         \4061 , \4062 , \4063 , \4064 , \4065 , \4066 , \4067 , \4068 , \4069 , \4070 ,
         \4071 , \4072 , \4073 , \4074 , \4075 , \4076 , \4077 , \4078 , \4079 , \4080 ,
         \4081 , \4082 , \4083 , \4084 , \4085 , \4086 , \4087 , \4088 , \4089 , \4090 ,
         \4091 , \4092 , \4093 , \4094 , \4095 , \4096 , \4097 , \4098 , \4099 , \4100 ,
         \4101 , \4102 , \4103 , \4104 , \4105 , \4106 , \4107 , \4108 , \4109 , \4110 ,
         \4111 , \4112 , \4113 , \4114 , \4115 , \4116 , \4117 , \4118 , \4119 , \4120 ,
         \4121 , \4122 , \4123 , \4124 , \4125 , \4126 , \4127 , \4128 , \4129 , \4130 ,
         \4131 , \4132 , \4133 , \4134 , \4135 , \4136 , \4137 , \4138 , \4139 , \4140 ,
         \4141 , \4142 , \4143 , \4144 , \4145 , \4146 , \4147 , \4148 , \4149 , \4150 ,
         \4151 , \4152 , \4153 , \4154 , \4155 , \4156 , \4157 , \4158 , \4159 , \4160 ,
         \4161 , \4162 , \4163 , \4164 , \4165 , \4166 , \4167 , \4168 , \4169 , \4170 ,
         \4171 , \4172 , \4173 , \4174 , \4175 , \4176 , \4177 , \4178 , \4179 , \4180 ,
         \4181 , \4182 , \4183 , \4184 , \4185 , \4186 , \4187 , \4188 , \4189 , \4190 ,
         \4191 , \4192 , \4193 , \4194 , \4195 , \4196 , \4197 , \4198 , \4199 , \4200 ,
         \4201 , \4202 , \4203 , \4204 , \4205 , \4206 , \4207 , \4208 , \4209 , \4210 ,
         \4211 , \4212 , \4213 , \4214 , \4215 , \4216 , \4217 , \4218 , \4219 , \4220 ,
         \4221 , \4222 , \4223 , \4224 , \4225 , \4226 , \4227 , \4228 , \4229 , \4230 ,
         \4231 , \4232 , \4233 , \4234 , \4235 , \4236 , \4237 , \4238 , \4239 , \4240 ,
         \4241 , \4242 , \4243 , \4244 , \4245 , \4246 , \4247 , \4248 , \4249 , \4250 ,
         \4251 , \4252 , \4253 , \4254 , \4255 , \4256 , \4257 , \4258 , \4259 , \4260 ,
         \4261 , \4262 , \4263 , \4264 , \4265 , \4266 , \4267 , \4268 , \4269 , \4270 ,
         \4271 , \4272 , \4273 , \4274 , \4275 , \4276 , \4277 , \4278 , \4279 , \4280 ,
         \4281 , \4282 , \4283 , \4284 , \4285 , \4286 , \4287 , \4288 , \4289 , \4290 ,
         \4291 , \4292 , \4293 , \4294 , \4295 , \4296 , \4297 , \4298 , \4299 , \4300 ,
         \4301 , \4302 , \4303 , \4304 , \4305 , \4306 , \4307 , \4308 , \4309 , \4310 ,
         \4311 , \4312 , \4313 , \4314 , \4315 , \4316 , \4317 , \4318 , \4319 , \4320 ,
         \4321 , \4322 , \4323 , \4324 , \4325 , \4326 , \4327 , \4328 , \4329 , \4330 ,
         \4331 , \4332 , \4333 , \4334 , \4335 , \4336 , \4337 , \4338 , \4339 , \4340 ,
         \4341 , \4342 , \4343 , \4344 , \4345 , \4346 , \4347 , \4348 , \4349 , \4350 ,
         \4351 , \4352 , \4353 , \4354 , \4355 , \4356 , \4357 , \4358 , \4359 , \4360 ,
         \4361 , \4362 , \4363 , \4364 , \4365 , \4366 , \4367 , \4368 , \4369 , \4370 ,
         \4371 , \4372 , \4373 , \4374 , \4375 , \4376 , \4377 , \4378 , \4379 , \4380 ,
         \4381 , \4382 , \4383 , \4384 , \4385 , \4386 , \4387 , \4388 , \4389 , \4390 ,
         \4391 , \4392 , \4393 , \4394 , \4395 , \4396 , \4397 , \4398 , \4399 , \4400 ,
         \4401 , \4402 , \4403 , \4404 , \4405 , \4406 , \4407 , \4408 , \4409 , \4410 ,
         \4411 , \4412 , \4413 , \4414 , \4415 , \4416 , \4417 , \4418 , \4419 , \4420 ,
         \4421 , \4422 , \4423 , \4424 , \4425 , \4426 , \4427 , \4428 , \4429 , \4430 ,
         \4431 , \4432 , \4433 , \4434 , \4435 , \4436 , \4437 , \4438 , \4439 , \4440 ,
         \4441 , \4442 , \4443 , \4444 , \4445 , \4446 , \4447 , \4448 , \4449 , \4450 ,
         \4451 , \4452 , \4453 , \4454 , \4455 , \4456 , \4457 , \4458 , \4459 , \4460 ,
         \4461 , \4462 , \4463 , \4464 , \4465 , \4466 , \4467 , \4468 , \4469 , \4470 ,
         \4471 , \4472 , \4473 , \4474 , \4475 , \4476 , \4477 , \4478 , \4479 , \4480 ,
         \4481 , \4482 , \4483 , \4484 , \4485 , \4486 , \4487 , \4488 , \4489 , \4490 ,
         \4491 , \4492 , \4493 , \4494 , \4495 , \4496 , \4497 , \4498 , \4499 , \4500 ,
         \4501 , \4502 , \4503 , \4504 , \4505 , \4506 , \4507 , \4508 , \4509 , \4510 ,
         \4511 , \4512 , \4513 , \4514 , \4515 , \4516 , \4517 , \4518 , \4519 , \4520 ,
         \4521 , \4522 , \4523 , \4524 , \4525 , \4526 , \4527 , \4528 , \4529 , \4530 ,
         \4531 , \4532 , \4533 , \4534 , \4535 , \4536 , \4537 , \4538 , \4539 , \4540 ,
         \4541 , \4542 , \4543 , \4544 , \4545 , \4546 , \4547 , \4548 , \4549 , \4550 ,
         \4551 , \4552 , \4553 , \4554 , \4555 , \4556 , \4557 , \4558 , \4559 , \4560 ,
         \4561 , \4562 , \4563 , \4564 , \4565 , \4566 , \4567 , \4568 , \4569 , \4570 ,
         \4571 , \4572 , \4573 , \4574 , \4575 , \4576 , \4577 , \4578 , \4579 , \4580 ,
         \4581 , \4582 , \4583 , \4584 , \4585 , \4586 , \4587 , \4588 , \4589 , \4590 ,
         \4591 , \4592 , \4593 , \4594 , \4595 , \4596 , \4597 , \4598 , \4599 , \4600 ,
         \4601 , \4602 , \4603 , \4604 , \4605 , \4606 , \4607 , \4608 , \4609 , \4610 ,
         \4611 , \4612 , \4613 , \4614 , \4615 , \4616 , \4617 , \4618 , \4619 , \4620 ,
         \4621 , \4622 , \4623 , \4624 , \4625 , \4626 , \4627 , \4628 , \4629 , \4630 ,
         \4631 , \4632 , \4633 , \4634 , \4635 , \4636 , \4637 , \4638 , \4639 , \4640 ,
         \4641 , \4642 , \4643 , \4644 , \4645 , \4646 , \4647 , \4648 , \4649 , \4650 ,
         \4651 , \4652 , \4653 , \4654 , \4655 , \4656 , \4657 , \4658 , \4659 , \4660 ,
         \4661 , \4662 , \4663 , \4664 , \4665 , \4666 , \4667 , \4668 , \4669 , \4670 ,
         \4671 , \4672 , \4673 , \4674 , \4675 , \4676 , \4677 , \4678 , \4679 , \4680 ,
         \4681 , \4682 , \4683 , \4684 , \4685 , \4686 , \4687 , \4688 , \4689 , \4690 ,
         \4691 , \4692 , \4693 , \4694 , \4695 , \4696 , \4697 , \4698 , \4699 , \4700 ,
         \4701 , \4702 , \4703 , \4704 , \4705 , \4706 , \4707 , \4708 , \4709 , \4710 ,
         \4711 , \4712 , \4713 , \4714 , \4715 , \4716 , \4717 , \4718 , \4719 , \4720 ,
         \4721 , \4722 , \4723 , \4724 , \4725 , \4726 , \4727 , \4728 , \4729 , \4730 ,
         \4731 , \4732 , \4733 , \4734 , \4735 , \4736 , \4737 , \4738 , \4739 , \4740 ,
         \4741 , \4742 , \4743 , \4744 , \4745 , \4746 , \4747 , \4748 , \4749 , \4750 ,
         \4751 , \4752 , \4753 , \4754 , \4755 , \4756 , \4757 , \4758 , \4759 , \4760 ,
         \4761 , \4762 , \4763 , \4764 , \4765 , \4766 , \4767 , \4768 , \4769 , \4770 ,
         \4771 , \4772 , \4773 , \4774 , \4775 , \4776 , \4777 , \4778 , \4779 , \4780 ,
         \4781 , \4782 , \4783 , \4784 , \4785 , \4786 , \4787 , \4788 , \4789 , \4790 ,
         \4791 , \4792 , \4793 , \4794 , \4795 , \4796 , \4797 , \4798 , \4799 , \4800 ,
         \4801 , \4802 , \4803 , \4804 , \4805 , \4806 , \4807 , \4808 , \4809 , \4810 ,
         \4811 , \4812 , \4813 , \4814 , \4815 , \4816 , \4817 , \4818 , \4819 , \4820 ,
         \4821 , \4822 , \4823 , \4824 , \4825 , \4826 , \4827 , \4828 , \4829 , \4830 ,
         \4831 , \4832 , \4833 , \4834 , \4835 , \4836 , \4837 , \4838 , \4839 , \4840 ,
         \4841 , \4842 , \4843 , \4844 , \4845 , \4846 , \4847 , \4848 , \4849 , \4850 ,
         \4851 , \4852 , \4853 , \4854 , \4855 , \4856 , \4857 , \4858 , \4859 , \4860 ,
         \4861 , \4862 , \4863 , \4864 , \4865 , \4866 , \4867 , \4868 , \4869 , \4870 ,
         \4871 , \4872 , \4873 , \4874 , \4875 , \4876 , \4877 , \4878 , \4879 , \4880 ,
         \4881 , \4882 , \4883 , \4884 , \4885 , \4886 , \4887 , \4888 , \4889 , \4890 ,
         \4891 , \4892 , \4893 , \4894 , \4895 , \4896 , \4897 , \4898 , \4899 , \4900 ,
         \4901 , \4902 , \4903 , \4904 , \4905 , \4906 , \4907 , \4908 , \4909 , \4910 ,
         \4911 , \4912 , \4913 , \4914 , \4915 , \4916 , \4917 , \4918 , \4919 , \4920 ,
         \4921 , \4922 , \4923 , \4924 , \4925 , \4926 , \4927 , \4928 , \4929 , \4930 ,
         \4931 , \4932 , \4933 , \4934 , \4935 , \4936 , \4937 , \4938 , \4939 , \4940 ,
         \4941 , \4942 , \4943 , \4944 , \4945 , \4946 , \4947 , \4948 , \4949 , \4950 ,
         \4951 , \4952 , \4953 , \4954 , \4955 , \4956 , \4957 , \4958 , \4959 , \4960 ,
         \4961 , \4962 , \4963 , \4964 , \4965 , \4966 , \4967 , \4968 , \4969 , \4970 ,
         \4971 , \4972 , \4973 , \4974 , \4975 , \4976 , \4977 , \4978 , \4979 , \4980 ,
         \4981 , \4982 , \4983 , \4984 , \4985 , \4986 , \4987 , \4988 , \4989 , \4990 ,
         \4991 , \4992 , \4993 , \4994 , \4995 , \4996 , \4997 , \4998 , \4999 , \5000 ,
         \5001 , \5002 , \5003 , \5004 , \5005 , \5006 , \5007 , \5008 , \5009 , \5010 ,
         \5011 , \5012 , \5013 , \5014 , \5015 , \5016 , \5017 , \5018 , \5019 , \5020 ,
         \5021 , \5022 , \5023 , \5024 , \5025 , \5026 , \5027 , \5028 , \5029 , \5030 ,
         \5031 , \5032 , \5033 , \5034 , \5035 , \5036 , \5037 , \5038 , \5039 , \5040 ,
         \5041 , \5042 , \5043 , \5044 , \5045 , \5046 , \5047 , \5048 , \5049 , \5050 ,
         \5051 , \5052 , \5053 , \5054 , \5055 , \5056 , \5057 , \5058 , \5059 , \5060 ,
         \5061 , \5062 , \5063 , \5064 , \5065 , \5066 , \5067 , \5068 , \5069 , \5070 ,
         \5071 , \5072 , \5073 , \5074 , \5075 , \5076 , \5077 , \5078 , \5079 , \5080 ,
         \5081 , \5082 , \5083 , \5084 , \5085 , \5086 , \5087 , \5088 , \5089 , \5090 ,
         \5091 , \5092 , \5093 , \5094 , \5095 , \5096 , \5097 , \5098 , \5099 , \5100 ,
         \5101 , \5102 , \5103 , \5104 , \5105 , \5106 , \5107 , \5108 , \5109 , \5110 ,
         \5111 , \5112 , \5113 , \5114 , \5115 , \5116 , \5117 , \5118 , \5119 , \5120 ,
         \5121 , \5122 , \5123 , \5124 , \5125 , \5126 , \5127 , \5128 , \5129 , \5130 ,
         \5131 , \5132 , \5133 , \5134 , \5135 , \5136 , \5137 , \5138 , \5139 , \5140 ,
         \5141 , \5142 , \5143 , \5144 , \5145 , \5146 , \5147 , \5148 , \5149 , \5150 ,
         \5151 , \5152 , \5153 , \5154 , \5155 , \5156 , \5157 , \5158 , \5159 , \5160 ,
         \5161 , \5162 , \5163 , \5164 , \5165 , \5166 , \5167 , \5168 , \5169 , \5170 ,
         \5171 , \5172 , \5173 , \5174 , \5175 , \5176 , \5177 , \5178 , \5179 , \5180 ,
         \5181 , \5182 , \5183 , \5184 , \5185 , \5186 , \5187 , \5188 , \5189 , \5190 ,
         \5191 , \5192 , \5193 , \5194 , \5195 , \5196 , \5197 , \5198 , \5199 , \5200 ,
         \5201 , \5202 , \5203 , \5204 , \5205 , \5206 , \5207 , \5208 , \5209 , \5210 ,
         \5211 , \5212 , \5213 , \5214 , \5215 , \5216 , \5217 , \5218 , \5219 , \5220 ,
         \5221 , \5222 , \5223 , \5224 , \5225 , \5226 , \5227 , \5228 , \5229 , \5230 ,
         \5231 , \5232 , \5233 , \5234 , \5235 , \5236 , \5237 , \5238 , \5239 , \5240 ,
         \5241 , \5242 , \5243 , \5244 , \5245 , \5246 , \5247 , \5248 , \5249 , \5250 ,
         \5251 , \5252 , \5253 , \5254 , \5255 , \5256 , \5257 , \5258 , \5259 , \5260 ,
         \5261 , \5262 , \5263 , \5264 , \5265 , \5266 , \5267 , \5268 , \5269 , \5270 ,
         \5271 , \5272 , \5273 , \5274 , \5275 , \5276 , \5277 , \5278 , \5279 , \5280 ,
         \5281 , \5282 , \5283 , \5284 , \5285 , \5286 , \5287 , \5288 , \5289 , \5290 ,
         \5291 , \5292 , \5293 , \5294 , \5295 , \5296 , \5297 , \5298 , \5299 , \5300 ,
         \5301 , \5302 , \5303 , \5304 , \5305 , \5306 , \5307 , \5308 , \5309 , \5310 ,
         \5311 , \5312 , \5313 , \5314 , \5315 , \5316 , \5317 , \5318 , \5319 , \5320 ,
         \5321 , \5322 , \5323 , \5324 , \5325 , \5326 , \5327 , \5328 , \5329 , \5330 ,
         \5331 , \5332 , \5333 , \5334 , \5335 , \5336 , \5337 , \5338 , \5339 , \5340 ,
         \5341 , \5342 , \5343 , \5344 , \5345 , \5346 , \5347 , \5348 , \5349 , \5350 ,
         \5351 , \5352 , \5353 , \5354 , \5355 , \5356 , \5357 , \5358 , \5359 , \5360 ,
         \5361 , \5362 , \5363 , \5364 , \5365 , \5366 , \5367 , \5368 , \5369 , \5370 ,
         \5371 , \5372 , \5373 , \5374 , \5375 , \5376 , \5377 , \5378 , \5379 , \5380 ,
         \5381 , \5382 , \5383 , \5384 , \5385 , \5386 , \5387 , \5388 , \5389 , \5390 ,
         \5391 , \5392 , \5393 , \5394 , \5395 , \5396 , \5397 , \5398 , \5399 , \5400 ,
         \5401 , \5402 , \5403 , \5404 , \5405 , \5406 , \5407 , \5408 , \5409 , \5410 ,
         \5411 , \5412 , \5413 , \5414 , \5415 , \5416 , \5417 , \5418 , \5419 , \5420 ,
         \5421 , \5422 , \5423 , \5424 , \5425 , \5426 , \5427 , \5428 , \5429 , \5430 ,
         \5431 , \5432 , \5433 , \5434 , \5435 , \5436 , \5437 , \5438 , \5439 , \5440 ,
         \5441 , \5442 , \5443 , \5444 , \5445 , \5446 , \5447 , \5448 , \5449 , \5450 ,
         \5451 , \5452 , \5453 , \5454 , \5455 , \5456 , \5457 , \5458 , \5459 , \5460 ,
         \5461 , \5462 , \5463 , \5464 , \5465 , \5466 , \5467 , \5468 , \5469 , \5470 ,
         \5471 , \5472 , \5473 , \5474 , \5475 , \5476 , \5477 , \5478 , \5479 , \5480 ,
         \5481 , \5482 , \5483 , \5484 , \5485 , \5486 , \5487 , \5488 , \5489 , \5490 ,
         \5491 , \5492 , \5493 , \5494 , \5495 , \5496 , \5497 , \5498 , \5499 , \5500 ,
         \5501 , \5502 , \5503 , \5504 , \5505 , \5506 , \5507 , \5508 , \5509 , \5510 ,
         \5511 , \5512 , \5513 , \5514 , \5515 , \5516 , \5517 , \5518 , \5519 , \5520 ,
         \5521 , \5522 , \5523 , \5524 , \5525 , \5526 , \5527 , \5528 , \5529 , \5530 ,
         \5531 , \5532 , \5533 , \5534 , \5535 , \5536 , \5537 , \5538 , \5539 , \5540 ,
         \5541 , \5542 , \5543 , \5544 , \5545 , \5546 , \5547 , \5548 , \5549 , \5550 ,
         \5551 , \5552 , \5553 , \5554 , \5555 , \5556 , \5557 , \5558 , \5559 , \5560 ,
         \5561 , \5562 , \5563 , \5564 , \5565 , \5566 , \5567 , \5568 , \5569 , \5570 ,
         \5571 , \5572 , \5573 , \5574 , \5575 , \5576 , \5577 , \5578 , \5579 , \5580 ,
         \5581 , \5582 , \5583 , \5584 , \5585 , \5586 , \5587 , \5588 , \5589 , \5590 ,
         \5591 , \5592 , \5593 , \5594 , \5595 , \5596 , \5597 , \5598 , \5599 , \5600 ,
         \5601 , \5602 , \5603 , \5604 , \5605 , \5606 , \5607 , \5608 , \5609 , \5610 ,
         \5611 , \5612 , \5613 , \5614 , \5615 , \5616 , \5617 , \5618 , \5619 , \5620 ,
         \5621 , \5622 , \5623 , \5624 , \5625 , \5626 , \5627 , \5628 , \5629 , \5630 ,
         \5631 , \5632 , \5633 , \5634 , \5635 , \5636 , \5637 , \5638 , \5639 , \5640 ,
         \5641 , \5642 , \5643 , \5644 , \5645 , \5646 , \5647 , \5648 , \5649 , \5650 ,
         \5651 , \5652 , \5653 , \5654 , \5655 , \5656 , \5657 , \5658 , \5659 , \5660 ,
         \5661 , \5662 , \5663 , \5664 , \5665 , \5666 , \5667 , \5668 , \5669 , \5670 ,
         \5671 , \5672 , \5673 , \5674 , \5675 , \5676 , \5677 , \5678 , \5679 , \5680 ,
         \5681 , \5682 , \5683 , \5684 , \5685 , \5686 , \5687 , \5688 , \5689 , \5690 ,
         \5691 , \5692 , \5693 , \5694 , \5695 , \5696 , \5697 , \5698 , \5699 , \5700 ,
         \5701 , \5702 , \5703 , \5704 , \5705 , \5706 , \5707 , \5708 , \5709 , \5710 ,
         \5711 , \5712 , \5713 , \5714 , \5715 , \5716 , \5717 , \5718 , \5719 , \5720 ,
         \5721 , \5722 , \5723 , \5724 , \5725 , \5726 , \5727 , \5728 , \5729 , \5730 ,
         \5731 , \5732 , \5733 , \5734 , \5735 , \5736 , \5737 , \5738 , \5739 , \5740 ,
         \5741 , \5742 , \5743 , \5744 , \5745 , \5746 , \5747 , \5748 , \5749 , \5750 ,
         \5751 , \5752 , \5753 , \5754 , \5755 , \5756 , \5757 , \5758 , \5759 , \5760 ,
         \5761 , \5762 , \5763 , \5764 , \5765 , \5766 , \5767 , \5768 , \5769 , \5770 ,
         \5771 , \5772 , \5773 , \5774 , \5775 , \5776 , \5777 , \5778 , \5779 , \5780 ,
         \5781 , \5782 , \5783 , \5784 , \5785 , \5786 , \5787 , \5788 , \5789 , \5790 ,
         \5791 , \5792 , \5793 , \5794 , \5795 , \5796 , \5797 , \5798 , \5799 , \5800 ,
         \5801 , \5802 , \5803 , \5804 , \5805 , \5806 , \5807 , \5808 , \5809 , \5810 ,
         \5811 , \5812 , \5813 , \5814 , \5815 , \5816 , \5817 , \5818 , \5819 , \5820 ,
         \5821 , \5822 , \5823 , \5824 , \5825 , \5826 , \5827 , \5828 , \5829 , \5830 ,
         \5831 , \5832 , \5833 , \5834 , \5835 , \5836 , \5837 , \5838 , \5839 , \5840 ,
         \5841 , \5842 , \5843 , \5844 , \5845 , \5846 , \5847 , \5848 , \5849 , \5850 ,
         \5851 , \5852 , \5853 , \5854 , \5855 , \5856 , \5857 , \5858 , \5859 , \5860 ,
         \5861 , \5862 , \5863 , \5864 , \5865 , \5866 , \5867 , \5868 , \5869 , \5870 ,
         \5871 , \5872 , \5873 , \5874 , \5875 , \5876 , \5877 , \5878 , \5879 , \5880 ,
         \5881 , \5882 , \5883 , \5884 , \5885 , \5886 , \5887 , \5888 , \5889 , \5890 ,
         \5891 , \5892 , \5893 , \5894 , \5895 , \5896 , \5897 , \5898 , \5899 , \5900 ,
         \5901 , \5902 , \5903 , \5904 , \5905 , \5906 , \5907 , \5908 , \5909 , \5910 ,
         \5911 , \5912 , \5913 , \5914 , \5915 , \5916 , \5917 , \5918 , \5919 , \5920 ,
         \5921 , \5922 , \5923 , \5924 , \5925 , \5926 , \5927 , \5928 , \5929 , \5930 ,
         \5931 , \5932 , \5933 , \5934 , \5935 , \5936 , \5937 , \5938 , \5939 , \5940 ,
         \5941 , \5942 , \5943 , \5944 , \5945 , \5946 , \5947 , \5948 , \5949 , \5950 ,
         \5951 , \5952 , \5953 , \5954 , \5955 , \5956 , \5957 , \5958 , \5959 , \5960 ,
         \5961 , \5962 , \5963 , \5964 , \5965 , \5966 , \5967 , \5968 , \5969 , \5970 ,
         \5971 , \5972 , \5973 , \5974 , \5975 , \5976 , \5977 , \5978 , \5979 , \5980 ,
         \5981 , \5982 , \5983 , \5984 , \5985 , \5986 , \5987 , \5988 , \5989 , \5990 ,
         \5991 , \5992 , \5993 , \5994 , \5995 , \5996 , \5997 , \5998 , \5999 , \6000 ,
         \6001 , \6002 , \6003 , \6004 , \6005 , \6006 , \6007 , \6008 , \6009 , \6010 ,
         \6011 , \6012 , \6013 , \6014 , \6015 , \6016 , \6017 , \6018 , \6019 , \6020 ,
         \6021 , \6022 , \6023 , \6024 , \6025 , \6026 , \6027 , \6028 , \6029 , \6030 ,
         \6031 , \6032 , \6033 , \6034 , \6035 , \6036 , \6037 , \6038 , \6039 , \6040 ,
         \6041 , \6042 , \6043 , \6044 , \6045 , \6046 , \6047 , \6048 , \6049 , \6050 ,
         \6051 , \6052 , \6053 , \6054 , \6055 , \6056 , \6057 , \6058 , \6059 , \6060 ,
         \6061 , \6062 , \6063 , \6064 , \6065 , \6066 , \6067 , \6068 , \6069 , \6070 ,
         \6071 , \6072 , \6073 , \6074 , \6075 , \6076 , \6077 , \6078 , \6079 , \6080 ,
         \6081 , \6082 , \6083 , \6084 , \6085 , \6086 , \6087 , \6088 , \6089 , \6090 ,
         \6091 , \6092 , \6093 , \6094 , \6095 , \6096 , \6097 , \6098 , \6099 , \6100 ,
         \6101 , \6102 , \6103 , \6104 , \6105 , \6106 , \6107 , \6108 , \6109 , \6110 ,
         \6111 , \6112 , \6113 , \6114 , \6115 , \6116 , \6117 , \6118 , \6119 , \6120 ,
         \6121 , \6122 , \6123 , \6124 , \6125 , \6126 , \6127 , \6128 , \6129 , \6130 ,
         \6131 , \6132 , \6133 , \6134 , \6135 , \6136 , \6137 , \6138 , \6139 , \6140 ,
         \6141 , \6142 , \6143 , \6144 , \6145 , \6146 , \6147 , \6148 , \6149 , \6150 ,
         \6151 , \6152 , \6153 , \6154 , \6155 , \6156 , \6157 , \6158 , \6159 , \6160 ,
         \6161 , \6162 , \6163 , \6164 , \6165 , \6166 , \6167 , \6168 , \6169 , \6170 ,
         \6171 , \6172 , \6173 , \6174 , \6175 , \6176 , \6177 , \6178 , \6179 , \6180 ,
         \6181 , \6182 , \6183 , \6184 , \6185 , \6186 , \6187 , \6188 , \6189 , \6190 ,
         \6191 , \6192 , \6193 , \6194 , \6195 , \6196 , \6197 , \6198 , \6199 , \6200 ,
         \6201 , \6202 , \6203 , \6204 , \6205 , \6206 , \6207 , \6208 , \6209 , \6210 ,
         \6211 , \6212 , \6213 , \6214 , \6215 , \6216 , \6217 , \6218 , \6219 , \6220 ,
         \6221 , \6222 , \6223 , \6224 , \6225 , \6226 , \6227 , \6228 , \6229 , \6230 ,
         \6231 , \6232 , \6233 , \6234 , \6235 , \6236 , \6237 , \6238 , \6239 , \6240 ,
         \6241 , \6242 , \6243 , \6244 , \6245 , \6246 , \6247 , \6248 , \6249 , \6250 ,
         \6251 , \6252 , \6253 , \6254 , \6255 , \6256 , \6257 , \6258 , \6259 , \6260 ,
         \6261 , \6262 , \6263 , \6264 , \6265 , \6266 , \6267 , \6268 , \6269 , \6270 ,
         \6271 , \6272 , \6273 , \6274 , \6275 , \6276 , \6277 , \6278 , \6279 , \6280 ,
         \6281 , \6282 , \6283 , \6284 , \6285 , \6286 , \6287 , \6288 , \6289 , \6290 ,
         \6291 , \6292 , \6293 , \6294 , \6295 , \6296 , \6297 , \6298 , \6299 , \6300 ,
         \6301 , \6302 , \6303 , \6304 , \6305 , \6306 , \6307 , \6308 , \6309 , \6310 ,
         \6311 , \6312 , \6313 , \6314 , \6315 , \6316 , \6317 , \6318 , \6319 , \6320 ,
         \6321 , \6322 , \6323 , \6324 , \6325 , \6326 , \6327 , \6328 , \6329 , \6330 ,
         \6331 , \6332 , \6333 , \6334 , \6335 , \6336 , \6337 , \6338 , \6339 , \6340 ,
         \6341 , \6342 , \6343 , \6344 , \6345 , \6346 , \6347 , \6348 , \6349 , \6350 ,
         \6351 , \6352 , \6353 , \6354 , \6355 , \6356 , \6357 , \6358 , \6359 , \6360 ,
         \6361 , \6362 , \6363 , \6364 , \6365 , \6366 , \6367 , \6368 , \6369 , \6370 ,
         \6371 , \6372 , \6373 , \6374 , \6375 , \6376 , \6377 , \6378 , \6379 , \6380 ,
         \6381 , \6382 , \6383 , \6384 , \6385 , \6386 , \6387 , \6388 , \6389 , \6390 ,
         \6391 , \6392 , \6393 , \6394 , \6395 , \6396 , \6397 , \6398 , \6399 , \6400 ,
         \6401 , \6402 , \6403 , \6404 , \6405 , \6406 , \6407 , \6408 , \6409 , \6410 ,
         \6411 , \6412 , \6413 , \6414 , \6415 , \6416 , \6417 , \6418 , \6419 , \6420 ,
         \6421 , \6422 , \6423 , \6424 , \6425 , \6426 , \6427 , \6428 , \6429 , \6430 ,
         \6431 , \6432 , \6433 , \6434 , \6435 , \6436 , \6437 , \6438 , \6439 , \6440 ,
         \6441 , \6442 , \6443 , \6444 , \6445 , \6446 , \6447 , \6448 , \6449 , \6450 ,
         \6451 , \6452 , \6453 , \6454 , \6455 , \6456 , \6457 , \6458 , \6459 , \6460 ,
         \6461 , \6462 , \6463 , \6464 , \6465 , \6466 , \6467 , \6468 , \6469 , \6470 ,
         \6471 , \6472 , \6473 , \6474 , \6475 , \6476 , \6477 , \6478 , \6479 , \6480 ,
         \6481 , \6482 , \6483 , \6484 , \6485 , \6486 , \6487 , \6488 , \6489 , \6490 ,
         \6491 , \6492 , \6493 , \6494 , \6495 , \6496 , \6497 , \6498 , \6499 , \6500 ,
         \6501 , \6502 , \6503 , \6504 , \6505 , \6506 , \6507 , \6508 , \6509 , \6510 ,
         \6511 , \6512 , \6513 , \6514 , \6515 , \6516 , \6517 , \6518 , \6519 , \6520 ,
         \6521 , \6522 , \6523 , \6524 , \6525 , \6526 , \6527 , \6528 , \6529 , \6530 ,
         \6531 , \6532 , \6533 , \6534 , \6535 , \6536 , \6537 , \6538 , \6539 , \6540 ,
         \6541 , \6542 , \6543 , \6544 , \6545 , \6546 , \6547 , \6548 , \6549 , \6550 ,
         \6551 , \6552 , \6553 , \6554 , \6555 , \6556 , \6557 , \6558 , \6559 , \6560 ,
         \6561 , \6562 , \6563 , \6564 , \6565 , \6566 , \6567 , \6568 , \6569 , \6570 ,
         \6571 , \6572 , \6573 , \6574 , \6575 , \6576 , \6577 , \6578 , \6579 , \6580 ,
         \6581 , \6582 , \6583 , \6584 , \6585 , \6586 , \6587 , \6588 , \6589 , \6590 ,
         \6591 , \6592 , \6593 , \6594 , \6595 , \6596 , \6597 , \6598 , \6599 , \6600 ,
         \6601 , \6602 , \6603 , \6604 , \6605 , \6606 , \6607 , \6608 , \6609 , \6610 ,
         \6611 , \6612 , \6613 , \6614 , \6615 , \6616 , \6617 , \6618 , \6619 , \6620 ,
         \6621 , \6622 , \6623 , \6624 , \6625 , \6626 , \6627 , \6628 , \6629 , \6630 ,
         \6631 , \6632 , \6633 , \6634 , \6635 , \6636 , \6637 , \6638 , \6639 , \6640 ,
         \6641 , \6642 , \6643 , \6644 , \6645 , \6646 , \6647 , \6648 , \6649 , \6650 ,
         \6651 , \6652 , \6653 , \6654 , \6655 , \6656 , \6657 , \6658 , \6659 , \6660 ,
         \6661 , \6662 , \6663 , \6664 , \6665 , \6666 , \6667 , \6668 , \6669 , \6670 ,
         \6671 , \6672 , \6673 , \6674 , \6675 , \6676 , \6677 , \6678 , \6679 , \6680 ,
         \6681 , \6682 , \6683 , \6684 , \6685 , \6686 , \6687 , \6688 , \6689 , \6690 ,
         \6691 , \6692 , \6693 , \6694 , \6695 , \6696 , \6697 , \6698 , \6699 , \6700 ,
         \6701 , \6702 , \6703 , \6704 , \6705 , \6706 , \6707 , \6708 , \6709 , \6710 ,
         \6711 , \6712 , \6713 , \6714 , \6715 , \6716 , \6717 , \6718 , \6719 , \6720 ,
         \6721 , \6722 , \6723 , \6724 , \6725 , \6726 , \6727 , \6728 , \6729 , \6730 ,
         \6731 , \6732 , \6733 , \6734 , \6735 , \6736 , \6737 , \6738 , \6739 , \6740 ,
         \6741 , \6742 , \6743 , \6744 , \6745 , \6746 , \6747 , \6748 , \6749 , \6750 ,
         \6751 , \6752 , \6753 , \6754 , \6755 , \6756 , \6757 , \6758 , \6759 , \6760 ,
         \6761 , \6762 , \6763 , \6764 , \6765 , \6766 , \6767 , \6768 , \6769 , \6770 ,
         \6771 , \6772 , \6773 , \6774 , \6775 , \6776 , \6777 , \6778 , \6779 , \6780 ,
         \6781 , \6782 , \6783 , \6784 , \6785 , \6786 , \6787 , \6788 , \6789 , \6790 ,
         \6791 , \6792 , \6793 , \6794 , \6795 , \6796 , \6797 , \6798 , \6799 , \6800 ,
         \6801 , \6802 , \6803 , \6804 , \6805 , \6806 , \6807 , \6808 , \6809 , \6810 ,
         \6811 , \6812 , \6813 , \6814 , \6815 , \6816 , \6817 , \6818 , \6819 , \6820 ,
         \6821 , \6822 , \6823 , \6824 , \6825 , \6826 , \6827 , \6828 , \6829 , \6830 ,
         \6831 , \6832 , \6833 , \6834 , \6835 , \6836 , \6837 , \6838 , \6839 , \6840 ,
         \6841 , \6842 , \6843 , \6844 , \6845 , \6846 , \6847 , \6848 , \6849 , \6850 ,
         \6851 , \6852 , \6853 , \6854 , \6855 , \6856 , \6857 , \6858 , \6859 , \6860 ,
         \6861 , \6862 , \6863 , \6864 , \6865 , \6866 , \6867 , \6868 , \6869 , \6870 ,
         \6871 , \6872 , \6873 , \6874 , \6875 , \6876 , \6877 , \6878 , \6879 , \6880 ,
         \6881 , \6882 , \6883 , \6884 , \6885 , \6886 , \6887 , \6888 , \6889 , \6890 ,
         \6891 , \6892 , \6893 , \6894 , \6895 , \6896 , \6897 , \6898 , \6899 , \6900 ,
         \6901 , \6902 , \6903 , \6904 , \6905 , \6906 , \6907 , \6908 , \6909 , \6910 ,
         \6911 , \6912 , \6913 , \6914 , \6915 , \6916 , \6917 , \6918 , \6919 , \6920 ,
         \6921 , \6922 , \6923 , \6924 , \6925 , \6926 , \6927 , \6928 , \6929 , \6930 ,
         \6931 , \6932 , \6933 , \6934 , \6935 , \6936 , \6937 , \6938 , \6939 , \6940 ,
         \6941 , \6942 , \6943 , \6944 , \6945 , \6946 , \6947 , \6948 , \6949 , \6950 ,
         \6951 , \6952 , \6953 , \6954 , \6955 , \6956 , \6957 , \6958 , \6959 , \6960 ,
         \6961 , \6962 , \6963 , \6964 , \6965 , \6966 , \6967 , \6968 , \6969 , \6970 ,
         \6971 , \6972 , \6973 , \6974 , \6975 , \6976 , \6977 , \6978 , \6979 , \6980 ,
         \6981 , \6982 , \6983 , \6984 , \6985 , \6986 , \6987 , \6988 , \6989 , \6990 ,
         \6991 , \6992 , \6993 , \6994 , \6995 , \6996 , \6997 , \6998 , \6999 , \7000 ,
         \7001 , \7002 , \7003 , \7004 , \7005 , \7006 , \7007 , \7008 , \7009 , \7010 ,
         \7011 , \7012 , \7013 , \7014 , \7015 , \7016 , \7017 , \7018 , \7019 , \7020 ,
         \7021 , \7022 , \7023 , \7024 , \7025 , \7026 , \7027 , \7028 , \7029 , \7030 ,
         \7031 , \7032 , \7033 , \7034 , \7035 , \7036 , \7037 , \7038 , \7039 , \7040 ,
         \7041 , \7042 , \7043 , \7044 , \7045 , \7046 , \7047 , \7048 , \7049 , \7050 ,
         \7051 , \7052 , \7053 , \7054 , \7055 , \7056 , \7057 , \7058 , \7059 , \7060 ,
         \7061 , \7062 , \7063 , \7064 , \7065 , \7066 , \7067 , \7068 , \7069 , \7070 ,
         \7071 , \7072 , \7073 , \7074 , \7075 , \7076 , \7077 , \7078 , \7079 , \7080 ,
         \7081 , \7082 , \7083 , \7084 , \7085 , \7086 , \7087 , \7088 , \7089 , \7090 ,
         \7091 , \7092 , \7093 , \7094 , \7095 , \7096 , \7097 , \7098 , \7099 , \7100 ,
         \7101 , \7102 , \7103 , \7104 , \7105 , \7106 , \7107 , \7108 , \7109 , \7110 ,
         \7111 , \7112 , \7113 , \7114 , \7115 , \7116 , \7117 , \7118 , \7119 , \7120 ,
         \7121 , \7122 , \7123 , \7124 , \7125 , \7126 , \7127 , \7128 , \7129 , \7130 ,
         \7131 , \7132 , \7133 , \7134 , \7135 , \7136 , \7137 , \7138 , \7139 , \7140 ,
         \7141 , \7142 , \7143 , \7144 , \7145 , \7146 , \7147 , \7148 , \7149 , \7150 ,
         \7151 , \7152 , \7153 , \7154 , \7155 , \7156 , \7157 , \7158 , \7159 , \7160 ,
         \7161 , \7162 , \7163 , \7164 , \7165 , \7166 , \7167 , \7168 , \7169 , \7170 ,
         \7171 , \7172 , \7173 , \7174 , \7175 , \7176 , \7177 , \7178 , \7179 , \7180 ,
         \7181 , \7182 , \7183 , \7184 , \7185 , \7186 , \7187 , \7188 , \7189 , \7190 ,
         \7191 , \7192 , \7193 , \7194 , \7195 , \7196 , \7197 , \7198 , \7199 , \7200 ,
         \7201 , \7202 , \7203 , \7204 , \7205 , \7206 , \7207 , \7208 , \7209 , \7210 ,
         \7211 , \7212 , \7213 , \7214 , \7215 , \7216 , \7217 , \7218 , \7219 , \7220 ,
         \7221 , \7222 , \7223 , \7224 , \7225 , \7226 , \7227 , \7228 , \7229 , \7230 ,
         \7231 , \7232 , \7233 , \7234 , \7235 , \7236 , \7237 , \7238 , \7239 , \7240 ,
         \7241 , \7242 , \7243 , \7244 , \7245 , \7246 , \7247 , \7248 , \7249 , \7250 ,
         \7251 , \7252 , \7253 , \7254 , \7255 , \7256 , \7257 , \7258 , \7259 , \7260 ,
         \7261 , \7262 , \7263 , \7264 , \7265 , \7266 , \7267 , \7268 , \7269 , \7270 ,
         \7271 , \7272 , \7273 , \7274 , \7275 , \7276 , \7277 , \7278 , \7279 , \7280 ,
         \7281 , \7282 , \7283 , \7284 , \7285 , \7286 , \7287 , \7288 , \7289 , \7290 ,
         \7291 , \7292 , \7293 , \7294 , \7295 , \7296 , \7297 , \7298 , \7299 , \7300 ,
         \7301 , \7302 , \7303 , \7304 , \7305 , \7306 , \7307 , \7308 , \7309 , \7310 ,
         \7311 , \7312 , \7313 , \7314 , \7315 , \7316 , \7317 , \7318 , \7319 , \7320 ,
         \7321 , \7322 , \7323 , \7324 , \7325 , \7326 , \7327 , \7328 , \7329 , \7330 ,
         \7331 , \7332 , \7333 , \7334 , \7335 , \7336 , \7337 , \7338 , \7339 , \7340 ,
         \7341 , \7342 , \7343 , \7344 , \7345 , \7346 , \7347 , \7348 , \7349 , \7350 ,
         \7351 , \7352 , \7353 , \7354 , \7355 , \7356 , \7357 , \7358 , \7359 , \7360 ,
         \7361 , \7362 , \7363 , \7364 , \7365 , \7366 , \7367 , \7368 , \7369 , \7370 ,
         \7371 , \7372 , \7373 , \7374 , \7375 , \7376 , \7377 , \7378 , \7379 , \7380 ,
         \7381 , \7382 , \7383 , \7384 , \7385 , \7386 , \7387 , \7388 , \7389 , \7390 ,
         \7391 , \7392 , \7393 , \7394 , \7395 , \7396 , \7397 , \7398 , \7399 , \7400 ,
         \7401 , \7402 , \7403 , \7404 , \7405 , \7406 , \7407 , \7408 , \7409 , \7410 ,
         \7411 , \7412 , \7413 , \7414 , \7415 , \7416 , \7417 , \7418 , \7419 , \7420 ,
         \7421 , \7422 , \7423 , \7424 , \7425 , \7426 , \7427 , \7428 , \7429 , \7430 ,
         \7431 , \7432 , \7433 , \7434 , \7435 , \7436 , \7437 , \7438 , \7439 , \7440 ,
         \7441 , \7442 , \7443 , \7444 , \7445 , \7446 , \7447 , \7448 , \7449 , \7450 ,
         \7451 , \7452 , \7453 , \7454 , \7455 , \7456 , \7457 , \7458 , \7459 , \7460 ,
         \7461 , \7462 , \7463 , \7464 , \7465 , \7466 , \7467 , \7468 , \7469 , \7470 ,
         \7471 , \7472 , \7473 , \7474 , \7475 , \7476 , \7477 , \7478 , \7479 , \7480 ,
         \7481 , \7482 , \7483 , \7484 , \7485 , \7486 , \7487 , \7488 , \7489 , \7490 ,
         \7491 , \7492 , \7493 , \7494 , \7495 , \7496 , \7497 , \7498 , \7499 , \7500 ,
         \7501 , \7502 , \7503 , \7504 , \7505 , \7506 , \7507 , \7508 , \7509 , \7510 ,
         \7511 , \7512 , \7513 , \7514 , \7515 , \7516 , \7517 , \7518 , \7519 , \7520 ,
         \7521 , \7522 , \7523 , \7524 , \7525 , \7526 , \7527 , \7528 , \7529 , \7530 ,
         \7531 , \7532 , \7533 , \7534 , \7535 , \7536 , \7537 , \7538 , \7539 , \7540 ,
         \7541 , \7542 , \7543 , \7544 , \7545 , \7546 , \7547 , \7548 , \7549 , \7550 ,
         \7551 , \7552 , \7553 , \7554 , \7555 , \7556 , \7557 , \7558 , \7559 , \7560 ,
         \7561 , \7562 , \7563 , \7564 , \7565 , \7566 , \7567 , \7568 , \7569 , \7570 ,
         \7571 , \7572 , \7573 , \7574 , \7575 , \7576 , \7577 , \7578 , \7579 , \7580 ,
         \7581 , \7582 , \7583 , \7584 , \7585 , \7586 , \7587 , \7588 , \7589 , \7590 ,
         \7591 , \7592 , \7593 , \7594 , \7595 , \7596 , \7597 , \7598 , \7599 , \7600 ,
         \7601 , \7602 , \7603 , \7604 , \7605 , \7606 , \7607 , \7608 , \7609 , \7610 ,
         \7611 , \7612 , \7613 , \7614 , \7615 , \7616 , \7617 , \7618 , \7619 , \7620 ,
         \7621 , \7622 , \7623 , \7624 , \7625 , \7626 , \7627 , \7628 , \7629 , \7630 ,
         \7631 , \7632 , \7633 , \7634 , \7635 , \7636 , \7637 , \7638 , \7639 , \7640 ,
         \7641 , \7642 , \7643 , \7644 , \7645 , \7646 , \7647 , \7648 , \7649 , \7650 ,
         \7651 , \7652 , \7653 , \7654 , \7655 , \7656 , \7657 , \7658 , \7659 , \7660 ,
         \7661 , \7662 , \7663 , \7664 , \7665 , \7666 , \7667 , \7668 , \7669 , \7670 ,
         \7671 , \7672 , \7673 , \7674 , \7675 , \7676 , \7677 , \7678 , \7679 , \7680 ,
         \7681 , \7682 , \7683 , \7684 , \7685 , \7686 , \7687 , \7688 , \7689 , \7690 ,
         \7691 , \7692 , \7693 , \7694 , \7695 , \7696 , \7697 , \7698 , \7699 , \7700 ,
         \7701 , \7702 , \7703 , \7704 , \7705 , \7706 , \7707 , \7708 , \7709 , \7710 ,
         \7711 , \7712 , \7713 , \7714 , \7715 , \7716 , \7717 , \7718 , \7719 , \7720 ,
         \7721 , \7722 , \7723 , \7724 , \7725 , \7726 , \7727 , \7728 , \7729 , \7730 ,
         \7731 , \7732 , \7733 , \7734 , \7735 , \7736 , \7737 , \7738 , \7739 , \7740 ,
         \7741 , \7742 , \7743 , \7744 , \7745 , \7746 , \7747 , \7748 , \7749 , \7750 ,
         \7751 , \7752 , \7753 , \7754 , \7755 , \7756 , \7757 , \7758 , \7759 , \7760 ,
         \7761 , \7762 , \7763 , \7764 , \7765 , \7766 , \7767 , \7768 , \7769 , \7770 ,
         \7771 , \7772 , \7773 , \7774 , \7775 , \7776 , \7777 , \7778 , \7779 , \7780 ,
         \7781 , \7782 , \7783 , \7784 , \7785 , \7786 , \7787 , \7788 , \7789 , \7790 ,
         \7791 , \7792 , \7793 , \7794 , \7795 , \7796 , \7797 , \7798 , \7799 , \7800 ,
         \7801 , \7802 , \7803 , \7804 , \7805 , \7806 , \7807 , \7808 , \7809 , \7810 ,
         \7811 , \7812 , \7813 , \7814 , \7815 , \7816 , \7817 , \7818 ;
buf \U$labaj798 ( R_41_7a88898, \7517 );
buf \U$labaj799 ( R_42_7a83a80, \7530 );
buf \U$labaj800 ( R_43_7a83bd0, \7551 );
buf \U$labaj801 ( R_44_7a87788, \7567 );
buf \U$labaj802 ( R_45_7a88be0, \7582 );
buf \U$labaj803 ( R_46_7a81ef0, \7597 );
buf \U$labaj804 ( R_47_7a889e8, \7609 );
buf \U$labaj805 ( R_48_7a84a40, \7612 );
buf \U$labaj806 ( R_49_7a882b0, \7638 );
buf \U$labaj807 ( R_4a_7a82c10, \7646 );
buf \U$labaj808 ( R_4b_7a82d60, \7657 );
buf \U$labaj809 ( R_4c_7a87b78, \7664 );
buf \U$labaj810 ( R_4d_7a84b90, \7687 );
buf \U$labaj811 ( R_4e_7a86f00, \7695 );
buf \U$labaj812 ( R_4f_7a84ce0, \7703 );
buf \U$labaj813 ( R_50_7a87440, \7715 );
buf \U$labaj814 ( R_51_7a88160, \7729 );
buf \U$labaj815 ( R_52_7a83d20, \7736 );
buf \U$labaj816 ( R_53_7a88c88, \7752 );
buf \U$labaj817 ( R_54_7a82040, \7759 );
buf \U$labaj818 ( R_55_7a84e30, \7769 );
buf \U$labaj819 ( R_56_7a876e0, \7776 );
buf \U$labaj820 ( R_57_7a87f68, \7789 );
buf \U$labaj821 ( R_58_7a82eb0, \7796 );
buf \U$labaj822 ( R_59_7a88dd8, \7799 );
buf \U$labaj823 ( R_5a_7a86e58, \7809 );
buf \U$labaj824 ( R_5b_7a83e70, \7818 );
not \U$1 ( \94 , RI8929640_33);
not \U$2 ( \95 , RI8929dc0_49);
nand \U$3 ( \96 , \94 , \95 );
not \U$4 ( \97 , \96 );
nand \U$5 ( \98 , RI8929730_35, RI8929eb0_51);
not \U$6 ( \99 , \98 );
not \U$7 ( \100 , RI8929fa0_53);
not \U$8 ( \101 , RI8929820_37);
nand \U$9 ( \102 , \100 , \101 );
not \U$10 ( \103 , \102 );
nand \U$11 ( \104 , RI8929910_39, RI892a090_55);
not \U$12 ( \105 , \104 );
not \U$13 ( \106 , RI8929a00_41);
not \U$14 ( \107 , RI892a180_57);
nand \U$15 ( \108 , \106 , \107 );
not \U$16 ( \109 , \108 );
not \U$17 ( \110 , RI8929a78_42);
not \U$18 ( \111 , RI892a1f8_58);
nand \U$19 ( \112 , \110 , \111 );
not \U$20 ( \113 , \112 );
not \U$21 ( \114 , RI8929af0_43);
not \U$22 ( \115 , RI892a270_59);
nand \U$23 ( \116 , \114 , \115 );
not \U$24 ( \117 , \116 );
not \U$25 ( \118 , RI892a2e8_60);
not \U$26 ( \119 , RI8929b68_44);
nand \U$27 ( \120 , \118 , \119 );
not \U$28 ( \121 , \120 );
nand \U$29 ( \122 , RI8929d48_48, RI892a4c8_64);
nor \U$30 ( \123 , RI8929cd0_47, RI892a450_63);
or \U$31 ( \124 , \122 , \123 );
nand \U$32 ( \125 , RI8929cd0_47, RI892a450_63);
nand \U$33 ( \126 , \124 , \125 );
and \U$34 ( \127 , RI8929c58_46, RI892a3d8_62);
or \U$35 ( \128 , \126 , \127 );
or \U$36 ( \129 , RI8929c58_46, RI892a3d8_62);
nand \U$37 ( \130 , \128 , \129 );
nand \U$38 ( \131 , RI8929be0_45, RI892a360_61);
and \U$39 ( \132 , \130 , \131 );
nor \U$40 ( \133 , RI8929be0_45, RI892a360_61);
nor \U$41 ( \134 , \132 , \133 );
not \U$42 ( \135 , \134 );
or \U$43 ( \136 , \121 , \135 );
nand \U$44 ( \137 , RI8929b68_44, RI892a2e8_60);
nand \U$45 ( \138 , \136 , \137 );
not \U$46 ( \139 , \138 );
or \U$47 ( \140 , \117 , \139 );
nand \U$48 ( \141 , RI8929af0_43, RI892a270_59);
nand \U$49 ( \142 , \140 , \141 );
not \U$50 ( \143 , \142 );
or \U$51 ( \144 , \113 , \143 );
nand \U$52 ( \145 , RI8929a78_42, RI892a1f8_58);
nand \U$53 ( \146 , \144 , \145 );
not \U$54 ( \147 , \146 );
or \U$55 ( \148 , \109 , \147 );
nand \U$56 ( \149 , RI8929a00_41, RI892a180_57);
nand \U$57 ( \150 , \148 , \149 );
not \U$58 ( \151 , RI8929988_40);
not \U$59 ( \152 , RI892a108_56);
nand \U$60 ( \153 , \151 , \152 );
and \U$61 ( \154 , \150 , \153 );
and \U$62 ( \155 , RI892a108_56, RI8929988_40);
nor \U$63 ( \156 , \154 , \155 );
not \U$64 ( \157 , \156 );
or \U$65 ( \158 , \105 , \157 );
not \U$66 ( \159 , RI8929910_39);
not \U$67 ( \160 , RI892a090_55);
nand \U$68 ( \161 , \159 , \160 );
nand \U$69 ( \162 , \158 , \161 );
nand \U$70 ( \163 , RI8929898_38, RI892a018_54);
and \U$71 ( \164 , \162 , \163 );
not \U$72 ( \165 , RI8929898_38);
not \U$73 ( \166 , RI892a018_54);
and \U$74 ( \167 , \165 , \166 );
nor \U$75 ( \168 , \164 , \167 );
not \U$76 ( \169 , \168 );
or \U$77 ( \170 , \103 , \169 );
nand \U$78 ( \171 , RI8929820_37, RI8929fa0_53);
nand \U$79 ( \172 , \170 , \171 );
not \U$80 ( \173 , RI89297a8_36);
not \U$81 ( \174 , RI8929f28_52);
nor \U$82 ( \175 , \173 , \174 );
or \U$83 ( \176 , \172 , \175 );
nand \U$84 ( \177 , \173 , \174 );
nand \U$85 ( \178 , \176 , \177 );
not \U$86 ( \179 , \178 );
or \U$87 ( \180 , \99 , \179 );
not \U$88 ( \181 , RI8929730_35);
not \U$89 ( \182 , RI8929eb0_51);
nand \U$90 ( \183 , \181 , \182 );
nand \U$91 ( \184 , \180 , \183 );
nand \U$92 ( \185 , RI89296b8_34, RI8929e38_50);
and \U$93 ( \186 , \184 , \185 );
nor \U$94 ( \187 , RI89296b8_34, RI8929e38_50);
nor \U$95 ( \188 , \186 , \187 );
not \U$96 ( \189 , \188 );
or \U$97 ( \190 , \97 , \189 );
nand \U$98 ( \191 , RI8929640_33, RI8929dc0_49);
nand \U$99 ( \192 , \190 , \191 );
not \U$100 ( \193 , \192 );
not \U$101 ( \194 , \193 );
not \U$102 ( \195 , RI8928b00_9);
xor \U$103 ( \196 , RI89293e8_28, RI8929460_29);
and \U$104 ( \197 , \196 , RI8928e48_16);
xor \U$105 ( \198 , RI8928ce0_13, RI8929550_31);
not \U$106 ( \199 , \198 );
not \U$107 ( \200 , RI8929550_31);
nor \U$108 ( \201 , \200 , RI89295c8_32);
not \U$109 ( \202 , \201 );
or \U$110 ( \203 , \199 , \202 );
xor \U$111 ( \204 , RI8928c68_12, RI8929550_31);
nand \U$112 ( \205 , \204 , RI89295c8_32);
nand \U$113 ( \206 , \203 , \205 );
xnor \U$114 ( \207 , \197 , \206 );
xor \U$115 ( \208 , RI8928dd0_15, RI8929460_29);
not \U$116 ( \209 , \208 );
not \U$117 ( \210 , RI8929460_29);
nor \U$118 ( \211 , RI89294d8_30, RI8929550_31);
not \U$119 ( \212 , \211 );
or \U$120 ( \213 , \210 , \212 );
not \U$121 ( \214 , RI8929460_29);
nand \U$122 ( \215 , \214 , RI8929550_31, RI89294d8_30);
nand \U$123 ( \216 , \213 , \215 );
not \U$124 ( \217 , \216 );
or \U$125 ( \218 , \209 , \217 );
xor \U$126 ( \219 , RI89294d8_30, RI8929550_31);
not \U$127 ( \220 , \219 );
not \U$128 ( \221 , \220 );
xor \U$129 ( \222 , RI8928d58_14, RI8929460_29);
nand \U$130 ( \223 , \221 , \222 );
nand \U$131 ( \224 , \218 , \223 );
not \U$132 ( \225 , \224 );
and \U$133 ( \226 , \207 , \225 );
not \U$134 ( \227 , \207 );
and \U$135 ( \228 , \227 , \224 );
nor \U$136 ( \229 , \226 , \228 );
xor \U$137 ( \230 , RI8928d58_14, RI8929550_31);
not \U$138 ( \231 , \230 );
not \U$139 ( \232 , \201 );
or \U$140 ( \233 , \231 , \232 );
nand \U$141 ( \234 , \198 , RI89295c8_32);
nand \U$142 ( \235 , \233 , \234 );
or \U$143 ( \236 , RI89294d8_30, RI8929550_31);
nand \U$144 ( \237 , \236 , RI8928e48_16);
not \U$145 ( \238 , \237 );
not \U$146 ( \239 , RI89294d8_30);
not \U$147 ( \240 , RI8929550_31);
or \U$148 ( \241 , \239 , \240 );
nand \U$149 ( \242 , \241 , RI8929460_29);
nor \U$150 ( \243 , \238 , \242 );
nand \U$151 ( \244 , \235 , \243 );
not \U$152 ( \245 , \244 );
nor \U$153 ( \246 , \229 , \245 );
or \U$154 ( \247 , \235 , \243 );
nand \U$155 ( \248 , \247 , \244 );
xor \U$156 ( \249 , RI8929460_29, RI8928e48_16);
and \U$157 ( \250 , \216 , \249 );
and \U$158 ( \251 , \221 , \208 );
nor \U$159 ( \252 , \250 , \251 );
nand \U$160 ( \253 , \248 , \252 );
xor \U$161 ( \254 , RI8928dd0_15, RI8929550_31);
not \U$162 ( \255 , \254 );
not \U$163 ( \256 , \201 );
or \U$164 ( \257 , \255 , \256 );
nand \U$165 ( \258 , \230 , RI89295c8_32);
nand \U$166 ( \259 , \257 , \258 );
nand \U$167 ( \260 , \221 , RI8928e48_16);
not \U$168 ( \261 , \260 );
nor \U$169 ( \262 , \259 , \261 );
not \U$170 ( \263 , RI89295c8_32);
not \U$171 ( \264 , \254 );
not \U$172 ( \265 , \264 );
or \U$173 ( \266 , \263 , \265 );
nand \U$174 ( \267 , RI8928e48_16, RI89295c8_32);
nand \U$175 ( \268 , \267 , RI8929550_31);
nor \U$176 ( \269 , \268 , RI8928e48_16);
nand \U$177 ( \270 , \266 , \269 );
or \U$178 ( \271 , \262 , \270 );
nand \U$179 ( \272 , \259 , \261 );
nand \U$180 ( \273 , \271 , \272 );
and \U$181 ( \274 , \253 , \273 );
nor \U$182 ( \275 , \248 , \252 );
nor \U$183 ( \276 , \274 , \275 );
or \U$184 ( \277 , \246 , \276 );
nand \U$185 ( \278 , \229 , \245 );
nand \U$186 ( \279 , \277 , \278 );
not \U$187 ( \280 , \279 );
xor \U$188 ( \281 , RI8928bf0_11, RI8929550_31);
not \U$189 ( \282 , \281 );
not \U$190 ( \283 , \282 );
not \U$191 ( \284 , RI89295c8_32);
not \U$192 ( \285 , \284 );
and \U$193 ( \286 , \283 , \285 );
not \U$194 ( \287 , RI8929550_31);
nor \U$195 ( \288 , \287 , RI89295c8_32);
buf \U$196 ( \289 , \288 );
and \U$197 ( \290 , \289 , \204 );
nor \U$198 ( \291 , \286 , \290 );
xor \U$199 ( \292 , RI8928e48_16, RI8929370_27);
not \U$200 ( \293 , \292 );
not \U$201 ( \294 , RI89293e8_28);
nand \U$202 ( \295 , \294 , RI8929370_27);
or \U$203 ( \296 , \295 , RI8929460_29);
not \U$204 ( \297 , RI8929370_27);
nand \U$205 ( \298 , \297 , RI89293e8_28, RI8929460_29);
nand \U$206 ( \299 , \296 , \298 );
buf \U$207 ( \300 , \299 );
not \U$208 ( \301 , \300 );
or \U$209 ( \302 , \293 , \301 );
xor \U$210 ( \303 , RI89293e8_28, RI8929460_29);
xor \U$211 ( \304 , RI8929370_27, RI8928dd0_15);
nand \U$212 ( \305 , \303 , \304 );
nand \U$213 ( \306 , \302 , \305 );
xor \U$214 ( \307 , \291 , \306 );
xor \U$215 ( \308 , RI8929460_29, RI89294d8_30);
nand \U$216 ( \309 , \308 , \222 );
or \U$217 ( \310 , \309 , \219 );
xor \U$218 ( \311 , RI8929460_29, RI8928ce0_13);
nand \U$219 ( \312 , \219 , \311 );
nand \U$220 ( \313 , \310 , \312 );
or \U$221 ( \314 , RI8928e48_16, RI89293e8_28);
nand \U$222 ( \315 , \314 , RI8929460_29);
nand \U$223 ( \316 , RI8928e48_16, RI89293e8_28);
and \U$224 ( \317 , \315 , \316 , RI8929370_27);
nor \U$225 ( \318 , \313 , \317 );
not \U$226 ( \319 , \318 );
nand \U$227 ( \320 , \313 , \317 );
nand \U$228 ( \321 , \319 , \320 );
xnor \U$229 ( \322 , \307 , \321 );
not \U$230 ( \323 , \206 );
not \U$231 ( \324 , \197 );
nand \U$232 ( \325 , \323 , \324 );
and \U$233 ( \326 , \325 , \224 );
not \U$234 ( \327 , \206 );
nor \U$235 ( \328 , \327 , \324 );
nor \U$236 ( \329 , \326 , \328 );
nand \U$237 ( \330 , \322 , \329 );
not \U$238 ( \331 , \330 );
or \U$239 ( \332 , \280 , \331 );
not \U$240 ( \333 , \329 );
not \U$241 ( \334 , \322 );
nand \U$242 ( \335 , \333 , \334 );
nand \U$243 ( \336 , \332 , \335 );
not \U$244 ( \337 , \336 );
not \U$245 ( \338 , \337 );
not \U$246 ( \339 , \281 );
not \U$247 ( \340 , \289 );
or \U$248 ( \341 , \339 , \340 );
not \U$249 ( \342 , RI8928b78_10);
and \U$250 ( \343 , RI8929550_31, \342 );
not \U$251 ( \344 , RI8929550_31);
and \U$252 ( \345 , \344 , RI8928b78_10);
or \U$253 ( \346 , \343 , \345 );
nand \U$254 ( \347 , \346 , RI89295c8_32);
nand \U$255 ( \348 , \341 , \347 );
not \U$256 ( \349 , \348 );
and \U$257 ( \350 , \320 , \349 );
not \U$258 ( \351 , \320 );
and \U$259 ( \352 , \351 , \348 );
nor \U$260 ( \353 , \350 , \352 );
not \U$261 ( \354 , \291 );
nor \U$262 ( \355 , \354 , \306 );
or \U$263 ( \356 , \355 , \321 );
not \U$264 ( \357 , \291 );
nand \U$265 ( \358 , \357 , \306 );
nand \U$266 ( \359 , \356 , \358 );
not \U$267 ( \360 , \359 );
xor \U$268 ( \361 , \353 , \360 );
not \U$269 ( \362 , \304 );
not \U$270 ( \363 , \300 );
or \U$271 ( \364 , \362 , \363 );
xor \U$272 ( \365 , RI8928d58_14, RI8929370_27);
nand \U$273 ( \366 , \365 , \303 );
nand \U$274 ( \367 , \364 , \366 );
xor \U$275 ( \368 , RI89292f8_26, RI8929370_27);
buf \U$276 ( \369 , \368 );
nand \U$277 ( \370 , \369 , RI8928e48_16);
xnor \U$278 ( \371 , \367 , \370 );
not \U$279 ( \372 , \311 );
not \U$280 ( \373 , \216 );
or \U$281 ( \374 , \372 , \373 );
not \U$282 ( \375 , RI8928c68_12);
not \U$283 ( \376 , RI8929460_29);
and \U$284 ( \377 , \375 , \376 );
and \U$285 ( \378 , RI8928c68_12, RI8929460_29);
nor \U$286 ( \379 , \377 , \378 );
nand \U$287 ( \380 , \221 , \379 );
nand \U$288 ( \381 , \374 , \380 );
buf \U$289 ( \382 , \381 );
and \U$290 ( \383 , \371 , \382 );
not \U$291 ( \384 , \371 );
not \U$292 ( \385 , \382 );
and \U$293 ( \386 , \384 , \385 );
nor \U$294 ( \387 , \383 , \386 );
xnor \U$295 ( \388 , \361 , \387 );
not \U$296 ( \389 , \388 );
or \U$297 ( \390 , \338 , \389 );
not \U$298 ( \391 , \381 );
xor \U$299 ( \392 , \391 , \353 );
xnor \U$300 ( \393 , \392 , \371 );
not \U$301 ( \394 , \393 );
nand \U$302 ( \395 , \394 , \360 );
not \U$303 ( \396 , \395 );
nand \U$304 ( \397 , \393 , \359 );
not \U$305 ( \398 , \397 );
or \U$306 ( \399 , \396 , \398 );
not \U$307 ( \400 , \337 );
nand \U$308 ( \401 , \399 , \400 );
nand \U$309 ( \402 , \390 , \401 );
not \U$310 ( \403 , \329 );
xor \U$311 ( \404 , \403 , \334 );
xnor \U$312 ( \405 , \404 , \279 );
not \U$313 ( \406 , \245 );
buf \U$314 ( \407 , \229 );
xor \U$315 ( \408 , \406 , \407 );
xnor \U$316 ( \409 , \408 , \276 );
not \U$317 ( \410 , \409 );
not \U$318 ( \411 , \275 );
nand \U$319 ( \412 , \411 , \253 );
xnor \U$320 ( \413 , \412 , \273 );
not \U$321 ( \414 , \413 );
not \U$322 ( \415 , \262 );
nand \U$323 ( \416 , \415 , \272 );
buf \U$324 ( \417 , \270 );
xor \U$325 ( \418 , \416 , \417 );
not \U$326 ( \419 , \418 );
or \U$327 ( \420 , \284 , \264 );
nand \U$328 ( \421 , \420 , \268 );
nand \U$329 ( \422 , \417 , \421 );
not \U$330 ( \423 , \422 );
not \U$331 ( \424 , \423 );
nand \U$332 ( \425 , \414 , \419 , \424 );
nor \U$333 ( \426 , \410 , \425 );
nand \U$334 ( \427 , \405 , \426 );
nor \U$335 ( \428 , \402 , \427 );
xor \U$336 ( \429 , RI8928e48_16, RI8929190_23);
not \U$337 ( \430 , \429 );
not \U$338 ( \431 , RI8929208_24);
not \U$339 ( \432 , RI8929190_23);
or \U$340 ( \433 , \431 , \432 );
or \U$341 ( \434 , RI8929190_23, RI8929208_24);
nand \U$342 ( \435 , \433 , \434 );
xor \U$343 ( \436 , RI8929208_24, RI8929280_25);
nor \U$344 ( \437 , \435 , \436 );
not \U$345 ( \438 , \437 );
or \U$346 ( \439 , \430 , \438 );
buf \U$347 ( \440 , \436 );
xor \U$348 ( \441 , RI8929190_23, RI8928dd0_15);
nand \U$349 ( \442 , \440 , \441 );
nand \U$350 ( \443 , \439 , \442 );
not \U$351 ( \444 , RI8929460_29);
not \U$352 ( \445 , \211 );
or \U$353 ( \446 , \444 , \445 );
nand \U$354 ( \447 , \446 , \215 );
xor \U$355 ( \448 , RI8928bf0_11, RI8929460_29);
and \U$356 ( \449 , \447 , \448 );
xor \U$357 ( \450 , RI8929460_29, RI8928b78_10);
and \U$358 ( \451 , \219 , \450 );
nor \U$359 ( \452 , \449 , \451 );
nand \U$360 ( \453 , \436 , RI8928e48_16);
not \U$361 ( \454 , \453 );
xor \U$362 ( \455 , RI8929550_31, RI8928b00_9);
not \U$363 ( \456 , \455 );
not \U$364 ( \457 , RI8929550_31);
nor \U$365 ( \458 , \457 , RI89295c8_32);
not \U$366 ( \459 , \458 );
or \U$367 ( \460 , \456 , \459 );
xor \U$368 ( \461 , RI8929550_31, RI8928a88_8);
nand \U$369 ( \462 , \461 , RI89295c8_32);
nand \U$370 ( \463 , \460 , \462 );
nor \U$371 ( \464 , \454 , \463 );
or \U$372 ( \465 , \452 , \464 );
buf \U$373 ( \466 , \463 );
not \U$374 ( \467 , \453 );
nand \U$375 ( \468 , \466 , \467 );
nand \U$376 ( \469 , \465 , \468 );
xor \U$377 ( \470 , \443 , \469 );
not \U$378 ( \471 , RI8929460_29);
nor \U$379 ( \472 , \471 , RI89293e8_28);
xor \U$380 ( \473 , RI8928bf0_11, RI8929370_27);
nand \U$381 ( \474 , \472 , \473 );
not \U$382 ( \475 , RI8929370_27);
nor \U$383 ( \476 , \475 , RI8929460_29);
xor \U$384 ( \477 , RI8928c68_12, RI8929370_27);
not \U$385 ( \478 , RI89293e8_28);
nand \U$386 ( \479 , \476 , \477 , \478 );
not \U$387 ( \480 , \298 );
nand \U$388 ( \481 , \480 , \477 );
not \U$389 ( \482 , RI8929460_29);
xor \U$390 ( \483 , RI8928bf0_11, RI8929370_27);
nand \U$391 ( \484 , \482 , \483 , RI89293e8_28);
nand \U$392 ( \485 , \474 , \479 , \481 , \484 );
or \U$393 ( \486 , RI8928e48_16, RI8929208_24);
nand \U$394 ( \487 , \486 , RI8929280_25);
nand \U$395 ( \488 , RI8928e48_16, RI8929208_24);
and \U$396 ( \489 , \487 , \488 , RI8929190_23);
xor \U$397 ( \490 , \485 , \489 );
and \U$398 ( \491 , \470 , \490 );
and \U$399 ( \492 , \443 , \469 );
or \U$400 ( \493 , \491 , \492 );
and \U$401 ( \494 , \437 , \441 );
xor \U$402 ( \495 , RI8929190_23, RI8928d58_14);
and \U$403 ( \496 , \495 , \436 );
nor \U$404 ( \497 , \494 , \496 );
not \U$405 ( \498 , \497 );
not \U$406 ( \499 , \498 );
xor \U$407 ( \500 , RI8928ce0_13, RI8929280_25);
not \U$408 ( \501 , \500 );
xor \U$409 ( \502 , RI8929280_25, RI89292f8_26);
not \U$410 ( \503 , \502 );
nor \U$411 ( \504 , \503 , \368 );
not \U$412 ( \505 , \504 );
or \U$413 ( \506 , \501 , \505 );
xor \U$414 ( \507 , RI8928c68_12, RI8929280_25);
nand \U$415 ( \508 , \507 , \368 );
nand \U$416 ( \509 , \506 , \508 );
not \U$417 ( \510 , \509 );
not \U$418 ( \511 , \510 );
or \U$419 ( \512 , \499 , \511 );
nand \U$420 ( \513 , \509 , \497 );
nand \U$421 ( \514 , \512 , \513 );
xor \U$422 ( \515 , RI8929460_29, RI8928b00_9);
not \U$423 ( \516 , \515 );
not \U$424 ( \517 , \216 );
or \U$425 ( \518 , \516 , \517 );
xor \U$426 ( \519 , RI8928a88_8, RI8929460_29);
nand \U$427 ( \520 , \221 , \519 );
nand \U$428 ( \521 , \518 , \520 );
xor \U$429 ( \522 , \514 , \521 );
xor \U$430 ( \523 , \493 , \522 );
xor \U$431 ( \524 , \443 , \469 );
xor \U$432 ( \525 , \524 , \490 );
not \U$433 ( \526 , \525 );
not \U$434 ( \527 , \220 );
xor \U$435 ( \528 , RI8929460_29, RI89294d8_30);
nand \U$436 ( \529 , \528 , \379 );
or \U$437 ( \530 , \527 , \529 );
nand \U$438 ( \531 , \448 , \219 );
nand \U$439 ( \532 , \530 , \531 );
or \U$440 ( \533 , RI8928e48_16, RI89292f8_26);
nand \U$441 ( \534 , \533 , RI8929370_27);
nand \U$442 ( \535 , RI8928e48_16, RI89292f8_26);
and \U$443 ( \536 , \534 , \535 , RI8929280_25);
and \U$444 ( \537 , \532 , \536 );
not \U$445 ( \538 , \537 );
xor \U$446 ( \539 , RI8928ce0_13, RI8929370_27);
not \U$447 ( \540 , \539 );
not \U$448 ( \541 , \299 );
or \U$449 ( \542 , \540 , \541 );
nand \U$450 ( \543 , \196 , \477 );
nand \U$451 ( \544 , \542 , \543 );
xor \U$452 ( \545 , RI8928dd0_15, RI8929280_25);
not \U$453 ( \546 , \545 );
not \U$454 ( \547 , \504 );
or \U$455 ( \548 , \546 , \547 );
xor \U$456 ( \549 , RI8928d58_14, RI8929280_25);
nand \U$457 ( \550 , \549 , \368 );
nand \U$458 ( \551 , \548 , \550 );
and \U$459 ( \552 , \544 , \551 );
not \U$460 ( \553 , \544 );
not \U$461 ( \554 , \551 );
and \U$462 ( \555 , \553 , \554 );
nor \U$463 ( \556 , \552 , \555 );
not \U$464 ( \557 , \556 );
or \U$465 ( \558 , \538 , \557 );
not \U$466 ( \559 , \554 );
nand \U$467 ( \560 , \559 , \544 );
nand \U$468 ( \561 , \558 , \560 );
not \U$469 ( \562 , \561 );
not \U$470 ( \563 , \461 );
not \U$471 ( \564 , \288 );
or \U$472 ( \565 , \563 , \564 );
xor \U$473 ( \566 , RI8929550_31, RI8928a10_7);
nand \U$474 ( \567 , \566 , RI89295c8_32);
nand \U$475 ( \568 , \565 , \567 );
not \U$476 ( \569 , \450 );
not \U$477 ( \570 , \447 );
or \U$478 ( \571 , \569 , \570 );
nand \U$479 ( \572 , \515 , \219 );
nand \U$480 ( \573 , \571 , \572 );
nor \U$481 ( \574 , \568 , \573 );
not \U$482 ( \575 , \574 );
nand \U$483 ( \576 , \573 , \568 );
nand \U$484 ( \577 , \575 , \576 );
not \U$485 ( \578 , \549 );
buf \U$486 ( \579 , \504 );
not \U$487 ( \580 , \579 );
or \U$488 ( \581 , \578 , \580 );
nand \U$489 ( \582 , \369 , \500 );
nand \U$490 ( \583 , \581 , \582 );
and \U$491 ( \584 , \577 , \583 );
not \U$492 ( \585 , \577 );
not \U$493 ( \586 , \583 );
and \U$494 ( \587 , \585 , \586 );
nor \U$495 ( \588 , \584 , \587 );
nand \U$496 ( \589 , \562 , \588 );
not \U$497 ( \590 , \589 );
or \U$498 ( \591 , \526 , \590 );
not \U$499 ( \592 , \588 );
nand \U$500 ( \593 , \561 , \592 );
nand \U$501 ( \594 , \591 , \593 );
not \U$502 ( \595 , \594 );
xor \U$503 ( \596 , \523 , \595 );
and \U$504 ( \597 , \485 , \489 );
buf \U$505 ( \598 , \574 );
or \U$506 ( \599 , \586 , \598 );
buf \U$507 ( \600 , \576 );
nand \U$508 ( \601 , \599 , \600 );
not \U$509 ( \602 , \601 );
xor \U$510 ( \603 , \597 , \602 );
not \U$511 ( \604 , RI8928a10_7);
not \U$512 ( \605 , \604 );
not \U$513 ( \606 , \289 );
or \U$514 ( \607 , \605 , \606 );
not \U$515 ( \608 , RI89295c8_32);
nor \U$516 ( \609 , \608 , RI8929550_31);
and \U$517 ( \610 , \609 , RI8928998_6);
nand \U$518 ( \611 , RI8929550_31, RI89295c8_32);
nor \U$519 ( \612 , \611 , RI8928998_6);
nor \U$520 ( \613 , \610 , \612 );
nand \U$521 ( \614 , \607 , \613 );
and \U$522 ( \615 , RI8929190_23, RI8929118_22);
not \U$523 ( \616 , RI8929190_23);
not \U$524 ( \617 , RI8929118_22);
and \U$525 ( \618 , \616 , \617 );
nor \U$526 ( \619 , \615 , \618 );
nand \U$527 ( \620 , \619 , RI8928e48_16);
not \U$528 ( \621 , \620 );
and \U$529 ( \622 , \614 , \621 );
not \U$530 ( \623 , \614 );
and \U$531 ( \624 , \623 , \620 );
nor \U$532 ( \625 , \622 , \624 );
not \U$533 ( \626 , \473 );
not \U$534 ( \627 , \300 );
or \U$535 ( \628 , \626 , \627 );
xor \U$536 ( \629 , RI8928b78_10, RI8929370_27);
nand \U$537 ( \630 , \303 , \629 );
nand \U$538 ( \631 , \628 , \630 );
and \U$539 ( \632 , \625 , \631 );
not \U$540 ( \633 , \625 );
not \U$541 ( \634 , \631 );
and \U$542 ( \635 , \633 , \634 );
nor \U$543 ( \636 , \632 , \635 );
xnor \U$544 ( \637 , \603 , \636 );
not \U$545 ( \638 , \637 );
xnor \U$546 ( \639 , \596 , \638 );
and \U$547 ( \640 , \561 , \588 );
not \U$548 ( \641 , \561 );
and \U$549 ( \642 , \641 , \592 );
nor \U$550 ( \643 , \640 , \642 );
not \U$551 ( \644 , \525 );
and \U$552 ( \645 , \643 , \644 );
not \U$553 ( \646 , \643 );
and \U$554 ( \647 , \646 , \525 );
nor \U$555 ( \648 , \645 , \647 );
not \U$556 ( \649 , \648 );
xor \U$557 ( \650 , \467 , \466 );
xnor \U$558 ( \651 , \650 , \452 );
and \U$559 ( \652 , RI89295c8_32, \455 );
not \U$560 ( \653 , RI89295c8_32);
not \U$561 ( \654 , RI8929550_31);
nor \U$562 ( \655 , \654 , RI8928b78_10);
and \U$563 ( \656 , \653 , \655 );
or \U$564 ( \657 , \652 , \656 );
xor \U$565 ( \658 , RI8928e48_16, RI8929280_25);
nand \U$566 ( \659 , \658 , \502 );
or \U$567 ( \660 , \659 , \368 );
nand \U$568 ( \661 , \368 , \545 );
nand \U$569 ( \662 , \660 , \661 );
and \U$570 ( \663 , \657 , \662 );
not \U$571 ( \664 , \657 );
not \U$572 ( \665 , \662 );
and \U$573 ( \666 , \664 , \665 );
nor \U$574 ( \667 , \663 , \666 );
not \U$575 ( \668 , \667 );
not \U$576 ( \669 , \365 );
not \U$577 ( \670 , \300 );
or \U$578 ( \671 , \669 , \670 );
nand \U$579 ( \672 , \303 , \539 );
nand \U$580 ( \673 , \671 , \672 );
not \U$581 ( \674 , \673 );
or \U$582 ( \675 , \668 , \674 );
not \U$583 ( \676 , \665 );
nand \U$584 ( \677 , \676 , \657 );
nand \U$585 ( \678 , \675 , \677 );
xor \U$586 ( \679 , \651 , \678 );
xor \U$587 ( \680 , \556 , \537 );
and \U$588 ( \681 , \679 , \680 );
and \U$589 ( \682 , \651 , \678 );
or \U$590 ( \683 , \681 , \682 );
not \U$591 ( \684 , \683 );
nand \U$592 ( \685 , \649 , \684 );
and \U$593 ( \686 , \639 , \685 );
not \U$594 ( \687 , \639 );
nor \U$595 ( \688 , \683 , \648 );
and \U$596 ( \689 , \687 , \688 );
nor \U$597 ( \690 , \686 , \689 );
xor \U$598 ( \691 , \532 , \536 );
not \U$599 ( \692 , \673 );
not \U$600 ( \693 , \667 );
not \U$601 ( \694 , \693 );
or \U$602 ( \695 , \692 , \694 );
not \U$603 ( \696 , \673 );
nand \U$604 ( \697 , \696 , \667 );
nand \U$605 ( \698 , \695 , \697 );
xor \U$606 ( \699 , \691 , \698 );
not \U$607 ( \700 , \367 );
nand \U$608 ( \701 , \700 , \370 );
and \U$609 ( \702 , \701 , \382 );
not \U$610 ( \703 , \367 );
nor \U$611 ( \704 , \703 , \370 );
nor \U$612 ( \705 , \702 , \704 );
xnor \U$613 ( \706 , \699 , \705 );
not \U$614 ( \707 , \706 );
nand \U$615 ( \708 , \320 , \349 );
not \U$616 ( \709 , \708 );
not \U$617 ( \710 , \387 );
or \U$618 ( \711 , \709 , \710 );
not \U$619 ( \712 , \320 );
nand \U$620 ( \713 , \712 , \348 );
nand \U$621 ( \714 , \711 , \713 );
not \U$622 ( \715 , \714 );
nand \U$623 ( \716 , \707 , \715 );
not \U$624 ( \717 , \716 );
not \U$625 ( \718 , \717 );
nand \U$626 ( \719 , \706 , \714 );
buf \U$627 ( \720 , \719 );
nand \U$628 ( \721 , \718 , \720 );
not \U$629 ( \722 , \336 );
not \U$630 ( \723 , \395 );
or \U$631 ( \724 , \722 , \723 );
nand \U$632 ( \725 , \724 , \397 );
and \U$633 ( \726 , \721 , \725 );
not \U$634 ( \727 , \721 );
not \U$635 ( \728 , \725 );
and \U$636 ( \729 , \727 , \728 );
nor \U$637 ( \730 , \726 , \729 );
nand \U$638 ( \731 , \395 , \336 );
nand \U$639 ( \732 , \731 , \719 , \397 );
or \U$640 ( \733 , \714 , \706 );
nand \U$641 ( \734 , \732 , \733 );
xor \U$642 ( \735 , \651 , \678 );
xor \U$643 ( \736 , \735 , \680 );
not \U$644 ( \737 , \705 );
not \U$645 ( \738 , \737 );
not \U$646 ( \739 , \691 );
not \U$647 ( \740 , \739 );
not \U$648 ( \741 , \698 );
or \U$649 ( \742 , \740 , \741 );
or \U$650 ( \743 , \698 , \739 );
nand \U$651 ( \744 , \742 , \743 );
not \U$652 ( \745 , \744 );
or \U$653 ( \746 , \738 , \745 );
not \U$654 ( \747 , \739 );
buf \U$655 ( \748 , \698 );
nand \U$656 ( \749 , \747 , \748 );
nand \U$657 ( \750 , \746 , \749 );
nand \U$658 ( \751 , \736 , \750 );
not \U$659 ( \752 , \751 );
nor \U$660 ( \753 , \736 , \750 );
nor \U$661 ( \754 , \752 , \753 );
xor \U$662 ( \755 , \734 , \754 );
nand \U$663 ( \756 , \428 , \690 , \730 , \755 );
not \U$664 ( \757 , \732 );
not \U$665 ( \758 , \736 );
not \U$666 ( \759 , \758 );
not \U$667 ( \760 , \750 );
not \U$668 ( \761 , \760 );
or \U$669 ( \762 , \759 , \761 );
nand \U$670 ( \763 , \762 , \716 );
not \U$671 ( \764 , \763 );
not \U$672 ( \765 , \764 );
or \U$673 ( \766 , \757 , \765 );
nand \U$674 ( \767 , \766 , \751 );
buf \U$675 ( \768 , \767 );
nand \U$676 ( \769 , \648 , \683 );
nand \U$677 ( \770 , \769 , \685 );
buf \U$678 ( \771 , \770 );
and \U$679 ( \772 , \768 , \771 );
not \U$680 ( \773 , \768 );
not \U$681 ( \774 , \771 );
and \U$682 ( \775 , \773 , \774 );
nor \U$683 ( \776 , \772 , \775 );
and \U$684 ( \777 , \756 , \776 );
not \U$685 ( \778 , \777 );
not \U$686 ( \779 , \778 );
or \U$687 ( \780 , \195 , \779 );
xnor \U$688 ( \781 , \637 , \523 );
buf \U$689 ( \782 , \595 );
nand \U$690 ( \783 , \781 , \782 );
not \U$691 ( \784 , \783 );
not \U$692 ( \785 , \395 );
not \U$693 ( \786 , \785 );
not \U$694 ( \787 , \719 );
or \U$695 ( \788 , \786 , \787 );
not \U$696 ( \789 , \336 );
nand \U$697 ( \790 , \789 , \719 , \397 );
nand \U$698 ( \791 , \788 , \790 );
nor \U$699 ( \792 , \784 , \791 , \688 , \763 );
nand \U$700 ( \793 , \783 , \685 );
and \U$701 ( \794 , \769 , \751 );
or \U$702 ( \795 , \793 , \794 );
or \U$703 ( \796 , \781 , \782 );
nand \U$704 ( \797 , \795 , \796 );
nor \U$705 ( \798 , \792 , \797 );
buf \U$706 ( \799 , \597 );
nor \U$707 ( \800 , \636 , \799 );
or \U$708 ( \801 , \800 , \602 );
nand \U$709 ( \802 , \636 , \799 );
nand \U$710 ( \803 , \801 , \802 );
not \U$711 ( \804 , \521 );
not \U$712 ( \805 , \514 );
or \U$713 ( \806 , \804 , \805 );
nand \U$714 ( \807 , \509 , \498 );
nand \U$715 ( \808 , \806 , \807 );
not \U$716 ( \809 , \634 );
nand \U$717 ( \810 , \809 , \625 );
nand \U$718 ( \811 , \614 , \621 );
nand \U$719 ( \812 , \810 , \811 );
xor \U$720 ( \813 , \808 , \812 );
not \U$721 ( \814 , \629 );
not \U$722 ( \815 , \300 );
or \U$723 ( \816 , \814 , \815 );
xor \U$724 ( \817 , RI8928b00_9, RI8929370_27);
nand \U$725 ( \818 , \303 , \817 );
nand \U$726 ( \819 , \816 , \818 );
not \U$727 ( \820 , \507 );
not \U$728 ( \821 , \579 );
or \U$729 ( \822 , \820 , \821 );
xor \U$730 ( \823 , RI8928bf0_11, RI8929280_25);
nand \U$731 ( \824 , \369 , \823 );
nand \U$732 ( \825 , \822 , \824 );
xor \U$733 ( \826 , \819 , \825 );
nor \U$734 ( \827 , \435 , \436 );
buf \U$735 ( \828 , \495 );
and \U$736 ( \829 , \827 , \828 );
xor \U$737 ( \830 , RI8929190_23, RI8928ce0_13);
and \U$738 ( \831 , \440 , \830 );
nor \U$739 ( \832 , \829 , \831 );
not \U$740 ( \833 , \832 );
not \U$741 ( \834 , RI8928998_6);
not \U$742 ( \835 , \834 );
not \U$743 ( \836 , \201 );
or \U$744 ( \837 , \835 , \836 );
not \U$745 ( \838 , \609 );
and \U$746 ( \839 , RI8928920_5, \838 );
not \U$747 ( \840 , RI8928920_5);
and \U$748 ( \841 , \840 , \611 );
or \U$749 ( \842 , \839 , \841 );
nand \U$750 ( \843 , \837 , \842 );
not \U$751 ( \844 , \843 );
and \U$752 ( \845 , \833 , \844 );
and \U$753 ( \846 , \832 , \843 );
nor \U$754 ( \847 , \845 , \846 );
xor \U$755 ( \848 , \826 , \847 );
not \U$756 ( \849 , \619 );
not \U$757 ( \850 , \849 );
xnor \U$758 ( \851 , RI8928dd0_15, RI89290a0_21);
not \U$759 ( \852 , \851 );
and \U$760 ( \853 , \850 , \852 );
not \U$761 ( \854 , RI89290a0_21);
nor \U$762 ( \855 , RI8928e48_16, RI8929118_22);
not \U$763 ( \856 , \855 );
or \U$764 ( \857 , \854 , \856 );
not \U$765 ( \858 , RI89290a0_21);
nand \U$766 ( \859 , \858 , RI8928e48_16, RI8929118_22);
nand \U$767 ( \860 , \857 , \859 );
and \U$768 ( \861 , \849 , \860 );
nor \U$769 ( \862 , \853 , \861 );
nand \U$770 ( \863 , RI8928e48_16, RI8929118_22);
nand \U$771 ( \864 , \863 , RI89290a0_21);
not \U$772 ( \865 , \864 );
or \U$773 ( \866 , RI8928e48_16, RI8929118_22);
nand \U$774 ( \867 , \866 , RI8929190_23);
nand \U$775 ( \868 , \865 , \867 );
and \U$776 ( \869 , \862 , \868 );
not \U$777 ( \870 , \862 );
not \U$778 ( \871 , \868 );
and \U$779 ( \872 , \870 , \871 );
nor \U$780 ( \873 , \869 , \872 );
not \U$781 ( \874 , \519 );
not \U$782 ( \875 , \216 );
or \U$783 ( \876 , \874 , \875 );
xor \U$784 ( \877 , RI8928a10_7, RI8929460_29);
nand \U$785 ( \878 , \221 , \877 );
nand \U$786 ( \879 , \876 , \878 );
and \U$787 ( \880 , \873 , \879 );
not \U$788 ( \881 , \873 );
not \U$789 ( \882 , \879 );
and \U$790 ( \883 , \881 , \882 );
nor \U$791 ( \884 , \880 , \883 );
and \U$792 ( \885 , \848 , \884 );
not \U$793 ( \886 , \848 );
not \U$794 ( \887 , \884 );
and \U$795 ( \888 , \886 , \887 );
nor \U$796 ( \889 , \885 , \888 );
and \U$797 ( \890 , \813 , \889 );
not \U$798 ( \891 , \813 );
not \U$799 ( \892 , \889 );
and \U$800 ( \893 , \891 , \892 );
nor \U$801 ( \894 , \890 , \893 );
xor \U$802 ( \895 , \803 , \894 );
buf \U$803 ( \896 , \522 );
buf \U$804 ( \897 , \493 );
or \U$805 ( \898 , \896 , \897 );
not \U$806 ( \899 , \898 );
not \U$807 ( \900 , \638 );
not \U$808 ( \901 , \900 );
or \U$809 ( \902 , \899 , \901 );
nand \U$810 ( \903 , \897 , \896 );
nand \U$811 ( \904 , \902 , \903 );
xor \U$812 ( \905 , \895 , \904 );
and \U$813 ( \906 , \798 , \905 );
not \U$814 ( \907 , \798 );
not \U$815 ( \908 , \905 );
and \U$816 ( \909 , \907 , \908 );
nor \U$817 ( \910 , \906 , \909 );
buf \U$818 ( \911 , \910 );
or \U$819 ( \912 , RI892a180_57, RI8928b00_9);
and \U$820 ( \913 , \911 , \912 );
not \U$821 ( \914 , RI8929cd0_47);
nor \U$822 ( \915 , \914 , RI8929d48_48);
not \U$823 ( \916 , \915 );
xor \U$824 ( \917 , RI89294d8_30, RI8929cd0_47);
not \U$825 ( \918 , \917 );
or \U$826 ( \919 , \916 , \918 );
xor \U$827 ( \920 , RI8929cd0_47, RI8929460_29);
nand \U$828 ( \921 , \920 , RI8929d48_48);
nand \U$829 ( \922 , \919 , \921 );
or \U$830 ( \923 , RI89295c8_32, RI8929c58_46);
nand \U$831 ( \924 , \923 , RI8929cd0_47);
nand \U$832 ( \925 , RI89295c8_32, RI8929c58_46);
and \U$833 ( \926 , \924 , \925 , RI8929be0_45);
nand \U$834 ( \927 , \922 , \926 );
not \U$835 ( \928 , \920 );
not \U$836 ( \929 , RI8929d48_48);
nand \U$837 ( \930 , \929 , RI8929cd0_47);
not \U$838 ( \931 , \930 );
not \U$839 ( \932 , \931 );
or \U$840 ( \933 , \928 , \932 );
xor \U$841 ( \934 , RI8929cd0_47, RI89293e8_28);
nand \U$842 ( \935 , \934 , RI8929d48_48);
nand \U$843 ( \936 , \933 , \935 );
not \U$844 ( \937 , \936 );
xnor \U$845 ( \938 , RI8929c58_46, RI8929cd0_47);
xor \U$846 ( \939 , RI8929be0_45, RI89294d8_30);
or \U$847 ( \940 , \938 , \939 );
xor \U$848 ( \941 , RI8929be0_45, RI8929c58_46);
not \U$849 ( \942 , \941 );
xor \U$850 ( \943 , RI8929550_31, RI8929be0_45);
not \U$851 ( \944 , \943 );
or \U$852 ( \945 , \942 , \944 );
xor \U$853 ( \946 , RI8929c58_46, RI8929cd0_47);
not \U$854 ( \947 , \946 );
nand \U$855 ( \948 , \945 , \947 );
nand \U$856 ( \949 , \940 , \948 );
xor \U$857 ( \950 , RI8929b68_44, RI8929be0_45);
nand \U$858 ( \951 , \950 , RI89295c8_32);
and \U$859 ( \952 , \949 , \951 );
not \U$860 ( \953 , \949 );
not \U$861 ( \954 , \951 );
and \U$862 ( \955 , \953 , \954 );
nor \U$863 ( \956 , \952 , \955 );
not \U$864 ( \957 , \956 );
or \U$865 ( \958 , \937 , \957 );
or \U$866 ( \959 , \956 , \936 );
nand \U$867 ( \960 , \958 , \959 );
xor \U$868 ( \961 , \927 , \960 );
or \U$869 ( \962 , \922 , \926 );
nand \U$870 ( \963 , \962 , \927 );
xor \U$871 ( \964 , RI89295c8_32, RI8929be0_45);
not \U$872 ( \965 , \964 );
not \U$873 ( \966 , \941 );
nor \U$874 ( \967 , \966 , \946 );
not \U$875 ( \968 , \967 );
or \U$876 ( \969 , \965 , \968 );
xor \U$877 ( \970 , RI8929c58_46, RI8929cd0_47);
nand \U$878 ( \971 , \970 , \943 );
nand \U$879 ( \972 , \969 , \971 );
not \U$880 ( \973 , \972 );
nand \U$881 ( \974 , \963 , \973 );
and \U$882 ( \975 , \970 , RI89295c8_32);
xor \U$883 ( \976 , RI8929cd0_47, RI8929550_31);
not \U$884 ( \977 , \976 );
not \U$885 ( \978 , \930 );
not \U$886 ( \979 , \978 );
or \U$887 ( \980 , \977 , \979 );
nand \U$888 ( \981 , \917 , RI8929d48_48);
nand \U$889 ( \982 , \980 , \981 );
nor \U$890 ( \983 , \975 , \982 );
not \U$891 ( \984 , \284 );
not \U$892 ( \985 , \978 );
or \U$893 ( \986 , \984 , \985 );
nand \U$894 ( \987 , \976 , RI8929d48_48);
nand \U$895 ( \988 , \986 , \987 );
nand \U$896 ( \989 , RI89295c8_32, RI8929d48_48);
and \U$897 ( \990 , \989 , RI8929cd0_47);
nand \U$898 ( \991 , \988 , \990 );
or \U$899 ( \992 , \983 , \991 );
nand \U$900 ( \993 , \975 , \982 );
nand \U$901 ( \994 , \992 , \993 );
and \U$902 ( \995 , \974 , \994 );
nor \U$903 ( \996 , \963 , \973 );
nor \U$904 ( \997 , \995 , \996 );
and \U$905 ( \998 , \961 , \997 );
and \U$906 ( \999 , \927 , \960 );
or \U$907 ( \1000 , \998 , \999 );
xor \U$908 ( \1001 , RI89295c8_32, RI8929af0_43);
not \U$909 ( \1002 , \1001 );
xnor \U$910 ( \1003 , RI8929af0_43, RI8929b68_44);
nor \U$911 ( \1004 , \1003 , \950 );
not \U$912 ( \1005 , \1004 );
or \U$913 ( \1006 , \1002 , \1005 );
buf \U$914 ( \1007 , \950 );
xor \U$915 ( \1008 , RI8929550_31, RI8929af0_43);
nand \U$916 ( \1009 , \1007 , \1008 );
nand \U$917 ( \1010 , \1006 , \1009 );
not \U$918 ( \1011 , \934 );
not \U$919 ( \1012 , \915 );
or \U$920 ( \1013 , \1011 , \1012 );
xor \U$921 ( \1014 , RI8929370_27, RI8929cd0_47);
nand \U$922 ( \1015 , \1014 , RI8929d48_48);
nand \U$923 ( \1016 , \1013 , \1015 );
or \U$924 ( \1017 , RI89295c8_32, RI8929b68_44);
nand \U$925 ( \1018 , \1017 , RI8929be0_45);
nand \U$926 ( \1019 , RI89295c8_32, RI8929b68_44);
and \U$927 ( \1020 , \1018 , \1019 , RI8929af0_43);
nand \U$928 ( \1021 , \1016 , \1020 );
not \U$929 ( \1022 , \1021 );
nor \U$930 ( \1023 , \1016 , \1020 );
nor \U$931 ( \1024 , \1022 , \1023 );
xor \U$932 ( \1025 , \1010 , \1024 );
not \U$933 ( \1026 , \939 );
not \U$934 ( \1027 , \967 );
or \U$935 ( \1028 , \1026 , \1027 );
not \U$936 ( \1029 , RI8929be0_45);
nand \U$937 ( \1030 , \1029 , RI8929460_29);
not \U$938 ( \1031 , \1030 );
not \U$939 ( \1032 , RI8929460_29);
nand \U$940 ( \1033 , \1032 , RI8929be0_45);
not \U$941 ( \1034 , \1033 );
or \U$942 ( \1035 , \1031 , \1034 );
nand \U$943 ( \1036 , \1035 , \970 );
nand \U$944 ( \1037 , \1028 , \1036 );
xor \U$945 ( \1038 , \1025 , \1037 );
buf \U$946 ( \1039 , \956 );
not \U$947 ( \1040 , \936 );
and \U$948 ( \1041 , \1039 , \1040 );
buf \U$949 ( \1042 , \949 );
and \U$950 ( \1043 , \1042 , \951 );
nor \U$951 ( \1044 , \1041 , \1043 );
nor \U$952 ( \1045 , \1038 , \1044 );
or \U$953 ( \1046 , \1000 , \1045 );
nand \U$954 ( \1047 , \1038 , \1044 );
nand \U$955 ( \1048 , \1046 , \1047 );
nand \U$956 ( \1049 , \1030 , \1033 );
not \U$957 ( \1050 , \1049 );
not \U$958 ( \1051 , \967 );
or \U$959 ( \1052 , \1050 , \1051 );
not \U$960 ( \1053 , RI8929be0_45);
nand \U$961 ( \1054 , \1053 , RI89293e8_28);
not \U$962 ( \1055 , \1054 );
not \U$963 ( \1056 , RI89293e8_28);
nand \U$964 ( \1057 , \1056 , RI8929be0_45);
not \U$965 ( \1058 , \1057 );
or \U$966 ( \1059 , \1055 , \1058 );
nand \U$967 ( \1060 , \1059 , \970 );
nand \U$968 ( \1061 , \1052 , \1060 );
not \U$969 ( \1062 , \1061 );
not \U$970 ( \1063 , \1014 );
not \U$971 ( \1064 , \915 );
or \U$972 ( \1065 , \1063 , \1064 );
xor \U$973 ( \1066 , RI89292f8_26, RI8929cd0_47);
nand \U$974 ( \1067 , \1066 , RI8929d48_48);
nand \U$975 ( \1068 , \1065 , \1067 );
xor \U$976 ( \1069 , RI8929a78_42, RI8929af0_43);
nand \U$977 ( \1070 , \1069 , RI89295c8_32);
xor \U$978 ( \1071 , \1068 , \1070 );
not \U$979 ( \1072 , \1071 );
or \U$980 ( \1073 , \1062 , \1072 );
or \U$981 ( \1074 , \1061 , \1071 );
nand \U$982 ( \1075 , \1073 , \1074 );
not \U$983 ( \1076 , \1021 );
not \U$984 ( \1077 , \1076 );
not \U$985 ( \1078 , \1008 );
buf \U$986 ( \1079 , \1004 );
not \U$987 ( \1080 , \1079 );
or \U$988 ( \1081 , \1078 , \1080 );
xor \U$989 ( \1082 , RI89294d8_30, RI8929af0_43);
nand \U$990 ( \1083 , \1007 , \1082 );
nand \U$991 ( \1084 , \1081 , \1083 );
not \U$992 ( \1085 , \1084 );
or \U$993 ( \1086 , \1077 , \1085 );
or \U$994 ( \1087 , \1084 , \1076 );
nand \U$995 ( \1088 , \1086 , \1087 );
nor \U$996 ( \1089 , \1075 , \1088 );
not \U$997 ( \1090 , \1089 );
nand \U$998 ( \1091 , \1075 , \1088 );
nand \U$999 ( \1092 , \1090 , \1091 );
xor \U$1000 ( \1093 , \1010 , \1024 );
and \U$1001 ( \1094 , \1093 , \1037 );
and \U$1002 ( \1095 , \1010 , \1024 );
or \U$1003 ( \1096 , \1094 , \1095 );
and \U$1004 ( \1097 , \1092 , \1096 );
or \U$1005 ( \1098 , \1048 , \1097 );
not \U$1006 ( \1099 , \1089 );
not \U$1007 ( \1100 , \1096 );
nand \U$1008 ( \1101 , \1099 , \1091 , \1100 );
nand \U$1009 ( \1102 , \1098 , \1101 );
buf \U$1010 ( \1103 , \1102 );
buf \U$1011 ( \1104 , \1103 );
not \U$1012 ( \1105 , \931 );
not \U$1013 ( \1106 , \1066 );
or \U$1014 ( \1107 , \1105 , \1106 );
xor \U$1015 ( \1108 , RI8929280_25, RI8929cd0_47);
nand \U$1016 ( \1109 , \1108 , RI8929d48_48);
nand \U$1017 ( \1110 , \1107 , \1109 );
not \U$1018 ( \1111 , \1110 );
or \U$1019 ( \1112 , RI89295c8_32, RI8929a78_42);
nand \U$1020 ( \1113 , \1112 , RI8929af0_43);
nand \U$1021 ( \1114 , RI89295c8_32, RI8929a78_42);
nand \U$1022 ( \1115 , \1113 , \1114 , RI8929a00_41);
nand \U$1023 ( \1116 , \1111 , \1115 );
not \U$1024 ( \1117 , \1115 );
nand \U$1025 ( \1118 , \1117 , \1110 );
nand \U$1026 ( \1119 , \1116 , \1118 );
not \U$1027 ( \1120 , \1068 );
nand \U$1028 ( \1121 , \1120 , \1070 );
not \U$1029 ( \1122 , \1121 );
not \U$1030 ( \1123 , \1061 );
or \U$1031 ( \1124 , \1122 , \1123 );
not \U$1032 ( \1125 , \1070 );
nand \U$1033 ( \1126 , \1125 , \1068 );
nand \U$1034 ( \1127 , \1124 , \1126 );
xor \U$1035 ( \1128 , \1119 , \1127 );
not \U$1036 ( \1129 , \1082 );
not \U$1037 ( \1130 , \1004 );
or \U$1038 ( \1131 , \1129 , \1130 );
xor \U$1039 ( \1132 , RI8929460_29, RI8929af0_43);
nand \U$1040 ( \1133 , \1007 , \1132 );
nand \U$1041 ( \1134 , \1131 , \1133 );
not \U$1042 ( \1135 , \1134 );
xor \U$1043 ( \1136 , RI8929a00_41, RI89295c8_32);
not \U$1044 ( \1137 , \1136 );
and \U$1045 ( \1138 , RI8929a78_42, RI8929a00_41);
not \U$1046 ( \1139 , RI8929a78_42);
and \U$1047 ( \1140 , \1139 , \106 );
nor \U$1048 ( \1141 , \1138 , \1140 );
not \U$1049 ( \1142 , \1141 );
nor \U$1050 ( \1143 , \1142 , \1069 );
not \U$1051 ( \1144 , \1143 );
or \U$1052 ( \1145 , \1137 , \1144 );
xor \U$1053 ( \1146 , RI8929a00_41, RI8929550_31);
nand \U$1054 ( \1147 , \1069 , \1146 );
nand \U$1055 ( \1148 , \1145 , \1147 );
not \U$1056 ( \1149 , \1148 );
not \U$1057 ( \1150 , \1149 );
or \U$1058 ( \1151 , \1135 , \1150 );
or \U$1059 ( \1152 , \1134 , \1149 );
nand \U$1060 ( \1153 , \1151 , \1152 );
nand \U$1061 ( \1154 , \1054 , \1057 );
not \U$1062 ( \1155 , \1154 );
buf \U$1063 ( \1156 , \967 );
not \U$1064 ( \1157 , \1156 );
or \U$1065 ( \1158 , \1155 , \1157 );
buf \U$1066 ( \1159 , \970 );
xor \U$1067 ( \1160 , RI8929370_27, RI8929be0_45);
nand \U$1068 ( \1161 , \1159 , \1160 );
nand \U$1069 ( \1162 , \1158 , \1161 );
xor \U$1070 ( \1163 , \1153 , \1162 );
xnor \U$1071 ( \1164 , \1128 , \1163 );
or \U$1072 ( \1165 , \1084 , \1076 );
not \U$1073 ( \1166 , \1165 );
not \U$1074 ( \1167 , \1075 );
or \U$1075 ( \1168 , \1166 , \1167 );
nand \U$1076 ( \1169 , \1084 , \1076 );
nand \U$1077 ( \1170 , \1168 , \1169 );
nand \U$1078 ( \1171 , \1164 , \1170 );
not \U$1079 ( \1172 , \1164 );
not \U$1080 ( \1173 , \1170 );
nand \U$1081 ( \1174 , \1172 , \1173 );
and \U$1082 ( \1175 , \1104 , \1171 , \1174 );
and \U$1083 ( \1176 , \1171 , \1174 );
nor \U$1084 ( \1177 , \1176 , \1104 );
nor \U$1085 ( \1178 , \1175 , \1177 );
not \U$1086 ( \1179 , \1178 );
buf \U$1087 ( \1180 , \730 );
not \U$1088 ( \1181 , \1180 );
and \U$1089 ( \1182 , \1179 , \1181 );
xor \U$1090 ( \1183 , RI8928d58_14, RI892a270_59);
not \U$1091 ( \1184 , \1183 );
xor \U$1092 ( \1185 , RI892a270_59, RI892a2e8_60);
not \U$1093 ( \1186 , \1185 );
xor \U$1094 ( \1187 , RI892a2e8_60, RI892a360_61);
nor \U$1095 ( \1188 , \1186 , \1187 );
not \U$1096 ( \1189 , \1188 );
or \U$1097 ( \1190 , \1184 , \1189 );
xor \U$1098 ( \1191 , RI8928ce0_13, RI892a270_59);
nand \U$1099 ( \1192 , \1187 , \1191 );
nand \U$1100 ( \1193 , \1190 , \1192 );
xor \U$1101 ( \1194 , RI892a180_57, RI8928e48_16);
not \U$1102 ( \1195 , \1194 );
not \U$1103 ( \1196 , RI892a1f8_58);
not \U$1104 ( \1197 , RI892a180_57);
or \U$1105 ( \1198 , \1196 , \1197 );
or \U$1106 ( \1199 , RI892a180_57, RI892a1f8_58);
nand \U$1107 ( \1200 , \1198 , \1199 );
xor \U$1108 ( \1201 , RI892a1f8_58, RI892a270_59);
nor \U$1109 ( \1202 , \1200 , \1201 );
buf \U$1110 ( \1203 , \1202 );
not \U$1111 ( \1204 , \1203 );
or \U$1112 ( \1205 , \1195 , \1204 );
not \U$1113 ( \1206 , \1201 );
not \U$1114 ( \1207 , \1206 );
xor \U$1115 ( \1208 , RI892a180_57, RI8928dd0_15);
nand \U$1116 ( \1209 , \1207 , \1208 );
nand \U$1117 ( \1210 , \1205 , \1209 );
and \U$1118 ( \1211 , \1193 , \1210 );
not \U$1119 ( \1212 , \1193 );
not \U$1120 ( \1213 , \1210 );
and \U$1121 ( \1214 , \1212 , \1213 );
nor \U$1122 ( \1215 , \1211 , \1214 );
xor \U$1123 ( \1216 , RI8928c68_12, RI892a360_61);
not \U$1124 ( \1217 , \1216 );
xor \U$1125 ( \1218 , RI892a3d8_62, RI892a360_61);
not \U$1126 ( \1219 , \1218 );
xor \U$1127 ( \1220 , RI892a3d8_62, RI892a450_63);
nor \U$1128 ( \1221 , \1219 , \1220 );
not \U$1129 ( \1222 , \1221 );
or \U$1130 ( \1223 , \1217 , \1222 );
buf \U$1131 ( \1224 , \1220 );
xor \U$1132 ( \1225 , RI8928bf0_11, RI892a360_61);
nand \U$1133 ( \1226 , \1224 , \1225 );
nand \U$1134 ( \1227 , \1223 , \1226 );
xnor \U$1135 ( \1228 , \1215 , \1227 );
not \U$1136 ( \1229 , \1228 );
xor \U$1137 ( \1230 , RI892a270_59, RI8928dd0_15);
and \U$1138 ( \1231 , \1188 , \1230 );
buf \U$1139 ( \1232 , \1187 );
and \U$1140 ( \1233 , \1232 , \1183 );
nor \U$1141 ( \1234 , \1231 , \1233 );
not \U$1142 ( \1235 , \1234 );
xor \U$1143 ( \1236 , RI892a450_63, RI8928c68_12);
not \U$1144 ( \1237 , \1236 );
not \U$1145 ( \1238 , RI892a450_63);
nor \U$1146 ( \1239 , \1238 , RI892a4c8_64);
not \U$1147 ( \1240 , \1239 );
or \U$1148 ( \1241 , \1237 , \1240 );
xor \U$1149 ( \1242 , RI8928bf0_11, RI892a450_63);
nand \U$1150 ( \1243 , \1242 , RI892a4c8_64);
nand \U$1151 ( \1244 , \1241 , \1243 );
or \U$1152 ( \1245 , RI8928e48_16, RI892a2e8_60);
nand \U$1153 ( \1246 , \1245 , RI892a360_61);
nand \U$1154 ( \1247 , RI8928e48_16, RI892a2e8_60);
and \U$1155 ( \1248 , \1246 , \1247 , RI892a270_59);
nand \U$1156 ( \1249 , \1244 , \1248 );
buf \U$1157 ( \1250 , \1249 );
not \U$1158 ( \1251 , \1250 );
or \U$1159 ( \1252 , \1235 , \1251 );
xor \U$1160 ( \1253 , RI8928ce0_13, RI892a360_61);
not \U$1161 ( \1254 , \1253 );
not \U$1162 ( \1255 , \1218 );
not \U$1163 ( \1256 , \1220 );
not \U$1164 ( \1257 , \1256 );
nor \U$1165 ( \1258 , \1255 , \1257 );
not \U$1166 ( \1259 , \1258 );
or \U$1167 ( \1260 , \1254 , \1259 );
nand \U$1168 ( \1261 , \1257 , \1216 );
nand \U$1169 ( \1262 , \1260 , \1261 );
not \U$1170 ( \1263 , \1239 );
not \U$1171 ( \1264 , \1242 );
or \U$1172 ( \1265 , \1263 , \1264 );
xor \U$1173 ( \1266 , RI8928b78_10, RI892a450_63);
nand \U$1174 ( \1267 , \1266 , RI892a4c8_64);
nand \U$1175 ( \1268 , \1265 , \1267 );
not \U$1176 ( \1269 , \1268 );
not \U$1177 ( \1270 , \1269 );
nand \U$1178 ( \1271 , \1201 , RI8928e48_16);
not \U$1179 ( \1272 , \1271 );
not \U$1180 ( \1273 , \1272 );
or \U$1181 ( \1274 , \1270 , \1273 );
nand \U$1182 ( \1275 , \1268 , \1271 );
nand \U$1183 ( \1276 , \1274 , \1275 );
xor \U$1184 ( \1277 , \1262 , \1276 );
nand \U$1185 ( \1278 , \1252 , \1277 );
or \U$1186 ( \1279 , \1234 , \1250 );
and \U$1187 ( \1280 , \1278 , \1279 );
xor \U$1188 ( \1281 , \1229 , \1280 );
not \U$1189 ( \1282 , \1269 );
not \U$1190 ( \1283 , \1271 );
and \U$1191 ( \1284 , \1282 , \1283 );
and \U$1192 ( \1285 , \1276 , \1262 );
nor \U$1193 ( \1286 , \1284 , \1285 );
not \U$1194 ( \1287 , \1286 );
not \U$1195 ( \1288 , \1266 );
not \U$1196 ( \1289 , RI892a450_63);
nor \U$1197 ( \1290 , \1289 , RI892a4c8_64);
buf \U$1198 ( \1291 , \1290 );
not \U$1199 ( \1292 , \1291 );
or \U$1200 ( \1293 , \1288 , \1292 );
xor \U$1201 ( \1294 , RI8928b00_9, RI892a450_63);
nand \U$1202 ( \1295 , \1294 , RI892a4c8_64);
nand \U$1203 ( \1296 , \1293 , \1295 );
or \U$1204 ( \1297 , RI8928e48_16, RI892a1f8_58);
nand \U$1205 ( \1298 , \1297 , RI892a270_59);
nand \U$1206 ( \1299 , RI8928e48_16, RI892a1f8_58);
and \U$1207 ( \1300 , \1298 , \1299 , RI892a180_57);
nand \U$1208 ( \1301 , \1296 , \1300 );
not \U$1209 ( \1302 , \1301 );
nor \U$1210 ( \1303 , \1296 , \1300 );
nor \U$1211 ( \1304 , \1302 , \1303 );
not \U$1212 ( \1305 , \1304 );
or \U$1213 ( \1306 , \1287 , \1305 );
or \U$1214 ( \1307 , \1304 , \1286 );
nand \U$1215 ( \1308 , \1306 , \1307 );
xor \U$1216 ( \1309 , \1281 , \1308 );
not \U$1217 ( \1310 , \1277 );
not \U$1218 ( \1311 , \1249 );
not \U$1219 ( \1312 , \1234 );
or \U$1220 ( \1313 , \1311 , \1312 );
or \U$1221 ( \1314 , \1250 , \1234 );
nand \U$1222 ( \1315 , \1313 , \1314 );
not \U$1223 ( \1316 , \1315 );
and \U$1224 ( \1317 , \1310 , \1316 );
and \U$1225 ( \1318 , \1277 , \1315 );
nor \U$1226 ( \1319 , \1317 , \1318 );
xor \U$1227 ( \1320 , RI8928e48_16, RI892a270_59);
nand \U$1228 ( \1321 , \1185 , \1320 );
not \U$1229 ( \1322 , \1321 );
not \U$1230 ( \1323 , \1187 );
and \U$1231 ( \1324 , \1322 , \1323 );
and \U$1232 ( \1325 , \1187 , \1230 );
nor \U$1233 ( \1326 , \1324 , \1325 );
xor \U$1234 ( \1327 , RI892a360_61, RI8928d58_14);
not \U$1235 ( \1328 , \1327 );
not \U$1236 ( \1329 , \1258 );
or \U$1237 ( \1330 , \1328 , \1329 );
nand \U$1238 ( \1331 , \1220 , \1253 );
nand \U$1239 ( \1332 , \1330 , \1331 );
not \U$1240 ( \1333 , \1332 );
xor \U$1241 ( \1334 , \1326 , \1333 );
or \U$1242 ( \1335 , \1244 , \1248 );
nand \U$1243 ( \1336 , \1335 , \1249 );
and \U$1244 ( \1337 , \1334 , \1336 );
and \U$1245 ( \1338 , \1326 , \1333 );
or \U$1246 ( \1339 , \1337 , \1338 );
nand \U$1247 ( \1340 , \1319 , \1339 );
not \U$1248 ( \1341 , \1340 );
xor \U$1249 ( \1342 , \1326 , \1333 );
xor \U$1250 ( \1343 , \1342 , \1336 );
not \U$1251 ( \1344 , RI892a450_63);
not \U$1252 ( \1345 , RI8928ce0_13);
not \U$1253 ( \1346 , \1345 );
or \U$1254 ( \1347 , \1344 , \1346 );
not \U$1255 ( \1348 , RI892a450_63);
nand \U$1256 ( \1349 , \1348 , RI8928ce0_13);
nand \U$1257 ( \1350 , \1347 , \1349 );
not \U$1258 ( \1351 , \1350 );
not \U$1259 ( \1352 , \1291 );
or \U$1260 ( \1353 , \1351 , \1352 );
nand \U$1261 ( \1354 , \1236 , RI892a4c8_64);
nand \U$1262 ( \1355 , \1353 , \1354 );
not \U$1263 ( \1356 , \1355 );
not \U$1264 ( \1357 , \1356 );
or \U$1265 ( \1358 , \1256 , \1327 );
not \U$1266 ( \1359 , \1218 );
xor \U$1267 ( \1360 , RI8928dd0_15, RI892a360_61);
not \U$1268 ( \1361 , \1360 );
or \U$1269 ( \1362 , \1359 , \1361 );
nand \U$1270 ( \1363 , \1362 , \1256 );
nand \U$1271 ( \1364 , \1358 , \1363 );
nand \U$1272 ( \1365 , \1187 , RI8928e48_16);
and \U$1273 ( \1366 , \1364 , \1365 );
not \U$1274 ( \1367 , \1364 );
not \U$1275 ( \1368 , \1365 );
and \U$1276 ( \1369 , \1367 , \1368 );
nor \U$1277 ( \1370 , \1366 , \1369 );
not \U$1278 ( \1371 , \1370 );
or \U$1279 ( \1372 , \1357 , \1371 );
not \U$1280 ( \1373 , \1368 );
nand \U$1281 ( \1374 , \1373 , \1364 );
nand \U$1282 ( \1375 , \1372 , \1374 );
nand \U$1283 ( \1376 , \1343 , \1375 );
not \U$1284 ( \1377 , \1376 );
xor \U$1285 ( \1378 , RI8928d58_14, RI892a450_63);
not \U$1286 ( \1379 , \1378 );
not \U$1287 ( \1380 , \1239 );
or \U$1288 ( \1381 , \1379 , \1380 );
nand \U$1289 ( \1382 , \1350 , RI892a4c8_64);
nand \U$1290 ( \1383 , \1381 , \1382 );
or \U$1291 ( \1384 , RI8928e48_16, RI892a3d8_62);
nand \U$1292 ( \1385 , \1384 , RI892a450_63);
nand \U$1293 ( \1386 , RI8928e48_16, RI892a3d8_62);
and \U$1294 ( \1387 , \1385 , \1386 , RI892a360_61);
nand \U$1295 ( \1388 , \1383 , \1387 );
not \U$1296 ( \1389 , \1388 );
not \U$1297 ( \1390 , \1355 );
not \U$1298 ( \1391 , \1370 );
or \U$1299 ( \1392 , \1390 , \1391 );
or \U$1300 ( \1393 , \1355 , \1370 );
nand \U$1301 ( \1394 , \1392 , \1393 );
not \U$1302 ( \1395 , \1394 );
or \U$1303 ( \1396 , \1389 , \1395 );
xor \U$1304 ( \1397 , RI8928e48_16, RI892a360_61);
not \U$1305 ( \1398 , \1397 );
not \U$1306 ( \1399 , \1258 );
or \U$1307 ( \1400 , \1398 , \1399 );
nand \U$1308 ( \1401 , \1257 , \1360 );
nand \U$1309 ( \1402 , \1400 , \1401 );
not \U$1310 ( \1403 , \1402 );
nor \U$1311 ( \1404 , \1383 , \1387 );
not \U$1312 ( \1405 , \1404 );
nand \U$1313 ( \1406 , \1405 , \1388 );
nand \U$1314 ( \1407 , \1403 , \1406 );
not \U$1315 ( \1408 , \1407 );
and \U$1316 ( \1409 , \1257 , RI8928e48_16);
xor \U$1317 ( \1410 , RI8928dd0_15, RI892a450_63);
not \U$1318 ( \1411 , \1410 );
not \U$1319 ( \1412 , \1239 );
or \U$1320 ( \1413 , \1411 , \1412 );
nand \U$1321 ( \1414 , \1378 , RI892a4c8_64);
nand \U$1322 ( \1415 , \1413 , \1414 );
nor \U$1323 ( \1416 , \1409 , \1415 );
not \U$1324 ( \1417 , RI8928e48_16);
not \U$1325 ( \1418 , \1417 );
not \U$1326 ( \1419 , \1291 );
or \U$1327 ( \1420 , \1418 , \1419 );
nand \U$1328 ( \1421 , \1410 , RI892a4c8_64);
nand \U$1329 ( \1422 , \1420 , \1421 );
nand \U$1330 ( \1423 , RI8928e48_16, RI892a4c8_64);
and \U$1331 ( \1424 , \1423 , RI892a450_63);
nand \U$1332 ( \1425 , \1422 , \1424 );
or \U$1333 ( \1426 , \1416 , \1425 );
nand \U$1334 ( \1427 , \1415 , \1409 );
nand \U$1335 ( \1428 , \1426 , \1427 );
not \U$1336 ( \1429 , \1428 );
or \U$1337 ( \1430 , \1408 , \1429 );
not \U$1338 ( \1431 , \1404 );
nand \U$1339 ( \1432 , \1431 , \1388 , \1402 );
nand \U$1340 ( \1433 , \1430 , \1432 );
nand \U$1341 ( \1434 , \1396 , \1433 );
not \U$1342 ( \1435 , \1394 );
not \U$1343 ( \1436 , \1388 );
nand \U$1344 ( \1437 , \1435 , \1436 );
nand \U$1345 ( \1438 , \1434 , \1437 );
not \U$1346 ( \1439 , \1438 );
or \U$1347 ( \1440 , \1377 , \1439 );
not \U$1348 ( \1441 , \1343 );
not \U$1349 ( \1442 , \1375 );
nand \U$1350 ( \1443 , \1441 , \1442 );
nand \U$1351 ( \1444 , \1440 , \1443 );
not \U$1352 ( \1445 , \1444 );
or \U$1353 ( \1446 , \1341 , \1445 );
not \U$1354 ( \1447 , \1319 );
not \U$1355 ( \1448 , \1339 );
nand \U$1356 ( \1449 , \1447 , \1448 );
nand \U$1357 ( \1450 , \1446 , \1449 );
buf \U$1358 ( \1451 , \1450 );
xor \U$1359 ( \1452 , \1309 , \1451 );
not \U$1360 ( \1453 , \402 );
or \U$1361 ( \1454 , \1452 , \1453 );
nor \U$1362 ( \1455 , RI89294d8_30, RI892a3d8_62);
not \U$1363 ( \1456 , \1455 );
not \U$1364 ( \1457 , \1456 );
nor \U$1365 ( \1458 , RI8929550_31, RI892a450_63);
nand \U$1366 ( \1459 , RI89295c8_32, RI892a4c8_64);
nor \U$1367 ( \1460 , \1458 , \1459 );
not \U$1368 ( \1461 , \1460 );
or \U$1369 ( \1462 , \1457 , \1461 );
and \U$1370 ( \1463 , RI8929550_31, RI892a450_63);
and \U$1371 ( \1464 , \1456 , \1463 );
and \U$1372 ( \1465 , RI89294d8_30, RI892a3d8_62);
nor \U$1373 ( \1466 , \1464 , \1465 );
nand \U$1374 ( \1467 , \1462 , \1466 );
and \U$1375 ( \1468 , RI8929460_29, RI892a360_61);
nor \U$1376 ( \1469 , \1467 , \1468 );
nor \U$1377 ( \1470 , RI8929460_29, RI892a360_61);
nor \U$1378 ( \1471 , RI89293e8_28, RI892a2e8_60);
or \U$1379 ( \1472 , \1470 , \1471 );
or \U$1380 ( \1473 , \1469 , \1472 );
nand \U$1381 ( \1474 , RI89293e8_28, RI892a2e8_60);
nand \U$1382 ( \1475 , \1473 , \1474 );
or \U$1383 ( \1476 , RI8929370_27, RI892a270_59);
and \U$1384 ( \1477 , \1475 , \1476 );
and \U$1385 ( \1478 , RI8929370_27, RI892a270_59);
nor \U$1386 ( \1479 , \1477 , \1478 );
nor \U$1387 ( \1480 , RI89292f8_26, RI892a1f8_58);
or \U$1388 ( \1481 , \1479 , \1480 );
nand \U$1389 ( \1482 , RI89292f8_26, RI892a1f8_58);
nand \U$1390 ( \1483 , \1481 , \1482 );
not \U$1391 ( \1484 , \1483 );
nor \U$1392 ( \1485 , RI8929280_25, RI892a180_57);
not \U$1393 ( \1486 , \1485 );
nand \U$1394 ( \1487 , RI8929280_25, RI892a180_57);
nand \U$1395 ( \1488 , \1486 , \1487 );
not \U$1396 ( \1489 , \1488 );
and \U$1397 ( \1490 , \1484 , \1489 );
and \U$1398 ( \1491 , \1483 , \1488 );
nor \U$1399 ( \1492 , \1490 , \1491 );
nor \U$1400 ( \1493 , \405 , \1492 );
nor \U$1401 ( \1494 , RI8928b78_10, RI8929a78_42);
not \U$1402 ( \1495 , \1494 );
not \U$1403 ( \1496 , \1495 );
nor \U$1404 ( \1497 , RI8928bf0_11, RI8929af0_43);
not \U$1405 ( \1498 , \1497 );
not \U$1406 ( \1499 , \1498 );
nor \U$1407 ( \1500 , RI8928c68_12, RI8929b68_44);
nor \U$1408 ( \1501 , RI8928ce0_13, RI8929be0_45);
nor \U$1409 ( \1502 , \1500 , \1501 );
not \U$1410 ( \1503 , \1502 );
nor \U$1411 ( \1504 , RI8928dd0_15, RI8929cd0_47);
nand \U$1412 ( \1505 , RI8928e48_16, RI8929d48_48);
or \U$1413 ( \1506 , \1504 , \1505 );
nand \U$1414 ( \1507 , RI8928dd0_15, RI8929cd0_47);
nand \U$1415 ( \1508 , \1506 , \1507 );
or \U$1416 ( \1509 , RI8928d58_14, RI8929c58_46);
and \U$1417 ( \1510 , \1508 , \1509 );
and \U$1418 ( \1511 , RI8928d58_14, RI8929c58_46);
nor \U$1419 ( \1512 , \1510 , \1511 );
nand \U$1420 ( \1513 , RI8928ce0_13, RI8929be0_45);
nand \U$1421 ( \1514 , \1512 , \1513 );
not \U$1422 ( \1515 , \1514 );
or \U$1423 ( \1516 , \1503 , \1515 );
nand \U$1424 ( \1517 , RI8928c68_12, RI8929b68_44);
nand \U$1425 ( \1518 , \1516 , \1517 );
not \U$1426 ( \1519 , \1518 );
or \U$1427 ( \1520 , \1499 , \1519 );
nand \U$1428 ( \1521 , RI8928bf0_11, RI8929af0_43);
nand \U$1429 ( \1522 , \1520 , \1521 );
not \U$1430 ( \1523 , \1522 );
or \U$1431 ( \1524 , \1496 , \1523 );
nand \U$1432 ( \1525 , RI8928b78_10, RI8929a78_42);
nand \U$1433 ( \1526 , \1524 , \1525 );
and \U$1434 ( \1527 , RI8928b00_9, RI8929a00_41);
nor \U$1435 ( \1528 , RI8928b00_9, RI8929a00_41);
nor \U$1436 ( \1529 , \1527 , \1528 );
not \U$1437 ( \1530 , \1529 );
and \U$1438 ( \1531 , \1526 , \1530 );
not \U$1439 ( \1532 , \1526 );
and \U$1440 ( \1533 , \1532 , \1529 );
nor \U$1441 ( \1534 , \1531 , \1533 );
or \U$1442 ( \1535 , \409 , \1534 );
and \U$1443 ( \1536 , \413 , RI892a180_57);
or \U$1444 ( \1537 , \419 , \106 );
not \U$1445 ( \1538 , RI8929280_25);
or \U$1446 ( \1539 , \422 , \1538 );
nand \U$1447 ( \1540 , \1537 , \1539 );
nor \U$1448 ( \1541 , \1536 , \1540 );
nand \U$1449 ( \1542 , \1535 , \1541 );
nor \U$1450 ( \1543 , \1493 , \1542 );
nand \U$1451 ( \1544 , \1454 , \1543 );
nor \U$1452 ( \1545 , \1182 , \1544 );
not \U$1453 ( \1546 , \770 );
xor \U$1454 ( \1547 , \767 , \1546 );
nand \U$1455 ( \1548 , \1547 , RI8929280_25);
not \U$1456 ( \1549 , \755 );
or \U$1457 ( \1550 , \106 , RI892a180_57);
or \U$1458 ( \1551 , \107 , RI8929a00_41);
nand \U$1459 ( \1552 , \1550 , \1551 );
nand \U$1460 ( \1553 , \1549 , \1552 );
not \U$1461 ( \1554 , \690 );
and \U$1462 ( \1555 , RI8929a00_41, RI8929280_25);
nand \U$1463 ( \1556 , \1554 , \1555 );
nand \U$1464 ( \1557 , \1545 , \1548 , \1553 , \1556 );
nor \U$1465 ( \1558 , \913 , \1557 );
nand \U$1466 ( \1559 , \780 , \1558 );
not \U$1467 ( \1560 , \1559 );
buf \U$1468 ( \1561 , \1560 );
not \U$1469 ( \1562 , \1561 );
not \U$1470 ( \1563 , \1562 );
or \U$1471 ( \1564 , \194 , \1563 );
or \U$1472 ( \1565 , \193 , \1562 );
nand \U$1473 ( \1566 , \1564 , \1565 );
not \U$1474 ( \1567 , \1566 );
not \U$1475 ( \1568 , RI8928b78_10);
not \U$1476 ( \1569 , \756 );
nor \U$1477 ( \1570 , \1569 , \910 );
not \U$1478 ( \1571 , \1570 );
not \U$1479 ( \1572 , \1571 );
or \U$1480 ( \1573 , \1568 , \1572 );
not \U$1481 ( \1574 , RI892a1f8_58);
buf \U$1482 ( \1575 , \910 );
not \U$1483 ( \1576 , \1575 );
or \U$1484 ( \1577 , \1574 , \1576 );
not \U$1485 ( \1578 , RI89292f8_26);
nor \U$1486 ( \1579 , \1578 , \110 );
nand \U$1487 ( \1580 , \1554 , \1579 );
nand \U$1488 ( \1581 , \1578 , \342 );
nand \U$1489 ( \1582 , \1547 , \1581 );
or \U$1490 ( \1583 , \110 , RI892a1f8_58);
or \U$1491 ( \1584 , \111 , RI8929a78_42);
nand \U$1492 ( \1585 , \1583 , \1584 );
nand \U$1493 ( \1586 , \1549 , \1585 );
not \U$1494 ( \1587 , \1180 );
not \U$1495 ( \1588 , \1097 );
nand \U$1496 ( \1589 , \1588 , \1101 );
buf \U$1497 ( \1590 , \1048 );
xnor \U$1498 ( \1591 , \1589 , \1590 );
and \U$1499 ( \1592 , \1587 , \1591 );
nand \U$1500 ( \1593 , \1479 , \1482 );
or \U$1501 ( \1594 , \1593 , \1480 );
not \U$1502 ( \1595 , \1482 );
nor \U$1503 ( \1596 , \1595 , \1480 );
or \U$1504 ( \1597 , \1479 , \1596 );
nand \U$1505 ( \1598 , \1594 , \1597 );
not \U$1506 ( \1599 , \1598 );
not \U$1507 ( \1600 , \405 );
not \U$1508 ( \1601 , \1600 );
or \U$1509 ( \1602 , \1599 , \1601 );
not \U$1510 ( \1603 , \1525 );
nor \U$1511 ( \1604 , \1603 , \1522 );
nand \U$1512 ( \1605 , \1604 , \1495 );
not \U$1513 ( \1606 , \1525 );
not \U$1514 ( \1607 , \1495 );
or \U$1515 ( \1608 , \1606 , \1607 );
nand \U$1516 ( \1609 , \1608 , \1522 );
nand \U$1517 ( \1610 , \1605 , \1609 );
not \U$1518 ( \1611 , \1610 );
not \U$1519 ( \1612 , \410 );
or \U$1520 ( \1613 , \1611 , \1612 );
and \U$1521 ( \1614 , \413 , RI892a1f8_58);
or \U$1522 ( \1615 , \419 , \110 );
or \U$1523 ( \1616 , \422 , \1578 );
nand \U$1524 ( \1617 , \1615 , \1616 );
nor \U$1525 ( \1618 , \1614 , \1617 );
nand \U$1526 ( \1619 , \1613 , \1618 );
not \U$1527 ( \1620 , \1619 );
nand \U$1528 ( \1621 , \1602 , \1620 );
not \U$1529 ( \1622 , \1621 );
xor \U$1530 ( \1623 , \1315 , \1448 );
xnor \U$1531 ( \1624 , \1623 , \1277 );
not \U$1532 ( \1625 , \1444 );
and \U$1533 ( \1626 , \1624 , \1625 );
not \U$1534 ( \1627 , \1624 );
and \U$1535 ( \1628 , \1627 , \1444 );
nor \U$1536 ( \1629 , \1626 , \1628 );
not \U$1537 ( \1630 , \1629 );
nand \U$1538 ( \1631 , \1630 , \402 );
nand \U$1539 ( \1632 , \1622 , \1631 );
nor \U$1540 ( \1633 , \1592 , \1632 );
and \U$1541 ( \1634 , \1580 , \1582 , \1586 , \1633 );
nand \U$1542 ( \1635 , \1577 , \1634 );
not \U$1543 ( \1636 , \1635 );
nand \U$1544 ( \1637 , \1573 , \1636 );
buf \U$1545 ( \1638 , \1569 );
and \U$1546 ( \1639 , \1638 , RI8928bf0_11);
not \U$1547 ( \1640 , RI8929370_27);
not \U$1548 ( \1641 , RI8928bf0_11);
nand \U$1549 ( \1642 , \1640 , \1641 );
nand \U$1550 ( \1643 , \1547 , \1642 );
not \U$1551 ( \1644 , \690 );
nand \U$1552 ( \1645 , \1644 , RI8929af0_43, RI8929370_27);
or \U$1553 ( \1646 , \114 , RI892a270_59);
or \U$1554 ( \1647 , \115 , RI8929af0_43);
nand \U$1555 ( \1648 , \1646 , \1647 );
nand \U$1556 ( \1649 , \1549 , \1648 );
not \U$1557 ( \1650 , \1180 );
buf \U$1558 ( \1651 , \1000 );
not \U$1559 ( \1652 , \1651 );
not \U$1560 ( \1653 , \1047 );
nor \U$1561 ( \1654 , \1653 , \1045 );
not \U$1562 ( \1655 , \1654 );
or \U$1563 ( \1656 , \1652 , \1655 );
or \U$1564 ( \1657 , \1654 , \1651 );
nand \U$1565 ( \1658 , \1656 , \1657 );
and \U$1566 ( \1659 , \1650 , \1658 );
not \U$1567 ( \1660 , \402 );
xor \U$1568 ( \1661 , \1441 , \1442 );
xor \U$1569 ( \1662 , \1661 , \1438 );
not \U$1570 ( \1663 , \1662 );
or \U$1571 ( \1664 , \1660 , \1663 );
not \U$1572 ( \1665 , \1478 );
nand \U$1573 ( \1666 , \1665 , \1476 );
not \U$1574 ( \1667 , \1666 );
not \U$1575 ( \1668 , \1470 );
and \U$1576 ( \1669 , \1467 , \1668 );
nor \U$1577 ( \1670 , \1669 , \1468 );
or \U$1578 ( \1671 , \1670 , \1471 );
nand \U$1579 ( \1672 , \1671 , \1474 );
not \U$1580 ( \1673 , \1672 );
or \U$1581 ( \1674 , \1667 , \1673 );
or \U$1582 ( \1675 , \1672 , \1666 );
nand \U$1583 ( \1676 , \1674 , \1675 );
and \U$1584 ( \1677 , \1600 , \1676 );
buf \U$1585 ( \1678 , \409 );
not \U$1586 ( \1679 , \1512 );
not \U$1587 ( \1680 , \1501 );
and \U$1588 ( \1681 , \1679 , \1680 );
not \U$1589 ( \1682 , \1513 );
nor \U$1590 ( \1683 , \1681 , \1682 );
or \U$1591 ( \1684 , \1683 , \1500 );
nand \U$1592 ( \1685 , \1684 , \1517 );
not \U$1593 ( \1686 , \1685 );
nand \U$1594 ( \1687 , \1498 , \1521 );
not \U$1595 ( \1688 , \1687 );
and \U$1596 ( \1689 , \1686 , \1688 );
and \U$1597 ( \1690 , \1685 , \1687 );
nor \U$1598 ( \1691 , \1689 , \1690 );
or \U$1599 ( \1692 , \1678 , \1691 );
and \U$1600 ( \1693 , \413 , RI892a270_59);
and \U$1601 ( \1694 , \418 , RI8929af0_43);
and \U$1602 ( \1695 , \423 , RI8929370_27);
nor \U$1603 ( \1696 , \1693 , \1694 , \1695 );
nand \U$1604 ( \1697 , \1692 , \1696 );
nor \U$1605 ( \1698 , \1677 , \1697 );
nand \U$1606 ( \1699 , \1664 , \1698 );
nor \U$1607 ( \1700 , \1659 , \1699 );
nand \U$1608 ( \1701 , \1643 , \1645 , \1649 , \1700 );
nor \U$1609 ( \1702 , \1639 , \1701 );
not \U$1610 ( \1703 , \1641 );
not \U$1611 ( \1704 , \115 );
or \U$1612 ( \1705 , \1703 , \1704 );
nand \U$1613 ( \1706 , \1705 , \1575 );
nand \U$1614 ( \1707 , \1702 , \1706 );
nor \U$1615 ( \1708 , \1637 , \1707 );
not \U$1616 ( \1709 , \1708 );
buf \U$1617 ( \1710 , \1707 );
nand \U$1618 ( \1711 , \1637 , \1710 );
nand \U$1619 ( \1712 , \1709 , \1711 );
buf \U$1620 ( \1713 , \1637 );
or \U$1621 ( \1714 , \1713 , \1560 );
not \U$1622 ( \1715 , \1559 );
nand \U$1623 ( \1716 , \1715 , \1637 );
nand \U$1624 ( \1717 , \1714 , \1716 );
and \U$1625 ( \1718 , \1712 , \1717 );
buf \U$1626 ( \1719 , \1718 );
not \U$1627 ( \1720 , \1719 );
or \U$1628 ( \1721 , \1567 , \1720 );
not \U$1629 ( \1722 , \1712 );
not \U$1630 ( \1723 , \1722 );
not \U$1631 ( \1724 , \1723 );
buf \U$1632 ( \1725 , \1715 );
not \U$1633 ( \1726 , \1725 );
buf \U$1634 ( \1727 , \1726 );
nand \U$1635 ( \1728 , \1724 , \1727 );
nand \U$1636 ( \1729 , \1721 , \1728 );
buf \U$1637 ( \1730 , \413 );
not \U$1638 ( \1731 , \1730 );
not \U$1639 ( \1732 , \911 );
nand \U$1640 ( \1733 , \1731 , \1732 );
and \U$1641 ( \1734 , \1733 , RI8929f28_52);
buf \U$1642 ( \1735 , \1547 );
nand \U$1643 ( \1736 , \1735 , RI89288a8_4);
and \U$1644 ( \1737 , \174 , RI89297a8_36);
and \U$1645 ( \1738 , \173 , RI8929f28_52);
nor \U$1646 ( \1739 , \1737 , \1738 );
not \U$1647 ( \1740 , \1739 );
not \U$1648 ( \1741 , \755 );
nand \U$1649 ( \1742 , \1740 , \1741 );
not \U$1650 ( \1743 , RI8929028_20);
nor \U$1651 ( \1744 , \174 , \1743 );
not \U$1652 ( \1745 , \1744 );
nand \U$1653 ( \1746 , \174 , \1743 );
nand \U$1654 ( \1747 , \1745 , \1746 );
not \U$1655 ( \1748 , RI89290a0_21);
not \U$1656 ( \1749 , RI8929fa0_53);
or \U$1657 ( \1750 , \1748 , \1749 );
nand \U$1658 ( \1751 , RI8929118_22, RI892a018_54);
not \U$1659 ( \1752 , \1751 );
nand \U$1660 ( \1753 , RI8929190_23, RI892a090_55);
not \U$1661 ( \1754 , \1753 );
nor \U$1662 ( \1755 , \1485 , \1480 );
not \U$1663 ( \1756 , \1755 );
not \U$1664 ( \1757 , \1593 );
or \U$1665 ( \1758 , \1756 , \1757 );
nand \U$1666 ( \1759 , \1758 , \1487 );
not \U$1667 ( \1760 , RI8929208_24);
nand \U$1668 ( \1761 , \1760 , \152 );
and \U$1669 ( \1762 , \1759 , \1761 );
and \U$1670 ( \1763 , RI8929208_24, RI892a108_56);
nor \U$1671 ( \1764 , \1762 , \1763 );
not \U$1672 ( \1765 , \1764 );
or \U$1673 ( \1766 , \1754 , \1765 );
not \U$1674 ( \1767 , RI8929190_23);
nand \U$1675 ( \1768 , \1767 , \160 );
nand \U$1676 ( \1769 , \1766 , \1768 );
not \U$1677 ( \1770 , \1769 );
or \U$1678 ( \1771 , \1752 , \1770 );
nand \U$1679 ( \1772 , \617 , \166 );
nand \U$1680 ( \1773 , \1771 , \1772 );
not \U$1681 ( \1774 , RI89290a0_21);
and \U$1682 ( \1775 , \1774 , \100 );
or \U$1683 ( \1776 , \1773 , \1775 );
nand \U$1684 ( \1777 , \1750 , \1776 );
xnor \U$1685 ( \1778 , \1747 , \1777 );
not \U$1686 ( \1779 , \405 );
nand \U$1687 ( \1780 , \1778 , \1779 );
not \U$1688 ( \1781 , RI89288a8_4);
nand \U$1689 ( \1782 , \173 , \1781 );
nand \U$1690 ( \1783 , RI89288a8_4, RI89297a8_36);
and \U$1691 ( \1784 , \1782 , \1783 );
not \U$1692 ( \1785 , \1784 );
nand \U$1693 ( \1786 , RI8928998_6, RI8929898_38);
nand \U$1694 ( \1787 , RI8928a10_7, RI8929910_39);
not \U$1695 ( \1788 , \1787 );
nor \U$1696 ( \1789 , \1528 , \1494 );
not \U$1697 ( \1790 , \1789 );
nor \U$1698 ( \1791 , RI8928a88_8, RI8929988_40);
nor \U$1699 ( \1792 , \1790 , \1497 , \1791 );
and \U$1700 ( \1793 , \1518 , \1792 );
nand \U$1701 ( \1794 , \1525 , \1521 );
and \U$1702 ( \1795 , \1789 , \1794 );
nor \U$1703 ( \1796 , \1795 , \1527 );
or \U$1704 ( \1797 , \1796 , \1791 );
nand \U$1705 ( \1798 , RI8928a88_8, RI8929988_40);
nand \U$1706 ( \1799 , \1797 , \1798 );
nor \U$1707 ( \1800 , \1793 , \1799 );
not \U$1708 ( \1801 , \1800 );
or \U$1709 ( \1802 , \1788 , \1801 );
nand \U$1710 ( \1803 , \159 , \604 );
nand \U$1711 ( \1804 , \1802 , \1803 );
and \U$1712 ( \1805 , \1786 , \1804 );
and \U$1713 ( \1806 , \165 , \834 );
nor \U$1714 ( \1807 , \1805 , \1806 );
not \U$1715 ( \1808 , RI8928920_5);
nand \U$1716 ( \1809 , \101 , \1808 );
and \U$1717 ( \1810 , \1807 , \1809 );
nor \U$1718 ( \1811 , \101 , \1808 );
nor \U$1719 ( \1812 , \1810 , \1811 );
not \U$1720 ( \1813 , \1812 );
or \U$1721 ( \1814 , \1785 , \1813 );
or \U$1722 ( \1815 , \1812 , \1784 );
nand \U$1723 ( \1816 , \1814 , \1815 );
buf \U$1724 ( \1817 , \410 );
buf \U$1725 ( \1818 , \1817 );
and \U$1726 ( \1819 , \1816 , \1818 );
and \U$1727 ( \1820 , \418 , RI89297a8_36);
nor \U$1728 ( \1821 , \1819 , \1820 );
nand \U$1729 ( \1822 , \1736 , \1742 , \1780 , \1821 );
nor \U$1730 ( \1823 , \1734 , \1822 );
xor \U$1731 ( \1824 , RI8929190_23, RI8929cd0_47);
not \U$1732 ( \1825 , \1824 );
not \U$1733 ( \1826 , \978 );
or \U$1734 ( \1827 , \1825 , \1826 );
xor \U$1735 ( \1828 , RI8929118_22, RI8929cd0_47);
nand \U$1736 ( \1829 , \1828 , RI8929d48_48);
nand \U$1737 ( \1830 , \1827 , \1829 );
not \U$1738 ( \1831 , \1830 );
xor \U$1739 ( \1832 , RI8929910_39, RI8929550_31);
not \U$1740 ( \1833 , \1832 );
not \U$1741 ( \1834 , RI8929988_40);
not \U$1742 ( \1835 , RI8929910_39);
or \U$1743 ( \1836 , \1834 , \1835 );
or \U$1744 ( \1837 , RI8929910_39, RI8929988_40);
nand \U$1745 ( \1838 , \1836 , \1837 );
xor \U$1746 ( \1839 , RI8929988_40, RI8929a00_41);
nor \U$1747 ( \1840 , \1838 , \1839 );
not \U$1748 ( \1841 , \1840 );
or \U$1749 ( \1842 , \1833 , \1841 );
buf \U$1750 ( \1843 , \1839 );
xor \U$1751 ( \1844 , RI89294d8_30, RI8929910_39);
nand \U$1752 ( \1845 , \1843 , \1844 );
nand \U$1753 ( \1846 , \1842 , \1845 );
not \U$1754 ( \1847 , \1846 );
or \U$1755 ( \1848 , \1831 , \1847 );
or \U$1756 ( \1849 , \1846 , \1830 );
xor \U$1757 ( \1850 , RI8929af0_43, RI8929370_27);
not \U$1758 ( \1851 , \1850 );
not \U$1759 ( \1852 , \1079 );
or \U$1760 ( \1853 , \1851 , \1852 );
xor \U$1761 ( \1854 , RI89292f8_26, RI8929af0_43);
nand \U$1762 ( \1855 , \1007 , \1854 );
nand \U$1763 ( \1856 , \1853 , \1855 );
nand \U$1764 ( \1857 , \1849 , \1856 );
nand \U$1765 ( \1858 , \1848 , \1857 );
and \U$1766 ( \1859 , RI8929cd0_47, RI89290a0_21);
not \U$1767 ( \1860 , RI8929cd0_47);
and \U$1768 ( \1861 , \1860 , \1774 );
nor \U$1769 ( \1862 , \1859 , \1861 );
and \U$1770 ( \1863 , RI8929d48_48, \1862 );
not \U$1771 ( \1864 , RI8929d48_48);
not \U$1772 ( \1865 , RI8929cd0_47);
nor \U$1773 ( \1866 , \1865 , RI8929118_22);
and \U$1774 ( \1867 , \1864 , \1866 );
or \U$1775 ( \1868 , \1863 , \1867 );
xor \U$1776 ( \1869 , RI89293e8_28, RI8929a00_41);
not \U$1777 ( \1870 , \1869 );
not \U$1778 ( \1871 , \1143 );
or \U$1779 ( \1872 , \1870 , \1871 );
xor \U$1780 ( \1873 , RI8929a78_42, RI8929af0_43);
xor \U$1781 ( \1874 , RI8929370_27, RI8929a00_41);
nand \U$1782 ( \1875 , \1873 , \1874 );
nand \U$1783 ( \1876 , \1872 , \1875 );
xor \U$1784 ( \1877 , \1868 , \1876 );
not \U$1785 ( \1878 , \1844 );
nor \U$1786 ( \1879 , \1839 , \1838 );
not \U$1787 ( \1880 , \1879 );
or \U$1788 ( \1881 , \1878 , \1880 );
xor \U$1789 ( \1882 , RI8929460_29, RI8929910_39);
nand \U$1790 ( \1883 , \1843 , \1882 );
nand \U$1791 ( \1884 , \1881 , \1883 );
xor \U$1792 ( \1885 , \1877 , \1884 );
xor \U$1793 ( \1886 , \1858 , \1885 );
xor \U$1794 ( \1887 , RI8929280_25, RI8929be0_45);
not \U$1795 ( \1888 , \1887 );
not \U$1796 ( \1889 , \967 );
or \U$1797 ( \1890 , \1888 , \1889 );
xor \U$1798 ( \1891 , RI8929be0_45, RI8929208_24);
nand \U$1799 ( \1892 , \970 , \1891 );
nand \U$1800 ( \1893 , \1890 , \1892 );
not \U$1801 ( \1894 , \1893 );
xor \U$1802 ( \1895 , RI8929898_38, RI8929910_39);
and \U$1803 ( \1896 , \1895 , RI89295c8_32);
xor \U$1804 ( \1897 , RI8929a00_41, RI8929460_29);
not \U$1805 ( \1898 , \1897 );
not \U$1806 ( \1899 , \1143 );
or \U$1807 ( \1900 , \1898 , \1899 );
nand \U$1808 ( \1901 , \1873 , \1869 );
nand \U$1809 ( \1902 , \1900 , \1901 );
not \U$1810 ( \1903 , \1902 );
xnor \U$1811 ( \1904 , \1896 , \1903 );
not \U$1812 ( \1905 , \1904 );
or \U$1813 ( \1906 , \1894 , \1905 );
not \U$1814 ( \1907 , \1903 );
nand \U$1815 ( \1908 , \1907 , \1896 );
nand \U$1816 ( \1909 , \1906 , \1908 );
xnor \U$1817 ( \1910 , \1886 , \1909 );
not \U$1818 ( \1911 , \1910 );
not \U$1819 ( \1912 , \1891 );
not \U$1820 ( \1913 , \967 );
or \U$1821 ( \1914 , \1912 , \1913 );
xor \U$1822 ( \1915 , RI8929be0_45, RI8929190_23);
nand \U$1823 ( \1916 , \970 , \1915 );
nand \U$1824 ( \1917 , \1914 , \1916 );
or \U$1825 ( \1918 , RI89295c8_32, RI8929898_38);
nand \U$1826 ( \1919 , \1918 , RI8929910_39);
nand \U$1827 ( \1920 , RI89295c8_32, RI8929898_38);
and \U$1828 ( \1921 , \1919 , \1920 , RI8929820_37);
nand \U$1829 ( \1922 , \1917 , \1921 );
not \U$1830 ( \1923 , \1922 );
nor \U$1831 ( \1924 , \1917 , \1921 );
nor \U$1832 ( \1925 , \1923 , \1924 );
not \U$1833 ( \1926 , \1079 );
not \U$1834 ( \1927 , \1926 );
and \U$1835 ( \1928 , \1927 , \1854 );
xor \U$1836 ( \1929 , RI8929af0_43, RI8929280_25);
and \U$1837 ( \1930 , \1007 , \1929 );
nor \U$1838 ( \1931 , \1928 , \1930 );
xor \U$1839 ( \1932 , RI89295c8_32, RI8929820_37);
not \U$1840 ( \1933 , \1932 );
not \U$1841 ( \1934 , \1895 );
xor \U$1842 ( \1935 , RI8929820_37, RI8929898_38);
nand \U$1843 ( \1936 , \1934 , \1935 );
not \U$1844 ( \1937 , \1936 );
not \U$1845 ( \1938 , \1937 );
or \U$1846 ( \1939 , \1933 , \1938 );
buf \U$1847 ( \1940 , \1895 );
xor \U$1848 ( \1941 , RI8929550_31, RI8929820_37);
nand \U$1849 ( \1942 , \1940 , \1941 );
nand \U$1850 ( \1943 , \1939 , \1942 );
not \U$1851 ( \1944 , \1943 );
and \U$1852 ( \1945 , \1931 , \1944 );
not \U$1853 ( \1946 , \1931 );
and \U$1854 ( \1947 , \1946 , \1943 );
nor \U$1855 ( \1948 , \1945 , \1947 );
xor \U$1856 ( \1949 , \1925 , \1948 );
xor \U$1857 ( \1950 , RI8929910_39, RI89295c8_32);
not \U$1858 ( \1951 , \1950 );
not \U$1859 ( \1952 , \1840 );
or \U$1860 ( \1953 , \1951 , \1952 );
nand \U$1861 ( \1954 , \1843 , \1832 );
nand \U$1862 ( \1955 , \1953 , \1954 );
xor \U$1863 ( \1956 , RI8929208_24, RI8929cd0_47);
not \U$1864 ( \1957 , \1956 );
not \U$1865 ( \1958 , \978 );
or \U$1866 ( \1959 , \1957 , \1958 );
nand \U$1867 ( \1960 , \1824 , RI8929d48_48);
nand \U$1868 ( \1961 , \1959 , \1960 );
and \U$1869 ( \1962 , \1955 , \1961 );
not \U$1870 ( \1963 , \1955 );
not \U$1871 ( \1964 , \1961 );
and \U$1872 ( \1965 , \1963 , \1964 );
xor \U$1873 ( \1966 , RI8929a00_41, RI89294d8_30);
not \U$1874 ( \1967 , \1966 );
nor \U$1875 ( \1968 , \1142 , \1069 );
not \U$1876 ( \1969 , \1968 );
or \U$1877 ( \1970 , \1967 , \1969 );
nand \U$1878 ( \1971 , \1873 , \1897 );
nand \U$1879 ( \1972 , \1970 , \1971 );
not \U$1880 ( \1973 , \1972 );
nor \U$1881 ( \1974 , \1965 , \1973 );
nor \U$1882 ( \1975 , \1962 , \1974 );
not \U$1883 ( \1976 , \1975 );
not \U$1884 ( \1977 , \1976 );
not \U$1885 ( \1978 , RI89295c8_32);
not \U$1886 ( \1979 , RI8929988_40);
or \U$1887 ( \1980 , \1978 , \1979 );
nand \U$1888 ( \1981 , \1980 , RI8929910_39);
not \U$1889 ( \1982 , \1981 );
or \U$1890 ( \1983 , RI89295c8_32, RI8929988_40);
nand \U$1891 ( \1984 , \1983 , RI8929a00_41);
nand \U$1892 ( \1985 , \1982 , \1984 );
not \U$1893 ( \1986 , \1985 );
xor \U$1894 ( \1987 , RI89292f8_26, RI8929be0_45);
not \U$1895 ( \1988 , \1987 );
not \U$1896 ( \1989 , \941 );
nor \U$1897 ( \1990 , \1989 , \970 );
not \U$1898 ( \1991 , \1990 );
or \U$1899 ( \1992 , \1988 , \1991 );
nand \U$1900 ( \1993 , \970 , \1887 );
nand \U$1901 ( \1994 , \1992 , \1993 );
nand \U$1902 ( \1995 , \1986 , \1994 );
xor \U$1903 ( \1996 , \1896 , \1903 );
xnor \U$1904 ( \1997 , \1996 , \1893 );
not \U$1905 ( \1998 , \1997 );
xor \U$1906 ( \1999 , \1995 , \1998 );
not \U$1907 ( \2000 , \1999 );
or \U$1908 ( \2001 , \1977 , \2000 );
not \U$1909 ( \2002 , \1995 );
nand \U$1910 ( \2003 , \2002 , \1997 );
nand \U$1911 ( \2004 , \2001 , \2003 );
nand \U$1912 ( \2005 , \1949 , \2004 );
not \U$1913 ( \2006 , \2005 );
or \U$1914 ( \2007 , \1911 , \2006 );
not \U$1915 ( \2008 , \1949 );
not \U$1916 ( \2009 , \2004 );
nand \U$1917 ( \2010 , \2008 , \2009 );
nand \U$1918 ( \2011 , \2007 , \2010 );
not \U$1919 ( \2012 , \2011 );
not \U$1920 ( \2013 , \1858 );
not \U$1921 ( \2014 , \2013 );
not \U$1922 ( \2015 , \1885 );
not \U$1923 ( \2016 , \2015 );
or \U$1924 ( \2017 , \2014 , \2016 );
nand \U$1925 ( \2018 , \2017 , \1909 );
not \U$1926 ( \2019 , \2013 );
nand \U$1927 ( \2020 , \2019 , \1885 );
nand \U$1928 ( \2021 , \2018 , \2020 );
not \U$1929 ( \2022 , \2021 );
and \U$1930 ( \2023 , \1927 , \1929 );
xor \U$1931 ( \2024 , RI8929af0_43, RI8929208_24);
and \U$1932 ( \2025 , \1007 , \2024 );
nor \U$1933 ( \2026 , \2023 , \2025 );
xor \U$1934 ( \2027 , \2026 , \1922 );
xor \U$1935 ( \2028 , \1868 , \1876 );
and \U$1936 ( \2029 , \2028 , \1884 );
and \U$1937 ( \2030 , \1868 , \1876 );
or \U$1938 ( \2031 , \2029 , \2030 );
xnor \U$1939 ( \2032 , \2027 , \2031 );
not \U$1940 ( \2033 , \2032 );
and \U$1941 ( \2034 , \2022 , \2033 );
and \U$1942 ( \2035 , \2021 , \2032 );
nor \U$1943 ( \2036 , \2034 , \2035 );
not \U$1944 ( \2037 , \2036 );
buf \U$1945 ( \2038 , \1931 );
nand \U$1946 ( \2039 , \2038 , \1944 );
not \U$1947 ( \2040 , \2039 );
not \U$1948 ( \2041 , \1925 );
or \U$1949 ( \2042 , \2040 , \2041 );
or \U$1950 ( \2043 , \2038 , \1944 );
nand \U$1951 ( \2044 , \2042 , \2043 );
not \U$1952 ( \2045 , \2044 );
not \U$1953 ( \2046 , \1915 );
not \U$1954 ( \2047 , \1156 );
or \U$1955 ( \2048 , \2046 , \2047 );
xor \U$1956 ( \2049 , RI8929be0_45, RI8929118_22);
nand \U$1957 ( \2050 , \1159 , \2049 );
nand \U$1958 ( \2051 , \2048 , \2050 );
xor \U$1959 ( \2052 , RI8929820_37, RI89297a8_36);
nand \U$1960 ( \2053 , \2052 , RI89295c8_32);
not \U$1961 ( \2054 , \2053 );
not \U$1962 ( \2055 , \1874 );
not \U$1963 ( \2056 , \1968 );
or \U$1964 ( \2057 , \2055 , \2056 );
xor \U$1965 ( \2058 , RI89292f8_26, RI8929a00_41);
nand \U$1966 ( \2059 , \1873 , \2058 );
nand \U$1967 ( \2060 , \2057 , \2059 );
not \U$1968 ( \2061 , \2060 );
or \U$1969 ( \2062 , \2054 , \2061 );
buf \U$1970 ( \2063 , \2053 );
or \U$1971 ( \2064 , \2060 , \2063 );
nand \U$1972 ( \2065 , \2062 , \2064 );
not \U$1973 ( \2066 , \2065 );
and \U$1974 ( \2067 , \2051 , \2066 );
not \U$1975 ( \2068 , \2051 );
and \U$1976 ( \2069 , \2068 , \2065 );
nor \U$1977 ( \2070 , \2067 , \2069 );
not \U$1978 ( \2071 , \2070 );
not \U$1979 ( \2072 , \2071 );
not \U$1980 ( \2073 , \1936 );
not \U$1981 ( \2074 , \1941 );
not \U$1982 ( \2075 , \2074 );
and \U$1983 ( \2076 , \2073 , \2075 );
xor \U$1984 ( \2077 , RI89294d8_30, RI8929820_37);
not \U$1985 ( \2078 , \2077 );
not \U$1986 ( \2079 , \1940 );
nor \U$1987 ( \2080 , \2078 , \2079 );
nor \U$1988 ( \2081 , \2076 , \2080 );
not \U$1989 ( \2082 , \2081 );
not \U$1990 ( \2083 , \1882 );
not \U$1991 ( \2084 , \1879 );
or \U$1992 ( \2085 , \2083 , \2084 );
xor \U$1993 ( \2086 , RI89293e8_28, RI8929910_39);
nand \U$1994 ( \2087 , \1843 , \2086 );
nand \U$1995 ( \2088 , \2085 , \2087 );
not \U$1996 ( \2089 , \2088 );
and \U$1997 ( \2090 , \931 , \1862 );
xor \U$1998 ( \2091 , RI8929028_20, RI8929cd0_47);
and \U$1999 ( \2092 , RI8929d48_48, \2091 );
nor \U$2000 ( \2093 , \2090 , \2092 );
not \U$2001 ( \2094 , \2093 );
or \U$2002 ( \2095 , \2089 , \2094 );
or \U$2003 ( \2096 , \2088 , \2093 );
nand \U$2004 ( \2097 , \2095 , \2096 );
not \U$2005 ( \2098 , \2097 );
or \U$2006 ( \2099 , \2082 , \2098 );
or \U$2007 ( \2100 , \2097 , \2081 );
nand \U$2008 ( \2101 , \2099 , \2100 );
not \U$2009 ( \2102 , \2101 );
not \U$2010 ( \2103 , \2102 );
or \U$2011 ( \2104 , \2072 , \2103 );
nand \U$2012 ( \2105 , \2101 , \2070 );
nand \U$2013 ( \2106 , \2104 , \2105 );
not \U$2014 ( \2107 , \2106 );
or \U$2015 ( \2108 , \2045 , \2107 );
or \U$2016 ( \2109 , \2106 , \2044 );
nand \U$2017 ( \2110 , \2108 , \2109 );
not \U$2018 ( \2111 , \2110 );
or \U$2019 ( \2112 , \2037 , \2111 );
or \U$2020 ( \2113 , \2110 , \2036 );
nand \U$2021 ( \2114 , \2112 , \2113 );
not \U$2022 ( \2115 , \2114 );
xor \U$2023 ( \2116 , \2012 , \2115 );
xor \U$2024 ( \2117 , \1949 , \1910 );
xnor \U$2025 ( \2118 , \2117 , \2009 );
xor \U$2026 ( \2119 , \1846 , \1830 );
xnor \U$2027 ( \2120 , \2119 , \1856 );
not \U$2028 ( \2121 , \2120 );
not \U$2029 ( \2122 , \1994 );
not \U$2030 ( \2123 , \1985 );
and \U$2031 ( \2124 , \2122 , \2123 );
and \U$2032 ( \2125 , \1985 , \1994 );
nor \U$2033 ( \2126 , \2124 , \2125 );
xor \U$2034 ( \2127 , RI89293e8_28, RI8929af0_43);
not \U$2035 ( \2128 , \2127 );
not \U$2036 ( \2129 , \1079 );
or \U$2037 ( \2130 , \2128 , \2129 );
nand \U$2038 ( \2131 , \1007 , \1850 );
nand \U$2039 ( \2132 , \2130 , \2131 );
not \U$2040 ( \2133 , \2132 );
and \U$2041 ( \2134 , \2126 , \2133 );
not \U$2042 ( \2135 , \2126 );
and \U$2043 ( \2136 , \2135 , \2132 );
nor \U$2044 ( \2137 , \2134 , \2136 );
and \U$2045 ( \2138 , \1839 , RI89295c8_32);
and \U$2046 ( \2139 , RI8929d48_48, \1956 );
not \U$2047 ( \2140 , RI8929d48_48);
not \U$2048 ( \2141 , RI8929cd0_47);
nor \U$2049 ( \2142 , \2141 , RI8929280_25);
and \U$2050 ( \2143 , \2140 , \2142 );
or \U$2051 ( \2144 , \2139 , \2143 );
xor \U$2052 ( \2145 , \2138 , \2144 );
not \U$2053 ( \2146 , \1146 );
not \U$2054 ( \2147 , \1968 );
or \U$2055 ( \2148 , \2146 , \2147 );
nand \U$2056 ( \2149 , \1873 , \1966 );
nand \U$2057 ( \2150 , \2148 , \2149 );
and \U$2058 ( \2151 , \2145 , \2150 );
and \U$2059 ( \2152 , \2138 , \2144 );
or \U$2060 ( \2153 , \2151 , \2152 );
nand \U$2061 ( \2154 , \2137 , \2153 );
not \U$2062 ( \2155 , \2133 );
not \U$2063 ( \2156 , \2126 );
nand \U$2064 ( \2157 , \2155 , \2156 );
nand \U$2065 ( \2158 , \2154 , \2157 );
nand \U$2066 ( \2159 , \2121 , \2158 );
not \U$2067 ( \2160 , \2159 );
xor \U$2068 ( \2161 , \1995 , \1975 );
xnor \U$2069 ( \2162 , \2161 , \1997 );
not \U$2070 ( \2163 , \2162 );
or \U$2071 ( \2164 , \2160 , \2163 );
nand \U$2072 ( \2165 , \2154 , \2157 , \2120 );
nand \U$2073 ( \2166 , \2164 , \2165 );
nor \U$2074 ( \2167 , \2118 , \2166 );
not \U$2075 ( \2168 , \2167 );
not \U$2076 ( \2169 , \2168 );
xor \U$2077 ( \2170 , \2158 , \2120 );
xor \U$2078 ( \2171 , \2170 , \2162 );
xor \U$2079 ( \2172 , \2132 , \2153 );
xnor \U$2080 ( \2173 , \2172 , \2156 );
buf \U$2081 ( \2174 , \2173 );
not \U$2082 ( \2175 , \1972 );
not \U$2083 ( \2176 , \1964 );
or \U$2084 ( \2177 , \2175 , \2176 );
nand \U$2085 ( \2178 , \1973 , \1961 );
nand \U$2086 ( \2179 , \2177 , \2178 );
and \U$2087 ( \2180 , \2179 , \1963 );
not \U$2088 ( \2181 , \2179 );
and \U$2089 ( \2182 , \2181 , \1955 );
nor \U$2090 ( \2183 , \2180 , \2182 );
not \U$2091 ( \2184 , \2183 );
not \U$2092 ( \2185 , \1132 );
not \U$2093 ( \2186 , \1079 );
or \U$2094 ( \2187 , \2185 , \2186 );
nand \U$2095 ( \2188 , \1007 , \2127 );
nand \U$2096 ( \2189 , \2187 , \2188 );
not \U$2097 ( \2190 , \2189 );
nand \U$2098 ( \2191 , \2190 , \1118 );
not \U$2099 ( \2192 , \2191 );
not \U$2100 ( \2193 , \1160 );
not \U$2101 ( \2194 , \1156 );
or \U$2102 ( \2195 , \2193 , \2194 );
nand \U$2103 ( \2196 , \1159 , \1987 );
nand \U$2104 ( \2197 , \2195 , \2196 );
not \U$2105 ( \2198 , \2197 );
or \U$2106 ( \2199 , \2192 , \2198 );
not \U$2107 ( \2200 , \1118 );
nand \U$2108 ( \2201 , \2200 , \2189 );
nand \U$2109 ( \2202 , \2199 , \2201 );
nand \U$2110 ( \2203 , \2184 , \2202 );
and \U$2111 ( \2204 , \2174 , \2203 );
nor \U$2112 ( \2205 , \2202 , \2184 );
nor \U$2113 ( \2206 , \2204 , \2205 );
nand \U$2114 ( \2207 , \2171 , \2206 );
nand \U$2115 ( \2208 , \1102 , \1171 );
xor \U$2116 ( \2209 , \2138 , \2144 );
xor \U$2117 ( \2210 , \2209 , \2150 );
not \U$2118 ( \2211 , \1162 );
not \U$2119 ( \2212 , \1153 );
or \U$2120 ( \2213 , \2211 , \2212 );
not \U$2121 ( \2214 , \1149 );
nand \U$2122 ( \2215 , \2214 , \1134 );
nand \U$2123 ( \2216 , \2213 , \2215 );
xor \U$2124 ( \2217 , \2210 , \2216 );
xor \U$2125 ( \2218 , \2189 , \2200 );
xor \U$2126 ( \2219 , \2218 , \2197 );
xnor \U$2127 ( \2220 , \2217 , \2219 );
not \U$2128 ( \2221 , \1119 );
and \U$2129 ( \2222 , \2221 , \1127 );
or \U$2130 ( \2223 , \2222 , \1163 );
or \U$2131 ( \2224 , \1127 , \2221 );
nand \U$2132 ( \2225 , \2223 , \2224 );
nand \U$2133 ( \2226 , \2220 , \2225 );
nand \U$2134 ( \2227 , \2208 , \2226 , \1174 );
nor \U$2135 ( \2228 , \2220 , \2225 );
not \U$2136 ( \2229 , \2173 );
and \U$2137 ( \2230 , \2202 , \2183 );
not \U$2138 ( \2231 , \2202 );
and \U$2139 ( \2232 , \2231 , \2184 );
nor \U$2140 ( \2233 , \2230 , \2232 );
not \U$2141 ( \2234 , \2233 );
or \U$2142 ( \2235 , \2229 , \2234 );
or \U$2143 ( \2236 , \2173 , \2233 );
nand \U$2144 ( \2237 , \2235 , \2236 );
not \U$2145 ( \2238 , \2219 );
not \U$2146 ( \2239 , \2238 );
not \U$2147 ( \2240 , \2210 );
not \U$2148 ( \2241 , \2216 );
xor \U$2149 ( \2242 , \2240 , \2241 );
not \U$2150 ( \2243 , \2242 );
or \U$2151 ( \2244 , \2239 , \2243 );
not \U$2152 ( \2245 , \2216 );
and \U$2153 ( \2246 , \2240 , \2245 );
not \U$2154 ( \2247 , \2246 );
nand \U$2155 ( \2248 , \2244 , \2247 );
nor \U$2156 ( \2249 , \2237 , \2248 );
nor \U$2157 ( \2250 , \2228 , \2249 );
nand \U$2158 ( \2251 , \2207 , \2227 , \2250 );
not \U$2159 ( \2252 , \2248 );
not \U$2160 ( \2253 , \2237 );
nor \U$2161 ( \2254 , \2252 , \2253 );
nand \U$2162 ( \2255 , \2207 , \2254 );
not \U$2163 ( \2256 , \2171 );
not \U$2164 ( \2257 , \2206 );
nand \U$2165 ( \2258 , \2256 , \2257 );
and \U$2166 ( \2259 , \2251 , \2255 , \2258 );
not \U$2167 ( \2260 , \2259 );
not \U$2168 ( \2261 , \2260 );
or \U$2169 ( \2262 , \2169 , \2261 );
nand \U$2170 ( \2263 , \2118 , \2166 );
nand \U$2171 ( \2264 , \2262 , \2263 );
xor \U$2172 ( \2265 , \2116 , \2264 );
not \U$2173 ( \2266 , \2265 );
not \U$2174 ( \2267 , \1587 );
not \U$2175 ( \2268 , \2267 );
and \U$2176 ( \2269 , \2266 , \2268 );
not \U$2177 ( \2270 , \1570 );
buf \U$2178 ( \2271 , \2270 );
and \U$2179 ( \2272 , \2271 , RI89288a8_4);
nor \U$2180 ( \2273 , \2269 , \2272 );
xnor \U$2181 ( \2274 , RI892a018_54, RI8929fa0_53);
xor \U$2182 ( \2275 , RI892a018_54, RI892a090_55);
nor \U$2183 ( \2276 , \2274 , \2275 );
xor \U$2184 ( \2277 , RI8929fa0_53, RI8928e48_16);
and \U$2185 ( \2278 , \2276 , \2277 );
xor \U$2186 ( \2279 , RI8929fa0_53, RI8928dd0_15);
and \U$2187 ( \2280 , \2275 , \2279 );
nor \U$2188 ( \2281 , \2278 , \2280 );
xor \U$2189 ( \2282 , RI8928b78_10, RI892a270_59);
not \U$2190 ( \2283 , \2282 );
xnor \U$2191 ( \2284 , RI892a270_59, RI892a2e8_60);
nor \U$2192 ( \2285 , \2284 , \1187 );
not \U$2193 ( \2286 , \2285 );
or \U$2194 ( \2287 , \2283 , \2286 );
xor \U$2195 ( \2288 , RI892a270_59, RI8928b00_9);
nand \U$2196 ( \2289 , \1232 , \2288 );
nand \U$2197 ( \2290 , \2287 , \2289 );
not \U$2198 ( \2291 , \2290 );
xor \U$2199 ( \2292 , \2281 , \2291 );
not \U$2200 ( \2293 , \2292 );
xor \U$2201 ( \2294 , RI8928a88_8, RI892a360_61);
not \U$2202 ( \2295 , \2294 );
not \U$2203 ( \2296 , \1221 );
or \U$2204 ( \2297 , \2295 , \2296 );
xor \U$2205 ( \2298 , RI892a360_61, RI8928a10_7);
nand \U$2206 ( \2299 , \1224 , \2298 );
nand \U$2207 ( \2300 , \2297 , \2299 );
or \U$2208 ( \2301 , RI8928e48_16, RI892a018_54);
nand \U$2209 ( \2302 , \2301 , RI892a090_55);
nand \U$2210 ( \2303 , RI8928e48_16, RI892a018_54);
and \U$2211 ( \2304 , \2302 , \2303 , RI8929fa0_53);
and \U$2212 ( \2305 , \2300 , \2304 );
not \U$2213 ( \2306 , \2305 );
not \U$2214 ( \2307 , \2304 );
nand \U$2215 ( \2308 , \1221 , \2294 );
nand \U$2216 ( \2309 , \2307 , \2308 , \2299 );
nand \U$2217 ( \2310 , \2306 , \2309 );
not \U$2218 ( \2311 , \2310 );
or \U$2219 ( \2312 , \2293 , \2311 );
or \U$2220 ( \2313 , \2310 , \2292 );
nand \U$2221 ( \2314 , \2312 , \2313 );
not \U$2222 ( \2315 , \2314 );
xor \U$2223 ( \2316 , RI892a450_63, RI8928a10_7);
not \U$2224 ( \2317 , \2316 );
not \U$2225 ( \2318 , \1291 );
or \U$2226 ( \2319 , \2317 , \2318 );
and \U$2227 ( \2320 , RI892a450_63, \834 );
not \U$2228 ( \2321 , RI892a450_63);
and \U$2229 ( \2322 , \2321 , RI8928998_6);
or \U$2230 ( \2323 , \2320 , \2322 );
nand \U$2231 ( \2324 , \2323 , RI892a4c8_64);
nand \U$2232 ( \2325 , \2319 , \2324 );
not \U$2233 ( \2326 , \2325 );
xor \U$2234 ( \2327 , RI8928dd0_15, RI892a090_55);
not \U$2235 ( \2328 , \2327 );
not \U$2236 ( \2329 , RI892a090_55);
not \U$2237 ( \2330 , RI892a108_56);
and \U$2238 ( \2331 , \2329 , \2330 );
and \U$2239 ( \2332 , RI892a090_55, RI892a108_56);
nor \U$2240 ( \2333 , \2331 , \2332 );
not \U$2241 ( \2334 , \2333 );
xor \U$2242 ( \2335 , RI892a108_56, RI892a180_57);
nor \U$2243 ( \2336 , \2334 , \2335 );
not \U$2244 ( \2337 , \2336 );
or \U$2245 ( \2338 , \2328 , \2337 );
not \U$2246 ( \2339 , RI892a180_57);
not \U$2247 ( \2340 , \152 );
or \U$2248 ( \2341 , \2339 , \2340 );
not \U$2249 ( \2342 , RI892a180_57);
nand \U$2250 ( \2343 , \2342 , RI892a108_56);
nand \U$2251 ( \2344 , \2341 , \2343 );
xor \U$2252 ( \2345 , RI8928d58_14, RI892a090_55);
nand \U$2253 ( \2346 , \2344 , \2345 );
nand \U$2254 ( \2347 , \2338 , \2346 );
not \U$2255 ( \2348 , \2347 );
or \U$2256 ( \2349 , \2326 , \2348 );
or \U$2257 ( \2350 , \2347 , \2325 );
xor \U$2258 ( \2351 , RI8928bf0_11, RI892a270_59);
not \U$2259 ( \2352 , \2351 );
not \U$2260 ( \2353 , \1188 );
or \U$2261 ( \2354 , \2352 , \2353 );
nand \U$2262 ( \2355 , \1187 , \2282 );
nand \U$2263 ( \2356 , \2354 , \2355 );
nand \U$2264 ( \2357 , \2350 , \2356 );
nand \U$2265 ( \2358 , \2349 , \2357 );
xor \U$2266 ( \2359 , RI892a180_57, RI8928ce0_13);
not \U$2267 ( \2360 , \2359 );
nor \U$2268 ( \2361 , \1201 , \1200 );
not \U$2269 ( \2362 , \2361 );
or \U$2270 ( \2363 , \2360 , \2362 );
xor \U$2271 ( \2364 , RI8928c68_12, RI892a180_57);
nand \U$2272 ( \2365 , \1201 , \2364 );
nand \U$2273 ( \2366 , \2363 , \2365 );
not \U$2274 ( \2367 , \2366 );
nand \U$2275 ( \2368 , \2275 , RI8928e48_16);
nor \U$2276 ( \2369 , \2367 , \2368 );
xor \U$2277 ( \2370 , RI892a360_61, RI8928b00_9);
not \U$2278 ( \2371 , \2370 );
not \U$2279 ( \2372 , \1221 );
or \U$2280 ( \2373 , \2371 , \2372 );
nand \U$2281 ( \2374 , \1224 , \2294 );
nand \U$2282 ( \2375 , \2373 , \2374 );
or \U$2283 ( \2376 , \2369 , \2375 );
not \U$2284 ( \2377 , \2366 );
nand \U$2285 ( \2378 , \2377 , \2368 );
nand \U$2286 ( \2379 , \2376 , \2378 );
xor \U$2287 ( \2380 , \2358 , \2379 );
not \U$2288 ( \2381 , \2364 );
not \U$2289 ( \2382 , \2361 );
or \U$2290 ( \2383 , \2381 , \2382 );
xor \U$2291 ( \2384 , RI8928bf0_11, RI892a180_57);
nand \U$2292 ( \2385 , \1207 , \2384 );
nand \U$2293 ( \2386 , \2383 , \2385 );
not \U$2294 ( \2387 , \2323 );
not \U$2295 ( \2388 , \1291 );
or \U$2296 ( \2389 , \2387 , \2388 );
xor \U$2297 ( \2390 , RI892a450_63, RI8928920_5);
nand \U$2298 ( \2391 , \2390 , RI892a4c8_64);
nand \U$2299 ( \2392 , \2389 , \2391 );
xor \U$2300 ( \2393 , \2386 , \2392 );
not \U$2301 ( \2394 , \2345 );
not \U$2302 ( \2395 , \2333 );
nor \U$2303 ( \2396 , \2395 , \2344 );
not \U$2304 ( \2397 , \2396 );
or \U$2305 ( \2398 , \2394 , \2397 );
xor \U$2306 ( \2399 , RI8928ce0_13, RI892a090_55);
nand \U$2307 ( \2400 , \2344 , \2399 );
nand \U$2308 ( \2401 , \2398 , \2400 );
xor \U$2309 ( \2402 , \2393 , \2401 );
xnor \U$2310 ( \2403 , \2380 , \2402 );
not \U$2311 ( \2404 , \2403 );
or \U$2312 ( \2405 , \2315 , \2404 );
not \U$2313 ( \2406 , \2403 );
not \U$2314 ( \2407 , \2314 );
nand \U$2315 ( \2408 , \2406 , \2407 );
nand \U$2316 ( \2409 , \2405 , \2408 );
xor \U$2317 ( \2410 , \2368 , \2366 );
xnor \U$2318 ( \2411 , \2410 , \2375 );
not \U$2319 ( \2412 , \2411 );
xor \U$2320 ( \2413 , RI892a450_63, RI8928a88_8);
not \U$2321 ( \2414 , \2413 );
not \U$2322 ( \2415 , \1291 );
or \U$2323 ( \2416 , \2414 , \2415 );
nand \U$2324 ( \2417 , \2316 , RI892a4c8_64);
nand \U$2325 ( \2418 , \2416 , \2417 );
xor \U$2326 ( \2419 , RI892a180_57, RI8928d58_14);
not \U$2327 ( \2420 , \2419 );
not \U$2328 ( \2421 , \2361 );
or \U$2329 ( \2422 , \2420 , \2421 );
nand \U$2330 ( \2423 , \1207 , \2359 );
nand \U$2331 ( \2424 , \2422 , \2423 );
or \U$2332 ( \2425 , \2418 , \2424 );
xor \U$2333 ( \2426 , RI892a090_55, RI8928e48_16);
not \U$2334 ( \2427 , \2426 );
not \U$2335 ( \2428 , \2396 );
or \U$2336 ( \2429 , \2427 , \2428 );
nand \U$2337 ( \2430 , \2344 , \2327 );
nand \U$2338 ( \2431 , \2429 , \2430 );
and \U$2339 ( \2432 , \2425 , \2431 );
and \U$2340 ( \2433 , \2424 , \2418 );
nor \U$2341 ( \2434 , \2432 , \2433 );
not \U$2342 ( \2435 , \2434 );
xor \U$2343 ( \2436 , RI892a360_61, RI8928b78_10);
not \U$2344 ( \2437 , \2436 );
not \U$2345 ( \2438 , \1221 );
or \U$2346 ( \2439 , \2437 , \2438 );
nand \U$2347 ( \2440 , \1257 , \2370 );
nand \U$2348 ( \2441 , \2439 , \2440 );
or \U$2349 ( \2442 , RI8928e48_16, RI892a108_56);
nand \U$2350 ( \2443 , \2442 , RI892a180_57);
nand \U$2351 ( \2444 , RI8928e48_16, RI892a108_56);
and \U$2352 ( \2445 , \2443 , \2444 , RI892a090_55);
and \U$2353 ( \2446 , \2441 , \2445 );
not \U$2354 ( \2447 , \2446 );
or \U$2355 ( \2448 , \2435 , \2447 );
or \U$2356 ( \2449 , \2434 , \2446 );
nand \U$2357 ( \2450 , \2448 , \2449 );
not \U$2358 ( \2451 , \2450 );
or \U$2359 ( \2452 , \2412 , \2451 );
not \U$2360 ( \2453 , \2434 );
nand \U$2361 ( \2454 , \2453 , \2446 );
nand \U$2362 ( \2455 , \2452 , \2454 );
not \U$2363 ( \2456 , \2455 );
xor \U$2364 ( \2457 , \2409 , \2456 );
xor \U$2365 ( \2458 , \2325 , \2347 );
xor \U$2366 ( \2459 , \2458 , \2356 );
not \U$2367 ( \2460 , \2411 );
not \U$2368 ( \2461 , \2450 );
not \U$2369 ( \2462 , \2461 );
or \U$2370 ( \2463 , \2460 , \2462 );
not \U$2371 ( \2464 , \2411 );
nand \U$2372 ( \2465 , \2464 , \2450 );
nand \U$2373 ( \2466 , \2463 , \2465 );
xor \U$2374 ( \2467 , \2459 , \2466 );
xor \U$2375 ( \2468 , RI8928c68_12, RI892a270_59);
not \U$2376 ( \2469 , \2468 );
not \U$2377 ( \2470 , \2285 );
or \U$2378 ( \2471 , \2469 , \2470 );
nand \U$2379 ( \2472 , \1232 , \2351 );
nand \U$2380 ( \2473 , \2471 , \2472 );
not \U$2381 ( \2474 , \2473 );
not \U$2382 ( \2475 , \1294 );
not \U$2383 ( \2476 , \1291 );
or \U$2384 ( \2477 , \2475 , \2476 );
nand \U$2385 ( \2478 , \2413 , RI892a4c8_64);
nand \U$2386 ( \2479 , \2477 , \2478 );
not \U$2387 ( \2480 , \2479 );
not \U$2388 ( \2481 , \1208 );
not \U$2389 ( \2482 , \1202 );
or \U$2390 ( \2483 , \2481 , \2482 );
nand \U$2391 ( \2484 , \2419 , \1201 );
nand \U$2392 ( \2485 , \2483 , \2484 );
nand \U$2393 ( \2486 , \2335 , RI8928e48_16);
or \U$2394 ( \2487 , \2485 , \2486 );
nand \U$2395 ( \2488 , \2485 , \2486 );
nand \U$2396 ( \2489 , \2487 , \2488 );
not \U$2397 ( \2490 , \2489 );
or \U$2398 ( \2491 , \2480 , \2490 );
not \U$2399 ( \2492 , \2486 );
nand \U$2400 ( \2493 , \2492 , \2485 );
nand \U$2401 ( \2494 , \2491 , \2493 );
not \U$2402 ( \2495 , \2494 );
not \U$2403 ( \2496 , \2495 );
or \U$2404 ( \2497 , \2474 , \2496 );
not \U$2405 ( \2498 , \2473 );
nand \U$2406 ( \2499 , \2498 , \2494 );
nand \U$2407 ( \2500 , \2497 , \2499 );
not \U$2408 ( \2501 , \2500 );
not \U$2409 ( \2502 , \2445 );
xor \U$2410 ( \2503 , \2441 , \2502 );
not \U$2411 ( \2504 , \2503 );
not \U$2412 ( \2505 , \2504 );
or \U$2413 ( \2506 , \2501 , \2505 );
nand \U$2414 ( \2507 , \2494 , \2473 );
nand \U$2415 ( \2508 , \2506 , \2507 );
and \U$2416 ( \2509 , \2467 , \2508 );
and \U$2417 ( \2510 , \2459 , \2466 );
or \U$2418 ( \2511 , \2509 , \2510 );
nand \U$2419 ( \2512 , \2457 , \2511 );
not \U$2420 ( \2513 , \2512 );
xor \U$2421 ( \2514 , \2459 , \2466 );
xor \U$2422 ( \2515 , \2514 , \2508 );
xor \U$2423 ( \2516 , \2424 , \2418 );
xor \U$2424 ( \2517 , \2516 , \2431 );
not \U$2425 ( \2518 , \2517 );
not \U$2426 ( \2519 , \1301 );
and \U$2427 ( \2520 , \1188 , \1191 );
and \U$2428 ( \2521 , \1187 , \2468 );
nor \U$2429 ( \2522 , \2520 , \2521 );
not \U$2430 ( \2523 , \2522 );
or \U$2431 ( \2524 , \2519 , \2523 );
not \U$2432 ( \2525 , \1225 );
not \U$2433 ( \2526 , \1221 );
or \U$2434 ( \2527 , \2525 , \2526 );
nand \U$2435 ( \2528 , \1257 , \2436 );
nand \U$2436 ( \2529 , \2527 , \2528 );
nand \U$2437 ( \2530 , \2524 , \2529 );
not \U$2438 ( \2531 , \1301 );
not \U$2439 ( \2532 , \2522 );
nand \U$2440 ( \2533 , \2531 , \2532 );
and \U$2441 ( \2534 , \2530 , \2533 );
nand \U$2442 ( \2535 , \2518 , \2534 );
not \U$2443 ( \2536 , \2535 );
not \U$2444 ( \2537 , \2503 );
not \U$2445 ( \2538 , \2500 );
or \U$2446 ( \2539 , \2537 , \2538 );
or \U$2447 ( \2540 , \2500 , \2503 );
nand \U$2448 ( \2541 , \2539 , \2540 );
not \U$2449 ( \2542 , \2541 );
or \U$2450 ( \2543 , \2536 , \2542 );
not \U$2451 ( \2544 , \2534 );
nand \U$2452 ( \2545 , \2544 , \2517 );
nand \U$2453 ( \2546 , \2543 , \2545 );
and \U$2454 ( \2547 , \2515 , \2546 );
xnor \U$2455 ( \2548 , \2517 , \2534 );
xor \U$2456 ( \2549 , \2541 , \2548 );
and \U$2457 ( \2550 , \1301 , \2532 );
not \U$2458 ( \2551 , \1301 );
and \U$2459 ( \2552 , \2551 , \2522 );
nor \U$2460 ( \2553 , \2550 , \2552 );
xnor \U$2461 ( \2554 , \2553 , \2529 );
not \U$2462 ( \2555 , \2554 );
and \U$2463 ( \2556 , \1215 , \1227 );
not \U$2464 ( \2557 , \1193 );
nor \U$2465 ( \2558 , \2557 , \1213 );
nor \U$2466 ( \2559 , \2556 , \2558 );
not \U$2467 ( \2560 , \2559 );
xor \U$2468 ( \2561 , \2489 , \2479 );
not \U$2469 ( \2562 , \2561 );
and \U$2470 ( \2563 , \2560 , \2562 );
and \U$2471 ( \2564 , \2559 , \2561 );
nor \U$2472 ( \2565 , \2563 , \2564 );
not \U$2473 ( \2566 , \2565 );
not \U$2474 ( \2567 , \2566 );
or \U$2475 ( \2568 , \2555 , \2567 );
not \U$2476 ( \2569 , \2559 );
nand \U$2477 ( \2570 , \2569 , \2561 );
nand \U$2478 ( \2571 , \2568 , \2570 );
nand \U$2479 ( \2572 , \2549 , \2571 );
not \U$2480 ( \2573 , \2572 );
nor \U$2481 ( \2574 , \2547 , \2573 );
not \U$2482 ( \2575 , \2574 );
not \U$2483 ( \2576 , \2554 );
not \U$2484 ( \2577 , \2576 );
not \U$2485 ( \2578 , \2566 );
or \U$2486 ( \2579 , \2577 , \2578 );
nand \U$2487 ( \2580 , \2565 , \2554 );
nand \U$2488 ( \2581 , \2579 , \2580 );
not \U$2489 ( \2582 , \2581 );
not \U$2490 ( \2583 , \1308 );
not \U$2491 ( \2584 , \1229 );
or \U$2492 ( \2585 , \2583 , \2584 );
not \U$2493 ( \2586 , \1286 );
nand \U$2494 ( \2587 , \2586 , \1304 );
nand \U$2495 ( \2588 , \2585 , \2587 );
not \U$2496 ( \2589 , \2588 );
nand \U$2497 ( \2590 , \2582 , \2589 );
not \U$2498 ( \2591 , \2590 );
not \U$2499 ( \2592 , \1308 );
not \U$2500 ( \2593 , \1228 );
and \U$2501 ( \2594 , \2592 , \2593 );
not \U$2502 ( \2595 , \1229 );
and \U$2503 ( \2596 , \2595 , \1308 );
nor \U$2504 ( \2597 , \2594 , \2596 );
not \U$2505 ( \2598 , \2597 );
not \U$2506 ( \2599 , \1280 );
or \U$2507 ( \2600 , \2598 , \2599 );
nand \U$2508 ( \2601 , \2600 , \1450 );
or \U$2509 ( \2602 , \1280 , \2597 );
nand \U$2510 ( \2603 , \2601 , \2602 );
not \U$2511 ( \2604 , \2603 );
or \U$2512 ( \2605 , \2591 , \2604 );
nand \U$2513 ( \2606 , \2581 , \2588 );
nand \U$2514 ( \2607 , \2605 , \2606 );
nor \U$2515 ( \2608 , \2549 , \2571 );
not \U$2516 ( \2609 , \2608 );
nand \U$2517 ( \2610 , \2607 , \2609 );
not \U$2518 ( \2611 , \2610 );
or \U$2519 ( \2612 , \2575 , \2611 );
nor \U$2520 ( \2613 , \2515 , \2546 );
not \U$2521 ( \2614 , \2613 );
nand \U$2522 ( \2615 , \2612 , \2614 );
not \U$2523 ( \2616 , \2615 );
or \U$2524 ( \2617 , \2513 , \2616 );
nor \U$2525 ( \2618 , \2457 , \2511 );
not \U$2526 ( \2619 , \2618 );
nand \U$2527 ( \2620 , \2617 , \2619 );
and \U$2528 ( \2621 , \2281 , \2291 );
or \U$2529 ( \2622 , \2310 , \2621 );
not \U$2530 ( \2623 , \2281 );
nand \U$2531 ( \2624 , \2623 , \2290 );
nand \U$2532 ( \2625 , \2622 , \2624 );
not \U$2533 ( \2626 , \2625 );
not \U$2534 ( \2627 , \2298 );
not \U$2535 ( \2628 , \1221 );
or \U$2536 ( \2629 , \2627 , \2628 );
xor \U$2537 ( \2630 , RI892a360_61, RI8928998_6);
nand \U$2538 ( \2631 , \1224 , \2630 );
nand \U$2539 ( \2632 , \2629 , \2631 );
not \U$2540 ( \2633 , \2384 );
not \U$2541 ( \2634 , \1203 );
or \U$2542 ( \2635 , \2633 , \2634 );
xor \U$2543 ( \2636 , RI8928b78_10, RI892a180_57);
nand \U$2544 ( \2637 , \1207 , \2636 );
nand \U$2545 ( \2638 , \2635 , \2637 );
not \U$2546 ( \2639 , RI8929f28_52);
not \U$2547 ( \2640 , \100 );
or \U$2548 ( \2641 , \2639 , \2640 );
not \U$2549 ( \2642 , RI8929f28_52);
nand \U$2550 ( \2643 , \2642 , RI8929fa0_53);
nand \U$2551 ( \2644 , \2641 , \2643 );
nand \U$2552 ( \2645 , \2644 , RI8928e48_16);
xnor \U$2553 ( \2646 , \2638 , \2645 );
xor \U$2554 ( \2647 , \2632 , \2646 );
not \U$2555 ( \2648 , \2647 );
not \U$2556 ( \2649 , \2648 );
and \U$2557 ( \2650 , \1291 , \2390 );
xor \U$2558 ( \2651 , RI892a450_63, RI89288a8_4);
and \U$2559 ( \2652 , \2651 , RI892a4c8_64);
nor \U$2560 ( \2653 , \2650 , \2652 );
not \U$2561 ( \2654 , \2653 );
not \U$2562 ( \2655 , \2399 );
not \U$2563 ( \2656 , \2336 );
or \U$2564 ( \2657 , \2655 , \2656 );
xor \U$2565 ( \2658 , RI8928c68_12, RI892a090_55);
nand \U$2566 ( \2659 , \2344 , \2658 );
nand \U$2567 ( \2660 , \2657 , \2659 );
not \U$2568 ( \2661 , \2660 );
or \U$2569 ( \2662 , \2654 , \2661 );
or \U$2570 ( \2663 , \2660 , \2653 );
nand \U$2571 ( \2664 , \2662 , \2663 );
not \U$2572 ( \2665 , \2664 );
and \U$2573 ( \2666 , \2276 , \2279 );
xor \U$2574 ( \2667 , RI8928d58_14, RI8929fa0_53);
and \U$2575 ( \2668 , \2667 , \2275 );
nor \U$2576 ( \2669 , \2666 , \2668 );
not \U$2577 ( \2670 , \2669 );
and \U$2578 ( \2671 , \2665 , \2670 );
and \U$2579 ( \2672 , \2664 , \2669 );
nor \U$2580 ( \2673 , \2671 , \2672 );
not \U$2581 ( \2674 , \2673 );
not \U$2582 ( \2675 , \2674 );
or \U$2583 ( \2676 , \2649 , \2675 );
not \U$2584 ( \2677 , \2647 );
or \U$2585 ( \2678 , \2674 , \2677 );
nand \U$2586 ( \2679 , \2676 , \2678 );
not \U$2587 ( \2680 , \2679 );
or \U$2588 ( \2681 , \2626 , \2680 );
or \U$2589 ( \2682 , \2625 , \2679 );
nand \U$2590 ( \2683 , \2681 , \2682 );
not \U$2591 ( \2684 , \2683 );
not \U$2592 ( \2685 , \2402 );
not \U$2593 ( \2686 , \2685 );
not \U$2594 ( \2687 , \2358 );
not \U$2595 ( \2688 , \2687 );
or \U$2596 ( \2689 , \2686 , \2688 );
not \U$2597 ( \2690 , \2358 );
not \U$2598 ( \2691 , \2402 );
or \U$2599 ( \2692 , \2690 , \2691 );
nand \U$2600 ( \2693 , \2692 , \2379 );
nand \U$2601 ( \2694 , \2689 , \2693 );
not \U$2602 ( \2695 , \2694 );
not \U$2603 ( \2696 , \2288 );
not \U$2604 ( \2697 , \2285 );
or \U$2605 ( \2698 , \2696 , \2697 );
xor \U$2606 ( \2699 , RI892a270_59, RI8928a88_8);
nand \U$2607 ( \2700 , \1232 , \2699 );
nand \U$2608 ( \2701 , \2698 , \2700 );
xor \U$2609 ( \2702 , \2701 , \2305 );
xor \U$2610 ( \2703 , \2386 , \2392 );
and \U$2611 ( \2704 , \2703 , \2401 );
and \U$2612 ( \2705 , \2386 , \2392 );
or \U$2613 ( \2706 , \2704 , \2705 );
xor \U$2614 ( \2707 , \2702 , \2706 );
not \U$2615 ( \2708 , \2707 );
and \U$2616 ( \2709 , \2695 , \2708 );
and \U$2617 ( \2710 , \2694 , \2707 );
nor \U$2618 ( \2711 , \2709 , \2710 );
not \U$2619 ( \2712 , \2711 );
or \U$2620 ( \2713 , \2684 , \2712 );
or \U$2621 ( \2714 , \2711 , \2683 );
nand \U$2622 ( \2715 , \2713 , \2714 );
not \U$2623 ( \2716 , \2314 );
not \U$2624 ( \2717 , \2403 );
or \U$2625 ( \2718 , \2716 , \2717 );
nand \U$2626 ( \2719 , \2718 , \2456 );
nand \U$2627 ( \2720 , \2408 , \2719 );
and \U$2628 ( \2721 , \2715 , \2720 );
not \U$2629 ( \2722 , \2721 );
or \U$2630 ( \2723 , \2720 , \2715 );
nand \U$2631 ( \2724 , \2722 , \2723 );
and \U$2632 ( \2725 , \2620 , \2724 );
not \U$2633 ( \2726 , \2620 );
not \U$2634 ( \2727 , \2724 );
and \U$2635 ( \2728 , \2726 , \2727 );
nor \U$2636 ( \2729 , \2725 , \2728 );
not \U$2637 ( \2730 , \1453 );
not \U$2638 ( \2731 , \2730 );
not \U$2639 ( \2732 , \2731 );
nand \U$2640 ( \2733 , \2729 , \2732 );
and \U$2641 ( \2734 , \776 , \424 );
not \U$2642 ( \2735 , \2734 );
not \U$2643 ( \2736 , \2735 );
not \U$2644 ( \2737 , \2736 );
not \U$2645 ( \2738 , \173 );
buf \U$2646 ( \2739 , \1644 );
nand \U$2647 ( \2740 , \2738 , \2739 );
not \U$2648 ( \2741 , \2740 );
or \U$2649 ( \2742 , \2737 , \2741 );
nand \U$2650 ( \2743 , \2742 , RI8929028_20);
nand \U$2651 ( \2744 , \1823 , \2273 , \2733 , \2743 );
not \U$2652 ( \2745 , \2744 );
not \U$2653 ( \2746 , \2745 );
buf \U$2654 ( \2747 , \1575 );
and \U$2655 ( \2748 , \2747 , RI8929fa0_53);
nand \U$2656 ( \2749 , \1735 , RI8928920_5);
or \U$2657 ( \2750 , \101 , RI8929fa0_53);
or \U$2658 ( \2751 , \100 , RI8929820_37);
nand \U$2659 ( \2752 , \2750 , \2751 );
nand \U$2660 ( \2753 , \1741 , \2752 );
xor \U$2661 ( \2754 , \1774 , \100 );
not \U$2662 ( \2755 , \2754 );
not \U$2663 ( \2756 , \1773 );
or \U$2664 ( \2757 , \2755 , \2756 );
or \U$2665 ( \2758 , \1773 , \2754 );
nand \U$2666 ( \2759 , \2757 , \2758 );
and \U$2667 ( \2760 , \2759 , \1779 );
not \U$2668 ( \2761 , \1807 );
and \U$2669 ( \2762 , \101 , RI8928920_5);
and \U$2670 ( \2763 , \1808 , RI8929820_37);
nor \U$2671 ( \2764 , \2762 , \2763 );
not \U$2672 ( \2765 , \2764 );
and \U$2673 ( \2766 , \2761 , \2765 );
and \U$2674 ( \2767 , \1807 , \2764 );
nor \U$2675 ( \2768 , \2766 , \2767 );
not \U$2676 ( \2769 , \1818 );
or \U$2677 ( \2770 , \2768 , \2769 );
and \U$2678 ( \2771 , \1730 , RI8929fa0_53);
and \U$2679 ( \2772 , \418 , RI8929820_37);
nor \U$2680 ( \2773 , \2771 , \2772 );
nand \U$2681 ( \2774 , \2770 , \2773 );
nor \U$2682 ( \2775 , \2760 , \2774 );
nand \U$2683 ( \2776 , \2749 , \2753 , \2775 );
nor \U$2684 ( \2777 , \2748 , \2776 );
not \U$2685 ( \2778 , \2270 );
not \U$2686 ( \2779 , \2778 );
nand \U$2687 ( \2780 , \2779 , RI8928920_5);
nand \U$2688 ( \2781 , \2739 , RI8929820_37);
not \U$2689 ( \2782 , \2781 );
not \U$2690 ( \2783 , \2736 );
or \U$2691 ( \2784 , \2782 , \2783 );
nand \U$2692 ( \2785 , \2784 , RI89290a0_21);
nand \U$2693 ( \2786 , \2619 , \2512 );
xor \U$2694 ( \2787 , \2786 , \2615 );
and \U$2695 ( \2788 , \2787 , \2732 );
not \U$2696 ( \2789 , \2260 );
nand \U$2697 ( \2790 , \2263 , \2168 );
xor \U$2698 ( \2791 , \2789 , \2790 );
nor \U$2699 ( \2792 , \2791 , \2267 );
nor \U$2700 ( \2793 , \2788 , \2792 );
nand \U$2701 ( \2794 , \2777 , \2780 , \2785 , \2793 );
not \U$2702 ( \2795 , \2794 );
and \U$2703 ( \2796 , \2746 , \2795 );
and \U$2704 ( \2797 , \2745 , \2794 );
nor \U$2705 ( \2798 , \2796 , \2797 );
not \U$2706 ( \2799 , \2798 );
not \U$2707 ( \2800 , \2799 );
not \U$2708 ( \2801 , \2800 );
not \U$2709 ( \2802 , \2801 );
xnor \U$2710 ( \2803 , \168 , \2752 );
not \U$2711 ( \2804 , \2803 );
nand \U$2712 ( \2805 , \911 , RI8929eb0_51);
nand \U$2713 ( \2806 , \2735 , RI8928fb0_19);
nand \U$2714 ( \2807 , \1554 , RI8928fb0_19);
and \U$2715 ( \2808 , \419 , \2807 );
nor \U$2716 ( \2809 , \2808 , \181 );
xor \U$2717 ( \2810 , RI8929730_35, RI8929eb0_51);
not \U$2718 ( \2811 , \2810 );
not \U$2719 ( \2812 , \1549 );
or \U$2720 ( \2813 , \2811 , \2812 );
nand \U$2721 ( \2814 , \1730 , RI8929eb0_51);
nand \U$2722 ( \2815 , \2813 , \2814 );
not \U$2723 ( \2816 , \1783 );
not \U$2724 ( \2817 , \1812 );
or \U$2725 ( \2818 , \2816 , \2817 );
nand \U$2726 ( \2819 , \2818 , \1782 );
not \U$2727 ( \2820 , \2819 );
and \U$2728 ( \2821 , RI8929730_35, RI8928830_3);
not \U$2729 ( \2822 , RI8929730_35);
not \U$2730 ( \2823 , RI8928830_3);
and \U$2731 ( \2824 , \2822 , \2823 );
nor \U$2732 ( \2825 , \2821 , \2824 );
not \U$2733 ( \2826 , \2825 );
and \U$2734 ( \2827 , \2820 , \2826 );
and \U$2735 ( \2828 , \2819 , \2825 );
nor \U$2736 ( \2829 , \2827 , \2828 );
nor \U$2737 ( \2830 , \2769 , \2829 );
nor \U$2738 ( \2831 , \2809 , \2815 , \2830 );
or \U$2739 ( \2832 , \1777 , \1744 );
nand \U$2740 ( \2833 , \2832 , \1746 );
not \U$2741 ( \2834 , RI8928fb0_19);
and \U$2742 ( \2835 , RI8929eb0_51, \2834 );
not \U$2743 ( \2836 , RI8929eb0_51);
and \U$2744 ( \2837 , \2836 , RI8928fb0_19);
nor \U$2745 ( \2838 , \2835 , \2837 );
xor \U$2746 ( \2839 , \2833 , \2838 );
nand \U$2747 ( \2840 , \2839 , \1779 );
and \U$2748 ( \2841 , \2805 , \2806 , \2831 , \2840 );
or \U$2749 ( \2842 , RI89295c8_32, RI89297a8_36);
nand \U$2750 ( \2843 , \2842 , RI8929820_37);
nand \U$2751 ( \2844 , RI89295c8_32, RI89297a8_36);
nand \U$2752 ( \2845 , \2843 , \2844 , RI8929730_35);
not \U$2753 ( \2846 , \2845 );
not \U$2754 ( \2847 , \2091 );
not \U$2755 ( \2848 , \931 );
or \U$2756 ( \2849 , \2847 , \2848 );
and \U$2757 ( \2850 , RI8929cd0_47, \2834 );
not \U$2758 ( \2851 , RI8929cd0_47);
and \U$2759 ( \2852 , \2851 , RI8928fb0_19);
or \U$2760 ( \2853 , \2850 , \2852 );
nand \U$2761 ( \2854 , \2853 , RI8929d48_48);
nand \U$2762 ( \2855 , \2849 , \2854 );
not \U$2763 ( \2856 , \2855 );
or \U$2764 ( \2857 , \2846 , \2856 );
or \U$2765 ( \2858 , \2855 , \2845 );
nand \U$2766 ( \2859 , \2857 , \2858 );
not \U$2767 ( \2860 , \2051 );
not \U$2768 ( \2861 , \2065 );
or \U$2769 ( \2862 , \2860 , \2861 );
not \U$2770 ( \2863 , \2063 );
nand \U$2771 ( \2864 , \2863 , \2060 );
nand \U$2772 ( \2865 , \2862 , \2864 );
xor \U$2773 ( \2866 , \2859 , \2865 );
not \U$2774 ( \2867 , \2081 );
not \U$2775 ( \2868 , \2867 );
not \U$2776 ( \2869 , \2097 );
or \U$2777 ( \2870 , \2868 , \2869 );
not \U$2778 ( \2871 , \2093 );
nand \U$2779 ( \2872 , \2871 , \2088 );
nand \U$2780 ( \2873 , \2870 , \2872 );
xor \U$2781 ( \2874 , \2866 , \2873 );
xor \U$2782 ( \2875 , RI89295c8_32, RI8929730_35);
not \U$2783 ( \2876 , \2875 );
not \U$2784 ( \2877 , RI8929730_35);
xor \U$2785 ( \2878 , RI89297a8_36, \2877 );
nor \U$2786 ( \2879 , \2878 , \2052 );
not \U$2787 ( \2880 , \2879 );
or \U$2788 ( \2881 , \2876 , \2880 );
xor \U$2789 ( \2882 , RI8929550_31, RI8929730_35);
nand \U$2790 ( \2883 , \2052 , \2882 );
nand \U$2791 ( \2884 , \2881 , \2883 );
not \U$2792 ( \2885 , \2077 );
not \U$2793 ( \2886 , \1937 );
or \U$2794 ( \2887 , \2885 , \2886 );
xor \U$2795 ( \2888 , RI8929460_29, RI8929820_37);
nand \U$2796 ( \2889 , \1940 , \2888 );
nand \U$2797 ( \2890 , \2887 , \2889 );
xor \U$2798 ( \2891 , \2884 , \2890 );
not \U$2799 ( \2892 , \2024 );
not \U$2800 ( \2893 , \1927 );
or \U$2801 ( \2894 , \2892 , \2893 );
xor \U$2802 ( \2895 , RI8929af0_43, RI8929190_23);
nand \U$2803 ( \2896 , \1007 , \2895 );
nand \U$2804 ( \2897 , \2894 , \2896 );
xor \U$2805 ( \2898 , \2891 , \2897 );
not \U$2806 ( \2899 , \2058 );
buf \U$2807 ( \2900 , \1968 );
not \U$2808 ( \2901 , \2900 );
or \U$2809 ( \2902 , \2899 , \2901 );
buf \U$2810 ( \2903 , \1873 );
xor \U$2811 ( \2904 , RI8929a00_41, RI8929280_25);
nand \U$2812 ( \2905 , \2903 , \2904 );
nand \U$2813 ( \2906 , \2902 , \2905 );
not \U$2814 ( \2907 , \2086 );
not \U$2815 ( \2908 , \1840 );
or \U$2816 ( \2909 , \2907 , \2908 );
xor \U$2817 ( \2910 , RI8929910_39, RI8929370_27);
nand \U$2818 ( \2911 , \1843 , \2910 );
nand \U$2819 ( \2912 , \2909 , \2911 );
xor \U$2820 ( \2913 , \2906 , \2912 );
not \U$2821 ( \2914 , \2049 );
not \U$2822 ( \2915 , \1156 );
or \U$2823 ( \2916 , \2914 , \2915 );
and \U$2824 ( \2917 , RI8929be0_45, RI89290a0_21);
not \U$2825 ( \2918 , RI8929be0_45);
and \U$2826 ( \2919 , \2918 , \1774 );
nor \U$2827 ( \2920 , \2917 , \2919 );
nand \U$2828 ( \2921 , \1159 , \2920 );
nand \U$2829 ( \2922 , \2916 , \2921 );
xor \U$2830 ( \2923 , \2913 , \2922 );
xor \U$2831 ( \2924 , \2898 , \2923 );
buf \U$2832 ( \2925 , \2026 );
not \U$2833 ( \2926 , \2925 );
not \U$2834 ( \2927 , \1922 );
or \U$2835 ( \2928 , \2926 , \2927 );
nand \U$2836 ( \2929 , \2928 , \2031 );
or \U$2837 ( \2930 , \1922 , \2925 );
nand \U$2838 ( \2931 , \2929 , \2930 );
xor \U$2839 ( \2932 , \2924 , \2931 );
xor \U$2840 ( \2933 , \2874 , \2932 );
nand \U$2841 ( \2934 , \2102 , \2070 );
not \U$2842 ( \2935 , \2934 );
not \U$2843 ( \2936 , \2044 );
or \U$2844 ( \2937 , \2935 , \2936 );
not \U$2845 ( \2938 , \2102 );
nand \U$2846 ( \2939 , \2938 , \2071 );
nand \U$2847 ( \2940 , \2937 , \2939 );
xor \U$2848 ( \2941 , \2933 , \2940 );
not \U$2849 ( \2942 , \2032 );
not \U$2850 ( \2943 , \2942 );
not \U$2851 ( \2944 , \2110 );
not \U$2852 ( \2945 , \2944 );
or \U$2853 ( \2946 , \2943 , \2945 );
not \U$2854 ( \2947 , \2032 );
not \U$2855 ( \2948 , \2110 );
or \U$2856 ( \2949 , \2947 , \2948 );
nand \U$2857 ( \2950 , \2949 , \2021 );
nand \U$2858 ( \2951 , \2946 , \2950 );
nor \U$2859 ( \2952 , \2941 , \2951 );
not \U$2860 ( \2953 , \2952 );
nand \U$2861 ( \2954 , \2941 , \2951 );
nand \U$2862 ( \2955 , \2953 , \2954 );
not \U$2863 ( \2956 , \2955 );
not \U$2864 ( \2957 , \2167 );
nand \U$2865 ( \2958 , \2114 , \2011 );
not \U$2866 ( \2959 , \2958 );
or \U$2867 ( \2960 , \2957 , \2959 );
nand \U$2868 ( \2961 , \2012 , \2115 );
nand \U$2869 ( \2962 , \2960 , \2961 );
not \U$2870 ( \2963 , \2962 );
nand \U$2871 ( \2964 , \2259 , \2958 , \2263 );
nand \U$2872 ( \2965 , \2963 , \2964 );
not \U$2873 ( \2966 , \2965 );
or \U$2874 ( \2967 , \2956 , \2966 );
or \U$2875 ( \2968 , \2965 , \2955 );
nand \U$2876 ( \2969 , \2967 , \2968 );
not \U$2877 ( \2970 , \2267 );
and \U$2878 ( \2971 , \2969 , \2970 );
not \U$2879 ( \2972 , \2651 );
not \U$2880 ( \2973 , \1291 );
or \U$2881 ( \2974 , \2972 , \2973 );
xor \U$2882 ( \2975 , RI8928830_3, RI892a450_63);
nand \U$2883 ( \2976 , \2975 , RI892a4c8_64);
nand \U$2884 ( \2977 , \2974 , \2976 );
not \U$2885 ( \2978 , \2977 );
or \U$2886 ( \2979 , RI8928e48_16, RI8929f28_52);
nand \U$2887 ( \2980 , \2979 , RI8929fa0_53);
nand \U$2888 ( \2981 , RI8928e48_16, RI8929f28_52);
nand \U$2889 ( \2982 , \2980 , \2981 , RI8929eb0_51);
not \U$2890 ( \2983 , \2982 );
and \U$2891 ( \2984 , \2978 , \2983 );
and \U$2892 ( \2985 , \2977 , \2982 );
nor \U$2893 ( \2986 , \2984 , \2985 );
not \U$2894 ( \2987 , \2632 );
not \U$2895 ( \2988 , \2646 );
or \U$2896 ( \2989 , \2987 , \2988 );
not \U$2897 ( \2990 , \2645 );
nand \U$2898 ( \2991 , \2990 , \2638 );
nand \U$2899 ( \2992 , \2989 , \2991 );
xor \U$2900 ( \2993 , \2986 , \2992 );
not \U$2901 ( \2994 , \2669 );
not \U$2902 ( \2995 , \2994 );
not \U$2903 ( \2996 , \2664 );
or \U$2904 ( \2997 , \2995 , \2996 );
not \U$2905 ( \2998 , \2653 );
nand \U$2906 ( \2999 , \2998 , \2660 );
nand \U$2907 ( \3000 , \2997 , \2999 );
xnor \U$2908 ( \3001 , \2993 , \3000 );
not \U$2909 ( \3002 , \2677 );
not \U$2910 ( \3003 , \3002 );
not \U$2911 ( \3004 , \2674 );
or \U$2912 ( \3005 , \3003 , \3004 );
not \U$2913 ( \3006 , \2677 );
not \U$2914 ( \3007 , \2673 );
or \U$2915 ( \3008 , \3006 , \3007 );
nand \U$2916 ( \3009 , \3008 , \2625 );
nand \U$2917 ( \3010 , \3005 , \3009 );
xor \U$2918 ( \3011 , \3001 , \3010 );
not \U$2919 ( \3012 , \2667 );
nor \U$2920 ( \3013 , \2275 , \2274 );
not \U$2921 ( \3014 , \3013 );
or \U$2922 ( \3015 , \3012 , \3014 );
xor \U$2923 ( \3016 , RI8929fa0_53, RI8928ce0_13);
nand \U$2924 ( \3017 , \2275 , \3016 );
nand \U$2925 ( \3018 , \3015 , \3017 );
xnor \U$2926 ( \3019 , RI8929f28_52, RI8929eb0_51);
nor \U$2927 ( \3020 , \2644 , \3019 );
xor \U$2928 ( \3021 , RI8929eb0_51, RI8928e48_16);
and \U$2929 ( \3022 , \3020 , \3021 );
xor \U$2930 ( \3023 , RI8929eb0_51, RI8928dd0_15);
and \U$2931 ( \3024 , \3023 , \2644 );
nor \U$2932 ( \3025 , \3022 , \3024 );
and \U$2933 ( \3026 , \3018 , \3025 );
not \U$2934 ( \3027 , \3018 );
not \U$2935 ( \3028 , \3025 );
and \U$2936 ( \3029 , \3027 , \3028 );
or \U$2937 ( \3030 , \3026 , \3029 );
not \U$2938 ( \3031 , \2699 );
not \U$2939 ( \3032 , \2285 );
or \U$2940 ( \3033 , \3031 , \3032 );
xnor \U$2941 ( \3034 , RI892a270_59, RI8928a10_7);
not \U$2942 ( \3035 , \3034 );
nand \U$2943 ( \3036 , \3035 , \1232 );
nand \U$2944 ( \3037 , \3033 , \3036 );
and \U$2945 ( \3038 , \3030 , \3037 );
not \U$2946 ( \3039 , \3030 );
not \U$2947 ( \3040 , \3037 );
and \U$2948 ( \3041 , \3039 , \3040 );
nor \U$2949 ( \3042 , \3038 , \3041 );
not \U$2950 ( \3043 , \2636 );
buf \U$2951 ( \3044 , \2361 );
not \U$2952 ( \3045 , \3044 );
or \U$2953 ( \3046 , \3043 , \3045 );
buf \U$2954 ( \3047 , \1201 );
xor \U$2955 ( \3048 , RI892a180_57, RI8928b00_9);
nand \U$2956 ( \3049 , \3047 , \3048 );
nand \U$2957 ( \3050 , \3046 , \3049 );
not \U$2958 ( \3051 , \2658 );
buf \U$2959 ( \3052 , \2396 );
not \U$2960 ( \3053 , \3052 );
or \U$2961 ( \3054 , \3051 , \3053 );
not \U$2962 ( \3055 , \2344 );
not \U$2963 ( \3056 , \3055 );
xor \U$2964 ( \3057 , RI892a090_55, RI8928bf0_11);
nand \U$2965 ( \3058 , \3056 , \3057 );
nand \U$2966 ( \3059 , \3054 , \3058 );
xor \U$2967 ( \3060 , \3050 , \3059 );
not \U$2968 ( \3061 , \2630 );
buf \U$2969 ( \3062 , \1221 );
not \U$2970 ( \3063 , \3062 );
or \U$2971 ( \3064 , \3061 , \3063 );
xnor \U$2972 ( \3065 , RI892a360_61, RI8928920_5);
not \U$2973 ( \3066 , \3065 );
nand \U$2974 ( \3067 , \3066 , \1257 );
nand \U$2975 ( \3068 , \3064 , \3067 );
xor \U$2976 ( \3069 , \3060 , \3068 );
xor \U$2977 ( \3070 , \3042 , \3069 );
xor \U$2978 ( \3071 , \2701 , \2305 );
and \U$2979 ( \3072 , \3071 , \2706 );
and \U$2980 ( \3073 , \2701 , \2305 );
or \U$2981 ( \3074 , \3072 , \3073 );
xor \U$2982 ( \3075 , \3070 , \3074 );
xor \U$2983 ( \3076 , \3011 , \3075 );
not \U$2984 ( \3077 , \3076 );
not \U$2985 ( \3078 , \2711 );
not \U$2986 ( \3079 , \3078 );
not \U$2987 ( \3080 , \2683 );
or \U$2988 ( \3081 , \3079 , \3080 );
not \U$2989 ( \3082 , \2707 );
nand \U$2990 ( \3083 , \3082 , \2694 );
nand \U$2991 ( \3084 , \3081 , \3083 );
nand \U$2992 ( \3085 , \3077 , \3084 );
not \U$2993 ( \3086 , \3084 );
nand \U$2994 ( \3087 , \3086 , \3076 );
and \U$2995 ( \3088 , \3085 , \3087 );
not \U$2996 ( \3089 , \3088 );
nand \U$2997 ( \3090 , \2610 , \2574 );
nor \U$2998 ( \3091 , \2721 , \2613 , \2618 );
and \U$2999 ( \3092 , \3090 , \3091 );
or \U$3000 ( \3093 , \2721 , \2512 );
nand \U$3001 ( \3094 , \3093 , \2723 );
nor \U$3002 ( \3095 , \3092 , \3094 );
not \U$3003 ( \3096 , \3095 );
or \U$3004 ( \3097 , \3089 , \3096 );
or \U$3005 ( \3098 , \3095 , \3088 );
nand \U$3006 ( \3099 , \3097 , \3098 );
and \U$3007 ( \3100 , \3099 , \2732 );
nor \U$3008 ( \3101 , \2971 , \3100 );
not \U$3009 ( \3102 , \777 );
not \U$3010 ( \3103 , \1732 );
or \U$3011 ( \3104 , \3102 , \3103 );
nand \U$3012 ( \3105 , \3104 , RI8928830_3);
nand \U$3013 ( \3106 , \2841 , \3101 , \3105 );
buf \U$3014 ( \3107 , \3106 );
not \U$3015 ( \3108 , \3107 );
not \U$3016 ( \3109 , \3108 );
buf \U$3017 ( \3110 , \3109 );
not \U$3018 ( \3111 , \3110 );
or \U$3019 ( \3112 , \2804 , \3111 );
not \U$3020 ( \3113 , \3106 );
buf \U$3021 ( \3114 , \3113 );
not \U$3022 ( \3115 , \3114 );
or \U$3023 ( \3116 , \3115 , \2803 );
nand \U$3024 ( \3117 , \3112 , \3116 );
not \U$3025 ( \3118 , \3117 );
or \U$3026 ( \3119 , \2802 , \3118 );
not \U$3027 ( \3120 , \3110 );
xor \U$3028 ( \3121 , \165 , \166 );
and \U$3029 ( \3122 , \162 , \3121 );
not \U$3030 ( \3123 , \162 );
not \U$3031 ( \3124 , \3121 );
and \U$3032 ( \3125 , \3123 , \3124 );
or \U$3033 ( \3126 , \3122 , \3125 );
not \U$3034 ( \3127 , \3126 );
not \U$3035 ( \3128 , \3127 );
and \U$3036 ( \3129 , \3120 , \3128 );
and \U$3037 ( \3130 , \3115 , \3127 );
nor \U$3038 ( \3131 , \3129 , \3130 );
not \U$3039 ( \3132 , \3131 );
not \U$3040 ( \3133 , \3113 );
not \U$3041 ( \3134 , \2745 );
or \U$3042 ( \3135 , \3133 , \3134 );
or \U$3043 ( \3136 , \3108 , \2745 );
nand \U$3044 ( \3137 , \3135 , \3136 );
not \U$3045 ( \3138 , \3137 );
nand \U$3046 ( \3139 , \3138 , \2798 );
not \U$3047 ( \3140 , \3139 );
not \U$3048 ( \3141 , \3140 );
not \U$3049 ( \3142 , \3141 );
nand \U$3050 ( \3143 , \3132 , \3142 );
nand \U$3051 ( \3144 , \3119 , \3143 );
xor \U$3052 ( \3145 , \1729 , \3144 );
xor \U$3053 ( \3146 , RI892a108_56, RI8929988_40);
and \U$3054 ( \3147 , \150 , \3146 );
not \U$3055 ( \3148 , \150 );
not \U$3056 ( \3149 , \3146 );
and \U$3057 ( \3150 , \3148 , \3149 );
or \U$3058 ( \3151 , \3147 , \3150 );
not \U$3059 ( \3152 , \3151 );
xor \U$3060 ( \3153 , \2874 , \2932 );
and \U$3061 ( \3154 , \3153 , \2940 );
and \U$3062 ( \3155 , \2874 , \2932 );
or \U$3063 ( \3156 , \3154 , \3155 );
not \U$3064 ( \3157 , \3156 );
xor \U$3065 ( \3158 , \2898 , \2923 );
and \U$3066 ( \3159 , \3158 , \2931 );
and \U$3067 ( \3160 , \2898 , \2923 );
or \U$3068 ( \3161 , \3159 , \3160 );
not \U$3069 ( \3162 , \3161 );
xor \U$3070 ( \3163 , \2906 , \2912 );
and \U$3071 ( \3164 , \3163 , \2922 );
and \U$3072 ( \3165 , \2906 , \2912 );
or \U$3073 ( \3166 , \3164 , \3165 );
not \U$3074 ( \3167 , \3166 );
not \U$3075 ( \3168 , \2920 );
not \U$3076 ( \3169 , \1156 );
or \U$3077 ( \3170 , \3168 , \3169 );
and \U$3078 ( \3171 , RI8929be0_45, RI8929028_20);
not \U$3079 ( \3172 , RI8929be0_45);
and \U$3080 ( \3173 , \3172 , \1743 );
nor \U$3081 ( \3174 , \3171 , \3173 );
nand \U$3082 ( \3175 , \1159 , \3174 );
nand \U$3083 ( \3176 , \3170 , \3175 );
not \U$3084 ( \3177 , \2853 );
not \U$3085 ( \3178 , \931 );
or \U$3086 ( \3179 , \3177 , \3178 );
xor \U$3087 ( \3180 , RI8928f38_18, RI8929cd0_47);
nand \U$3088 ( \3181 , \3180 , RI8929d48_48);
nand \U$3089 ( \3182 , \3179 , \3181 );
and \U$3090 ( \3183 , RI8929730_35, RI89296b8_34);
not \U$3091 ( \3184 , RI8929730_35);
not \U$3092 ( \3185 , RI89296b8_34);
and \U$3093 ( \3186 , \3184 , \3185 );
nor \U$3094 ( \3187 , \3183 , \3186 );
and \U$3095 ( \3188 , \3187 , RI89295c8_32);
xor \U$3096 ( \3189 , \3182 , \3188 );
xnor \U$3097 ( \3190 , \3176 , \3189 );
not \U$3098 ( \3191 , \3190 );
or \U$3099 ( \3192 , \3167 , \3191 );
or \U$3100 ( \3193 , \3190 , \3166 );
nand \U$3101 ( \3194 , \3192 , \3193 );
not \U$3102 ( \3195 , \3194 );
xor \U$3103 ( \3196 , \2884 , \2890 );
and \U$3104 ( \3197 , \3196 , \2897 );
and \U$3105 ( \3198 , \2884 , \2890 );
or \U$3106 ( \3199 , \3197 , \3198 );
not \U$3107 ( \3200 , \3199 );
not \U$3108 ( \3201 , \3200 );
and \U$3109 ( \3202 , \3195 , \3201 );
and \U$3110 ( \3203 , \3194 , \3200 );
nor \U$3111 ( \3204 , \3202 , \3203 );
not \U$3112 ( \3205 , \3204 );
or \U$3113 ( \3206 , \3162 , \3205 );
or \U$3114 ( \3207 , \3204 , \3161 );
nand \U$3115 ( \3208 , \3206 , \3207 );
not \U$3116 ( \3209 , \3208 );
not \U$3117 ( \3210 , \2845 );
nand \U$3118 ( \3211 , \3210 , \2855 );
not \U$3119 ( \3212 , \3211 );
and \U$3120 ( \3213 , \2879 , \2882 );
xor \U$3121 ( \3214 , RI8929730_35, RI89294d8_30);
and \U$3122 ( \3215 , \3214 , \2052 );
nor \U$3123 ( \3216 , \3213 , \3215 );
not \U$3124 ( \3217 , \3216 );
not \U$3125 ( \3218 , \2888 );
not \U$3126 ( \3219 , \1937 );
or \U$3127 ( \3220 , \3218 , \3219 );
xor \U$3128 ( \3221 , RI8929820_37, RI89293e8_28);
nand \U$3129 ( \3222 , \1940 , \3221 );
nand \U$3130 ( \3223 , \3220 , \3222 );
not \U$3131 ( \3224 , \3223 );
or \U$3132 ( \3225 , \3217 , \3224 );
or \U$3133 ( \3226 , \3223 , \3216 );
nand \U$3134 ( \3227 , \3225 , \3226 );
not \U$3135 ( \3228 , \3227 );
or \U$3136 ( \3229 , \3212 , \3228 );
or \U$3137 ( \3230 , \3227 , \3211 );
nand \U$3138 ( \3231 , \3229 , \3230 );
not \U$3139 ( \3232 , \3231 );
not \U$3140 ( \3233 , \2910 );
not \U$3141 ( \3234 , \1840 );
or \U$3142 ( \3235 , \3233 , \3234 );
xor \U$3143 ( \3236 , RI8929910_39, RI89292f8_26);
nand \U$3144 ( \3237 , \1843 , \3236 );
nand \U$3145 ( \3238 , \3235 , \3237 );
not \U$3146 ( \3239 , \3238 );
not \U$3147 ( \3240 , \2903 );
not \U$3148 ( \3241 , \3240 );
xnor \U$3149 ( \3242 , RI8929a00_41, RI8929208_24);
not \U$3150 ( \3243 , \3242 );
and \U$3151 ( \3244 , \3241 , \3243 );
and \U$3152 ( \3245 , \2900 , \2904 );
nor \U$3153 ( \3246 , \3244 , \3245 );
not \U$3154 ( \3247 , \3246 );
or \U$3155 ( \3248 , \3239 , \3247 );
or \U$3156 ( \3249 , \3238 , \3246 );
nand \U$3157 ( \3250 , \3248 , \3249 );
not \U$3158 ( \3251 , \3250 );
not \U$3159 ( \3252 , \2895 );
not \U$3160 ( \3253 , \1927 );
or \U$3161 ( \3254 , \3252 , \3253 );
xor \U$3162 ( \3255 , RI8929af0_43, RI8929118_22);
nand \U$3163 ( \3256 , \1007 , \3255 );
nand \U$3164 ( \3257 , \3254 , \3256 );
not \U$3165 ( \3258 , \3257 );
not \U$3166 ( \3259 , \3258 );
and \U$3167 ( \3260 , \3251 , \3259 );
and \U$3168 ( \3261 , \3250 , \3258 );
nor \U$3169 ( \3262 , \3260 , \3261 );
not \U$3170 ( \3263 , \3262 );
or \U$3171 ( \3264 , \3232 , \3263 );
or \U$3172 ( \3265 , \3262 , \3231 );
nand \U$3173 ( \3266 , \3264 , \3265 );
xor \U$3174 ( \3267 , \2859 , \2865 );
and \U$3175 ( \3268 , \3267 , \2873 );
and \U$3176 ( \3269 , \2859 , \2865 );
or \U$3177 ( \3270 , \3268 , \3269 );
xnor \U$3178 ( \3271 , \3266 , \3270 );
not \U$3179 ( \3272 , \3271 );
and \U$3180 ( \3273 , \3209 , \3272 );
and \U$3181 ( \3274 , \3208 , \3271 );
nor \U$3182 ( \3275 , \3273 , \3274 );
nand \U$3183 ( \3276 , \3157 , \3275 );
not \U$3184 ( \3277 , \3276 );
not \U$3185 ( \3278 , \2952 );
not \U$3186 ( \3279 , \3278 );
nand \U$3187 ( \3280 , \2963 , \2964 );
not \U$3188 ( \3281 , \3280 );
or \U$3189 ( \3282 , \3279 , \3281 );
nand \U$3190 ( \3283 , \3282 , \2954 );
not \U$3191 ( \3284 , \3283 );
or \U$3192 ( \3285 , \3277 , \3284 );
not \U$3193 ( \3286 , \3275 );
nand \U$3194 ( \3287 , \3286 , \3156 );
nand \U$3195 ( \3288 , \3285 , \3287 );
not \U$3196 ( \3289 , \3288 );
not \U$3197 ( \3290 , \3270 );
not \U$3198 ( \3291 , \3266 );
or \U$3199 ( \3292 , \3290 , \3291 );
not \U$3200 ( \3293 , \3262 );
nand \U$3201 ( \3294 , \3293 , \3231 );
nand \U$3202 ( \3295 , \3292 , \3294 );
not \U$3203 ( \3296 , \3295 );
not \U$3204 ( \3297 , \3199 );
not \U$3205 ( \3298 , \3194 );
or \U$3206 ( \3299 , \3297 , \3298 );
not \U$3207 ( \3300 , \3190 );
nand \U$3208 ( \3301 , \3300 , \3166 );
nand \U$3209 ( \3302 , \3299 , \3301 );
not \U$3210 ( \3303 , \3302 );
and \U$3211 ( \3304 , \3296 , \3303 );
and \U$3212 ( \3305 , \3295 , \3302 );
nor \U$3213 ( \3306 , \3304 , \3305 );
not \U$3214 ( \3307 , \3187 );
and \U$3215 ( \3308 , RI8929550_31, RI8929640_33);
nor \U$3216 ( \3309 , RI8929550_31, RI8929640_33);
nor \U$3217 ( \3310 , \3308 , \3309 );
or \U$3218 ( \3311 , \3307 , \3310 );
and \U$3219 ( \3312 , RI89296b8_34, RI89295c8_32);
not \U$3220 ( \3313 , RI89296b8_34);
and \U$3221 ( \3314 , \3313 , RI8929640_33);
nor \U$3222 ( \3315 , \3312 , \3314 );
and \U$3223 ( \3316 , RI89295c8_32, RI8929640_33);
or \U$3224 ( \3317 , \3315 , \3316 );
nand \U$3225 ( \3318 , \3317 , \3307 );
nand \U$3226 ( \3319 , \3311 , \3318 );
not \U$3227 ( \3320 , \3236 );
not \U$3228 ( \3321 , \1840 );
or \U$3229 ( \3322 , \3320 , \3321 );
xor \U$3230 ( \3323 , RI8929280_25, RI8929910_39);
nand \U$3231 ( \3324 , \1843 , \3323 );
nand \U$3232 ( \3325 , \3322 , \3324 );
xor \U$3233 ( \3326 , \3319 , \3325 );
not \U$3234 ( \3327 , \3255 );
not \U$3235 ( \3328 , \1927 );
or \U$3236 ( \3329 , \3327 , \3328 );
and \U$3237 ( \3330 , \114 , RI89290a0_21);
and \U$3238 ( \3331 , \1774 , RI8929af0_43);
nor \U$3239 ( \3332 , \3330 , \3331 );
not \U$3240 ( \3333 , \3332 );
nand \U$3241 ( \3334 , \3333 , \1007 );
nand \U$3242 ( \3335 , \3329 , \3334 );
xnor \U$3243 ( \3336 , \3326 , \3335 );
and \U$3244 ( \3337 , \2879 , \3214 );
xor \U$3245 ( \3338 , RI8929730_35, RI8929460_29);
and \U$3246 ( \3339 , \2052 , \3338 );
nor \U$3247 ( \3340 , \3337 , \3339 );
not \U$3248 ( \3341 , \3242 );
not \U$3249 ( \3342 , \3341 );
not \U$3250 ( \3343 , \2900 );
or \U$3251 ( \3344 , \3342 , \3343 );
xor \U$3252 ( \3345 , RI8929190_23, RI8929a00_41);
nand \U$3253 ( \3346 , \2903 , \3345 );
nand \U$3254 ( \3347 , \3344 , \3346 );
xor \U$3255 ( \3348 , \3340 , \3347 );
not \U$3256 ( \3349 , \3180 );
not \U$3257 ( \3350 , \931 );
or \U$3258 ( \3351 , \3349 , \3350 );
and \U$3259 ( \3352 , RI8929cd0_47, RI8928ec0_17);
not \U$3260 ( \3353 , RI8929cd0_47);
not \U$3261 ( \3354 , RI8928ec0_17);
and \U$3262 ( \3355 , \3353 , \3354 );
nor \U$3263 ( \3356 , \3352 , \3355 );
nand \U$3264 ( \3357 , \3356 , RI8929d48_48);
nand \U$3265 ( \3358 , \3351 , \3357 );
not \U$3266 ( \3359 , \3358 );
or \U$3267 ( \3360 , RI89295c8_32, RI89296b8_34);
nand \U$3268 ( \3361 , \3360 , RI8929730_35);
nand \U$3269 ( \3362 , RI89295c8_32, RI89296b8_34);
and \U$3270 ( \3363 , \3361 , \3362 , RI8929640_33);
not \U$3271 ( \3364 , \3363 );
and \U$3272 ( \3365 , \3359 , \3364 );
and \U$3273 ( \3366 , \3358 , \3363 );
nor \U$3274 ( \3367 , \3365 , \3366 );
xor \U$3275 ( \3368 , \3348 , \3367 );
xor \U$3276 ( \3369 , \3336 , \3368 );
and \U$3277 ( \3370 , \3250 , \3257 );
not \U$3278 ( \3371 , \3246 );
and \U$3279 ( \3372 , \3238 , \3371 );
nor \U$3280 ( \3373 , \3370 , \3372 );
xnor \U$3281 ( \3374 , \3369 , \3373 );
not \U$3282 ( \3375 , \3189 );
not \U$3283 ( \3376 , \3176 );
or \U$3284 ( \3377 , \3375 , \3376 );
nand \U$3285 ( \3378 , \3182 , \3188 );
nand \U$3286 ( \3379 , \3377 , \3378 );
not \U$3287 ( \3380 , \3174 );
not \U$3288 ( \3381 , \1156 );
or \U$3289 ( \3382 , \3380 , \3381 );
and \U$3290 ( \3383 , RI8929be0_45, \2834 );
not \U$3291 ( \3384 , RI8929be0_45);
and \U$3292 ( \3385 , \3384 , RI8928fb0_19);
nor \U$3293 ( \3386 , \3383 , \3385 );
not \U$3294 ( \3387 , \3386 );
nand \U$3295 ( \3388 , \3387 , \1159 );
nand \U$3296 ( \3389 , \3382 , \3388 );
not \U$3297 ( \3390 , \3221 );
or \U$3298 ( \3391 , \1936 , \3390 );
and \U$3299 ( \3392 , RI8929370_27, \101 );
not \U$3300 ( \3393 , RI8929370_27);
and \U$3301 ( \3394 , \3393 , RI8929820_37);
nor \U$3302 ( \3395 , \3392 , \3394 );
or \U$3303 ( \3396 , \2079 , \3395 );
nand \U$3304 ( \3397 , \3391 , \3396 );
xnor \U$3305 ( \3398 , \3389 , \3397 );
xor \U$3306 ( \3399 , \3379 , \3398 );
not \U$3307 ( \3400 , \3211 );
nand \U$3308 ( \3401 , \3400 , \3227 );
not \U$3309 ( \3402 , \3216 );
nand \U$3310 ( \3403 , \3402 , \3223 );
and \U$3311 ( \3404 , \3401 , \3403 );
xor \U$3312 ( \3405 , \3399 , \3404 );
and \U$3313 ( \3406 , \3374 , \3405 );
not \U$3314 ( \3407 , \3374 );
not \U$3315 ( \3408 , \3405 );
and \U$3316 ( \3409 , \3407 , \3408 );
nor \U$3317 ( \3410 , \3406 , \3409 );
xnor \U$3318 ( \3411 , \3306 , \3410 );
not \U$3319 ( \3412 , \3411 );
not \U$3320 ( \3413 , \3271 );
not \U$3321 ( \3414 , \3413 );
not \U$3322 ( \3415 , \3208 );
or \U$3323 ( \3416 , \3414 , \3415 );
not \U$3324 ( \3417 , \3204 );
nand \U$3325 ( \3418 , \3417 , \3161 );
nand \U$3326 ( \3419 , \3416 , \3418 );
not \U$3327 ( \3420 , \3419 );
or \U$3328 ( \3421 , \3412 , \3420 );
or \U$3329 ( \3422 , \3419 , \3411 );
nand \U$3330 ( \3423 , \3421 , \3422 );
not \U$3331 ( \3424 , \3423 );
and \U$3332 ( \3425 , \3289 , \3424 );
and \U$3333 ( \3426 , \3288 , \3423 );
nor \U$3334 ( \3427 , \3425 , \3426 );
buf \U$3335 ( \3428 , \2267 );
nor \U$3336 ( \3429 , \3427 , \3428 );
not \U$3337 ( \3430 , \1779 );
nand \U$3338 ( \3431 , RI8928fb0_19, RI8929eb0_51);
not \U$3339 ( \3432 , \3431 );
not \U$3340 ( \3433 , \2833 );
or \U$3341 ( \3434 , \3432 , \3433 );
nand \U$3342 ( \3435 , \182 , \2834 );
nand \U$3343 ( \3436 , \3434 , \3435 );
nand \U$3344 ( \3437 , RI8928f38_18, RI8929e38_50);
and \U$3345 ( \3438 , \3436 , \3437 );
not \U$3346 ( \3439 , RI8928f38_18);
not \U$3347 ( \3440 , RI8929e38_50);
and \U$3348 ( \3441 , \3439 , \3440 );
nor \U$3349 ( \3442 , \3438 , \3441 );
and \U$3350 ( \3443 , \95 , RI8928ec0_17);
and \U$3351 ( \3444 , \3354 , RI8929dc0_49);
nor \U$3352 ( \3445 , \3443 , \3444 );
xor \U$3353 ( \3446 , \3442 , \3445 );
nor \U$3354 ( \3447 , \3430 , \3446 );
nand \U$3355 ( \3448 , \1554 , RI8929640_33);
not \U$3356 ( \3449 , \3448 );
not \U$3357 ( \3450 , \2734 );
or \U$3358 ( \3451 , \3449 , \3450 );
nand \U$3359 ( \3452 , \3451 , RI8928ec0_17);
and \U$3360 ( \3453 , \95 , RI8929640_33);
and \U$3361 ( \3454 , \94 , RI8929dc0_49);
nor \U$3362 ( \3455 , \3453 , \3454 );
not \U$3363 ( \3456 , \3455 );
not \U$3364 ( \3457 , \3456 );
not \U$3365 ( \3458 , \1741 );
or \U$3366 ( \3459 , \3457 , \3458 );
nand \U$3367 ( \3460 , \418 , RI8929640_33);
nand \U$3368 ( \3461 , \3459 , \3460 );
not \U$3369 ( \3462 , RI8928740_1);
nor \U$3370 ( \3463 , \776 , \3462 );
nor \U$3371 ( \3464 , \3461 , \3463 );
nand \U$3372 ( \3465 , \3452 , \3464 );
nor \U$3373 ( \3466 , \3447 , \3465 );
not \U$3374 ( \3467 , \1730 );
nand \U$3375 ( \3468 , \3467 , \1732 );
nand \U$3376 ( \3469 , \3468 , RI8929dc0_49);
nand \U$3377 ( \3470 , \2271 , RI8928740_1);
or \U$3378 ( \3471 , \3462 , RI8929640_33);
or \U$3379 ( \3472 , \94 , RI8928740_1);
nand \U$3380 ( \3473 , \3471 , \3472 );
nand \U$3381 ( \3474 , RI89287b8_2, RI89296b8_34);
not \U$3382 ( \3475 , \3474 );
nand \U$3383 ( \3476 , RI8928830_3, RI8929730_35);
not \U$3384 ( \3477 , \3476 );
not \U$3385 ( \3478 , \2819 );
or \U$3386 ( \3479 , \3477 , \3478 );
nand \U$3387 ( \3480 , \181 , \2823 );
nand \U$3388 ( \3481 , \3479 , \3480 );
not \U$3389 ( \3482 , \3481 );
or \U$3390 ( \3483 , \3475 , \3482 );
not \U$3391 ( \3484 , RI89287b8_2);
nand \U$3392 ( \3485 , \3185 , \3484 );
nand \U$3393 ( \3486 , \3483 , \3485 );
xnor \U$3394 ( \3487 , \3473 , \3486 );
nand \U$3395 ( \3488 , \3487 , \1818 );
nand \U$3396 ( \3489 , \3466 , \3469 , \3470 , \3488 );
nor \U$3397 ( \3490 , \3429 , \3489 );
xor \U$3398 ( \3491 , \3042 , \3069 );
and \U$3399 ( \3492 , \3491 , \3074 );
and \U$3400 ( \3493 , \3042 , \3069 );
or \U$3401 ( \3494 , \3492 , \3493 );
xor \U$3402 ( \3495 , \3050 , \3059 );
and \U$3403 ( \3496 , \3495 , \3068 );
and \U$3404 ( \3497 , \3050 , \3059 );
or \U$3405 ( \3498 , \3496 , \3497 );
not \U$3406 ( \3499 , \3037 );
not \U$3407 ( \3500 , \3030 );
or \U$3408 ( \3501 , \3499 , \3500 );
nand \U$3409 ( \3502 , \3028 , \3018 );
nand \U$3410 ( \3503 , \3501 , \3502 );
xor \U$3411 ( \3504 , \3498 , \3503 );
not \U$3412 ( \3505 , \3062 );
or \U$3413 ( \3506 , \3505 , \3065 );
not \U$3414 ( \3507 , \1257 );
and \U$3415 ( \3508 , RI892a360_61, \1781 );
not \U$3416 ( \3509 , RI892a360_61);
and \U$3417 ( \3510 , \3509 , RI89288a8_4);
nor \U$3418 ( \3511 , \3508 , \3510 );
or \U$3419 ( \3512 , \3507 , \3511 );
nand \U$3420 ( \3513 , \3506 , \3512 );
not \U$3421 ( \3514 , \3513 );
xnor \U$3422 ( \3515 , RI89287b8_2, RI892a450_63);
not \U$3423 ( \3516 , \3515 );
not \U$3424 ( \3517 , RI892a4c8_64);
not \U$3425 ( \3518 , \3517 );
and \U$3426 ( \3519 , \3516 , \3518 );
and \U$3427 ( \3520 , \1291 , \2975 );
nor \U$3428 ( \3521 , \3519 , \3520 );
and \U$3429 ( \3522 , RI8929eb0_51, RI8929e38_50);
not \U$3430 ( \3523 , RI8929eb0_51);
and \U$3431 ( \3524 , \3523 , \3440 );
nor \U$3432 ( \3525 , \3522 , \3524 );
and \U$3433 ( \3526 , \3525 , RI8928e48_16);
and \U$3434 ( \3527 , \3521 , \3526 );
not \U$3435 ( \3528 , \3521 );
not \U$3436 ( \3529 , \3526 );
and \U$3437 ( \3530 , \3528 , \3529 );
nor \U$3438 ( \3531 , \3527 , \3530 );
not \U$3439 ( \3532 , \3531 );
or \U$3440 ( \3533 , \3514 , \3532 );
or \U$3441 ( \3534 , \3531 , \3513 );
nand \U$3442 ( \3535 , \3533 , \3534 );
xor \U$3443 ( \3536 , \3504 , \3535 );
xor \U$3444 ( \3537 , \3494 , \3536 );
not \U$3445 ( \3538 , \3057 );
not \U$3446 ( \3539 , \3052 );
or \U$3447 ( \3540 , \3538 , \3539 );
xnor \U$3448 ( \3541 , RI8928b78_10, RI892a090_55);
or \U$3449 ( \3542 , \3055 , \3541 );
nand \U$3450 ( \3543 , \3540 , \3542 );
not \U$3451 ( \3544 , \3048 );
not \U$3452 ( \3545 , \3044 );
or \U$3453 ( \3546 , \3544 , \3545 );
xnor \U$3454 ( \3547 , RI892a180_57, RI8928a88_8);
not \U$3455 ( \3548 , \3547 );
nand \U$3456 ( \3549 , \3548 , \3047 );
nand \U$3457 ( \3550 , \3546 , \3549 );
xor \U$3458 ( \3551 , \3543 , \3550 );
not \U$3459 ( \3552 , \2285 );
or \U$3460 ( \3553 , \3552 , \3034 );
not \U$3461 ( \3554 , \1232 );
and \U$3462 ( \3555 , RI892a270_59, \834 );
not \U$3463 ( \3556 , RI892a270_59);
and \U$3464 ( \3557 , \3556 , RI8928998_6);
nor \U$3465 ( \3558 , \3555 , \3557 );
or \U$3466 ( \3559 , \3554 , \3558 );
nand \U$3467 ( \3560 , \3553 , \3559 );
xor \U$3468 ( \3561 , \3551 , \3560 );
xor \U$3469 ( \3562 , RI8929fa0_53, RI8928c68_12);
and \U$3470 ( \3563 , \2275 , \3562 );
and \U$3471 ( \3564 , \3013 , \3016 );
nor \U$3472 ( \3565 , \3563 , \3564 );
not \U$3473 ( \3566 , \3565 );
not \U$3474 ( \3567 , \2644 );
xor \U$3475 ( \3568 , RI8929eb0_51, RI8928d58_14);
not \U$3476 ( \3569 , \3568 );
or \U$3477 ( \3570 , \3567 , \3569 );
nand \U$3478 ( \3571 , \3020 , \3023 );
nand \U$3479 ( \3572 , \3570 , \3571 );
not \U$3480 ( \3573 , \3572 );
or \U$3481 ( \3574 , \3566 , \3573 );
or \U$3482 ( \3575 , \3565 , \3572 );
nand \U$3483 ( \3576 , \3574 , \3575 );
not \U$3484 ( \3577 , \3576 );
not \U$3485 ( \3578 , \2982 );
nand \U$3486 ( \3579 , \3578 , \2977 );
not \U$3487 ( \3580 , \3579 );
or \U$3488 ( \3581 , \3577 , \3580 );
or \U$3489 ( \3582 , \3576 , \3579 );
nand \U$3490 ( \3583 , \3581 , \3582 );
xor \U$3491 ( \3584 , \3561 , \3583 );
not \U$3492 ( \3585 , \2992 );
buf \U$3493 ( \3586 , \2986 );
nand \U$3494 ( \3587 , \3585 , \3586 );
and \U$3495 ( \3588 , \3587 , \3000 );
nor \U$3496 ( \3589 , \3585 , \3586 );
nor \U$3497 ( \3590 , \3588 , \3589 );
not \U$3498 ( \3591 , \3590 );
and \U$3499 ( \3592 , \3584 , \3591 );
not \U$3500 ( \3593 , \3584 );
and \U$3501 ( \3594 , \3593 , \3590 );
nor \U$3502 ( \3595 , \3592 , \3594 );
and \U$3503 ( \3596 , \3537 , \3595 );
and \U$3504 ( \3597 , \3494 , \3536 );
or \U$3505 ( \3598 , \3596 , \3597 );
not \U$3506 ( \3599 , \3598 );
xor \U$3507 ( \3600 , \3543 , \3550 );
and \U$3508 ( \3601 , \3600 , \3560 );
and \U$3509 ( \3602 , \3543 , \3550 );
nor \U$3510 ( \3603 , \3601 , \3602 );
not \U$3511 ( \3604 , \3603 );
not \U$3512 ( \3605 , \3576 );
not \U$3513 ( \3606 , \3579 );
not \U$3514 ( \3607 , \3606 );
or \U$3515 ( \3608 , \3605 , \3607 );
not \U$3516 ( \3609 , \3565 );
nand \U$3517 ( \3610 , \3609 , \3572 );
nand \U$3518 ( \3611 , \3608 , \3610 );
and \U$3519 ( \3612 , RI8928dd0_15, RI8929dc0_49);
not \U$3520 ( \3613 , RI8928dd0_15);
and \U$3521 ( \3614 , \3613 , \95 );
nor \U$3522 ( \3615 , \3612 , \3614 );
and \U$3523 ( \3616 , \3525 , \3615 );
not \U$3524 ( \3617 , \3525 );
not \U$3525 ( \3618 , RI8929dc0_49);
nor \U$3526 ( \3619 , RI8928e48_16, RI8929e38_50);
not \U$3527 ( \3620 , \3619 );
or \U$3528 ( \3621 , \3618 , \3620 );
nand \U$3529 ( \3622 , RI8928e48_16, RI8929e38_50);
not \U$3530 ( \3623 , \3622 );
nand \U$3531 ( \3624 , \3623 , \95 );
nand \U$3532 ( \3625 , \3621 , \3624 );
and \U$3533 ( \3626 , \3617 , \3625 );
nor \U$3534 ( \3627 , \3616 , \3626 );
not \U$3535 ( \3628 , \3627 );
not \U$3536 ( \3629 , \3562 );
not \U$3537 ( \3630 , \2276 );
or \U$3538 ( \3631 , \3629 , \3630 );
xor \U$3539 ( \3632 , RI8928bf0_11, RI8929fa0_53);
nand \U$3540 ( \3633 , \2275 , \3632 );
nand \U$3541 ( \3634 , \3631 , \3633 );
not \U$3542 ( \3635 , \3634 );
or \U$3543 ( \3636 , \3628 , \3635 );
or \U$3544 ( \3637 , \3627 , \3634 );
nand \U$3545 ( \3638 , \3636 , \3637 );
not \U$3546 ( \3639 , \3044 );
or \U$3547 ( \3640 , \3639 , \3547 );
not \U$3548 ( \3641 , \3047 );
xnor \U$3549 ( \3642 , RI892a180_57, RI8928a10_7);
or \U$3550 ( \3643 , \3641 , \3642 );
nand \U$3551 ( \3644 , \3640 , \3643 );
or \U$3552 ( \3645 , \3638 , \3644 );
nand \U$3553 ( \3646 , \3638 , \3644 );
nand \U$3554 ( \3647 , \3645 , \3646 );
and \U$3555 ( \3648 , \3611 , \3647 );
not \U$3556 ( \3649 , \3611 );
not \U$3557 ( \3650 , \3647 );
and \U$3558 ( \3651 , \3649 , \3650 );
nor \U$3559 ( \3652 , \3648 , \3651 );
not \U$3560 ( \3653 , \3652 );
or \U$3561 ( \3654 , \3604 , \3653 );
or \U$3562 ( \3655 , \3603 , \3652 );
nand \U$3563 ( \3656 , \3654 , \3655 );
not \U$3564 ( \3657 , \3584 );
not \U$3565 ( \3658 , \3591 );
or \U$3566 ( \3659 , \3657 , \3658 );
nand \U$3567 ( \3660 , \3561 , \3583 );
nand \U$3568 ( \3661 , \3659 , \3660 );
xor \U$3569 ( \3662 , \3656 , \3661 );
not \U$3570 ( \3663 , \3521 );
not \U$3571 ( \3664 , \3529 );
and \U$3572 ( \3665 , \3663 , \3664 );
not \U$3573 ( \3666 , \3531 );
and \U$3574 ( \3667 , \3666 , \3513 );
nor \U$3575 ( \3668 , \3665 , \3667 );
not \U$3576 ( \3669 , \3511 );
not \U$3577 ( \3670 , \3669 );
not \U$3578 ( \3671 , \3062 );
or \U$3579 ( \3672 , \3670 , \3671 );
and \U$3580 ( \3673 , RI892a360_61, RI8928830_3);
not \U$3581 ( \3674 , RI892a360_61);
and \U$3582 ( \3675 , \3674 , \2823 );
nor \U$3583 ( \3676 , \3673 , \3675 );
nand \U$3584 ( \3677 , \1257 , \3676 );
nand \U$3585 ( \3678 , \3672 , \3677 );
not \U$3586 ( \3679 , \3052 );
or \U$3587 ( \3680 , \3679 , \3541 );
xnor \U$3588 ( \3681 , RI892a090_55, RI8928b00_9);
or \U$3589 ( \3682 , \3055 , \3681 );
nand \U$3590 ( \3683 , \3680 , \3682 );
and \U$3591 ( \3684 , \3678 , \3683 );
not \U$3592 ( \3685 , \3678 );
not \U$3593 ( \3686 , \3683 );
and \U$3594 ( \3687 , \3685 , \3686 );
nor \U$3595 ( \3688 , \3684 , \3687 );
xor \U$3596 ( \3689 , \3668 , \3688 );
or \U$3597 ( \3690 , RI8928e48_16, RI8929e38_50);
nand \U$3598 ( \3691 , \3690 , RI8929eb0_51);
nand \U$3599 ( \3692 , \3691 , \3622 , RI8929dc0_49);
and \U$3600 ( \3693 , \3020 , \3568 );
xor \U$3601 ( \3694 , RI8929eb0_51, RI8928ce0_13);
and \U$3602 ( \3695 , \2644 , \3694 );
nor \U$3603 ( \3696 , \3693 , \3695 );
xor \U$3604 ( \3697 , \3692 , \3696 );
not \U$3605 ( \3698 , \1291 );
or \U$3606 ( \3699 , \3698 , \3515 );
and \U$3607 ( \3700 , RI892a450_63, \3462 );
not \U$3608 ( \3701 , RI892a450_63);
and \U$3609 ( \3702 , \3701 , RI8928740_1);
nor \U$3610 ( \3703 , \3700 , \3702 );
or \U$3611 ( \3704 , \3517 , \3703 );
nand \U$3612 ( \3705 , \3699 , \3704 );
xnor \U$3613 ( \3706 , \3697 , \3705 );
or \U$3614 ( \3707 , \3552 , \3558 );
and \U$3615 ( \3708 , \115 , RI8928920_5);
and \U$3616 ( \3709 , \1808 , RI892a270_59);
nor \U$3617 ( \3710 , \3708 , \3709 );
or \U$3618 ( \3711 , \3554 , \3710 );
nand \U$3619 ( \3712 , \3707 , \3711 );
xor \U$3620 ( \3713 , \3706 , \3712 );
xor \U$3621 ( \3714 , \3689 , \3713 );
xor \U$3622 ( \3715 , \3498 , \3503 );
and \U$3623 ( \3716 , \3715 , \3535 );
and \U$3624 ( \3717 , \3498 , \3503 );
or \U$3625 ( \3718 , \3716 , \3717 );
not \U$3626 ( \3719 , \3718 );
and \U$3627 ( \3720 , \3714 , \3719 );
not \U$3628 ( \3721 , \3714 );
and \U$3629 ( \3722 , \3721 , \3718 );
nor \U$3630 ( \3723 , \3720 , \3722 );
xnor \U$3631 ( \3724 , \3662 , \3723 );
not \U$3632 ( \3725 , \3724 );
or \U$3633 ( \3726 , \3599 , \3725 );
or \U$3634 ( \3727 , \3724 , \3598 );
nand \U$3635 ( \3728 , \3726 , \3727 );
not \U$3636 ( \3729 , \3728 );
xor \U$3637 ( \3730 , \3494 , \3536 );
xor \U$3638 ( \3731 , \3730 , \3595 );
xor \U$3639 ( \3732 , \3001 , \3010 );
and \U$3640 ( \3733 , \3732 , \3075 );
and \U$3641 ( \3734 , \3001 , \3010 );
or \U$3642 ( \3735 , \3733 , \3734 );
or \U$3643 ( \3736 , \3731 , \3735 );
not \U$3644 ( \3737 , \3736 );
buf \U$3645 ( \3738 , \3087 );
and \U$3646 ( \3739 , \3095 , \3738 );
not \U$3647 ( \3740 , \3085 );
nor \U$3648 ( \3741 , \3739 , \3740 );
not \U$3649 ( \3742 , \3741 );
or \U$3650 ( \3743 , \3737 , \3742 );
nand \U$3651 ( \3744 , \3731 , \3735 );
nand \U$3652 ( \3745 , \3743 , \3744 );
not \U$3653 ( \3746 , \3745 );
or \U$3654 ( \3747 , \3729 , \3746 );
not \U$3655 ( \3748 , \3745 );
not \U$3656 ( \3749 , \3728 );
and \U$3657 ( \3750 , \3748 , \3749 );
not \U$3658 ( \3751 , \2732 );
nor \U$3659 ( \3752 , \3750 , \3751 );
nand \U$3660 ( \3753 , \3747 , \3752 );
nand \U$3661 ( \3754 , \3490 , \3753 );
buf \U$3662 ( \3755 , \3754 );
not \U$3663 ( \3756 , \3755 );
or \U$3664 ( \3757 , \3152 , \3756 );
or \U$3665 ( \3758 , \3755 , \3151 );
nand \U$3666 ( \3759 , \3757 , \3758 );
not \U$3667 ( \3760 , \3759 );
not \U$3668 ( \3761 , \3753 );
buf \U$3669 ( \3762 , \1733 );
and \U$3670 ( \3763 , \3762 , RI8929e38_50);
nand \U$3671 ( \3764 , \2739 , RI89296b8_34);
and \U$3672 ( \3765 , \3764 , \2736 );
nor \U$3673 ( \3766 , \3765 , \3439 );
nor \U$3674 ( \3767 , \3763 , \3766 );
not \U$3675 ( \3768 , \3428 );
nand \U$3676 ( \3769 , \3276 , \3287 );
buf \U$3677 ( \3770 , \3283 );
xnor \U$3678 ( \3771 , \3769 , \3770 );
nand \U$3679 ( \3772 , \3768 , \3771 );
not \U$3680 ( \3773 , RI89287b8_2);
not \U$3681 ( \3774 , \1575 );
nand \U$3682 ( \3775 , \3774 , \777 );
not \U$3683 ( \3776 , \3775 );
or \U$3684 ( \3777 , \3773 , \3776 );
xor \U$3685 ( \3778 , \3439 , \3440 );
not \U$3686 ( \3779 , \3778 );
not \U$3687 ( \3780 , \3436 );
or \U$3688 ( \3781 , \3779 , \3780 );
or \U$3689 ( \3782 , \3436 , \3778 );
nand \U$3690 ( \3783 , \3781 , \3782 );
nand \U$3691 ( \3784 , \3783 , \1779 );
nand \U$3692 ( \3785 , \3777 , \3784 );
and \U$3693 ( \3786 , \3440 , RI89296b8_34);
and \U$3694 ( \3787 , \3185 , RI8929e38_50);
nor \U$3695 ( \3788 , \3786 , \3787 );
not \U$3696 ( \3789 , \3788 );
nand \U$3697 ( \3790 , \1741 , \3789 );
and \U$3698 ( \3791 , \3185 , RI89287b8_2);
and \U$3699 ( \3792 , \3484 , RI89296b8_34);
nor \U$3700 ( \3793 , \3791 , \3792 );
xor \U$3701 ( \3794 , \3793 , \3481 );
nand \U$3702 ( \3795 , \3794 , \1818 );
nand \U$3703 ( \3796 , \418 , RI89296b8_34);
nand \U$3704 ( \3797 , \3790 , \3795 , \3796 );
nor \U$3705 ( \3798 , \3785 , \3797 );
nand \U$3706 ( \3799 , \3736 , \3744 );
not \U$3707 ( \3800 , \3799 );
buf \U$3708 ( \3801 , \3741 );
not \U$3709 ( \3802 , \3801 );
or \U$3710 ( \3803 , \3800 , \3802 );
or \U$3711 ( \3804 , \3801 , \3799 );
nand \U$3712 ( \3805 , \3803 , \3804 );
nand \U$3713 ( \3806 , \3805 , \2732 );
nand \U$3714 ( \3807 , \3767 , \3772 , \3798 , \3806 );
not \U$3715 ( \3808 , \3807 );
nand \U$3716 ( \3809 , \3761 , \3114 , \3808 );
not \U$3717 ( \3810 , \3490 );
nand \U$3718 ( \3811 , \3808 , \3810 , \3114 );
nand \U$3719 ( \3812 , \3109 , \3490 , \3807 , \3753 );
nand \U$3720 ( \3813 , \3809 , \3811 , \3812 );
buf \U$3721 ( \3814 , \3813 );
buf \U$3722 ( \3815 , \3814 );
not \U$3723 ( \3816 , \3815 );
or \U$3724 ( \3817 , \3760 , \3816 );
or \U$3725 ( \3818 , \159 , RI892a090_55);
or \U$3726 ( \3819 , \160 , RI8929910_39);
nand \U$3727 ( \3820 , \3818 , \3819 );
xnor \U$3728 ( \3821 , \156 , \3820 );
not \U$3729 ( \3822 , \3821 );
buf \U$3730 ( \3823 , \3755 );
xnor \U$3731 ( \3824 , \3822 , \3823 );
not \U$3732 ( \3825 , \3107 );
not \U$3733 ( \3826 , \3825 );
not \U$3734 ( \3827 , \3808 );
or \U$3735 ( \3828 , \3826 , \3827 );
not \U$3736 ( \3829 , \3825 );
nand \U$3737 ( \3830 , \3829 , \3807 );
nand \U$3738 ( \3831 , \3828 , \3830 );
not \U$3739 ( \3832 , \3831 );
buf \U$3740 ( \3833 , \3832 );
nand \U$3741 ( \3834 , \3824 , \3833 );
nand \U$3742 ( \3835 , \3817 , \3834 );
xor \U$3743 ( \3836 , \3145 , \3835 );
buf \U$3744 ( \3837 , \3836 );
not \U$3745 ( \3838 , \3837 );
and \U$3746 ( \3839 , \142 , \1585 );
not \U$3747 ( \3840 , \142 );
not \U$3748 ( \3841 , \1585 );
and \U$3749 ( \3842 , \3840 , \3841 );
or \U$3750 ( \3843 , \3839 , \3842 );
not \U$3751 ( \3844 , \3843 );
and \U$3752 ( \3845 , \3823 , \3844 );
not \U$3753 ( \3846 , \3845 );
not \U$3754 ( \3847 , RI8928c68_12);
not \U$3755 ( \3848 , \3775 );
or \U$3756 ( \3849 , \3847 , \3848 );
and \U$3757 ( \3850 , \1575 , RI892a2e8_60);
not \U$3758 ( \3851 , RI89293e8_28);
not \U$3759 ( \3852 , RI8929b68_44);
not \U$3760 ( \3853 , \1554 );
or \U$3761 ( \3854 , \3852 , \3853 );
nand \U$3762 ( \3855 , \3854 , \776 );
not \U$3763 ( \3856 , \3855 );
or \U$3764 ( \3857 , \3851 , \3856 );
or \U$3765 ( \3858 , \119 , RI892a2e8_60);
or \U$3766 ( \3859 , \118 , RI8929b68_44);
nand \U$3767 ( \3860 , \3858 , \3859 );
and \U$3768 ( \3861 , \1741 , \3860 );
xor \U$3769 ( \3862 , \927 , \960 );
xor \U$3770 ( \3863 , \3862 , \997 );
or \U$3771 ( \3864 , \2267 , \3863 );
not \U$3772 ( \3865 , \1433 );
not \U$3773 ( \3866 , \3865 );
and \U$3774 ( \3867 , \1394 , \1388 );
not \U$3775 ( \3868 , \1437 );
nor \U$3776 ( \3869 , \3867 , \3868 );
not \U$3777 ( \3870 , \3869 );
or \U$3778 ( \3871 , \3866 , \3870 );
or \U$3779 ( \3872 , \3869 , \3865 );
nand \U$3780 ( \3873 , \3871 , \3872 );
not \U$3781 ( \3874 , \3873 );
not \U$3782 ( \3875 , \402 );
or \U$3783 ( \3876 , \3874 , \3875 );
not \U$3784 ( \3877 , \1474 );
nor \U$3785 ( \3878 , \3877 , \1471 );
not \U$3786 ( \3879 , \3878 );
not \U$3787 ( \3880 , \1670 );
or \U$3788 ( \3881 , \3879 , \3880 );
or \U$3789 ( \3882 , \1670 , \3878 );
nand \U$3790 ( \3883 , \3881 , \3882 );
and \U$3791 ( \3884 , \3883 , \1600 );
not \U$3792 ( \3885 , \1517 );
nor \U$3793 ( \3886 , \3885 , \1500 );
not \U$3794 ( \3887 , \3886 );
not \U$3795 ( \3888 , \1683 );
or \U$3796 ( \3889 , \3887 , \3888 );
or \U$3797 ( \3890 , \1683 , \3886 );
nand \U$3798 ( \3891 , \3889 , \3890 );
not \U$3799 ( \3892 , \3891 );
not \U$3800 ( \3893 , \410 );
or \U$3801 ( \3894 , \3892 , \3893 );
and \U$3802 ( \3895 , \413 , RI892a2e8_60);
or \U$3803 ( \3896 , \419 , \119 );
or \U$3804 ( \3897 , \424 , \478 );
nand \U$3805 ( \3898 , \3896 , \3897 );
nor \U$3806 ( \3899 , \3895 , \3898 );
nand \U$3807 ( \3900 , \3894 , \3899 );
nor \U$3808 ( \3901 , \3884 , \3900 );
nand \U$3809 ( \3902 , \3876 , \3901 );
not \U$3810 ( \3903 , \3902 );
nand \U$3811 ( \3904 , \3864 , \3903 );
nor \U$3812 ( \3905 , \3861 , \3904 );
nand \U$3813 ( \3906 , \3857 , \3905 );
nor \U$3814 ( \3907 , \3850 , \3906 );
nand \U$3815 ( \3908 , \3849 , \3907 );
not \U$3816 ( \3909 , RI8928ce0_13);
not \U$3817 ( \3910 , \1571 );
or \U$3818 ( \3911 , \3909 , \3910 );
and \U$3819 ( \3912 , \1575 , RI892a360_61);
not \U$3820 ( \3913 , \996 );
nand \U$3821 ( \3914 , \3913 , \974 );
xnor \U$3822 ( \3915 , \994 , \3914 );
not \U$3823 ( \3916 , \1180 );
and \U$3824 ( \3917 , \3915 , \3916 );
nand \U$3825 ( \3918 , \1432 , \1407 );
xnor \U$3826 ( \3919 , \1428 , \3918 );
not \U$3827 ( \3920 , \3919 );
not \U$3828 ( \3921 , \402 );
or \U$3829 ( \3922 , \3920 , \3921 );
not \U$3830 ( \3923 , \1668 );
not \U$3831 ( \3924 , \1469 );
or \U$3832 ( \3925 , \3923 , \3924 );
or \U$3833 ( \3926 , \1468 , \1470 );
nand \U$3834 ( \3927 , \3926 , \1467 );
nand \U$3835 ( \3928 , \3925 , \3927 );
and \U$3836 ( \3929 , \1600 , \3928 );
not \U$3837 ( \3930 , \1514 );
and \U$3838 ( \3931 , \3930 , \1680 );
nand \U$3839 ( \3932 , \1680 , \1513 );
and \U$3840 ( \3933 , \1679 , \3932 );
nor \U$3841 ( \3934 , \3931 , \3933 );
or \U$3842 ( \3935 , \1678 , \3934 );
and \U$3843 ( \3936 , \413 , RI892a360_61);
and \U$3844 ( \3937 , \418 , RI8929be0_45);
and \U$3845 ( \3938 , \423 , RI8929460_29);
nor \U$3846 ( \3939 , \3936 , \3937 , \3938 );
nand \U$3847 ( \3940 , \3935 , \3939 );
nor \U$3848 ( \3941 , \3929 , \3940 );
nand \U$3849 ( \3942 , \3922 , \3941 );
nor \U$3850 ( \3943 , \3917 , \3942 );
and \U$3851 ( \3944 , RI892a360_61, RI8929be0_45);
not \U$3852 ( \3945 , RI892a360_61);
not \U$3853 ( \3946 , RI8929be0_45);
and \U$3854 ( \3947 , \3945 , \3946 );
nor \U$3855 ( \3948 , \3944 , \3947 );
nand \U$3856 ( \3949 , \1549 , \3948 );
not \U$3857 ( \3950 , RI8929460_29);
nor \U$3858 ( \3951 , \3950 , \3946 );
nand \U$3859 ( \3952 , \1644 , \3951 );
nand \U$3860 ( \3953 , \3950 , \1345 );
nand \U$3861 ( \3954 , \1547 , \3953 );
nand \U$3862 ( \3955 , \3943 , \3949 , \3952 , \3954 );
nor \U$3863 ( \3956 , \3912 , \3955 );
nand \U$3864 ( \3957 , \3911 , \3956 );
xor \U$3865 ( \3958 , \3908 , \3957 );
not \U$3866 ( \3959 , \3958 );
not \U$3867 ( \3960 , \3908 );
not \U$3868 ( \3961 , \3960 );
and \U$3869 ( \3962 , \1710 , \3961 );
not \U$3870 ( \3963 , \1710 );
and \U$3871 ( \3964 , \3963 , \3960 );
nor \U$3872 ( \3965 , \3962 , \3964 );
nand \U$3873 ( \3966 , \3959 , \3965 );
not \U$3874 ( \3967 , \3966 );
not \U$3875 ( \3968 , \192 );
not \U$3876 ( \3969 , \1710 );
not \U$3877 ( \3970 , \3969 );
or \U$3878 ( \3971 , \3968 , \3970 );
or \U$3879 ( \3972 , \192 , \3969 );
nand \U$3880 ( \3973 , \3971 , \3972 );
nand \U$3881 ( \3974 , \3967 , \3973 );
buf \U$3882 ( \3975 , \3958 );
buf \U$3883 ( \3976 , \3975 );
buf \U$3884 ( \3977 , \1710 );
nand \U$3885 ( \3978 , \3976 , \3977 );
and \U$3886 ( \3979 , \3974 , \3978 );
nand \U$3887 ( \3980 , \3846 , \3979 );
not \U$3888 ( \3981 , \3980 );
not \U$3889 ( \3982 , \3126 );
buf \U$3890 ( \3983 , \2794 );
not \U$3891 ( \3984 , \3983 );
not \U$3892 ( \3985 , \3984 );
or \U$3893 ( \3986 , \3982 , \3985 );
not \U$3894 ( \3987 , \3983 );
or \U$3895 ( \3988 , \3987 , \3126 );
nand \U$3896 ( \3989 , \3986 , \3988 );
not \U$3897 ( \3990 , \3989 );
not \U$3898 ( \3991 , \1730 );
not \U$3899 ( \3992 , \3991 );
not \U$3900 ( \3993 , \2747 );
not \U$3901 ( \3994 , \3993 );
or \U$3902 ( \3995 , \3992 , \3994 );
nand \U$3903 ( \3996 , \3995 , RI892a018_54);
nand \U$3904 ( \3997 , \2779 , RI8928998_6);
not \U$3905 ( \3998 , \2228 );
not \U$3906 ( \3999 , \3998 );
buf \U$3907 ( \4000 , \2227 );
not \U$3908 ( \4001 , \4000 );
or \U$3909 ( \4002 , \3999 , \4001 );
not \U$3910 ( \4003 , \2254 );
nand \U$3911 ( \4004 , \4002 , \4003 );
buf \U$3912 ( \4005 , \2249 );
not \U$3913 ( \4006 , \4005 );
nand \U$3914 ( \4007 , \4004 , \4006 );
nand \U$3915 ( \4008 , \2258 , \2207 );
not \U$3916 ( \4009 , \4008 );
and \U$3917 ( \4010 , \4007 , \4009 );
nor \U$3918 ( \4011 , \4010 , \2267 );
not \U$3919 ( \4012 , \4011 );
nand \U$3920 ( \4013 , \4004 , \4008 , \4006 );
not \U$3921 ( \4014 , \4013 );
or \U$3922 ( \4015 , \4012 , \4014 );
and \U$3923 ( \4016 , \1741 , \3121 );
and \U$3924 ( \4017 , RI8929118_22, RI892a018_54);
not \U$3925 ( \4018 , RI8929118_22);
and \U$3926 ( \4019 , \4018 , \166 );
nor \U$3927 ( \4020 , \4017 , \4019 );
xor \U$3928 ( \4021 , \1769 , \4020 );
not \U$3929 ( \4022 , \1779 );
or \U$3930 ( \4023 , \4021 , \4022 );
xor \U$3931 ( \4024 , \165 , \834 );
not \U$3932 ( \4025 , \4024 );
not \U$3933 ( \4026 , \1804 );
or \U$3934 ( \4027 , \4025 , \4026 );
or \U$3935 ( \4028 , \1804 , \4024 );
nand \U$3936 ( \4029 , \4027 , \4028 );
and \U$3937 ( \4030 , \1818 , \4029 );
and \U$3938 ( \4031 , RI8929898_38, \418 );
nor \U$3939 ( \4032 , \4030 , \4031 );
nand \U$3940 ( \4033 , \4023 , \4032 );
nor \U$3941 ( \4034 , \4016 , \4033 );
nand \U$3942 ( \4035 , \4015 , \4034 );
not \U$3943 ( \4036 , RI8928998_6);
not \U$3944 ( \4037 , \1735 );
or \U$3945 ( \4038 , \4036 , \4037 );
not \U$3946 ( \4039 , \2613 );
nand \U$3947 ( \4040 , \2515 , \2546 );
nand \U$3948 ( \4041 , \4039 , \4040 );
not \U$3949 ( \4042 , \4041 );
buf \U$3950 ( \4043 , \2610 );
nand \U$3951 ( \4044 , \4043 , \2572 );
and \U$3952 ( \4045 , \4042 , \4044 );
nor \U$3953 ( \4046 , \4045 , \2731 );
nand \U$3954 ( \4047 , \4043 , \4041 , \2572 );
nand \U$3955 ( \4048 , \4046 , \4047 );
nand \U$3956 ( \4049 , \4038 , \4048 );
nor \U$3957 ( \4050 , \4035 , \4049 );
not \U$3958 ( \4051 , RI8929898_38);
not \U$3959 ( \4052 , \2739 );
or \U$3960 ( \4053 , \4051 , \4052 );
nand \U$3961 ( \4054 , \4053 , \2736 );
nand \U$3962 ( \4055 , \4054 , RI8929118_22);
nand \U$3963 ( \4056 , \3996 , \3997 , \4050 , \4055 );
not \U$3964 ( \4057 , \4056 );
not \U$3965 ( \4058 , \4057 );
not \U$3966 ( \4059 , RI8928a10_7);
not \U$3967 ( \4060 , \1571 );
or \U$3968 ( \4061 , \4059 , \4060 );
and \U$3969 ( \4062 , \911 , RI892a090_55);
not \U$3970 ( \4063 , \2608 );
nand \U$3971 ( \4064 , \4063 , \2572 );
not \U$3972 ( \4065 , \4064 );
not \U$3973 ( \4066 , \2607 );
and \U$3974 ( \4067 , \4065 , \4066 );
and \U$3975 ( \4068 , \4064 , \2607 );
nor \U$3976 ( \4069 , \4067 , \4068 );
not \U$3977 ( \4070 , \4069 );
not \U$3978 ( \4071 , \2731 );
and \U$3979 ( \4072 , \4070 , \4071 );
and \U$3980 ( \4073 , \1549 , \3820 );
nor \U$3981 ( \4074 , \4072 , \4073 );
not \U$3982 ( \4075 , RI8929190_23);
not \U$3983 ( \4076 , \690 );
not \U$3984 ( \4077 , \4076 );
or \U$3985 ( \4078 , \4075 , \4077 );
nand \U$3986 ( \4079 , \4078 , \419 );
nand \U$3987 ( \4080 , \4079 , RI8929910_39);
not \U$3988 ( \4081 , \4005 );
nand \U$3989 ( \4082 , \4081 , \4003 );
not \U$3990 ( \4083 , \4082 );
nand \U$3991 ( \4084 , \4000 , \3998 );
not \U$3992 ( \4085 , \4084 );
or \U$3993 ( \4086 , \4083 , \4085 );
or \U$3994 ( \4087 , \4084 , \4082 );
nand \U$3995 ( \4088 , \4086 , \4087 );
not \U$3996 ( \4089 , \730 );
buf \U$3997 ( \4090 , \4089 );
and \U$3998 ( \4091 , \4088 , \4090 );
and \U$3999 ( \4092 , \1768 , \1753 );
xnor \U$4000 ( \4093 , \4092 , \1764 );
not \U$4001 ( \4094 , \4093 );
not \U$4002 ( \4095 , \1779 );
or \U$4003 ( \4096 , \4094 , \4095 );
and \U$4004 ( \4097 , \1803 , \1787 );
not \U$4005 ( \4098 , \4097 );
not \U$4006 ( \4099 , \1800 );
or \U$4007 ( \4100 , \4098 , \4099 );
or \U$4008 ( \4101 , \1800 , \4097 );
nand \U$4009 ( \4102 , \4100 , \4101 );
and \U$4010 ( \4103 , \1817 , \4102 );
or \U$4011 ( \4104 , \3991 , \160 );
or \U$4012 ( \4105 , \424 , \1767 );
nand \U$4013 ( \4106 , \4104 , \4105 );
nor \U$4014 ( \4107 , \4103 , \4106 );
nand \U$4015 ( \4108 , \4096 , \4107 );
nor \U$4016 ( \4109 , \4091 , \4108 );
not \U$4017 ( \4110 , RI8928a10_7);
nand \U$4018 ( \4111 , \4110 , \1767 );
nand \U$4019 ( \4112 , \4111 , \1547 );
nand \U$4020 ( \4113 , \4074 , \4080 , \4109 , \4112 );
nor \U$4021 ( \4114 , \4062 , \4113 );
nand \U$4022 ( \4115 , \4061 , \4114 );
buf \U$4023 ( \4116 , \4115 );
not \U$4024 ( \4117 , \4116 );
not \U$4025 ( \4118 , \4117 );
or \U$4026 ( \4119 , \4058 , \4118 );
not \U$4027 ( \4120 , \4115 );
not \U$4028 ( \4121 , \4120 );
nand \U$4029 ( \4122 , \4056 , \4121 );
nand \U$4030 ( \4123 , \4119 , \4122 );
not \U$4031 ( \4124 , \4057 );
not \U$4032 ( \4125 , \2794 );
or \U$4033 ( \4126 , \4124 , \4125 );
and \U$4034 ( \4127 , \3996 , \3997 , \4050 , \4055 );
or \U$4035 ( \4128 , \3983 , \4127 );
nand \U$4036 ( \4129 , \4126 , \4128 );
nand \U$4037 ( \4130 , \4123 , \4129 );
not \U$4038 ( \4131 , \4130 );
not \U$4039 ( \4132 , \4131 );
or \U$4040 ( \4133 , \3990 , \4132 );
not \U$4041 ( \4134 , \4123 );
buf \U$4042 ( \4135 , \4134 );
not \U$4043 ( \4136 , \2803 );
buf \U$4044 ( \4137 , \3983 );
not \U$4045 ( \4138 , \4137 );
or \U$4046 ( \4139 , \4136 , \4138 );
not \U$4047 ( \4140 , \3984 );
or \U$4048 ( \4141 , \4140 , \2803 );
nand \U$4049 ( \4142 , \4139 , \4141 );
nand \U$4050 ( \4143 , \4135 , \4142 );
nand \U$4051 ( \4144 , \4133 , \4143 );
not \U$4052 ( \4145 , \4144 );
and \U$4053 ( \4146 , \1712 , \1717 );
not \U$4054 ( \4147 , \4146 );
and \U$4055 ( \4148 , \184 , \3789 );
not \U$4056 ( \4149 , \184 );
and \U$4057 ( \4150 , \4149 , \3788 );
nor \U$4058 ( \4151 , \4148 , \4150 );
not \U$4059 ( \4152 , \4151 );
not \U$4060 ( \4153 , \1725 );
not \U$4061 ( \4154 , \4153 );
or \U$4062 ( \4155 , \4152 , \4154 );
or \U$4063 ( \4156 , \4153 , \4151 );
nand \U$4064 ( \4157 , \4155 , \4156 );
not \U$4065 ( \4158 , \4157 );
or \U$4066 ( \4159 , \4147 , \4158 );
buf \U$4067 ( \4160 , \1712 );
not \U$4068 ( \4161 , \4160 );
and \U$4069 ( \4162 , \188 , \3455 );
not \U$4070 ( \4163 , \188 );
and \U$4071 ( \4164 , \4163 , \3456 );
nor \U$4072 ( \4165 , \4162 , \4164 );
not \U$4073 ( \4166 , \4165 );
not \U$4074 ( \4167 , \1725 );
not \U$4075 ( \4168 , \4167 );
or \U$4076 ( \4169 , \4166 , \4168 );
not \U$4077 ( \4170 , \1725 );
not \U$4078 ( \4171 , \4165 );
not \U$4079 ( \4172 , \4171 );
or \U$4080 ( \4173 , \4170 , \4172 );
nand \U$4081 ( \4174 , \4169 , \4173 );
nand \U$4082 ( \4175 , \4161 , \4174 );
nand \U$4083 ( \4176 , \4159 , \4175 );
xnor \U$4084 ( \4177 , \172 , \1739 );
not \U$4085 ( \4178 , \4177 );
not \U$4086 ( \4179 , \4178 );
not \U$4087 ( \4180 , \4121 );
not \U$4088 ( \4181 , \4180 );
not \U$4089 ( \4182 , \4181 );
or \U$4090 ( \4183 , \4179 , \4182 );
buf \U$4091 ( \4184 , \4116 );
or \U$4092 ( \4185 , \4178 , \4184 );
nand \U$4093 ( \4186 , \4183 , \4185 );
not \U$4094 ( \4187 , \4186 );
not \U$4095 ( \4188 , RI8928a88_8);
not \U$4096 ( \4189 , \1571 );
or \U$4097 ( \4190 , \4188 , \4189 );
and \U$4098 ( \4191 , \1575 , RI892a108_56);
and \U$4099 ( \4192 , \1549 , \3146 );
not \U$4100 ( \4193 , \4089 );
not \U$4101 ( \4194 , \2228 );
nand \U$4102 ( \4195 , \4194 , \2226 );
not \U$4103 ( \4196 , \4195 );
not \U$4104 ( \4197 , \1164 );
not \U$4105 ( \4198 , \1170 );
or \U$4106 ( \4199 , \4197 , \4198 );
not \U$4107 ( \4200 , \1174 );
or \U$4108 ( \4201 , \4200 , \1103 );
nand \U$4109 ( \4202 , \4199 , \4201 );
not \U$4110 ( \4203 , \4202 );
or \U$4111 ( \4204 , \4196 , \4203 );
or \U$4112 ( \4205 , \4195 , \4202 );
nand \U$4113 ( \4206 , \4204 , \4205 );
not \U$4114 ( \4207 , \4206 );
or \U$4115 ( \4208 , \4193 , \4207 );
not \U$4116 ( \4209 , \2588 );
not \U$4117 ( \4210 , \2581 );
or \U$4118 ( \4211 , \4209 , \4210 );
or \U$4119 ( \4212 , \2581 , \2588 );
nand \U$4120 ( \4213 , \4211 , \4212 );
not \U$4121 ( \4214 , \4213 );
not \U$4122 ( \4215 , \2603 );
or \U$4123 ( \4216 , \4214 , \4215 );
buf \U$4124 ( \4217 , \2603 );
or \U$4125 ( \4218 , \4213 , \4217 );
nand \U$4126 ( \4219 , \4216 , \4218 );
nand \U$4127 ( \4220 , \4219 , \402 );
nand \U$4128 ( \4221 , \4208 , \4220 );
nor \U$4129 ( \4222 , \4192 , \4221 );
or \U$4130 ( \4223 , \690 , \1760 );
nand \U$4131 ( \4224 , \4223 , \419 );
nand \U$4132 ( \4225 , \4224 , RI8929988_40);
not \U$4133 ( \4226 , RI8928a88_8);
nand \U$4134 ( \4227 , \4226 , \1760 );
nand \U$4135 ( \4228 , \1547 , \4227 );
not \U$4136 ( \4229 , \1791 );
nand \U$4137 ( \4230 , \4229 , \1798 );
not \U$4138 ( \4231 , \4230 );
or \U$4139 ( \4232 , \1604 , \1790 );
not \U$4140 ( \4233 , \1527 );
nand \U$4141 ( \4234 , \4232 , \4233 );
not \U$4142 ( \4235 , \4234 );
or \U$4143 ( \4236 , \4231 , \4235 );
or \U$4144 ( \4237 , \4234 , \4230 );
nand \U$4145 ( \4238 , \4236 , \4237 );
and \U$4146 ( \4239 , \4238 , \1817 );
or \U$4147 ( \4240 , \3991 , \152 );
or \U$4148 ( \4241 , \424 , \1760 );
nand \U$4149 ( \4242 , \4240 , \4241 );
nor \U$4150 ( \4243 , \4239 , \4242 );
not \U$4151 ( \4244 , \1763 );
nand \U$4152 ( \4245 , \4244 , \1761 );
not \U$4153 ( \4246 , \4245 );
not \U$4154 ( \4247 , \1759 );
or \U$4155 ( \4248 , \4246 , \4247 );
or \U$4156 ( \4249 , \1759 , \4245 );
nand \U$4157 ( \4250 , \4248 , \4249 );
nand \U$4158 ( \4251 , \1779 , \4250 );
and \U$4159 ( \4252 , \4243 , \4251 );
nand \U$4160 ( \4253 , \4222 , \4225 , \4228 , \4252 );
nor \U$4161 ( \4254 , \4191 , \4253 );
nand \U$4162 ( \4255 , \4190 , \4254 );
not \U$4163 ( \4256 , \4255 );
and \U$4164 ( \4257 , \4256 , \1559 );
not \U$4165 ( \4258 , \4256 );
and \U$4166 ( \4259 , \4258 , \1715 );
nor \U$4167 ( \4260 , \4257 , \4259 );
not \U$4168 ( \4261 , \4256 );
not \U$4169 ( \4262 , \4115 );
or \U$4170 ( \4263 , \4261 , \4262 );
or \U$4171 ( \4264 , \4256 , \4115 );
nand \U$4172 ( \4265 , \4263 , \4264 );
nand \U$4173 ( \4266 , \4260 , \4265 );
not \U$4174 ( \4267 , \4266 );
not \U$4175 ( \4268 , \4267 );
or \U$4176 ( \4269 , \4187 , \4268 );
not \U$4177 ( \4270 , \4260 );
buf \U$4178 ( \4271 , \4270 );
or \U$4179 ( \4272 , \178 , \2810 );
nand \U$4180 ( \4273 , \178 , \2810 );
and \U$4181 ( \4274 , \4272 , \4273 );
not \U$4182 ( \4275 , \4274 );
not \U$4183 ( \4276 , \4115 );
buf \U$4184 ( \4277 , \4276 );
not \U$4185 ( \4278 , \4277 );
not \U$4186 ( \4279 , \4278 );
or \U$4187 ( \4280 , \4275 , \4279 );
or \U$4188 ( \4281 , \4274 , \4184 );
nand \U$4189 ( \4282 , \4280 , \4281 );
nand \U$4190 ( \4283 , \4271 , \4282 );
nand \U$4191 ( \4284 , \4269 , \4283 );
xor \U$4192 ( \4285 , \4176 , \4284 );
not \U$4193 ( \4286 , \4285 );
or \U$4194 ( \4287 , \4145 , \4286 );
nand \U$4195 ( \4288 , \4176 , \4284 );
nand \U$4196 ( \4289 , \4287 , \4288 );
not \U$4197 ( \4290 , \4289 );
or \U$4198 ( \4291 , \3981 , \4290 );
not \U$4199 ( \4292 , \3979 );
nand \U$4200 ( \4293 , \4292 , \3845 );
nand \U$4201 ( \4294 , \4291 , \4293 );
not \U$4202 ( \4295 , \4294 );
nand \U$4203 ( \4296 , \3838 , \4295 );
not \U$4204 ( \4297 , \4296 );
not \U$4205 ( \4298 , \3814 );
not \U$4206 ( \4299 , \3843 );
not \U$4207 ( \4300 , \3755 );
or \U$4208 ( \4301 , \4299 , \4300 );
buf \U$4209 ( \4302 , \3754 );
not \U$4210 ( \4303 , \4302 );
not \U$4211 ( \4304 , \4303 );
or \U$4212 ( \4305 , \4304 , \3843 );
nand \U$4213 ( \4306 , \4301 , \4305 );
not \U$4214 ( \4307 , \4306 );
or \U$4215 ( \4308 , \4298 , \4307 );
not \U$4216 ( \4309 , \3832 );
not \U$4217 ( \4310 , \4309 );
and \U$4218 ( \4311 , \146 , \1552 );
not \U$4219 ( \4312 , \146 );
not \U$4220 ( \4313 , \1552 );
and \U$4221 ( \4314 , \4312 , \4313 );
or \U$4222 ( \4315 , \4311 , \4314 );
not \U$4223 ( \4316 , \4315 );
not \U$4224 ( \4317 , \3755 );
or \U$4225 ( \4318 , \4316 , \4317 );
or \U$4226 ( \4319 , \4304 , \4315 );
nand \U$4227 ( \4320 , \4318 , \4319 );
nand \U$4228 ( \4321 , \4310 , \4320 );
nand \U$4229 ( \4322 , \4308 , \4321 );
and \U$4230 ( \4323 , \138 , \1648 );
not \U$4231 ( \4324 , \138 );
not \U$4232 ( \4325 , \1648 );
and \U$4233 ( \4326 , \4324 , \4325 );
or \U$4234 ( \4327 , \4323 , \4326 );
not \U$4235 ( \4328 , \4327 );
nand \U$4236 ( \4329 , \4304 , \4328 );
not \U$4237 ( \4330 , \4329 );
nor \U$4238 ( \4331 , \4322 , \4330 );
not \U$4239 ( \4332 , \3107 );
buf \U$4240 ( \4333 , \4332 );
not \U$4241 ( \4334 , \4333 );
and \U$4242 ( \4335 , \3822 , \4334 );
not \U$4243 ( \4336 , \3822 );
and \U$4244 ( \4337 , \4336 , \4333 );
nor \U$4245 ( \4338 , \4335 , \4337 );
not \U$4246 ( \4339 , \4338 );
not \U$4247 ( \4340 , \2800 );
and \U$4248 ( \4341 , \4339 , \4340 );
not \U$4249 ( \4342 , \3141 );
and \U$4250 ( \4343 , \3151 , \4333 );
not \U$4251 ( \4344 , \3151 );
and \U$4252 ( \4345 , \4344 , \4334 );
nor \U$4253 ( \4346 , \4343 , \4345 );
and \U$4254 ( \4347 , \4342 , \4346 );
nor \U$4255 ( \4348 , \4341 , \4347 );
buf \U$4256 ( \4349 , \4348 );
or \U$4257 ( \4350 , \4331 , \4349 );
nand \U$4258 ( \4351 , \4322 , \4330 );
nand \U$4259 ( \4352 , \4350 , \4351 );
not \U$4260 ( \4353 , \4352 );
not \U$4261 ( \4354 , \4266 );
buf \U$4262 ( \4355 , \4354 );
not \U$4263 ( \4356 , \4355 );
not \U$4264 ( \4357 , \4282 );
or \U$4265 ( \4358 , \4356 , \4357 );
not \U$4266 ( \4359 , \4151 );
not \U$4267 ( \4360 , \4277 );
not \U$4268 ( \4361 , \4360 );
or \U$4269 ( \4362 , \4359 , \4361 );
or \U$4270 ( \4363 , \4360 , \4151 );
nand \U$4271 ( \4364 , \4362 , \4363 );
nand \U$4272 ( \4365 , \4271 , \4364 );
nand \U$4273 ( \4366 , \4358 , \4365 );
not \U$4274 ( \4367 , \4174 );
not \U$4275 ( \4368 , \1719 );
or \U$4276 ( \4369 , \4367 , \4368 );
nand \U$4277 ( \4370 , \1724 , \1566 );
nand \U$4278 ( \4371 , \4369 , \4370 );
xor \U$4279 ( \4372 , \4366 , \4371 );
buf \U$4280 ( \4373 , \3958 );
not \U$4281 ( \4374 , \4373 );
not \U$4282 ( \4375 , \4374 );
buf \U$4283 ( \4376 , \3966 );
not \U$4284 ( \4377 , \4376 );
or \U$4285 ( \4378 , \4375 , \4377 );
nand \U$4286 ( \4379 , \4378 , \3977 );
xor \U$4287 ( \4380 , \4372 , \4379 );
not \U$4288 ( \4381 , \4380 );
or \U$4289 ( \4382 , \4353 , \4381 );
not \U$4290 ( \4383 , \2800 );
not \U$4291 ( \4384 , \3131 );
and \U$4292 ( \4385 , \4383 , \4384 );
not \U$4293 ( \4386 , \3141 );
not \U$4294 ( \4387 , \4338 );
and \U$4295 ( \4388 , \4386 , \4387 );
nor \U$4296 ( \4389 , \4385 , \4388 );
not \U$4297 ( \4390 , \4142 );
not \U$4298 ( \4391 , \4130 );
not \U$4299 ( \4392 , \4391 );
or \U$4300 ( \4393 , \4390 , \4392 );
not \U$4301 ( \4394 , \4178 );
not \U$4302 ( \4395 , \3983 );
not \U$4303 ( \4396 , \4395 );
not \U$4304 ( \4397 , \4396 );
or \U$4305 ( \4398 , \4394 , \4397 );
or \U$4306 ( \4399 , \4137 , \4178 );
nand \U$4307 ( \4400 , \4398 , \4399 );
nand \U$4308 ( \4401 , \4135 , \4400 );
nand \U$4309 ( \4402 , \4393 , \4401 );
not \U$4310 ( \4403 , \4402 );
xor \U$4311 ( \4404 , \4389 , \4403 );
not \U$4312 ( \4405 , \3833 );
not \U$4313 ( \4406 , \4405 );
not \U$4314 ( \4407 , \3759 );
not \U$4315 ( \4408 , \4407 );
and \U$4316 ( \4409 , \4406 , \4408 );
and \U$4317 ( \4410 , \4320 , \3815 );
nor \U$4318 ( \4411 , \4409 , \4410 );
xor \U$4319 ( \4412 , \4404 , \4411 );
nand \U$4320 ( \4413 , \4382 , \4412 );
or \U$4321 ( \4414 , \4352 , \4380 );
nand \U$4322 ( \4415 , \4413 , \4414 );
not \U$4323 ( \4416 , \4415 );
not \U$4324 ( \4417 , \4416 );
or \U$4325 ( \4418 , \4297 , \4417 );
nand \U$4326 ( \4419 , \4294 , \3837 );
nand \U$4327 ( \4420 , \4418 , \4419 );
xor \U$4328 ( \4421 , \4389 , \4403 );
and \U$4329 ( \4422 , \4421 , \4411 );
and \U$4330 ( \4423 , \4389 , \4403 );
or \U$4331 ( \4424 , \4422 , \4423 );
not \U$4332 ( \4425 , \4424 );
not \U$4333 ( \4426 , \4425 );
xor \U$4334 ( \4427 , \4366 , \4371 );
and \U$4335 ( \4428 , \4427 , \4379 );
and \U$4336 ( \4429 , \4366 , \4371 );
or \U$4337 ( \4430 , \4428 , \4429 );
not \U$4338 ( \4431 , \4430 );
not \U$4339 ( \4432 , \4364 );
not \U$4340 ( \4433 , \4355 );
or \U$4341 ( \4434 , \4432 , \4433 );
not \U$4342 ( \4435 , \4172 );
not \U$4343 ( \4436 , \4360 );
or \U$4344 ( \4437 , \4435 , \4436 );
not \U$4345 ( \4438 , \4184 );
not \U$4346 ( \4439 , \4438 );
or \U$4347 ( \4440 , \4439 , \4172 );
nand \U$4348 ( \4441 , \4437 , \4440 );
nand \U$4349 ( \4442 , \4271 , \4441 );
nand \U$4350 ( \4443 , \4434 , \4442 );
not \U$4351 ( \4444 , \4315 );
nand \U$4352 ( \4445 , \3823 , \4444 );
nor \U$4353 ( \4446 , \4443 , \4445 );
not \U$4354 ( \4447 , \4446 );
nand \U$4355 ( \4448 , \4443 , \4445 );
nand \U$4356 ( \4449 , \4447 , \4448 );
not \U$4357 ( \4450 , \4449 );
not \U$4358 ( \4451 , \4400 );
not \U$4359 ( \4452 , \4391 );
or \U$4360 ( \4453 , \4451 , \4452 );
not \U$4361 ( \4454 , \4395 );
not \U$4362 ( \4455 , \4274 );
and \U$4363 ( \4456 , \4454 , \4455 );
not \U$4364 ( \4457 , \4137 );
and \U$4365 ( \4458 , \4457 , \4274 );
nor \U$4366 ( \4459 , \4456 , \4458 );
nand \U$4367 ( \4460 , \4135 , \4459 );
nand \U$4368 ( \4461 , \4453 , \4460 );
not \U$4369 ( \4462 , \4461 );
and \U$4370 ( \4463 , \4450 , \4462 );
and \U$4371 ( \4464 , \4449 , \4461 );
nor \U$4372 ( \4465 , \4463 , \4464 );
not \U$4373 ( \4466 , \4465 );
or \U$4374 ( \4467 , \4431 , \4466 );
or \U$4375 ( \4468 , \4465 , \4430 );
nand \U$4376 ( \4469 , \4467 , \4468 );
not \U$4377 ( \4470 , \4469 );
or \U$4378 ( \4471 , \4426 , \4470 );
not \U$4379 ( \4472 , \4465 );
nand \U$4380 ( \4473 , \4472 , \4430 );
nand \U$4381 ( \4474 , \4471 , \4473 );
not \U$4382 ( \4475 , \4474 );
xor \U$4383 ( \4476 , \4420 , \4475 );
not \U$4384 ( \4477 , \4459 );
buf \U$4385 ( \4478 , \4391 );
not \U$4386 ( \4479 , \4478 );
or \U$4387 ( \4480 , \4477 , \4479 );
not \U$4388 ( \4481 , \4457 );
buf \U$4389 ( \4482 , \4151 );
not \U$4390 ( \4483 , \4482 );
and \U$4391 ( \4484 , \4481 , \4483 );
and \U$4392 ( \4485 , \4457 , \4482 );
nor \U$4393 ( \4486 , \4484 , \4485 );
nand \U$4394 ( \4487 , \4135 , \4486 );
nand \U$4395 ( \4488 , \4480 , \4487 );
not \U$4396 ( \4489 , \4448 );
not \U$4397 ( \4490 , \4461 );
or \U$4398 ( \4491 , \4489 , \4490 );
not \U$4399 ( \4492 , \4446 );
nand \U$4400 ( \4493 , \4491 , \4492 );
not \U$4401 ( \4494 , \4493 );
xor \U$4402 ( \4495 , \4488 , \4494 );
not \U$4403 ( \4496 , \3824 );
not \U$4404 ( \4497 , \3815 );
or \U$4405 ( \4498 , \4496 , \4497 );
not \U$4406 ( \4499 , \3127 );
not \U$4407 ( \4500 , \3823 );
or \U$4408 ( \4501 , \4499 , \4500 );
or \U$4409 ( \4502 , \3823 , \3127 );
nand \U$4410 ( \4503 , \4501 , \4502 );
nand \U$4411 ( \4504 , \4503 , \3833 );
nand \U$4412 ( \4505 , \4498 , \4504 );
not \U$4413 ( \4506 , \3151 );
nand \U$4414 ( \4507 , \3823 , \4506 );
xnor \U$4415 ( \4508 , \4505 , \4507 );
xor \U$4416 ( \4509 , \4495 , \4508 );
xor \U$4417 ( \4510 , \1729 , \3144 );
and \U$4418 ( \4511 , \4510 , \3835 );
and \U$4419 ( \4512 , \1729 , \3144 );
or \U$4420 ( \4513 , \4511 , \4512 );
xor \U$4421 ( \4514 , \4443 , \4513 );
not \U$4422 ( \4515 , \4355 );
not \U$4423 ( \4516 , \4441 );
or \U$4424 ( \4517 , \4515 , \4516 );
not \U$4425 ( \4518 , \193 );
not \U$4426 ( \4519 , \4277 );
not \U$4427 ( \4520 , \4519 );
or \U$4428 ( \4521 , \4518 , \4520 );
or \U$4429 ( \4522 , \4519 , \193 );
nand \U$4430 ( \4523 , \4521 , \4522 );
nand \U$4431 ( \4524 , \4523 , \4271 );
nand \U$4432 ( \4525 , \4517 , \4524 );
not \U$4433 ( \4526 , \1717 );
not \U$4434 ( \4527 , \4526 );
not \U$4435 ( \4528 , \1723 );
or \U$4436 ( \4529 , \4527 , \4528 );
nand \U$4437 ( \4530 , \4529 , \1727 );
nor \U$4438 ( \4531 , \4525 , \4530 );
not \U$4439 ( \4532 , \4531 );
nand \U$4440 ( \4533 , \4525 , \4530 );
nand \U$4441 ( \4534 , \4532 , \4533 );
xor \U$4442 ( \4535 , \3110 , \4178 );
not \U$4443 ( \4536 , \4535 );
not \U$4444 ( \4537 , \2800 );
and \U$4445 ( \4538 , \4536 , \4537 );
not \U$4446 ( \4539 , \4386 );
not \U$4447 ( \4540 , \4539 );
and \U$4448 ( \4541 , \4540 , \3117 );
nor \U$4449 ( \4542 , \4538 , \4541 );
xor \U$4450 ( \4543 , \4534 , \4542 );
xor \U$4451 ( \4544 , \4514 , \4543 );
xnor \U$4452 ( \4545 , \4509 , \4544 );
buf \U$4453 ( \4546 , \4545 );
xnor \U$4454 ( \4547 , \4476 , \4546 );
not \U$4455 ( \4548 , \4416 );
not \U$4456 ( \4549 , \3836 );
not \U$4457 ( \4550 , \4295 );
or \U$4458 ( \4551 , \4549 , \4550 );
or \U$4459 ( \4552 , \4295 , \3836 );
nand \U$4460 ( \4553 , \4551 , \4552 );
not \U$4461 ( \4554 , \4553 );
not \U$4462 ( \4555 , \4554 );
or \U$4463 ( \4556 , \4548 , \4555 );
nand \U$4464 ( \4557 , \4553 , \4415 );
nand \U$4465 ( \4558 , \4556 , \4557 );
buf \U$4466 ( \4559 , \4558 );
xor \U$4467 ( \4560 , \4469 , \4424 );
not \U$4468 ( \4561 , \4560 );
or \U$4469 ( \4562 , \4559 , \4561 );
not \U$4470 ( \4563 , RI8928dd0_15);
not \U$4471 ( \4564 , \2270 );
or \U$4472 ( \4565 , \4563 , \4564 );
nand \U$4473 ( \4566 , \1575 , RI892a450_63);
not \U$4474 ( \4567 , \988 );
not \U$4475 ( \4568 , \990 );
and \U$4476 ( \4569 , \4567 , \4568 );
not \U$4477 ( \4570 , \991 );
nor \U$4478 ( \4571 , \4569 , \4570 );
and \U$4479 ( \4572 , \1650 , \4571 );
or \U$4480 ( \4573 , \1422 , \1424 );
nand \U$4481 ( \4574 , \4573 , \1425 );
not \U$4482 ( \4575 , \4574 );
not \U$4483 ( \4576 , \4575 );
not \U$4484 ( \4577 , \402 );
or \U$4485 ( \4578 , \4576 , \4577 );
not \U$4486 ( \4579 , \1459 );
nor \U$4487 ( \4580 , \1463 , \1458 );
not \U$4488 ( \4581 , \4580 );
or \U$4489 ( \4582 , \4579 , \4581 );
or \U$4490 ( \4583 , \4580 , \1459 );
nand \U$4491 ( \4584 , \4582 , \4583 );
not \U$4492 ( \4585 , \4584 );
not \U$4493 ( \4586 , \1600 );
or \U$4494 ( \4587 , \4585 , \4586 );
not \U$4495 ( \4588 , \1505 );
not \U$4496 ( \4589 , \1507 );
nor \U$4497 ( \4590 , \4589 , \1504 );
not \U$4498 ( \4591 , \4590 );
or \U$4499 ( \4592 , \4588 , \4591 );
or \U$4500 ( \4593 , \4590 , \1505 );
nand \U$4501 ( \4594 , \4592 , \4593 );
and \U$4502 ( \4595 , \410 , \4594 );
not \U$4503 ( \4596 , RI892a450_63);
not \U$4504 ( \4597 , \413 );
or \U$4505 ( \4598 , \4596 , \4597 );
and \U$4506 ( \4599 , \418 , RI8929cd0_47);
and \U$4507 ( \4600 , \423 , RI8929550_31);
nor \U$4508 ( \4601 , \4599 , \4600 );
nand \U$4509 ( \4602 , \4598 , \4601 );
nor \U$4510 ( \4603 , \4595 , \4602 );
nand \U$4511 ( \4604 , \4587 , \4603 );
not \U$4512 ( \4605 , \4604 );
nand \U$4513 ( \4606 , \4578 , \4605 );
nor \U$4514 ( \4607 , \4572 , \4606 );
and \U$4515 ( \4608 , RI8929cd0_47, RI8929550_31);
nand \U$4516 ( \4609 , \4076 , \4608 );
xor \U$4517 ( \4610 , RI8929cd0_47, RI892a450_63);
nand \U$4518 ( \4611 , \1549 , \4610 );
nand \U$4519 ( \4612 , \4607 , \4609 , \4611 );
not \U$4520 ( \4613 , RI8928dd0_15);
not \U$4521 ( \4614 , RI8929550_31);
and \U$4522 ( \4615 , \4613 , \4614 );
nor \U$4523 ( \4616 , \4615 , \776 );
nor \U$4524 ( \4617 , \4612 , \4616 );
nand \U$4525 ( \4618 , \4566 , \4617 );
not \U$4526 ( \4619 , \4618 );
nand \U$4527 ( \4620 , \4565 , \4619 );
buf \U$4528 ( \4621 , \4620 );
not \U$4529 ( \4622 , \4621 );
not \U$4530 ( \4623 , RI8928d58_14);
not \U$4531 ( \4624 , \2270 );
or \U$4532 ( \4625 , \4623 , \4624 );
and \U$4533 ( \4626 , RI892a3d8_62, \1575 );
not \U$4534 ( \4627 , RI8928d58_14);
not \U$4535 ( \4628 , RI89294d8_30);
nand \U$4536 ( \4629 , \4627 , \4628 );
nand \U$4537 ( \4630 , \1547 , \4629 );
and \U$4538 ( \4631 , RI892a3d8_62, RI8929c58_46);
not \U$4539 ( \4632 , RI892a3d8_62);
not \U$4540 ( \4633 , RI8929c58_46);
and \U$4541 ( \4634 , \4632 , \4633 );
nor \U$4542 ( \4635 , \4631 , \4634 );
nand \U$4543 ( \4636 , \1549 , \4635 );
nor \U$4544 ( \4637 , \4628 , \4633 );
nand \U$4545 ( \4638 , \1644 , \4637 );
not \U$4546 ( \4639 , \993 );
or \U$4547 ( \4640 , \4639 , \983 , \4570 );
nand \U$4548 ( \4641 , \4570 , \983 );
nand \U$4549 ( \4642 , \4640 , \4641 );
not \U$4550 ( \4643 , \4642 );
not \U$4551 ( \4644 , \3916 );
or \U$4552 ( \4645 , \4643 , \4644 );
not \U$4553 ( \4646 , \1425 );
not \U$4554 ( \4647 , \1427 );
nor \U$4555 ( \4648 , \4647 , \1416 );
not \U$4556 ( \4649 , \4648 );
or \U$4557 ( \4650 , \4646 , \4649 );
or \U$4558 ( \4651 , \4648 , \1425 );
nand \U$4559 ( \4652 , \4650 , \4651 );
not \U$4560 ( \4653 , \4652 );
not \U$4561 ( \4654 , \402 );
or \U$4562 ( \4655 , \4653 , \4654 );
not \U$4563 ( \4656 , \405 );
nor \U$4564 ( \4657 , \1460 , \1463 );
not \U$4565 ( \4658 , \4657 );
not \U$4566 ( \4659 , \1456 );
nor \U$4567 ( \4660 , \4659 , \1465 );
not \U$4568 ( \4661 , \4660 );
and \U$4569 ( \4662 , \4658 , \4661 );
and \U$4570 ( \4663 , \4657 , \4660 );
nor \U$4571 ( \4664 , \4662 , \4663 );
not \U$4572 ( \4665 , \4664 );
and \U$4573 ( \4666 , \4656 , \4665 );
not \U$4574 ( \4667 , \1511 );
nand \U$4575 ( \4668 , \4667 , \1509 );
not \U$4576 ( \4669 , \4668 );
not \U$4577 ( \4670 , \1508 );
or \U$4578 ( \4671 , \4669 , \4670 );
or \U$4579 ( \4672 , \4668 , \1508 );
nand \U$4580 ( \4673 , \4671 , \4672 );
not \U$4581 ( \4674 , \4673 );
not \U$4582 ( \4675 , \1817 );
or \U$4583 ( \4676 , \4674 , \4675 );
and \U$4584 ( \4677 , \1730 , RI892a3d8_62);
or \U$4585 ( \4678 , \419 , \4633 );
or \U$4586 ( \4679 , \424 , \4628 );
nand \U$4587 ( \4680 , \4678 , \4679 );
nor \U$4588 ( \4681 , \4677 , \4680 );
nand \U$4589 ( \4682 , \4676 , \4681 );
nor \U$4590 ( \4683 , \4666 , \4682 );
nand \U$4591 ( \4684 , \4655 , \4683 );
not \U$4592 ( \4685 , \4684 );
nand \U$4593 ( \4686 , \4645 , \4685 );
not \U$4594 ( \4687 , \4686 );
nand \U$4595 ( \4688 , \4630 , \4636 , \4638 , \4687 );
nor \U$4596 ( \4689 , \4626 , \4688 );
nand \U$4597 ( \4690 , \4625 , \4689 );
not \U$4598 ( \4691 , \4690 );
nand \U$4599 ( \4692 , \4622 , \4691 );
nand \U$4600 ( \4693 , \4621 , \4690 );
and \U$4601 ( \4694 , \4692 , \4693 );
not \U$4602 ( \4695 , \4694 );
not \U$4603 ( \4696 , \4695 );
not \U$4604 ( \4697 , \4696 );
buf \U$4605 ( \4698 , \3957 );
not \U$4606 ( \4699 , \4698 );
not \U$4607 ( \4700 , \4699 );
not \U$4608 ( \4701 , \4700 );
buf \U$4609 ( \4702 , \4701 );
not \U$4610 ( \4703 , \4702 );
not \U$4611 ( \4704 , \4703 );
or \U$4612 ( \4705 , \4697 , \4704 );
or \U$4613 ( \4706 , \4693 , \4698 );
not \U$4614 ( \4707 , \4690 );
not \U$4615 ( \4708 , \4621 );
nand \U$4616 ( \4709 , \4707 , \4708 , \4698 );
nand \U$4617 ( \4710 , \4706 , \4709 );
buf \U$4618 ( \4711 , \4710 );
not \U$4619 ( \4712 , \4698 );
not \U$4620 ( \4713 , \4712 );
not \U$4621 ( \4714 , \4713 );
not \U$4622 ( \4715 , \192 );
and \U$4623 ( \4716 , \4714 , \4715 );
and \U$4624 ( \4717 , \4698 , \192 );
nor \U$4625 ( \4718 , \4716 , \4717 );
nand \U$4626 ( \4719 , \4711 , \4718 );
nand \U$4627 ( \4720 , \4705 , \4719 );
not \U$4628 ( \4721 , \4720 );
not \U$4629 ( \4722 , \3814 );
and \U$4630 ( \4723 , \4327 , \3755 );
not \U$4631 ( \4724 , \4327 );
and \U$4632 ( \4725 , \4724 , \4303 );
or \U$4633 ( \4726 , \4723 , \4725 );
not \U$4634 ( \4727 , \4726 );
or \U$4635 ( \4728 , \4722 , \4727 );
nand \U$4636 ( \4729 , \4306 , \4310 );
nand \U$4637 ( \4730 , \4728 , \4729 );
not \U$4638 ( \4731 , \4730 );
or \U$4639 ( \4732 , \4721 , \4731 );
not \U$4640 ( \4733 , \4444 );
not \U$4641 ( \4734 , \4333 );
or \U$4642 ( \4735 , \4733 , \4734 );
or \U$4643 ( \4736 , \3114 , \4444 );
nand \U$4644 ( \4737 , \4735 , \4736 );
not \U$4645 ( \4738 , \4737 );
not \U$4646 ( \4739 , \3140 );
or \U$4647 ( \4740 , \4738 , \4739 );
nand \U$4648 ( \4741 , \4346 , \2799 );
nand \U$4649 ( \4742 , \4740 , \4741 );
not \U$4650 ( \4743 , \4742 );
nand \U$4651 ( \4744 , \4732 , \4743 );
not \U$4652 ( \4745 , \4730 );
not \U$4653 ( \4746 , \4720 );
nand \U$4654 ( \4747 , \4745 , \4746 );
nand \U$4655 ( \4748 , \4744 , \4747 );
not \U$4656 ( \4749 , \4144 );
xor \U$4657 ( \4750 , \4285 , \4749 );
xor \U$4658 ( \4751 , \4748 , \4750 );
xor \U$4659 ( \4752 , \4329 , \4348 );
xnor \U$4660 ( \4753 , \4752 , \4322 );
and \U$4661 ( \4754 , \4751 , \4753 );
and \U$4662 ( \4755 , \4748 , \4750 );
or \U$4663 ( \4756 , \4754 , \4755 );
not \U$4664 ( \4757 , \4756 );
not \U$4665 ( \4758 , \4757 );
not \U$4666 ( \4759 , \3973 );
not \U$4667 ( \4760 , \3958 );
or \U$4668 ( \4761 , \4759 , \4760 );
not \U$4669 ( \4762 , \3958 );
not \U$4670 ( \4763 , \4762 );
not \U$4671 ( \4764 , \1710 );
not \U$4672 ( \4765 , \4165 );
or \U$4673 ( \4766 , \4764 , \4765 );
or \U$4674 ( \4767 , \3977 , \4165 );
nand \U$4675 ( \4768 , \4766 , \4767 );
nand \U$4676 ( \4769 , \3965 , \4768 );
or \U$4677 ( \4770 , \4763 , \4769 );
nand \U$4678 ( \4771 , \4761 , \4770 );
not \U$4679 ( \4772 , \4266 );
not \U$4680 ( \4773 , \4772 );
not \U$4681 ( \4774 , \2803 );
not \U$4682 ( \4775 , \4120 );
not \U$4683 ( \4776 , \4775 );
or \U$4684 ( \4777 , \4774 , \4776 );
or \U$4685 ( \4778 , \4116 , \2803 );
nand \U$4686 ( \4779 , \4777 , \4778 );
not \U$4687 ( \4780 , \4779 );
or \U$4688 ( \4781 , \4773 , \4780 );
nand \U$4689 ( \4782 , \4186 , \4271 );
nand \U$4690 ( \4783 , \4781 , \4782 );
xor \U$4691 ( \4784 , \4771 , \4783 );
not \U$4692 ( \4785 , \4690 );
not \U$4693 ( \4786 , \4695 );
or \U$4694 ( \4787 , \4785 , \4786 );
nand \U$4695 ( \4788 , \4787 , \4703 );
and \U$4696 ( \4789 , \4784 , \4788 );
and \U$4697 ( \4790 , \4771 , \4783 );
or \U$4698 ( \4791 , \4789 , \4790 );
xor \U$4699 ( \4792 , \3979 , \4791 );
xnor \U$4700 ( \4793 , \134 , \3860 );
nor \U$4701 ( \4794 , \4303 , \4793 );
not \U$4702 ( \4795 , \4274 );
not \U$4703 ( \4796 , \4153 );
or \U$4704 ( \4797 , \4795 , \4796 );
not \U$4705 ( \4798 , \1561 );
or \U$4706 ( \4799 , \4798 , \4274 );
nand \U$4707 ( \4800 , \4797 , \4799 );
not \U$4708 ( \4801 , \4800 );
not \U$4709 ( \4802 , \1719 );
or \U$4710 ( \4803 , \4801 , \4802 );
nand \U$4711 ( \4804 , \4161 , \4157 );
nand \U$4712 ( \4805 , \4803 , \4804 );
xor \U$4713 ( \4806 , \4794 , \4805 );
and \U$4714 ( \4807 , \3821 , \4137 );
not \U$4715 ( \4808 , \3821 );
and \U$4716 ( \4809 , \4808 , \3987 );
nor \U$4717 ( \4810 , \4807 , \4809 );
not \U$4718 ( \4811 , \4810 );
not \U$4719 ( \4812 , \4131 );
or \U$4720 ( \4813 , \4811 , \4812 );
buf \U$4721 ( \4814 , \4123 );
not \U$4722 ( \4815 , \4814 );
nand \U$4723 ( \4816 , \4815 , \3989 );
nand \U$4724 ( \4817 , \4813 , \4816 );
and \U$4725 ( \4818 , \4806 , \4817 );
and \U$4726 ( \4819 , \4794 , \4805 );
or \U$4727 ( \4820 , \4818 , \4819 );
and \U$4728 ( \4821 , \4792 , \4820 );
and \U$4729 ( \4822 , \3979 , \4791 );
or \U$4730 ( \4823 , \4821 , \4822 );
not \U$4731 ( \4824 , \4823 );
not \U$4732 ( \4825 , \4289 );
not \U$4733 ( \4826 , \4825 );
not \U$4734 ( \4827 , \3845 );
not \U$4735 ( \4828 , \4292 );
or \U$4736 ( \4829 , \4827 , \4828 );
or \U$4737 ( \4830 , \4292 , \3845 );
nand \U$4738 ( \4831 , \4829 , \4830 );
not \U$4739 ( \4832 , \4831 );
and \U$4740 ( \4833 , \4826 , \4832 );
and \U$4741 ( \4834 , \4825 , \4831 );
nor \U$4742 ( \4835 , \4833 , \4834 );
not \U$4743 ( \4836 , \4835 );
nand \U$4744 ( \4837 , \4824 , \4836 );
not \U$4745 ( \4838 , \4837 );
or \U$4746 ( \4839 , \4758 , \4838 );
nand \U$4747 ( \4840 , \4835 , \4823 );
nand \U$4748 ( \4841 , \4839 , \4840 );
nand \U$4749 ( \4842 , \4562 , \4841 );
nand \U$4750 ( \4843 , \4559 , \4561 );
nand \U$4751 ( \4844 , \4842 , \4843 );
or \U$4752 ( \4845 , \4547 , \4844 );
not \U$4753 ( \4846 , \4420 );
not \U$4754 ( \4847 , \4475 );
not \U$4755 ( \4848 , \4545 );
or \U$4756 ( \4849 , \4847 , \4848 );
or \U$4757 ( \4850 , \4545 , \4475 );
nand \U$4758 ( \4851 , \4849 , \4850 );
not \U$4759 ( \4852 , \4851 );
or \U$4760 ( \4853 , \4846 , \4852 );
nand \U$4761 ( \4854 , \4546 , \4474 );
nand \U$4762 ( \4855 , \4853 , \4854 );
not \U$4763 ( \4856 , \4855 );
not \U$4764 ( \4857 , \4535 );
not \U$4765 ( \4858 , \4857 );
not \U$4766 ( \4859 , \4540 );
or \U$4767 ( \4860 , \4858 , \4859 );
not \U$4768 ( \4861 , \4274 );
and \U$4769 ( \4862 , \4861 , \3110 );
not \U$4770 ( \4863 , \4861 );
not \U$4771 ( \4864 , \3110 );
and \U$4772 ( \4865 , \4863 , \4864 );
nor \U$4773 ( \4866 , \4862 , \4865 );
nand \U$4774 ( \4867 , \2801 , \4866 );
nand \U$4775 ( \4868 , \4860 , \4867 );
not \U$4776 ( \4869 , \4355 );
not \U$4777 ( \4870 , \4523 );
or \U$4778 ( \4871 , \4869 , \4870 );
nand \U$4779 ( \4872 , \4271 , \4519 );
nand \U$4780 ( \4873 , \4871 , \4872 );
xnor \U$4781 ( \4874 , \4868 , \4873 );
not \U$4782 ( \4875 , \4488 );
not \U$4783 ( \4876 , \4508 );
or \U$4784 ( \4877 , \4875 , \4876 );
not \U$4785 ( \4878 , \4507 );
nand \U$4786 ( \4879 , \4878 , \4505 );
nand \U$4787 ( \4880 , \4877 , \4879 );
xor \U$4788 ( \4881 , \4874 , \4880 );
xor \U$4789 ( \4882 , \4507 , \4488 );
xor \U$4790 ( \4883 , \4882 , \4505 );
nand \U$4791 ( \4884 , \4883 , \4494 );
not \U$4792 ( \4885 , \4884 );
not \U$4793 ( \4886 , \4544 );
or \U$4794 ( \4887 , \4885 , \4886 );
not \U$4795 ( \4888 , \4883 );
nand \U$4796 ( \4889 , \4888 , \4493 );
nand \U$4797 ( \4890 , \4887 , \4889 );
xor \U$4798 ( \4891 , \4881 , \4890 );
not \U$4799 ( \4892 , \4891 );
nand \U$4800 ( \4893 , \3823 , \3821 );
not \U$4801 ( \4894 , \4486 );
not \U$4802 ( \4895 , \4478 );
or \U$4803 ( \4896 , \4894 , \4895 );
and \U$4804 ( \4897 , \4172 , \4137 );
not \U$4805 ( \4898 , \4172 );
and \U$4806 ( \4899 , \4898 , \4457 );
or \U$4807 ( \4900 , \4897 , \4899 );
nand \U$4808 ( \4901 , \4135 , \4900 );
nand \U$4809 ( \4902 , \4896 , \4901 );
xor \U$4810 ( \4903 , \4893 , \4902 );
not \U$4811 ( \4904 , \4503 );
buf \U$4812 ( \4905 , \3815 );
not \U$4813 ( \4906 , \4905 );
or \U$4814 ( \4907 , \4904 , \4906 );
not \U$4815 ( \4908 , \2803 );
not \U$4816 ( \4909 , \3823 );
or \U$4817 ( \4910 , \4908 , \4909 );
or \U$4818 ( \4911 , \3823 , \2803 );
nand \U$4819 ( \4912 , \4910 , \4911 );
nand \U$4820 ( \4913 , \4912 , \3833 );
nand \U$4821 ( \4914 , \4907 , \4913 );
xnor \U$4822 ( \4915 , \4903 , \4914 );
and \U$4823 ( \4916 , \4533 , \4542 );
nor \U$4824 ( \4917 , \4916 , \4531 );
nor \U$4825 ( \4918 , \4915 , \4917 );
not \U$4826 ( \4919 , \4918 );
nand \U$4827 ( \4920 , \4915 , \4917 );
nand \U$4828 ( \4921 , \4919 , \4920 );
not \U$4829 ( \4922 , \4921 );
xor \U$4830 ( \4923 , \4443 , \4513 );
and \U$4831 ( \4924 , \4923 , \4543 );
and \U$4832 ( \4925 , \4443 , \4513 );
or \U$4833 ( \4926 , \4924 , \4925 );
not \U$4834 ( \4927 , \4926 );
and \U$4835 ( \4928 , \4922 , \4927 );
and \U$4836 ( \4929 , \4921 , \4926 );
nor \U$4837 ( \4930 , \4928 , \4929 );
not \U$4838 ( \4931 , \4930 );
and \U$4839 ( \4932 , \4892 , \4931 );
and \U$4840 ( \4933 , \4930 , \4891 );
nor \U$4841 ( \4934 , \4932 , \4933 );
nand \U$4842 ( \4935 , \4856 , \4934 );
not \U$4843 ( \4936 , \4874 );
not \U$4844 ( \4937 , \4880 );
or \U$4845 ( \4938 , \4936 , \4937 );
not \U$4846 ( \4939 , \4873 );
not \U$4847 ( \4940 , \4857 );
not \U$4848 ( \4941 , \4540 );
or \U$4849 ( \4942 , \4940 , \4941 );
nand \U$4850 ( \4943 , \4942 , \4867 );
nand \U$4851 ( \4944 , \4939 , \4943 );
nand \U$4852 ( \4945 , \4938 , \4944 );
not \U$4853 ( \4946 , \4918 );
nand \U$4854 ( \4947 , \4946 , \4926 );
nand \U$4855 ( \4948 , \4947 , \4920 );
not \U$4856 ( \4949 , \4948 );
xor \U$4857 ( \4950 , \4945 , \4949 );
not \U$4858 ( \4951 , \4866 );
not \U$4859 ( \4952 , \4540 );
or \U$4860 ( \4953 , \4951 , \4952 );
not \U$4861 ( \4954 , \4482 );
and \U$4862 ( \4955 , \4954 , \3110 );
not \U$4863 ( \4956 , \4954 );
and \U$4864 ( \4957 , \4956 , \4864 );
nor \U$4865 ( \4958 , \4955 , \4957 );
nand \U$4866 ( \4959 , \2801 , \4958 );
nand \U$4867 ( \4960 , \4953 , \4959 );
not \U$4868 ( \4961 , \4873 );
nand \U$4869 ( \4962 , \3823 , \3126 );
not \U$4870 ( \4963 , \4962 );
or \U$4871 ( \4964 , \4961 , \4963 );
or \U$4872 ( \4965 , \4873 , \4962 );
nand \U$4873 ( \4966 , \4964 , \4965 );
xor \U$4874 ( \4967 , \4960 , \4966 );
not \U$4875 ( \4968 , \4912 );
not \U$4876 ( \4969 , \4905 );
or \U$4877 ( \4970 , \4968 , \4969 );
not \U$4878 ( \4971 , \4178 );
not \U$4879 ( \4972 , \3823 );
or \U$4880 ( \4973 , \4971 , \4972 );
buf \U$4881 ( \4974 , \3823 );
or \U$4882 ( \4975 , \4974 , \4178 );
nand \U$4883 ( \4976 , \4973 , \4975 );
nand \U$4884 ( \4977 , \3833 , \4976 );
nand \U$4885 ( \4978 , \4970 , \4977 );
not \U$4886 ( \4979 , \4978 );
not \U$4887 ( \4980 , \4900 );
not \U$4888 ( \4981 , \4478 );
or \U$4889 ( \4982 , \4980 , \4981 );
not \U$4890 ( \4983 , \192 );
not \U$4891 ( \4984 , \4457 );
or \U$4892 ( \4985 , \4983 , \4984 );
or \U$4893 ( \4986 , \4457 , \192 );
nand \U$4894 ( \4987 , \4985 , \4986 );
nand \U$4895 ( \4988 , \4135 , \4987 );
nand \U$4896 ( \4989 , \4982 , \4988 );
not \U$4897 ( \4990 , \4355 );
not \U$4898 ( \4991 , \4271 );
and \U$4899 ( \4992 , \4990 , \4991 );
nor \U$4900 ( \4993 , \4992 , \4277 );
xor \U$4901 ( \4994 , \4989 , \4993 );
not \U$4902 ( \4995 , \4994 );
or \U$4903 ( \4996 , \4979 , \4995 );
or \U$4904 ( \4997 , \4994 , \4978 );
nand \U$4905 ( \4998 , \4996 , \4997 );
xor \U$4906 ( \4999 , \4967 , \4998 );
not \U$4907 ( \5000 , \4893 );
xor \U$4908 ( \5001 , \5000 , \4914 );
and \U$4909 ( \5002 , \5001 , \4902 );
and \U$4910 ( \5003 , \5000 , \4914 );
nor \U$4911 ( \5004 , \5002 , \5003 );
xnor \U$4912 ( \5005 , \4999 , \5004 );
xor \U$4913 ( \5006 , \4950 , \5005 );
not \U$4914 ( \5007 , \4930 );
and \U$4915 ( \5008 , \5007 , \4891 );
and \U$4916 ( \5009 , \4881 , \4890 );
nor \U$4917 ( \5010 , \5008 , \5009 );
nand \U$4918 ( \5011 , \5006 , \5010 );
and \U$4919 ( \5012 , \4845 , \4935 , \5011 );
not \U$4920 ( \5013 , \4998 );
not \U$4921 ( \5014 , \5004 );
or \U$4922 ( \5015 , \5014 , \4967 );
not \U$4923 ( \5016 , \5015 );
or \U$4924 ( \5017 , \5013 , \5016 );
nand \U$4925 ( \5018 , \5014 , \4967 );
nand \U$4926 ( \5019 , \5017 , \5018 );
not \U$4927 ( \5020 , \4974 );
nor \U$4928 ( \5021 , \5020 , \2803 );
not \U$4929 ( \5022 , \4958 );
not \U$4930 ( \5023 , \4539 );
not \U$4931 ( \5024 , \5023 );
or \U$4932 ( \5025 , \5022 , \5024 );
xnor \U$4933 ( \5026 , \3110 , \4172 );
nand \U$4934 ( \5027 , \2801 , \5026 );
nand \U$4935 ( \5028 , \5025 , \5027 );
xor \U$4936 ( \5029 , \5021 , \5028 );
not \U$4937 ( \5030 , \4976 );
not \U$4938 ( \5031 , \4905 );
or \U$4939 ( \5032 , \5030 , \5031 );
xor \U$4940 ( \5033 , \4861 , \4974 );
nand \U$4941 ( \5034 , \3833 , \5033 );
nand \U$4942 ( \5035 , \5032 , \5034 );
xor \U$4943 ( \5036 , \5029 , \5035 );
not \U$4944 ( \5037 , \4993 );
or \U$4945 ( \5038 , \4978 , \5037 );
nand \U$4946 ( \5039 , \5038 , \4989 );
nand \U$4947 ( \5040 , \4978 , \5037 );
and \U$4948 ( \5041 , \5039 , \5040 );
not \U$4949 ( \5042 , \4987 );
not \U$4950 ( \5043 , \4478 );
or \U$4951 ( \5044 , \5042 , \5043 );
not \U$4952 ( \5045 , \4457 );
nand \U$4953 ( \5046 , \5045 , \4135 );
nand \U$4954 ( \5047 , \5044 , \5046 );
not \U$4955 ( \5048 , \5047 );
not \U$4956 ( \5049 , \4960 );
not \U$4957 ( \5050 , \4966 );
or \U$4958 ( \5051 , \5049 , \5050 );
not \U$4959 ( \5052 , \4962 );
nand \U$4960 ( \5053 , \5052 , \4873 );
nand \U$4961 ( \5054 , \5051 , \5053 );
xor \U$4962 ( \5055 , \5048 , \5054 );
xnor \U$4963 ( \5056 , \5041 , \5055 );
xor \U$4964 ( \5057 , \5036 , \5056 );
xor \U$4965 ( \5058 , \5019 , \5057 );
not \U$4966 ( \5059 , \5058 );
not \U$4967 ( \5060 , \4949 );
xor \U$4968 ( \5061 , \4945 , \5005 );
nand \U$4969 ( \5062 , \5060 , \5061 );
nand \U$4970 ( \5063 , \5005 , \4945 );
nand \U$4971 ( \5064 , \5059 , \5062 , \5063 );
and \U$4972 ( \5065 , \5036 , \5056 );
or \U$4973 ( \5066 , \5019 , \5065 );
or \U$4974 ( \5067 , \5056 , \5036 );
nand \U$4975 ( \5068 , \5066 , \5067 );
nand \U$4976 ( \5069 , \4974 , \4177 );
not \U$4977 ( \5070 , \193 );
xnor \U$4978 ( \5071 , \5070 , \4864 );
and \U$4979 ( \5072 , \5071 , \2801 );
and \U$4980 ( \5073 , \5023 , \5026 );
nor \U$4981 ( \5074 , \5072 , \5073 );
not \U$4982 ( \5075 , \5074 );
and \U$4983 ( \5076 , \5069 , \5075 );
not \U$4984 ( \5077 , \5069 );
and \U$4985 ( \5078 , \5077 , \5074 );
or \U$4986 ( \5079 , \5076 , \5078 );
not \U$4987 ( \5080 , \5079 );
or \U$4988 ( \5081 , \4478 , \4135 );
and \U$4989 ( \5082 , \5081 , \4137 );
not \U$4990 ( \5083 , \5082 );
and \U$4991 ( \5084 , \5080 , \5083 );
and \U$4992 ( \5085 , \5079 , \5082 );
nor \U$4993 ( \5086 , \5084 , \5085 );
xor \U$4994 ( \5087 , \5021 , \5028 );
and \U$4995 ( \5088 , \5087 , \5035 );
and \U$4996 ( \5089 , \5021 , \5028 );
nor \U$4997 ( \5090 , \5088 , \5089 );
not \U$4998 ( \5091 , \5048 );
not \U$4999 ( \5092 , \5033 );
not \U$5000 ( \5093 , \4905 );
or \U$5001 ( \5094 , \5092 , \5093 );
not \U$5002 ( \5095 , \4482 );
not \U$5003 ( \5096 , \4974 );
or \U$5004 ( \5097 , \5095 , \5096 );
or \U$5005 ( \5098 , \4974 , \4482 );
nand \U$5006 ( \5099 , \5097 , \5098 );
nand \U$5007 ( \5100 , \3833 , \5099 );
nand \U$5008 ( \5101 , \5094 , \5100 );
not \U$5009 ( \5102 , \5101 );
or \U$5010 ( \5103 , \5091 , \5102 );
or \U$5011 ( \5104 , \5101 , \5048 );
nand \U$5012 ( \5105 , \5103 , \5104 );
xor \U$5013 ( \5106 , \5090 , \5105 );
xor \U$5014 ( \5107 , \5086 , \5106 );
not \U$5015 ( \5108 , \5041 );
and \U$5016 ( \5109 , \5108 , \5055 );
and \U$5017 ( \5110 , \5048 , \5054 );
nor \U$5018 ( \5111 , \5109 , \5110 );
xor \U$5019 ( \5112 , \5107 , \5111 );
nand \U$5020 ( \5113 , \5068 , \5112 );
buf \U$5021 ( \5114 , \5113 );
xor \U$5022 ( \5115 , \5086 , \5106 );
and \U$5023 ( \5116 , \5115 , \5111 );
and \U$5024 ( \5117 , \5086 , \5106 );
or \U$5025 ( \5118 , \5116 , \5117 );
not \U$5026 ( \5119 , \5079 );
or \U$5027 ( \5120 , \5119 , \5082 );
not \U$5028 ( \5121 , \5069 );
nand \U$5029 ( \5122 , \5121 , \5075 );
nand \U$5030 ( \5123 , \5120 , \5122 );
not \U$5031 ( \5124 , \5123 );
not \U$5032 ( \5125 , \3833 );
xor \U$5033 ( \5126 , \4171 , \4974 );
not \U$5034 ( \5127 , \5126 );
or \U$5035 ( \5128 , \5125 , \5127 );
nand \U$5036 ( \5129 , \4905 , \5099 );
nand \U$5037 ( \5130 , \5128 , \5129 );
and \U$5038 ( \5131 , \4861 , \4974 );
not \U$5039 ( \5132 , \2800 );
not \U$5040 ( \5133 , \4864 );
and \U$5041 ( \5134 , \5132 , \5133 );
and \U$5042 ( \5135 , \5071 , \5023 );
nor \U$5043 ( \5136 , \5134 , \5135 );
xor \U$5044 ( \5137 , \5131 , \5136 );
xnor \U$5045 ( \5138 , \5130 , \5137 );
not \U$5046 ( \5139 , \5138 );
or \U$5047 ( \5140 , \5124 , \5139 );
or \U$5048 ( \5141 , \5138 , \5123 );
nand \U$5049 ( \5142 , \5140 , \5141 );
not \U$5050 ( \5143 , \5142 );
xor \U$5051 ( \5144 , \5021 , \5028 );
and \U$5052 ( \5145 , \5144 , \5035 );
and \U$5053 ( \5146 , \5021 , \5028 );
or \U$5054 ( \5147 , \5145 , \5146 );
and \U$5055 ( \5148 , \5147 , \5105 );
and \U$5056 ( \5149 , \5101 , \5047 );
nor \U$5057 ( \5150 , \5148 , \5149 );
not \U$5058 ( \5151 , \5150 );
and \U$5059 ( \5152 , \5143 , \5151 );
and \U$5060 ( \5153 , \5142 , \5150 );
nor \U$5061 ( \5154 , \5152 , \5153 );
nand \U$5062 ( \5155 , \5118 , \5154 );
not \U$5063 ( \5156 , \5155 );
not \U$5064 ( \5157 , \5023 );
not \U$5065 ( \5158 , \2801 );
and \U$5066 ( \5159 , \5157 , \5158 );
nor \U$5067 ( \5160 , \5159 , \4864 );
nand \U$5068 ( \5161 , \4974 , \4954 );
xor \U$5069 ( \5162 , \5160 , \5161 );
and \U$5070 ( \5163 , \4905 , \5126 );
xor \U$5071 ( \5164 , \4974 , \5070 );
and \U$5072 ( \5165 , \5164 , \3833 );
nor \U$5073 ( \5166 , \5163 , \5165 );
xor \U$5074 ( \5167 , \5162 , \5166 );
not \U$5075 ( \5168 , \5167 );
not \U$5076 ( \5169 , \5136 );
not \U$5077 ( \5170 , \5169 );
and \U$5078 ( \5171 , \5131 , \5136 );
not \U$5079 ( \5172 , \5171 );
nand \U$5080 ( \5173 , \5137 , \5130 );
nand \U$5081 ( \5174 , \5172 , \5173 );
not \U$5082 ( \5175 , \5174 );
not \U$5083 ( \5176 , \5175 );
or \U$5084 ( \5177 , \5170 , \5176 );
nand \U$5085 ( \5178 , \5174 , \5136 );
nand \U$5086 ( \5179 , \5177 , \5178 );
not \U$5087 ( \5180 , \5179 );
or \U$5088 ( \5181 , \5168 , \5180 );
or \U$5089 ( \5182 , \5167 , \5179 );
nand \U$5090 ( \5183 , \5181 , \5182 );
not \U$5091 ( \5184 , \5150 );
not \U$5092 ( \5185 , \5184 );
not \U$5093 ( \5186 , \5142 );
or \U$5094 ( \5187 , \5185 , \5186 );
not \U$5095 ( \5188 , \5138 );
nand \U$5096 ( \5189 , \5188 , \5123 );
nand \U$5097 ( \5190 , \5187 , \5189 );
nor \U$5098 ( \5191 , \5183 , \5190 );
nor \U$5099 ( \5192 , \5156 , \5191 );
and \U$5100 ( \5193 , \5012 , \5064 , \5114 , \5192 );
not \U$5101 ( \5194 , \5193 );
not \U$5102 ( \5195 , \4841 );
not \U$5103 ( \5196 , \4560 );
not \U$5104 ( \5197 , \4558 );
or \U$5105 ( \5198 , \5196 , \5197 );
or \U$5106 ( \5199 , \4560 , \4558 );
nand \U$5107 ( \5200 , \5198 , \5199 );
not \U$5108 ( \5201 , \5200 );
or \U$5109 ( \5202 , \5195 , \5201 );
or \U$5110 ( \5203 , \4841 , \5200 );
nand \U$5111 ( \5204 , \5202 , \5203 );
xor \U$5112 ( \5205 , \4380 , \4352 );
xor \U$5113 ( \5206 , \5205 , \4412 );
not \U$5114 ( \5207 , \4823 );
not \U$5115 ( \5208 , \4836 );
or \U$5116 ( \5209 , \5207 , \5208 );
not \U$5117 ( \5210 , \4823 );
nand \U$5118 ( \5211 , \5210 , \4835 );
nand \U$5119 ( \5212 , \5209 , \5211 );
and \U$5120 ( \5213 , \5212 , \4756 );
not \U$5121 ( \5214 , \5212 );
and \U$5122 ( \5215 , \5214 , \4757 );
nor \U$5123 ( \5216 , \5213 , \5215 );
xor \U$5124 ( \5217 , \5206 , \5216 );
not \U$5125 ( \5218 , \3127 );
not \U$5126 ( \5219 , \4116 );
or \U$5127 ( \5220 , \5218 , \5219 );
not \U$5128 ( \5221 , \4276 );
or \U$5129 ( \5222 , \5221 , \3127 );
nand \U$5130 ( \5223 , \5220 , \5222 );
not \U$5131 ( \5224 , \5223 );
not \U$5132 ( \5225 , \4266 );
not \U$5133 ( \5226 , \5225 );
or \U$5134 ( \5227 , \5224 , \5226 );
nand \U$5135 ( \5228 , \4779 , \4270 );
nand \U$5136 ( \5229 , \5227 , \5228 );
buf \U$5137 ( \5230 , \5229 );
not \U$5138 ( \5231 , \5230 );
not \U$5139 ( \5232 , \3977 );
and \U$5140 ( \5233 , \4151 , \5232 );
not \U$5141 ( \5234 , \4151 );
buf \U$5142 ( \5235 , \1710 );
and \U$5143 ( \5236 , \5234 , \5235 );
nor \U$5144 ( \5237 , \5233 , \5236 );
not \U$5145 ( \5238 , \5237 );
not \U$5146 ( \5239 , \3967 );
or \U$5147 ( \5240 , \5238 , \5239 );
nand \U$5148 ( \5241 , \4768 , \4373 );
nand \U$5149 ( \5242 , \5240 , \5241 );
not \U$5150 ( \5243 , \5242 );
or \U$5151 ( \5244 , \5231 , \5243 );
or \U$5152 ( \5245 , \5242 , \5230 );
and \U$5153 ( \5246 , \4178 , \4153 );
not \U$5154 ( \5247 , \4178 );
not \U$5155 ( \5248 , \4170 );
and \U$5156 ( \5249 , \5247 , \5248 );
or \U$5157 ( \5250 , \5246 , \5249 );
not \U$5158 ( \5251 , \5250 );
not \U$5159 ( \5252 , \4146 );
or \U$5160 ( \5253 , \5251 , \5252 );
nand \U$5161 ( \5254 , \1722 , \4800 );
nand \U$5162 ( \5255 , \5253 , \5254 );
nand \U$5163 ( \5256 , \5245 , \5255 );
nand \U$5164 ( \5257 , \5244 , \5256 );
not \U$5165 ( \5258 , \5257 );
xor \U$5166 ( \5259 , \4771 , \4783 );
xor \U$5167 ( \5260 , \5259 , \4788 );
not \U$5168 ( \5261 , \5260 );
or \U$5169 ( \5262 , \5258 , \5261 );
or \U$5170 ( \5263 , \5257 , \5260 );
xor \U$5171 ( \5264 , \130 , \3948 );
not \U$5172 ( \5265 , \5264 );
nand \U$5173 ( \5266 , \3755 , \5265 );
not \U$5174 ( \5267 , \5266 );
and \U$5175 ( \5268 , \3844 , \4333 );
not \U$5176 ( \5269 , \3844 );
and \U$5177 ( \5270 , \5269 , \3110 );
or \U$5178 ( \5271 , \5268 , \5270 );
not \U$5179 ( \5272 , \5271 );
not \U$5180 ( \5273 , \3140 );
or \U$5181 ( \5274 , \5272 , \5273 );
nand \U$5182 ( \5275 , \2799 , \4737 );
nand \U$5183 ( \5276 , \5274 , \5275 );
not \U$5184 ( \5277 , \5276 );
not \U$5185 ( \5278 , \5277 );
or \U$5186 ( \5279 , \5267 , \5278 );
and \U$5187 ( \5280 , \4506 , \3984 );
not \U$5188 ( \5281 , \4506 );
and \U$5189 ( \5282 , \5281 , \4137 );
or \U$5190 ( \5283 , \5280 , \5282 );
not \U$5191 ( \5284 , \5283 );
not \U$5192 ( \5285 , \4391 );
or \U$5193 ( \5286 , \5284 , \5285 );
not \U$5194 ( \5287 , \4814 );
nand \U$5195 ( \5288 , \5287 , \4810 );
nand \U$5196 ( \5289 , \5286 , \5288 );
nand \U$5197 ( \5290 , \5279 , \5289 );
not \U$5198 ( \5291 , \5266 );
nand \U$5199 ( \5292 , \5291 , \5276 );
nand \U$5200 ( \5293 , \5290 , \5292 );
nand \U$5201 ( \5294 , \5263 , \5293 );
nand \U$5202 ( \5295 , \5262 , \5294 );
not \U$5203 ( \5296 , \5295 );
xor \U$5204 ( \5297 , \3979 , \4791 );
xor \U$5205 ( \5298 , \5297 , \4820 );
not \U$5206 ( \5299 , \5298 );
nand \U$5207 ( \5300 , \5296 , \5299 );
xor \U$5208 ( \5301 , \4748 , \4750 );
xor \U$5209 ( \5302 , \5301 , \4753 );
not \U$5210 ( \5303 , \5302 );
and \U$5211 ( \5304 , \5300 , \5303 );
nor \U$5212 ( \5305 , \5296 , \5299 );
nor \U$5213 ( \5306 , \5304 , \5305 );
and \U$5214 ( \5307 , \5217 , \5306 );
and \U$5215 ( \5308 , \5206 , \5216 );
or \U$5216 ( \5309 , \5307 , \5308 );
nand \U$5217 ( \5310 , \5204 , \5309 );
xor \U$5218 ( \5311 , \5257 , \5260 );
xor \U$5219 ( \5312 , \5311 , \5293 );
not \U$5220 ( \5313 , \5312 );
xor \U$5221 ( \5314 , \5229 , \5255 );
xnor \U$5222 ( \5315 , \5314 , \5242 );
not \U$5223 ( \5316 , \5315 );
and \U$5224 ( \5317 , \3821 , \4775 );
not \U$5225 ( \5318 , \3821 );
and \U$5226 ( \5319 , \5318 , \4276 );
nor \U$5227 ( \5320 , \5317 , \5319 );
not \U$5228 ( \5321 , \5320 );
nand \U$5229 ( \5322 , \4260 , \4265 );
not \U$5230 ( \5323 , \5322 );
not \U$5231 ( \5324 , \5323 );
or \U$5232 ( \5325 , \5321 , \5324 );
nand \U$5233 ( \5326 , \5223 , \4270 );
nand \U$5234 ( \5327 , \5325 , \5326 );
buf \U$5235 ( \5328 , \5327 );
not \U$5236 ( \5329 , \5328 );
not \U$5237 ( \5330 , \4274 );
not \U$5238 ( \5331 , \5235 );
or \U$5239 ( \5332 , \5330 , \5331 );
or \U$5240 ( \5333 , \5235 , \4274 );
nand \U$5241 ( \5334 , \5332 , \5333 );
not \U$5242 ( \5335 , \5334 );
nand \U$5243 ( \5336 , \4762 , \3965 );
not \U$5244 ( \5337 , \5336 );
not \U$5245 ( \5338 , \5337 );
or \U$5246 ( \5339 , \5335 , \5338 );
nand \U$5247 ( \5340 , \5237 , \3975 );
nand \U$5248 ( \5341 , \5339 , \5340 );
buf \U$5249 ( \5342 , \5341 );
not \U$5250 ( \5343 , \5342 );
or \U$5251 ( \5344 , \5329 , \5343 );
or \U$5252 ( \5345 , \5342 , \5328 );
not \U$5253 ( \5346 , \4718 );
not \U$5254 ( \5347 , \4696 );
or \U$5255 ( \5348 , \5346 , \5347 );
not \U$5256 ( \5349 , \4172 );
not \U$5257 ( \5350 , \4713 );
or \U$5258 ( \5351 , \5349 , \5350 );
not \U$5259 ( \5352 , \4699 );
or \U$5260 ( \5353 , \5352 , \4172 );
nand \U$5261 ( \5354 , \5351 , \5353 );
nand \U$5262 ( \5355 , \4711 , \5354 );
nand \U$5263 ( \5356 , \5348 , \5355 );
nand \U$5264 ( \5357 , \5345 , \5356 );
nand \U$5265 ( \5358 , \5344 , \5357 );
nand \U$5266 ( \5359 , \5316 , \5358 );
not \U$5267 ( \5360 , \5359 );
nand \U$5268 ( \5361 , \3490 , \3753 );
xnor \U$5269 ( \5362 , \126 , \4635 );
not \U$5270 ( \5363 , \5362 );
nand \U$5271 ( \5364 , \5361 , \5363 );
not \U$5272 ( \5365 , \5364 );
and \U$5273 ( \5366 , \4315 , \3984 );
not \U$5274 ( \5367 , \4315 );
and \U$5275 ( \5368 , \5367 , \4137 );
nor \U$5276 ( \5369 , \5366 , \5368 );
not \U$5277 ( \5370 , \5369 );
not \U$5278 ( \5371 , \4131 );
or \U$5279 ( \5372 , \5370 , \5371 );
not \U$5280 ( \5373 , \4814 );
nand \U$5281 ( \5374 , \5373 , \5283 );
nand \U$5282 ( \5375 , \5372 , \5374 );
xor \U$5283 ( \5376 , \5365 , \5375 );
not \U$5284 ( \5377 , \5264 );
not \U$5285 ( \5378 , \5361 );
or \U$5286 ( \5379 , \5377 , \5378 );
or \U$5287 ( \5380 , \4302 , \5264 );
nand \U$5288 ( \5381 , \5379 , \5380 );
not \U$5289 ( \5382 , \5381 );
not \U$5290 ( \5383 , \3814 );
or \U$5291 ( \5384 , \5382 , \5383 );
not \U$5292 ( \5385 , \4793 );
not \U$5293 ( \5386 , \4302 );
or \U$5294 ( \5387 , \5385 , \5386 );
not \U$5295 ( \5388 , \3755 );
not \U$5296 ( \5389 , \5388 );
or \U$5297 ( \5390 , \5389 , \4793 );
nand \U$5298 ( \5391 , \5387 , \5390 );
nand \U$5299 ( \5392 , \5391 , \3833 );
nand \U$5300 ( \5393 , \5384 , \5392 );
and \U$5301 ( \5394 , \5376 , \5393 );
and \U$5302 ( \5395 , \5365 , \5375 );
or \U$5303 ( \5396 , \5394 , \5395 );
not \U$5304 ( \5397 , \5396 );
not \U$5305 ( \5398 , \5397 );
or \U$5306 ( \5399 , \5360 , \5398 );
or \U$5307 ( \5400 , \5358 , \5316 );
nand \U$5308 ( \5401 , \5399 , \5400 );
not \U$5309 ( \5402 , \5401 );
and \U$5310 ( \5403 , \5313 , \5402 );
and \U$5311 ( \5404 , \5401 , \5312 );
nor \U$5312 ( \5405 , \5403 , \5404 );
not \U$5313 ( \5406 , \5405 );
not \U$5314 ( \5407 , \5406 );
not \U$5315 ( \5408 , \4746 );
not \U$5316 ( \5409 , \5408 );
buf \U$5317 ( \5410 , \4621 );
buf \U$5318 ( \5411 , \5410 );
not \U$5319 ( \5412 , \2803 );
not \U$5320 ( \5413 , \1562 );
or \U$5321 ( \5414 , \5412 , \5413 );
or \U$5322 ( \5415 , \1562 , \2803 );
nand \U$5323 ( \5416 , \5414 , \5415 );
not \U$5324 ( \5417 , \5416 );
not \U$5325 ( \5418 , \1719 );
or \U$5326 ( \5419 , \5417 , \5418 );
nand \U$5327 ( \5420 , \1722 , \5250 );
nand \U$5328 ( \5421 , \5419 , \5420 );
not \U$5329 ( \5422 , \5421 );
and \U$5330 ( \5423 , \5411 , \5422 );
not \U$5331 ( \5424 , \5423 );
not \U$5332 ( \5425 , \3815 );
not \U$5333 ( \5426 , \5391 );
or \U$5334 ( \5427 , \5425 , \5426 );
nand \U$5335 ( \5428 , \3833 , \4726 );
nand \U$5336 ( \5429 , \5427 , \5428 );
nand \U$5337 ( \5430 , \5424 , \5429 );
not \U$5338 ( \5431 , \5430 );
or \U$5339 ( \5432 , \5409 , \5431 );
not \U$5340 ( \5433 , \5429 );
nand \U$5341 ( \5434 , \5433 , \5423 );
nand \U$5342 ( \5435 , \5432 , \5434 );
not \U$5343 ( \5436 , \5435 );
buf \U$5344 ( \5437 , \4730 );
not \U$5345 ( \5438 , \5437 );
not \U$5346 ( \5439 , \4746 );
not \U$5347 ( \5440 , \4742 );
or \U$5348 ( \5441 , \5439 , \5440 );
or \U$5349 ( \5442 , \4742 , \4746 );
nand \U$5350 ( \5443 , \5441 , \5442 );
not \U$5351 ( \5444 , \5443 );
or \U$5352 ( \5445 , \5438 , \5444 );
or \U$5353 ( \5446 , \5443 , \5437 );
nand \U$5354 ( \5447 , \5445 , \5446 );
not \U$5355 ( \5448 , \5447 );
xor \U$5356 ( \5449 , \4794 , \4805 );
xor \U$5357 ( \5450 , \5449 , \4817 );
not \U$5358 ( \5451 , \5450 );
and \U$5359 ( \5452 , \5448 , \5451 );
and \U$5360 ( \5453 , \5447 , \5450 );
nor \U$5361 ( \5454 , \5452 , \5453 );
not \U$5362 ( \5455 , \5454 );
or \U$5363 ( \5456 , \5436 , \5455 );
or \U$5364 ( \5457 , \5435 , \5454 );
nand \U$5365 ( \5458 , \5456 , \5457 );
not \U$5366 ( \5459 , \5458 );
or \U$5367 ( \5460 , \5407 , \5459 );
not \U$5368 ( \5461 , \5312 );
nand \U$5369 ( \5462 , \5461 , \5401 );
nand \U$5370 ( \5463 , \5460 , \5462 );
not \U$5371 ( \5464 , \5463 );
not \U$5372 ( \5465 , \5435 );
not \U$5373 ( \5466 , \5454 );
not \U$5374 ( \5467 , \5466 );
or \U$5375 ( \5468 , \5465 , \5467 );
not \U$5376 ( \5469 , \5450 );
nand \U$5377 ( \5470 , \5469 , \5447 );
nand \U$5378 ( \5471 , \5468 , \5470 );
not \U$5379 ( \5472 , \5471 );
not \U$5380 ( \5473 , \5295 );
not \U$5381 ( \5474 , \5298 );
or \U$5382 ( \5475 , \5473 , \5474 );
or \U$5383 ( \5476 , \5295 , \5298 );
nand \U$5384 ( \5477 , \5475 , \5476 );
not \U$5385 ( \5478 , \5477 );
not \U$5386 ( \5479 , \5478 );
not \U$5387 ( \5480 , \5302 );
not \U$5388 ( \5481 , \5480 );
or \U$5389 ( \5482 , \5479 , \5481 );
nand \U$5390 ( \5483 , \5302 , \5477 );
nand \U$5391 ( \5484 , \5482 , \5483 );
not \U$5392 ( \5485 , \5484 );
not \U$5393 ( \5486 , \5485 );
or \U$5394 ( \5487 , \5472 , \5486 );
not \U$5395 ( \5488 , \5471 );
nand \U$5396 ( \5489 , \5488 , \5484 );
nand \U$5397 ( \5490 , \5487 , \5489 );
not \U$5398 ( \5491 , \5490 );
or \U$5399 ( \5492 , \5464 , \5491 );
not \U$5400 ( \5493 , \5478 );
not \U$5401 ( \5494 , \5480 );
or \U$5402 ( \5495 , \5493 , \5494 );
nand \U$5403 ( \5496 , \5495 , \5483 );
nand \U$5404 ( \5497 , \5496 , \5471 );
nand \U$5405 ( \5498 , \5492 , \5497 );
xor \U$5406 ( \5499 , \5206 , \5216 );
xor \U$5407 ( \5500 , \5499 , \5306 );
nand \U$5408 ( \5501 , \5498 , \5500 );
nand \U$5409 ( \5502 , \5310 , \5501 );
not \U$5410 ( \5503 , \5502 );
not \U$5411 ( \5504 , \5503 );
not \U$5412 ( \5505 , \5463 );
not \U$5413 ( \5506 , \5490 );
not \U$5414 ( \5507 , \5506 );
or \U$5415 ( \5508 , \5505 , \5507 );
not \U$5416 ( \5509 , \5463 );
nand \U$5417 ( \5510 , \5509 , \5490 );
nand \U$5418 ( \5511 , \5508 , \5510 );
xnor \U$5419 ( \5512 , \4327 , \3115 );
and \U$5420 ( \5513 , \4540 , \5512 );
not \U$5421 ( \5514 , \5271 );
nor \U$5422 ( \5515 , \5514 , \2800 );
nor \U$5423 ( \5516 , \5513 , \5515 );
not \U$5424 ( \5517 , \5516 );
not \U$5425 ( \5518 , \3127 );
not \U$5426 ( \5519 , \1562 );
or \U$5427 ( \5520 , \5518 , \5519 );
or \U$5428 ( \5521 , \4167 , \3127 );
nand \U$5429 ( \5522 , \5520 , \5521 );
not \U$5430 ( \5523 , \5522 );
not \U$5431 ( \5524 , \1719 );
or \U$5432 ( \5525 , \5523 , \5524 );
nand \U$5433 ( \5526 , \1724 , \5416 );
nand \U$5434 ( \5527 , \5525 , \5526 );
not \U$5435 ( \5528 , \5527 );
not \U$5436 ( \5529 , \4267 );
not \U$5437 ( \5530 , \3151 );
not \U$5438 ( \5531 , \4116 );
or \U$5439 ( \5532 , \5530 , \5531 );
not \U$5440 ( \5533 , \4120 );
or \U$5441 ( \5534 , \5533 , \3151 );
nand \U$5442 ( \5535 , \5532 , \5534 );
not \U$5443 ( \5536 , \5535 );
or \U$5444 ( \5537 , \5529 , \5536 );
buf \U$5445 ( \5538 , \5320 );
nand \U$5446 ( \5539 , \5538 , \4271 );
nand \U$5447 ( \5540 , \5537 , \5539 );
not \U$5448 ( \5541 , \5540 );
not \U$5449 ( \5542 , \4151 );
not \U$5450 ( \5543 , \4698 );
or \U$5451 ( \5544 , \5542 , \5543 );
not \U$5452 ( \5545 , \4698 );
not \U$5453 ( \5546 , \5545 );
or \U$5454 ( \5547 , \5546 , \4151 );
nand \U$5455 ( \5548 , \5544 , \5547 );
not \U$5456 ( \5549 , \5548 );
not \U$5457 ( \5550 , \4711 );
or \U$5458 ( \5551 , \5549 , \5550 );
nand \U$5459 ( \5552 , \5354 , \4696 );
nand \U$5460 ( \5553 , \5551 , \5552 );
not \U$5461 ( \5554 , \5553 );
xor \U$5462 ( \5555 , \5541 , \5554 );
nand \U$5463 ( \5556 , \5528 , \5555 );
and \U$5464 ( \5557 , \5541 , \5554 );
not \U$5465 ( \5558 , \5557 );
nand \U$5466 ( \5559 , \5517 , \5556 , \5558 );
xor \U$5467 ( \5560 , \5266 , \5276 );
xor \U$5468 ( \5561 , \5560 , \5289 );
xor \U$5469 ( \5562 , \5559 , \5561 );
xor \U$5470 ( \5563 , \5408 , \5423 );
xnor \U$5471 ( \5564 , \5563 , \5429 );
and \U$5472 ( \5565 , \5562 , \5564 );
and \U$5473 ( \5566 , \5559 , \5561 );
nor \U$5474 ( \5567 , \5565 , \5566 );
not \U$5475 ( \5568 , \5567 );
not \U$5476 ( \5569 , \5397 );
not \U$5477 ( \5570 , \5358 );
not \U$5478 ( \5571 , \5315 );
or \U$5479 ( \5572 , \5570 , \5571 );
or \U$5480 ( \5573 , \5358 , \5315 );
nand \U$5481 ( \5574 , \5572 , \5573 );
not \U$5482 ( \5575 , \5574 );
or \U$5483 ( \5576 , \5569 , \5575 );
or \U$5484 ( \5577 , \5574 , \5397 );
nand \U$5485 ( \5578 , \5576 , \5577 );
xor \U$5486 ( \5579 , \4177 , \3977 );
not \U$5487 ( \5580 , \5579 );
not \U$5488 ( \5581 , \3967 );
or \U$5489 ( \5582 , \5580 , \5581 );
nand \U$5490 ( \5583 , \4375 , \5334 );
nand \U$5491 ( \5584 , \5582 , \5583 );
not \U$5492 ( \5585 , \5584 );
not \U$5493 ( \5586 , \3813 );
not \U$5494 ( \5587 , \5362 );
not \U$5495 ( \5588 , \5361 );
not \U$5496 ( \5589 , \5588 );
or \U$5497 ( \5590 , \5587 , \5589 );
nand \U$5498 ( \5591 , \5590 , \5364 );
not \U$5499 ( \5592 , \5591 );
not \U$5500 ( \5593 , \5592 );
or \U$5501 ( \5594 , \5586 , \5593 );
nand \U$5502 ( \5595 , \3832 , \5381 );
nand \U$5503 ( \5596 , \5594 , \5595 );
xor \U$5504 ( \5597 , \122 , \4610 );
not \U$5505 ( \5598 , \5597 );
nand \U$5506 ( \5599 , \4304 , \5598 );
not \U$5507 ( \5600 , \5599 );
and \U$5508 ( \5601 , \5596 , \5600 );
not \U$5509 ( \5602 , \5596 );
and \U$5510 ( \5603 , \5602 , \5599 );
nor \U$5511 ( \5604 , \5601 , \5603 );
not \U$5512 ( \5605 , \5604 );
or \U$5513 ( \5606 , \5585 , \5605 );
buf \U$5514 ( \5607 , \5596 );
nand \U$5515 ( \5608 , \5607 , \5600 );
nand \U$5516 ( \5609 , \5606 , \5608 );
not \U$5517 ( \5610 , \5609 );
xor \U$5518 ( \5611 , \5327 , \5341 );
xnor \U$5519 ( \5612 , \5611 , \5356 );
not \U$5520 ( \5613 , \5612 );
xor \U$5521 ( \5614 , \5411 , \5422 );
not \U$5522 ( \5615 , \5614 );
nand \U$5523 ( \5616 , \5613 , \5615 );
buf \U$5524 ( \5617 , \5616 );
and \U$5525 ( \5618 , \5610 , \5617 );
not \U$5526 ( \5619 , \5614 );
nor \U$5527 ( \5620 , \5619 , \5613 );
nor \U$5528 ( \5621 , \5618 , \5620 );
nand \U$5529 ( \5622 , \5578 , \5621 );
not \U$5530 ( \5623 , \5622 );
not \U$5531 ( \5624 , \5516 );
not \U$5532 ( \5625 , \5556 );
nor \U$5533 ( \5626 , \5625 , \5557 );
not \U$5534 ( \5627 , \5626 );
or \U$5535 ( \5628 , \5624 , \5627 );
not \U$5536 ( \5629 , \5558 );
not \U$5537 ( \5630 , \5556 );
or \U$5538 ( \5631 , \5629 , \5630 );
nand \U$5539 ( \5632 , \5631 , \5517 );
nand \U$5540 ( \5633 , \5628 , \5632 );
not \U$5541 ( \5634 , \5633 );
not \U$5542 ( \5635 , \5634 );
xor \U$5543 ( \5636 , \5365 , \5375 );
xor \U$5544 ( \5637 , \5636 , \5393 );
not \U$5545 ( \5638 , \5637 );
not \U$5546 ( \5639 , \5638 );
or \U$5547 ( \5640 , \5635 , \5639 );
not \U$5548 ( \5641 , \5637 );
not \U$5549 ( \5642 , \5633 );
or \U$5550 ( \5643 , \5641 , \5642 );
and \U$5551 ( \5644 , \2779 , RI8928e48_16);
not \U$5552 ( \5645 , RI892a4c8_64);
not \U$5553 ( \5646 , \1575 );
or \U$5554 ( \5647 , \5645 , \5646 );
not \U$5555 ( \5648 , \1644 );
not \U$5556 ( \5649 , \4090 );
nand \U$5557 ( \5650 , \5648 , \5649 );
not \U$5558 ( \5651 , \989 );
and \U$5559 ( \5652 , \5650 , \5651 );
and \U$5560 ( \5653 , RI8928e48_16, \2730 );
or \U$5561 ( \5654 , \405 , RI89295c8_32);
nand \U$5562 ( \5655 , \5654 , \3991 );
nor \U$5563 ( \5656 , \5653 , \5655 );
or \U$5564 ( \5657 , \5656 , \3517 );
or \U$5565 ( \5658 , \405 , RI892a4c8_64);
nand \U$5566 ( \5659 , \5658 , \424 );
and \U$5567 ( \5660 , \5659 , RI89295c8_32);
not \U$5568 ( \5661 , \1817 );
and \U$5569 ( \5662 , RI8929d48_48, \1417 );
not \U$5570 ( \5663 , RI8929d48_48);
and \U$5571 ( \5664 , \5663 , RI8928e48_16);
nor \U$5572 ( \5665 , \5662 , \5664 );
or \U$5573 ( \5666 , \5661 , \5665 );
not \U$5574 ( \5667 , RI8929d48_48);
or \U$5575 ( \5668 , \419 , \5667 );
nand \U$5576 ( \5669 , \5666 , \5668 );
nor \U$5577 ( \5670 , \5660 , \5669 );
nand \U$5578 ( \5671 , \5657 , \5670 );
nor \U$5579 ( \5672 , \5652 , \5671 );
and \U$5580 ( \5673 , RI8929d48_48, RI892a4c8_64);
not \U$5581 ( \5674 , RI8929d48_48);
and \U$5582 ( \5675 , \5674 , \3517 );
nor \U$5583 ( \5676 , \5673 , \5675 );
nand \U$5584 ( \5677 , \1741 , \5676 );
nand \U$5585 ( \5678 , \1417 , \284 );
nand \U$5586 ( \5679 , \5678 , \1547 );
and \U$5587 ( \5680 , \5672 , \5677 , \5679 );
nand \U$5588 ( \5681 , \5647 , \5680 );
nor \U$5589 ( \5682 , \5644 , \5681 );
and \U$5590 ( \5683 , \4621 , \5682 );
buf \U$5591 ( \5684 , \5683 );
not \U$5592 ( \5685 , \193 );
buf \U$5593 ( \5686 , \4621 );
not \U$5594 ( \5687 , \5686 );
or \U$5595 ( \5688 , \5685 , \5687 );
or \U$5596 ( \5689 , \5410 , \193 );
nand \U$5597 ( \5690 , \5688 , \5689 );
nand \U$5598 ( \5691 , \5684 , \5690 );
not \U$5599 ( \5692 , \5682 );
buf \U$5600 ( \5693 , \5692 );
nand \U$5601 ( \5694 , \5411 , \5693 );
nand \U$5602 ( \5695 , \5691 , \5694 );
and \U$5603 ( \5696 , \3843 , \3984 );
not \U$5604 ( \5697 , \3843 );
and \U$5605 ( \5698 , \5697 , \4137 );
nor \U$5606 ( \5699 , \5696 , \5698 );
not \U$5607 ( \5700 , \5699 );
not \U$5608 ( \5701 , \4131 );
or \U$5609 ( \5702 , \5700 , \5701 );
nand \U$5610 ( \5703 , \4135 , \5369 );
nand \U$5611 ( \5704 , \5702 , \5703 );
xor \U$5612 ( \5705 , \5695 , \5704 );
not \U$5613 ( \5706 , \4793 );
not \U$5614 ( \5707 , \3115 );
or \U$5615 ( \5708 , \5706 , \5707 );
or \U$5616 ( \5709 , \3110 , \4793 );
nand \U$5617 ( \5710 , \5708 , \5709 );
not \U$5618 ( \5711 , \5710 );
not \U$5619 ( \5712 , \3142 );
or \U$5620 ( \5713 , \5711 , \5712 );
nand \U$5621 ( \5714 , \2801 , \5512 );
nand \U$5622 ( \5715 , \5713 , \5714 );
and \U$5623 ( \5716 , \5705 , \5715 );
and \U$5624 ( \5717 , \5695 , \5704 );
or \U$5625 ( \5718 , \5716 , \5717 );
not \U$5626 ( \5719 , \5718 );
nand \U$5627 ( \5720 , \5643 , \5719 );
nand \U$5628 ( \5721 , \5640 , \5720 );
not \U$5629 ( \5722 , \5721 );
or \U$5630 ( \5723 , \5623 , \5722 );
not \U$5631 ( \5724 , \5578 );
not \U$5632 ( \5725 , \5621 );
nand \U$5633 ( \5726 , \5724 , \5725 );
nand \U$5634 ( \5727 , \5723 , \5726 );
not \U$5635 ( \5728 , \5727 );
or \U$5636 ( \5729 , \5568 , \5728 );
or \U$5637 ( \5730 , \5727 , \5567 );
nand \U$5638 ( \5731 , \5729 , \5730 );
not \U$5639 ( \5732 , \5731 );
not \U$5640 ( \5733 , \5405 );
not \U$5641 ( \5734 , \5458 );
and \U$5642 ( \5735 , \5733 , \5734 );
and \U$5643 ( \5736 , \5458 , \5405 );
nor \U$5644 ( \5737 , \5735 , \5736 );
not \U$5645 ( \5738 , \5737 );
not \U$5646 ( \5739 , \5738 );
or \U$5647 ( \5740 , \5732 , \5739 );
not \U$5648 ( \5741 , \5567 );
nand \U$5649 ( \5742 , \5741 , \5727 );
nand \U$5650 ( \5743 , \5740 , \5742 );
nand \U$5651 ( \5744 , \5511 , \5743 );
not \U$5652 ( \5745 , \5744 );
not \U$5653 ( \5746 , \5745 );
not \U$5654 ( \5747 , \5731 );
not \U$5655 ( \5748 , \5737 );
and \U$5656 ( \5749 , \5747 , \5748 );
and \U$5657 ( \5750 , \5737 , \5731 );
nor \U$5658 ( \5751 , \5749 , \5750 );
not \U$5659 ( \5752 , \5751 );
xnor \U$5660 ( \5753 , \5597 , \3755 );
not \U$5661 ( \5754 , \5753 );
not \U$5662 ( \5755 , \3814 );
or \U$5663 ( \5756 , \5754 , \5755 );
not \U$5664 ( \5757 , \5591 );
nand \U$5665 ( \5758 , \5757 , \3832 );
nand \U$5666 ( \5759 , \5756 , \5758 );
not \U$5667 ( \5760 , \4328 );
not \U$5668 ( \5761 , \3987 );
or \U$5669 ( \5762 , \5760 , \5761 );
or \U$5670 ( \5763 , \3984 , \4328 );
nand \U$5671 ( \5764 , \5762 , \5763 );
not \U$5672 ( \5765 , \5764 );
not \U$5673 ( \5766 , \4131 );
or \U$5674 ( \5767 , \5765 , \5766 );
nand \U$5675 ( \5768 , \4134 , \5699 );
nand \U$5676 ( \5769 , \5767 , \5768 );
nand \U$5677 ( \5770 , \5759 , \5769 );
and \U$5678 ( \5771 , \5264 , \3825 );
not \U$5679 ( \5772 , \5264 );
and \U$5680 ( \5773 , \5772 , \3115 );
nor \U$5681 ( \5774 , \5771 , \5773 );
not \U$5682 ( \5775 , \5774 );
not \U$5683 ( \5776 , \3140 );
or \U$5684 ( \5777 , \5775 , \5776 );
nand \U$5685 ( \5778 , \2799 , \5710 );
nand \U$5686 ( \5779 , \5777 , \5778 );
nand \U$5687 ( \5780 , \5759 , \5779 );
nand \U$5688 ( \5781 , \5779 , \5769 );
nand \U$5689 ( \5782 , \5770 , \5780 , \5781 );
not \U$5690 ( \5783 , \5782 );
and \U$5691 ( \5784 , \3822 , \5248 );
not \U$5692 ( \5785 , \3822 );
and \U$5693 ( \5786 , \5785 , \4798 );
nor \U$5694 ( \5787 , \5784 , \5786 );
not \U$5695 ( \5788 , \5787 );
not \U$5696 ( \5789 , \1719 );
or \U$5697 ( \5790 , \5788 , \5789 );
nand \U$5698 ( \5791 , \4161 , \5522 );
nand \U$5699 ( \5792 , \5790 , \5791 );
not \U$5700 ( \5793 , \5792 );
not \U$5701 ( \5794 , \5579 );
not \U$5702 ( \5795 , \3958 );
or \U$5703 ( \5796 , \5794 , \5795 );
not \U$5704 ( \5797 , \2803 );
not \U$5705 ( \5798 , \1710 );
or \U$5706 ( \5799 , \5797 , \5798 );
or \U$5707 ( \5800 , \3977 , \2803 );
nand \U$5708 ( \5801 , \5799 , \5800 );
nand \U$5709 ( \5802 , \4762 , \5801 , \3965 );
nand \U$5710 ( \5803 , \5796 , \5802 );
not \U$5711 ( \5804 , \4315 );
not \U$5712 ( \5805 , \4775 );
or \U$5713 ( \5806 , \5804 , \5805 );
or \U$5714 ( \5807 , \5533 , \4315 );
nand \U$5715 ( \5808 , \5806 , \5807 );
not \U$5716 ( \5809 , \5808 );
not \U$5717 ( \5810 , \5225 );
or \U$5718 ( \5811 , \5809 , \5810 );
nand \U$5719 ( \5812 , \5535 , \4270 );
nand \U$5720 ( \5813 , \5811 , \5812 );
and \U$5721 ( \5814 , \5803 , \5813 );
not \U$5722 ( \5815 , \5803 );
not \U$5723 ( \5816 , \5813 );
and \U$5724 ( \5817 , \5815 , \5816 );
nor \U$5725 ( \5818 , \5814 , \5817 );
not \U$5726 ( \5819 , \5818 );
or \U$5727 ( \5820 , \5793 , \5819 );
nand \U$5728 ( \5821 , \5813 , \5803 );
nand \U$5729 ( \5822 , \5820 , \5821 );
not \U$5730 ( \5823 , \5822 );
and \U$5731 ( \5824 , \4621 , \5682 );
not \U$5732 ( \5825 , \5824 );
not \U$5733 ( \5826 , \4165 );
not \U$5734 ( \5827 , \5686 );
or \U$5735 ( \5828 , \5826 , \5827 );
or \U$5736 ( \5829 , \5410 , \4165 );
nand \U$5737 ( \5830 , \5828 , \5829 );
not \U$5738 ( \5831 , \5830 );
or \U$5739 ( \5832 , \5825 , \5831 );
nand \U$5740 ( \5833 , \5690 , \5693 );
nand \U$5741 ( \5834 , \5832 , \5833 );
not \U$5742 ( \5835 , \5834 );
not \U$5743 ( \5836 , \5835 );
buf \U$5744 ( \5837 , \5676 );
buf \U$5745 ( \5838 , \5837 );
buf \U$5746 ( \5839 , \5838 );
nand \U$5747 ( \5840 , \5836 , \5389 , \5839 );
not \U$5748 ( \5841 , \5840 );
buf \U$5749 ( \5842 , \5838 );
and \U$5750 ( \5843 , \4302 , \5842 );
nand \U$5751 ( \5844 , \5843 , \5835 );
not \U$5752 ( \5845 , \5839 );
not \U$5753 ( \5846 , \3755 );
or \U$5754 ( \5847 , \5845 , \5846 );
nand \U$5755 ( \5848 , \5847 , \5834 );
and \U$5756 ( \5849 , \5844 , \5848 );
not \U$5757 ( \5850 , \4694 );
not \U$5758 ( \5851 , \5850 );
not \U$5759 ( \5852 , \5851 );
not \U$5760 ( \5853 , \5548 );
or \U$5761 ( \5854 , \5852 , \5853 );
and \U$5762 ( \5855 , \4274 , \4699 );
not \U$5763 ( \5856 , \4274 );
and \U$5764 ( \5857 , \5856 , \4698 );
or \U$5765 ( \5858 , \5855 , \5857 );
not \U$5766 ( \5859 , \5858 );
nand \U$5767 ( \5860 , \5859 , \4711 );
nand \U$5768 ( \5861 , \5854 , \5860 );
not \U$5769 ( \5862 , \5861 );
nor \U$5770 ( \5863 , \5849 , \5862 );
nor \U$5771 ( \5864 , \5841 , \5863 );
not \U$5772 ( \5865 , \5864 );
or \U$5773 ( \5866 , \5823 , \5865 );
not \U$5774 ( \5867 , \5840 );
not \U$5775 ( \5868 , \5863 );
not \U$5776 ( \5869 , \5868 );
or \U$5777 ( \5870 , \5867 , \5869 );
not \U$5778 ( \5871 , \5822 );
nand \U$5779 ( \5872 , \5870 , \5871 );
nand \U$5780 ( \5873 , \5866 , \5872 );
not \U$5781 ( \5874 , \5873 );
or \U$5782 ( \5875 , \5783 , \5874 );
not \U$5783 ( \5876 , \5840 );
not \U$5784 ( \5877 , \5868 );
or \U$5785 ( \5878 , \5876 , \5877 );
nand \U$5786 ( \5879 , \5878 , \5822 );
nand \U$5787 ( \5880 , \5875 , \5879 );
not \U$5788 ( \5881 , \5880 );
not \U$5789 ( \5882 , \5881 );
not \U$5790 ( \5883 , \5555 );
not \U$5791 ( \5884 , \5527 );
and \U$5792 ( \5885 , \5883 , \5884 );
and \U$5793 ( \5886 , \5555 , \5527 );
nor \U$5794 ( \5887 , \5885 , \5886 );
not \U$5795 ( \5888 , \5887 );
xor \U$5796 ( \5889 , \5599 , \5596 );
xor \U$5797 ( \5890 , \5889 , \5584 );
not \U$5798 ( \5891 , \5890 );
not \U$5799 ( \5892 , \5891 );
or \U$5800 ( \5893 , \5888 , \5892 );
not \U$5801 ( \5894 , \5887 );
not \U$5802 ( \5895 , \5894 );
not \U$5803 ( \5896 , \5890 );
or \U$5804 ( \5897 , \5895 , \5896 );
xor \U$5805 ( \5898 , \5695 , \5704 );
xor \U$5806 ( \5899 , \5898 , \5715 );
nand \U$5807 ( \5900 , \5897 , \5899 );
nand \U$5808 ( \5901 , \5893 , \5900 );
not \U$5809 ( \5902 , \5901 );
not \U$5810 ( \5903 , \5902 );
or \U$5811 ( \5904 , \5882 , \5903 );
not \U$5812 ( \5905 , \5901 );
not \U$5813 ( \5906 , \5880 );
or \U$5814 ( \5907 , \5905 , \5906 );
not \U$5815 ( \5908 , \5614 );
not \U$5816 ( \5909 , \5612 );
or \U$5817 ( \5910 , \5908 , \5909 );
nand \U$5818 ( \5911 , \5910 , \5616 );
and \U$5819 ( \5912 , \5911 , \5609 );
not \U$5820 ( \5913 , \5911 );
and \U$5821 ( \5914 , \5913 , \5610 );
nor \U$5822 ( \5915 , \5912 , \5914 );
buf \U$5823 ( \5916 , \5915 );
nand \U$5824 ( \5917 , \5907 , \5916 );
nand \U$5825 ( \5918 , \5904 , \5917 );
xor \U$5826 ( \5919 , \5564 , \5562 );
nor \U$5827 ( \5920 , \5918 , \5919 );
nand \U$5828 ( \5921 , \5726 , \5622 );
buf \U$5829 ( \5922 , \5721 );
xor \U$5830 ( \5923 , \5921 , \5922 );
or \U$5831 ( \5924 , \5920 , \5923 );
nand \U$5832 ( \5925 , \5918 , \5919 );
nand \U$5833 ( \5926 , \5924 , \5925 );
nand \U$5834 ( \5927 , \5752 , \5926 );
nand \U$5835 ( \5928 , \5746 , \5927 );
nor \U$5836 ( \5929 , \5504 , \5928 );
not \U$5837 ( \5930 , \5929 );
xor \U$5838 ( \5931 , \5919 , \5918 );
xnor \U$5839 ( \5932 , \5931 , \5923 );
xor \U$5840 ( \5933 , \5718 , \5637 );
xor \U$5841 ( \5934 , \5933 , \5633 );
not \U$5842 ( \5935 , \5934 );
xor \U$5843 ( \5936 , \5818 , \5792 );
not \U$5844 ( \5937 , \5838 );
and \U$5845 ( \5938 , \5388 , \5937 );
not \U$5846 ( \5939 , \5388 );
and \U$5847 ( \5940 , \5939 , \5839 );
nor \U$5848 ( \5941 , \5938 , \5940 );
not \U$5849 ( \5942 , \5941 );
not \U$5850 ( \5943 , \3814 );
or \U$5851 ( \5944 , \5942 , \5943 );
nand \U$5852 ( \5945 , \3833 , \5753 );
nand \U$5853 ( \5946 , \5944 , \5945 );
not \U$5854 ( \5947 , \5946 );
buf \U$5855 ( \5948 , \5801 );
and \U$5856 ( \5949 , \3976 , \5948 );
and \U$5857 ( \5950 , \3127 , \5235 );
not \U$5858 ( \5951 , \3127 );
and \U$5859 ( \5952 , \5951 , \5232 );
nor \U$5860 ( \5953 , \5950 , \5952 );
not \U$5861 ( \5954 , \5953 );
and \U$5862 ( \5955 , \4377 , \5954 );
nor \U$5863 ( \5956 , \5949 , \5955 );
not \U$5864 ( \5957 , \5956 );
not \U$5865 ( \5958 , \4793 );
not \U$5866 ( \5959 , \3983 );
or \U$5867 ( \5960 , \5958 , \5959 );
or \U$5868 ( \5961 , \4137 , \4793 );
nand \U$5869 ( \5962 , \5960 , \5961 );
not \U$5870 ( \5963 , \5962 );
not \U$5871 ( \5964 , \4391 );
or \U$5872 ( \5965 , \5963 , \5964 );
nand \U$5873 ( \5966 , \4134 , \5764 );
nand \U$5874 ( \5967 , \5965 , \5966 );
not \U$5875 ( \5968 , \5967 );
or \U$5876 ( \5969 , \5957 , \5968 );
or \U$5877 ( \5970 , \5967 , \5956 );
nand \U$5878 ( \5971 , \5969 , \5970 );
not \U$5879 ( \5972 , \5971 );
or \U$5880 ( \5973 , \5947 , \5972 );
not \U$5881 ( \5974 , \5956 );
nand \U$5882 ( \5975 , \5974 , \5967 );
nand \U$5883 ( \5976 , \5973 , \5975 );
xor \U$5884 ( \5977 , \5936 , \5976 );
xor \U$5885 ( \5978 , \5779 , \5769 );
xor \U$5886 ( \5979 , \5978 , \5759 );
and \U$5887 ( \5980 , \5977 , \5979 );
and \U$5888 ( \5981 , \5936 , \5976 );
or \U$5889 ( \5982 , \5980 , \5981 );
not \U$5890 ( \5983 , \5982 );
not \U$5891 ( \5984 , \4695 );
not \U$5892 ( \5985 , \5858 );
and \U$5893 ( \5986 , \5984 , \5985 );
and \U$5894 ( \5987 , \4178 , \4698 );
not \U$5895 ( \5988 , \4178 );
and \U$5896 ( \5989 , \5988 , \5545 );
or \U$5897 ( \5990 , \5987 , \5989 );
and \U$5898 ( \5991 , \5990 , \4711 );
nor \U$5899 ( \5992 , \5986 , \5991 );
not \U$5900 ( \5993 , \5992 );
not \U$5901 ( \5994 , \5993 );
not \U$5902 ( \5995 , \3843 );
not \U$5903 ( \5996 , \4181 );
or \U$5904 ( \5997 , \5995 , \5996 );
or \U$5905 ( \5998 , \4278 , \3843 );
nand \U$5906 ( \5999 , \5997 , \5998 );
not \U$5907 ( \6000 , \5999 );
not \U$5908 ( \6001 , \4354 );
or \U$5909 ( \6002 , \6000 , \6001 );
nand \U$5910 ( \6003 , \5808 , \4271 );
nand \U$5911 ( \6004 , \6002 , \6003 );
not \U$5912 ( \6005 , \6004 );
or \U$5913 ( \6006 , \5994 , \6005 );
not \U$5914 ( \6007 , \5992 );
not \U$5915 ( \6008 , \6004 );
not \U$5916 ( \6009 , \6008 );
or \U$5917 ( \6010 , \6007 , \6009 );
not \U$5918 ( \6011 , \3151 );
not \U$5919 ( \6012 , \1727 );
or \U$5920 ( \6013 , \6011 , \6012 );
or \U$5921 ( \6014 , \1727 , \3151 );
nand \U$5922 ( \6015 , \6013 , \6014 );
not \U$5923 ( \6016 , \6015 );
not \U$5924 ( \6017 , \1719 );
or \U$5925 ( \6018 , \6016 , \6017 );
nand \U$5926 ( \6019 , \4161 , \5787 );
nand \U$5927 ( \6020 , \6018 , \6019 );
nand \U$5928 ( \6021 , \6010 , \6020 );
nand \U$5929 ( \6022 , \6006 , \6021 );
not \U$5930 ( \6023 , \6022 );
not \U$5931 ( \6024 , \3825 );
not \U$5932 ( \6025 , \3808 );
or \U$5933 ( \6026 , \6024 , \6025 );
nand \U$5934 ( \6027 , \6026 , \5842 );
and \U$5935 ( \6028 , \6027 , \3755 , \3830 );
not \U$5936 ( \6029 , \5683 );
not \U$5937 ( \6030 , \4151 );
buf \U$5938 ( \6031 , \5686 );
not \U$5939 ( \6032 , \6031 );
or \U$5940 ( \6033 , \6030 , \6032 );
or \U$5941 ( \6034 , \6031 , \4151 );
nand \U$5942 ( \6035 , \6033 , \6034 );
not \U$5943 ( \6036 , \6035 );
or \U$5944 ( \6037 , \6029 , \6036 );
nand \U$5945 ( \6038 , \5693 , \5830 );
nand \U$5946 ( \6039 , \6037 , \6038 );
nand \U$5947 ( \6040 , \6028 , \6039 );
buf \U$5948 ( \6041 , \6040 );
not \U$5949 ( \6042 , \6041 );
xor \U$5950 ( \6043 , \5834 , \5843 );
xnor \U$5951 ( \6044 , \6043 , \5862 );
not \U$5952 ( \6045 , \6044 );
or \U$5953 ( \6046 , \6042 , \6045 );
or \U$5954 ( \6047 , \6044 , \6041 );
nand \U$5955 ( \6048 , \6046 , \6047 );
not \U$5956 ( \6049 , \6048 );
or \U$5957 ( \6050 , \6023 , \6049 );
not \U$5958 ( \6051 , \6041 );
nand \U$5959 ( \6052 , \6051 , \6044 );
nand \U$5960 ( \6053 , \6050 , \6052 );
not \U$5961 ( \6054 , \5873 );
not \U$5962 ( \6055 , \5782 );
not \U$5963 ( \6056 , \6055 );
and \U$5964 ( \6057 , \6054 , \6056 );
and \U$5965 ( \6058 , \5873 , \6055 );
nor \U$5966 ( \6059 , \6057 , \6058 );
xnor \U$5967 ( \6060 , \6053 , \6059 );
not \U$5968 ( \6061 , \6060 );
or \U$5969 ( \6062 , \5983 , \6061 );
not \U$5970 ( \6063 , \6059 );
nand \U$5971 ( \6064 , \6063 , \6053 );
nand \U$5972 ( \6065 , \6062 , \6064 );
not \U$5973 ( \6066 , \6065 );
or \U$5974 ( \6067 , \5935 , \6066 );
not \U$5975 ( \6068 , \5880 );
not \U$5976 ( \6069 , \5915 );
or \U$5977 ( \6070 , \6068 , \6069 );
or \U$5978 ( \6071 , \5880 , \5915 );
nand \U$5979 ( \6072 , \6070 , \6071 );
and \U$5980 ( \6073 , \6072 , \5901 );
not \U$5981 ( \6074 , \6072 );
and \U$5982 ( \6075 , \6074 , \5902 );
nor \U$5983 ( \6076 , \6073 , \6075 );
not \U$5984 ( \6077 , \6076 );
nand \U$5985 ( \6078 , \6067 , \6077 );
or \U$5986 ( \6079 , \6065 , \5934 );
nand \U$5987 ( \6080 , \6078 , \6079 );
nand \U$5988 ( \6081 , \5932 , \6080 );
xor \U$5989 ( \6082 , \5934 , \6076 );
xnor \U$5990 ( \6083 , \6082 , \6065 );
xor \U$5991 ( \6084 , \5887 , \5899 );
xnor \U$5992 ( \6085 , \6084 , \5891 );
buf \U$5993 ( \6086 , \6085 );
not \U$5994 ( \6087 , \6086 );
xor \U$5995 ( \6088 , \6053 , \6059 );
xor \U$5996 ( \6089 , \6088 , \5982 );
not \U$5997 ( \6090 , \6089 );
or \U$5998 ( \6091 , \6087 , \6090 );
or \U$5999 ( \6092 , \6089 , \6086 );
xor \U$6000 ( \6093 , \5936 , \5976 );
xor \U$6001 ( \6094 , \6093 , \5979 );
not \U$6002 ( \6095 , \6094 );
xor \U$6003 ( \6096 , \6040 , \6022 );
xnor \U$6004 ( \6097 , \6096 , \6044 );
not \U$6005 ( \6098 , \4274 );
not \U$6006 ( \6099 , \6031 );
or \U$6007 ( \6100 , \6098 , \6099 );
or \U$6008 ( \6101 , \4274 , \5411 );
nand \U$6009 ( \6102 , \6100 , \6101 );
not \U$6010 ( \6103 , \6102 );
not \U$6011 ( \6104 , \5684 );
or \U$6012 ( \6105 , \6103 , \6104 );
nand \U$6013 ( \6106 , \6035 , \5693 );
nand \U$6014 ( \6107 , \6105 , \6106 );
buf \U$6015 ( \6108 , \6107 );
not \U$6016 ( \6109 , \6108 );
nor \U$6017 ( \6110 , \4309 , \5937 );
not \U$6018 ( \6111 , \6110 );
or \U$6019 ( \6112 , \6109 , \6111 );
or \U$6020 ( \6113 , \6108 , \6110 );
and \U$6021 ( \6114 , \2803 , \5545 );
not \U$6022 ( \6115 , \2803 );
and \U$6023 ( \6116 , \6115 , \4700 );
nor \U$6024 ( \6117 , \6114 , \6116 );
not \U$6025 ( \6118 , \6117 );
not \U$6026 ( \6119 , \4711 );
or \U$6027 ( \6120 , \6118 , \6119 );
not \U$6028 ( \6121 , \4695 );
nand \U$6029 ( \6122 , \6121 , \5990 );
nand \U$6030 ( \6123 , \6120 , \6122 );
nand \U$6031 ( \6124 , \6113 , \6123 );
nand \U$6032 ( \6125 , \6112 , \6124 );
not \U$6033 ( \6126 , \6125 );
xor \U$6034 ( \6127 , \6039 , \6028 );
not \U$6035 ( \6128 , \3115 );
not \U$6036 ( \6129 , \5363 );
and \U$6037 ( \6130 , \6128 , \6129 );
and \U$6038 ( \6131 , \4334 , \5363 );
nor \U$6039 ( \6132 , \6130 , \6131 );
not \U$6040 ( \6133 , \6132 );
not \U$6041 ( \6134 , \3140 );
or \U$6042 ( \6135 , \6133 , \6134 );
nand \U$6043 ( \6136 , \2799 , \5774 );
nand \U$6044 ( \6137 , \6135 , \6136 );
not \U$6045 ( \6138 , \6137 );
xnor \U$6046 ( \6139 , \6127 , \6138 );
not \U$6047 ( \6140 , \6139 );
or \U$6048 ( \6141 , \6126 , \6140 );
not \U$6049 ( \6142 , \6138 );
xor \U$6050 ( \6143 , \6039 , \6028 );
nand \U$6051 ( \6144 , \6142 , \6143 );
nand \U$6052 ( \6145 , \6141 , \6144 );
and \U$6053 ( \6146 , \6097 , \6145 );
not \U$6054 ( \6147 , \6097 );
not \U$6055 ( \6148 , \6145 );
and \U$6056 ( \6149 , \6147 , \6148 );
nor \U$6057 ( \6150 , \6146 , \6149 );
not \U$6058 ( \6151 , \6150 );
or \U$6059 ( \6152 , \6095 , \6151 );
nand \U$6060 ( \6153 , \6097 , \6145 );
nand \U$6061 ( \6154 , \6152 , \6153 );
not \U$6062 ( \6155 , \6154 );
nand \U$6063 ( \6156 , \6092 , \6155 );
nand \U$6064 ( \6157 , \6091 , \6156 );
nand \U$6065 ( \6158 , \6083 , \6157 );
and \U$6066 ( \6159 , \6081 , \6158 );
xor \U$6067 ( \6160 , \6085 , \6155 );
xnor \U$6068 ( \6161 , \6160 , \6089 );
xnor \U$6069 ( \6162 , \6139 , \6125 );
not \U$6070 ( \6163 , \6162 );
not \U$6071 ( \6164 , \6163 );
not \U$6072 ( \6165 , \3108 );
not \U$6073 ( \6166 , \5598 );
and \U$6074 ( \6167 , \6165 , \6166 );
and \U$6075 ( \6168 , \3114 , \5598 );
nor \U$6076 ( \6169 , \6167 , \6168 );
not \U$6077 ( \6170 , \6169 );
not \U$6078 ( \6171 , \6170 );
not \U$6079 ( \6172 , \3142 );
or \U$6080 ( \6173 , \6171 , \6172 );
nand \U$6081 ( \6174 , \2801 , \6132 );
nand \U$6082 ( \6175 , \6173 , \6174 );
not \U$6083 ( \6176 , \6175 );
not \U$6084 ( \6177 , \5684 );
not \U$6085 ( \6178 , \4178 );
not \U$6086 ( \6179 , \4621 );
not \U$6087 ( \6180 , \6179 );
buf \U$6088 ( \6181 , \6180 );
not \U$6089 ( \6182 , \6181 );
or \U$6090 ( \6183 , \6178 , \6182 );
or \U$6091 ( \6184 , \6181 , \4178 );
nand \U$6092 ( \6185 , \6183 , \6184 );
not \U$6093 ( \6186 , \6185 );
or \U$6094 ( \6187 , \6177 , \6186 );
nand \U$6095 ( \6188 , \6102 , \5693 );
nand \U$6096 ( \6189 , \6187 , \6188 );
not \U$6097 ( \6190 , \5837 );
not \U$6098 ( \6191 , \6190 );
not \U$6099 ( \6192 , \3983 );
not \U$6100 ( \6193 , \6192 );
or \U$6101 ( \6194 , \6191 , \6193 );
not \U$6102 ( \6195 , \2745 );
nand \U$6103 ( \6196 , \6194 , \6195 );
nand \U$6104 ( \6197 , \3983 , \5837 );
and \U$6105 ( \6198 , \6196 , \4334 , \6197 );
nand \U$6106 ( \6199 , \6189 , \6198 );
not \U$6107 ( \6200 , \4134 );
or \U$6108 ( \6201 , \6200 , \5962 );
not \U$6109 ( \6202 , \4129 );
not \U$6110 ( \6203 , \5265 );
not \U$6111 ( \6204 , \6192 );
or \U$6112 ( \6205 , \6203 , \6204 );
or \U$6113 ( \6206 , \3987 , \5265 );
nand \U$6114 ( \6207 , \6205 , \6206 );
not \U$6115 ( \6208 , \6207 );
or \U$6116 ( \6209 , \6202 , \6208 );
nand \U$6117 ( \6210 , \6209 , \4814 );
nand \U$6118 ( \6211 , \6201 , \6210 );
xor \U$6119 ( \6212 , \6199 , \6211 );
and \U$6120 ( \6213 , \6176 , \6212 );
and \U$6121 ( \6214 , \6199 , \6211 );
nor \U$6122 ( \6215 , \6213 , \6214 );
not \U$6123 ( \6216 , \6215 );
or \U$6124 ( \6217 , \6164 , \6216 );
not \U$6125 ( \6218 , \6215 );
not \U$6126 ( \6219 , \6218 );
not \U$6127 ( \6220 , \6162 );
or \U$6128 ( \6221 , \6219 , \6220 );
not \U$6129 ( \6222 , \4793 );
not \U$6130 ( \6223 , \4775 );
not \U$6131 ( \6224 , \6223 );
not \U$6132 ( \6225 , \6224 );
or \U$6133 ( \6226 , \6222 , \6225 );
or \U$6134 ( \6227 , \6224 , \4793 );
nand \U$6135 ( \6228 , \6226 , \6227 );
not \U$6136 ( \6229 , \6228 );
not \U$6137 ( \6230 , \4772 );
or \U$6138 ( \6231 , \6229 , \6230 );
xor \U$6139 ( \6232 , \4327 , \4277 );
nand \U$6140 ( \6233 , \4271 , \6232 );
nand \U$6141 ( \6234 , \6231 , \6233 );
not \U$6142 ( \6235 , \3843 );
not \U$6143 ( \6236 , \1727 );
or \U$6144 ( \6237 , \6235 , \6236 );
or \U$6145 ( \6238 , \4167 , \3843 );
nand \U$6146 ( \6239 , \6237 , \6238 );
not \U$6147 ( \6240 , \6239 );
not \U$6148 ( \6241 , \1719 );
or \U$6149 ( \6242 , \6240 , \6241 );
not \U$6150 ( \6243 , \4315 );
not \U$6151 ( \6244 , \1562 );
or \U$6152 ( \6245 , \6243 , \6244 );
or \U$6153 ( \6246 , \1562 , \4315 );
nand \U$6154 ( \6247 , \6245 , \6246 );
nand \U$6155 ( \6248 , \6247 , \4161 );
nand \U$6156 ( \6249 , \6242 , \6248 );
xor \U$6157 ( \6250 , \6234 , \6249 );
not \U$6158 ( \6251 , \4698 );
not \U$6159 ( \6252 , \3127 );
and \U$6160 ( \6253 , \6251 , \6252 );
buf \U$6161 ( \6254 , \4698 );
and \U$6162 ( \6255 , \6254 , \3127 );
nor \U$6163 ( \6256 , \6253 , \6255 );
not \U$6164 ( \6257 , \6256 );
not \U$6165 ( \6258 , \6257 );
not \U$6166 ( \6259 , \4711 );
or \U$6167 ( \6260 , \6258 , \6259 );
nand \U$6168 ( \6261 , \4696 , \6117 );
nand \U$6169 ( \6262 , \6260 , \6261 );
and \U$6170 ( \6263 , \6250 , \6262 );
and \U$6171 ( \6264 , \6234 , \6249 );
or \U$6172 ( \6265 , \6263 , \6264 );
not \U$6173 ( \6266 , \6265 );
not \U$6174 ( \6267 , \6266 );
not \U$6175 ( \6268 , \4267 );
not \U$6176 ( \6269 , \6232 );
or \U$6177 ( \6270 , \6268 , \6269 );
nand \U$6178 ( \6271 , \5999 , \4271 );
nand \U$6179 ( \6272 , \6270 , \6271 );
not \U$6180 ( \6273 , \6247 );
not \U$6181 ( \6274 , \1719 );
or \U$6182 ( \6275 , \6273 , \6274 );
nand \U$6183 ( \6276 , \6015 , \4161 );
nand \U$6184 ( \6277 , \6275 , \6276 );
xor \U$6185 ( \6278 , \6272 , \6277 );
not \U$6186 ( \6279 , \3822 );
not \U$6187 ( \6280 , \5235 );
or \U$6188 ( \6281 , \6279 , \6280 );
or \U$6189 ( \6282 , \5235 , \3822 );
nand \U$6190 ( \6283 , \6281 , \6282 );
not \U$6191 ( \6284 , \6283 );
not \U$6192 ( \6285 , \3967 );
or \U$6193 ( \6286 , \6284 , \6285 );
not \U$6194 ( \6287 , \5953 );
nand \U$6195 ( \6288 , \6287 , \3976 );
nand \U$6196 ( \6289 , \6286 , \6288 );
xor \U$6197 ( \6290 , \6278 , \6289 );
not \U$6198 ( \6291 , \6290 );
not \U$6199 ( \6292 , \6291 );
or \U$6200 ( \6293 , \6267 , \6292 );
not \U$6201 ( \6294 , \6265 );
not \U$6202 ( \6295 , \6290 );
or \U$6203 ( \6296 , \6294 , \6295 );
xor \U$6204 ( \6297 , \6107 , \6123 );
xnor \U$6205 ( \6298 , \6297 , \6110 );
nand \U$6206 ( \6299 , \6296 , \6298 );
nand \U$6207 ( \6300 , \6293 , \6299 );
not \U$6208 ( \6301 , \6300 );
nand \U$6209 ( \6302 , \6221 , \6301 );
nand \U$6210 ( \6303 , \6217 , \6302 );
not \U$6211 ( \6304 , \5946 );
not \U$6212 ( \6305 , \6304 );
buf \U$6213 ( \6306 , \5971 );
not \U$6214 ( \6307 , \6306 );
or \U$6215 ( \6308 , \6305 , \6307 );
or \U$6216 ( \6309 , \6306 , \6304 );
nand \U$6217 ( \6310 , \6308 , \6309 );
not \U$6218 ( \6311 , \6310 );
xor \U$6219 ( \6312 , \6272 , \6277 );
and \U$6220 ( \6313 , \6312 , \6289 );
and \U$6221 ( \6314 , \6272 , \6277 );
or \U$6222 ( \6315 , \6313 , \6314 );
not \U$6223 ( \6316 , \6315 );
and \U$6224 ( \6317 , \5992 , \6008 );
not \U$6225 ( \6318 , \5992 );
and \U$6226 ( \6319 , \6318 , \6004 );
or \U$6227 ( \6320 , \6317 , \6319 );
xor \U$6228 ( \6321 , \6320 , \6020 );
not \U$6229 ( \6322 , \6321 );
or \U$6230 ( \6323 , \6316 , \6322 );
or \U$6231 ( \6324 , \6321 , \6315 );
nand \U$6232 ( \6325 , \6323 , \6324 );
not \U$6233 ( \6326 , \6325 );
or \U$6234 ( \6327 , \6311 , \6326 );
not \U$6235 ( \6328 , \6321 );
nand \U$6236 ( \6329 , \6328 , \6315 );
nand \U$6237 ( \6330 , \6327 , \6329 );
and \U$6238 ( \6331 , \6303 , \6330 );
not \U$6239 ( \6332 , \6303 );
not \U$6240 ( \6333 , \6330 );
and \U$6241 ( \6334 , \6332 , \6333 );
nor \U$6242 ( \6335 , \6331 , \6334 );
not \U$6243 ( \6336 , \6335 );
not \U$6244 ( \6337 , \6150 );
not \U$6245 ( \6338 , \6094 );
not \U$6246 ( \6339 , \6338 );
or \U$6247 ( \6340 , \6337 , \6339 );
or \U$6248 ( \6341 , \6338 , \6150 );
nand \U$6249 ( \6342 , \6340 , \6341 );
not \U$6250 ( \6343 , \6342 );
or \U$6251 ( \6344 , \6336 , \6343 );
nand \U$6252 ( \6345 , \6303 , \6330 );
nand \U$6253 ( \6346 , \6344 , \6345 );
nand \U$6254 ( \6347 , \6161 , \6346 );
not \U$6255 ( \6348 , \6310 );
not \U$6256 ( \6349 , \6325 );
or \U$6257 ( \6350 , \6348 , \6349 );
or \U$6258 ( \6351 , \6325 , \6310 );
nand \U$6259 ( \6352 , \6350 , \6351 );
not \U$6260 ( \6353 , \6352 );
xor \U$6261 ( \6354 , \6215 , \6300 );
xnor \U$6262 ( \6355 , \6354 , \6162 );
not \U$6263 ( \6356 , \6355 );
or \U$6264 ( \6357 , \6353 , \6356 );
not \U$6265 ( \6358 , \5362 );
not \U$6266 ( \6359 , \4137 );
or \U$6267 ( \6360 , \6358 , \6359 );
or \U$6268 ( \6361 , \4396 , \5362 );
nand \U$6269 ( \6362 , \6360 , \6361 );
not \U$6270 ( \6363 , \6362 );
not \U$6271 ( \6364 , \4131 );
or \U$6272 ( \6365 , \6363 , \6364 );
nand \U$6273 ( \6366 , \5287 , \6207 );
nand \U$6274 ( \6367 , \6365 , \6366 );
not \U$6275 ( \6368 , \6367 );
buf \U$6276 ( \6369 , \2798 );
or \U$6277 ( \6370 , \6169 , \6369 );
buf \U$6278 ( \6371 , \5837 );
and \U$6279 ( \6372 , \6371 , \4332 );
not \U$6280 ( \6373 , \6371 );
not \U$6281 ( \6374 , \4332 );
and \U$6282 ( \6375 , \6373 , \6374 );
nor \U$6283 ( \6376 , \6372 , \6375 );
nor \U$6284 ( \6377 , \6376 , \3137 );
nand \U$6285 ( \6378 , \6369 , \6377 );
nand \U$6286 ( \6379 , \6370 , \6378 );
not \U$6287 ( \6380 , \6379 );
not \U$6288 ( \6381 , \3151 );
not \U$6289 ( \6382 , \5235 );
or \U$6290 ( \6383 , \6381 , \6382 );
or \U$6291 ( \6384 , \5235 , \3151 );
nand \U$6292 ( \6385 , \6383 , \6384 );
not \U$6293 ( \6386 , \6385 );
not \U$6294 ( \6387 , \3967 );
or \U$6295 ( \6388 , \6386 , \6387 );
nand \U$6296 ( \6389 , \4373 , \6283 );
nand \U$6297 ( \6390 , \6388 , \6389 );
not \U$6298 ( \6391 , \6390 );
not \U$6299 ( \6392 , \6391 );
or \U$6300 ( \6393 , \6380 , \6392 );
not \U$6301 ( \6394 , \6379 );
nand \U$6302 ( \6395 , \6390 , \6394 );
nand \U$6303 ( \6396 , \6393 , \6395 );
not \U$6304 ( \6397 , \6396 );
or \U$6305 ( \6398 , \6368 , \6397 );
nand \U$6306 ( \6399 , \6390 , \6379 );
nand \U$6307 ( \6400 , \6398 , \6399 );
not \U$6308 ( \6401 , \6400 );
not \U$6309 ( \6402 , \6175 );
not \U$6310 ( \6403 , \6212 );
or \U$6311 ( \6404 , \6402 , \6403 );
or \U$6312 ( \6405 , \6212 , \6175 );
nand \U$6313 ( \6406 , \6404 , \6405 );
buf \U$6314 ( \6407 , \6406 );
nand \U$6315 ( \6408 , \6401 , \6407 );
not \U$6316 ( \6409 , \6408 );
not \U$6317 ( \6410 , \4772 );
not \U$6318 ( \6411 , \6410 );
not \U$6319 ( \6412 , \4181 );
not \U$6320 ( \6413 , \5264 );
and \U$6321 ( \6414 , \6412 , \6413 );
and \U$6322 ( \6415 , \6224 , \5264 );
nor \U$6323 ( \6416 , \6414 , \6415 );
not \U$6324 ( \6417 , \6416 );
and \U$6325 ( \6418 , \6411 , \6417 );
and \U$6326 ( \6419 , \6228 , \4271 );
nor \U$6327 ( \6420 , \6418 , \6419 );
not \U$6328 ( \6421 , \6420 );
not \U$6329 ( \6422 , \4315 );
not \U$6330 ( \6423 , \5235 );
or \U$6331 ( \6424 , \6422 , \6423 );
or \U$6332 ( \6425 , \3977 , \4315 );
nand \U$6333 ( \6426 , \6424 , \6425 );
not \U$6334 ( \6427 , \6426 );
not \U$6335 ( \6428 , \3967 );
or \U$6336 ( \6429 , \6427 , \6428 );
nand \U$6337 ( \6430 , \3976 , \6385 );
nand \U$6338 ( \6431 , \6429 , \6430 );
or \U$6339 ( \6432 , \6421 , \6431 );
not \U$6340 ( \6433 , \5684 );
not \U$6341 ( \6434 , \2803 );
not \U$6342 ( \6435 , \5411 );
or \U$6343 ( \6436 , \6434 , \6435 );
or \U$6344 ( \6437 , \6181 , \2803 );
nand \U$6345 ( \6438 , \6436 , \6437 );
not \U$6346 ( \6439 , \6438 );
or \U$6347 ( \6440 , \6433 , \6439 );
nand \U$6348 ( \6441 , \6185 , \5693 );
nand \U$6349 ( \6442 , \6440 , \6441 );
nand \U$6350 ( \6443 , \6432 , \6442 );
nand \U$6351 ( \6444 , \6431 , \6421 );
nand \U$6352 ( \6445 , \6443 , \6444 );
not \U$6353 ( \6446 , \6445 );
xor \U$6354 ( \6447 , \6198 , \6189 );
not \U$6355 ( \6448 , \6447 );
not \U$6356 ( \6449 , \5937 );
not \U$6357 ( \6450 , \2798 );
nand \U$6358 ( \6451 , \6449 , \6450 );
not \U$6359 ( \6452 , \5850 );
not \U$6360 ( \6453 , \6256 );
and \U$6361 ( \6454 , \6452 , \6453 );
not \U$6362 ( \6455 , \3822 );
not \U$6363 ( \6456 , \6254 );
or \U$6364 ( \6457 , \6455 , \6456 );
or \U$6365 ( \6458 , \6254 , \3822 );
nand \U$6366 ( \6459 , \6457 , \6458 );
and \U$6367 ( \6460 , \4711 , \6459 );
nor \U$6368 ( \6461 , \6454 , \6460 );
xor \U$6369 ( \6462 , \6451 , \6461 );
not \U$6370 ( \6463 , \4327 );
not \U$6371 ( \6464 , \1562 );
or \U$6372 ( \6465 , \6463 , \6464 );
or \U$6373 ( \6466 , \1727 , \4327 );
nand \U$6374 ( \6467 , \6465 , \6466 );
and \U$6375 ( \6468 , \1719 , \6467 );
and \U$6376 ( \6469 , \1722 , \6239 );
nor \U$6377 ( \6470 , \6468 , \6469 );
and \U$6378 ( \6471 , \6462 , \6470 );
and \U$6379 ( \6472 , \6451 , \6461 );
or \U$6380 ( \6473 , \6471 , \6472 );
not \U$6381 ( \6474 , \6473 );
or \U$6382 ( \6475 , \6448 , \6474 );
or \U$6383 ( \6476 , \6473 , \6447 );
nand \U$6384 ( \6477 , \6475 , \6476 );
not \U$6385 ( \6478 , \6477 );
or \U$6386 ( \6479 , \6446 , \6478 );
not \U$6387 ( \6480 , \6473 );
nand \U$6388 ( \6481 , \6480 , \6447 );
nand \U$6389 ( \6482 , \6479 , \6481 );
not \U$6390 ( \6483 , \6482 );
or \U$6391 ( \6484 , \6409 , \6483 );
not \U$6392 ( \6485 , \6407 );
nand \U$6393 ( \6486 , \6485 , \6400 );
nand \U$6394 ( \6487 , \6484 , \6486 );
buf \U$6395 ( \6488 , \6487 );
nand \U$6396 ( \6489 , \6357 , \6488 );
not \U$6397 ( \6490 , \6352 );
not \U$6398 ( \6491 , \6355 );
nand \U$6399 ( \6492 , \6490 , \6491 );
nand \U$6400 ( \6493 , \6489 , \6492 );
not \U$6401 ( \6494 , \6493 );
not \U$6402 ( \6495 , \6494 );
not \U$6403 ( \6496 , \6335 );
nand \U$6404 ( \6497 , \6496 , \6342 );
not \U$6405 ( \6498 , \6342 );
nand \U$6406 ( \6499 , \6498 , \6335 );
nand \U$6407 ( \6500 , \6497 , \6499 );
nand \U$6408 ( \6501 , \6495 , \6500 );
and \U$6409 ( \6502 , \6347 , \6501 );
nor \U$6410 ( \6503 , \6161 , \6346 );
nor \U$6411 ( \6504 , \6502 , \6503 );
and \U$6412 ( \6505 , \6159 , \6504 );
nor \U$6413 ( \6506 , \6083 , \6157 );
not \U$6414 ( \6507 , \6506 );
not \U$6415 ( \6508 , \6081 );
or \U$6416 ( \6509 , \6507 , \6508 );
not \U$6417 ( \6510 , \5932 );
nand \U$6418 ( \6511 , \6510 , \6078 , \6079 );
nand \U$6419 ( \6512 , \6509 , \6511 );
nor \U$6420 ( \6513 , \6505 , \6512 );
not \U$6421 ( \6514 , \6513 );
not \U$6422 ( \6515 , \6514 );
or \U$6423 ( \6516 , \5930 , \6515 );
and \U$6424 ( \6517 , \5927 , \6081 );
and \U$6425 ( \6518 , \5744 , \6158 );
not \U$6426 ( \6519 , \5693 );
not \U$6427 ( \6520 , \3843 );
not \U$6428 ( \6521 , \6179 );
not \U$6429 ( \6522 , \6521 );
or \U$6430 ( \6523 , \6520 , \6522 );
or \U$6431 ( \6524 , \6521 , \3843 );
nand \U$6432 ( \6525 , \6523 , \6524 );
not \U$6433 ( \6526 , \6525 );
or \U$6434 ( \6527 , \6519 , \6526 );
and \U$6435 ( \6528 , \4327 , \6179 );
not \U$6436 ( \6529 , \4327 );
and \U$6437 ( \6530 , \6529 , \5410 );
nor \U$6438 ( \6531 , \6528 , \6530 );
nand \U$6439 ( \6532 , \6531 , \5683 );
nand \U$6440 ( \6533 , \6527 , \6532 );
not \U$6441 ( \6534 , \6533 );
nand \U$6442 ( \6535 , \1722 , \5842 );
not \U$6443 ( \6536 , \6535 );
or \U$6444 ( \6537 , \6534 , \6536 );
or \U$6445 ( \6538 , \6535 , \6533 );
nand \U$6446 ( \6539 , \6537 , \6538 );
xnor \U$6447 ( \6540 , \4793 , \5352 );
not \U$6448 ( \6541 , \6540 );
not \U$6449 ( \6542 , \4696 );
or \U$6450 ( \6543 , \6541 , \6542 );
not \U$6451 ( \6544 , \5264 );
not \U$6452 ( \6545 , \4700 );
or \U$6453 ( \6546 , \6544 , \6545 );
or \U$6454 ( \6547 , \6254 , \5264 );
nand \U$6455 ( \6548 , \6546 , \6547 );
nand \U$6456 ( \6549 , \4711 , \6548 );
nand \U$6457 ( \6550 , \6543 , \6549 );
xor \U$6458 ( \6551 , \6539 , \6550 );
not \U$6459 ( \6552 , \6551 );
not \U$6460 ( \6553 , \5597 );
not \U$6461 ( \6554 , \5235 );
or \U$6462 ( \6555 , \6553 , \6554 );
or \U$6463 ( \6556 , \3977 , \5597 );
nand \U$6464 ( \6557 , \6555 , \6556 );
not \U$6465 ( \6558 , \6557 );
not \U$6466 ( \6559 , \3967 );
or \U$6467 ( \6560 , \6558 , \6559 );
xnor \U$6468 ( \6561 , \5362 , \5235 );
nand \U$6469 ( \6562 , \4373 , \6561 );
nand \U$6470 ( \6563 , \6560 , \6562 );
not \U$6471 ( \6564 , \5693 );
not \U$6472 ( \6565 , \6531 );
or \U$6473 ( \6566 , \6564 , \6565 );
not \U$6474 ( \6567 , \4793 );
not \U$6475 ( \6568 , \4708 );
not \U$6476 ( \6569 , \6568 );
or \U$6477 ( \6570 , \6567 , \6569 );
or \U$6478 ( \6571 , \6180 , \4793 );
nand \U$6479 ( \6572 , \6570 , \6571 );
nand \U$6480 ( \6573 , \6572 , \5824 );
nand \U$6481 ( \6574 , \6566 , \6573 );
nand \U$6482 ( \6575 , \4699 , \6190 );
and \U$6483 ( \6576 , \6575 , \3961 );
not \U$6484 ( \6577 , \5837 );
not \U$6485 ( \6578 , \4698 );
or \U$6486 ( \6579 , \6577 , \6578 );
nand \U$6487 ( \6580 , \6579 , \5235 );
nor \U$6488 ( \6581 , \6576 , \6580 );
nand \U$6489 ( \6582 , \6574 , \6581 );
not \U$6490 ( \6583 , \6582 );
nand \U$6491 ( \6584 , \6563 , \6583 );
not \U$6492 ( \6585 , \6584 );
not \U$6493 ( \6586 , \6585 );
and \U$6494 ( \6587 , \6552 , \6586 );
nor \U$6495 ( \6588 , \6563 , \6583 );
buf \U$6496 ( \6589 , \6588 );
nor \U$6497 ( \6590 , \6587 , \6589 );
not \U$6498 ( \6591 , \5683 );
not \U$6499 ( \6592 , \6525 );
or \U$6500 ( \6593 , \6591 , \6592 );
not \U$6501 ( \6594 , \4315 );
not \U$6502 ( \6595 , \6521 );
or \U$6503 ( \6596 , \6594 , \6595 );
or \U$6504 ( \6597 , \6521 , \4315 );
nand \U$6505 ( \6598 , \6596 , \6597 );
nand \U$6506 ( \6599 , \6598 , \5693 );
nand \U$6507 ( \6600 , \6593 , \6599 );
not \U$6508 ( \6601 , \1708 );
and \U$6509 ( \6602 , \6601 , \5837 );
not \U$6510 ( \6603 , \5235 );
not \U$6511 ( \6604 , \1713 );
or \U$6512 ( \6605 , \6603 , \6604 );
nand \U$6513 ( \6606 , \6605 , \4798 );
nor \U$6514 ( \6607 , \6602 , \6606 );
xor \U$6515 ( \6608 , \6600 , \6607 );
not \U$6516 ( \6609 , \6550 );
not \U$6517 ( \6610 , \6539 );
or \U$6518 ( \6611 , \6609 , \6610 );
not \U$6519 ( \6612 , \6535 );
nand \U$6520 ( \6613 , \6612 , \6533 );
nand \U$6521 ( \6614 , \6611 , \6613 );
xor \U$6522 ( \6615 , \6608 , \6614 );
not \U$6523 ( \6616 , \6561 );
not \U$6524 ( \6617 , \5337 );
or \U$6525 ( \6618 , \6616 , \6617 );
not \U$6526 ( \6619 , \1710 );
not \U$6527 ( \6620 , \5264 );
and \U$6528 ( \6621 , \6619 , \6620 );
and \U$6529 ( \6622 , \5235 , \5264 );
nor \U$6530 ( \6623 , \6621 , \6622 );
not \U$6531 ( \6624 , \6623 );
nand \U$6532 ( \6625 , \6624 , \4763 );
nand \U$6533 ( \6626 , \6618 , \6625 );
and \U$6534 ( \6627 , \4167 , \5838 );
nor \U$6535 ( \6628 , \4170 , \6371 );
nor \U$6536 ( \6629 , \6627 , \6628 );
not \U$6537 ( \6630 , \6629 );
not \U$6538 ( \6631 , \1719 );
or \U$6539 ( \6632 , \6630 , \6631 );
and \U$6540 ( \6633 , \5597 , \1561 );
not \U$6541 ( \6634 , \5597 );
and \U$6542 ( \6635 , \6634 , \1726 );
nor \U$6543 ( \6636 , \6633 , \6635 );
nand \U$6544 ( \6637 , \4161 , \6636 );
nand \U$6545 ( \6638 , \6632 , \6637 );
xor \U$6546 ( \6639 , \6626 , \6638 );
not \U$6547 ( \6640 , \6540 );
not \U$6548 ( \6641 , \4711 );
or \U$6549 ( \6642 , \6640 , \6641 );
not \U$6550 ( \6643 , \4327 );
not \U$6551 ( \6644 , \6254 );
or \U$6552 ( \6645 , \6643 , \6644 );
or \U$6553 ( \6646 , \6254 , \4327 );
nand \U$6554 ( \6647 , \6645 , \6646 );
nand \U$6555 ( \6648 , \4696 , \6647 );
nand \U$6556 ( \6649 , \6642 , \6648 );
xor \U$6557 ( \6650 , \6639 , \6649 );
xor \U$6558 ( \6651 , \6615 , \6650 );
xor \U$6559 ( \6652 , \6590 , \6651 );
not \U$6560 ( \6653 , \3967 );
buf \U$6561 ( \6654 , \5837 );
xor \U$6562 ( \6655 , \6654 , \3977 );
not \U$6563 ( \6656 , \6655 );
or \U$6564 ( \6657 , \6653 , \6656 );
nand \U$6565 ( \6658 , \3976 , \6557 );
nand \U$6566 ( \6659 , \6657 , \6658 );
not \U$6567 ( \6660 , \6659 );
not \U$6568 ( \6661 , \6660 );
not \U$6569 ( \6662 , \5362 );
not \U$6570 ( \6663 , \4698 );
or \U$6571 ( \6664 , \6662 , \6663 );
not \U$6572 ( \6665 , \4712 );
or \U$6573 ( \6666 , \6665 , \5362 );
nand \U$6574 ( \6667 , \6664 , \6666 );
not \U$6575 ( \6668 , \6667 );
not \U$6576 ( \6669 , \4711 );
or \U$6577 ( \6670 , \6668 , \6669 );
nand \U$6578 ( \6671 , \5851 , \6548 );
nand \U$6579 ( \6672 , \6670 , \6671 );
not \U$6580 ( \6673 , \6672 );
nor \U$6581 ( \6674 , \6574 , \6581 );
not \U$6582 ( \6675 , \6674 );
nand \U$6583 ( \6676 , \6675 , \6582 );
xor \U$6584 ( \6677 , \6673 , \6676 );
not \U$6585 ( \6678 , \6677 );
not \U$6586 ( \6679 , \6678 );
or \U$6587 ( \6680 , \6661 , \6679 );
nand \U$6588 ( \6681 , \6677 , \6659 );
nand \U$6589 ( \6682 , \6680 , \6681 );
nand \U$6590 ( \6683 , \4763 , \5838 );
not \U$6591 ( \6684 , \6683 );
not \U$6592 ( \6685 , \5683 );
not \U$6593 ( \6686 , \5264 );
not \U$6594 ( \6687 , \5686 );
or \U$6595 ( \6688 , \6686 , \6687 );
or \U$6596 ( \6689 , \5410 , \5264 );
nand \U$6597 ( \6690 , \6688 , \6689 );
not \U$6598 ( \6691 , \6690 );
or \U$6599 ( \6692 , \6685 , \6691 );
nand \U$6600 ( \6693 , \6572 , \5693 );
nand \U$6601 ( \6694 , \6692 , \6693 );
buf \U$6602 ( \6695 , \6694 );
nand \U$6603 ( \6696 , \6684 , \6695 );
not \U$6604 ( \6697 , \6696 );
not \U$6605 ( \6698 , \5597 );
not \U$6606 ( \6699 , \4713 );
or \U$6607 ( \6700 , \6698 , \6699 );
or \U$6608 ( \6701 , \6665 , \5597 );
nand \U$6609 ( \6702 , \6700 , \6701 );
not \U$6610 ( \6703 , \6702 );
not \U$6611 ( \6704 , \4711 );
or \U$6612 ( \6705 , \6703 , \6704 );
nand \U$6613 ( \6706 , \5851 , \6667 );
nand \U$6614 ( \6707 , \6705 , \6706 );
not \U$6615 ( \6708 , \6707 );
not \U$6616 ( \6709 , \6708 );
or \U$6617 ( \6710 , \6697 , \6709 );
not \U$6618 ( \6711 , \6695 );
nand \U$6619 ( \6712 , \6711 , \6683 );
nand \U$6620 ( \6713 , \6710 , \6712 );
nand \U$6621 ( \6714 , \6682 , \6713 );
not \U$6622 ( \6715 , \6371 );
not \U$6623 ( \6716 , \4699 );
or \U$6624 ( \6717 , \6715 , \6716 );
or \U$6625 ( \6718 , \4701 , \6371 );
nand \U$6626 ( \6719 , \6717 , \6718 );
not \U$6627 ( \6720 , \6719 );
not \U$6628 ( \6721 , \4711 );
or \U$6629 ( \6722 , \6720 , \6721 );
nand \U$6630 ( \6723 , \5851 , \6702 );
nand \U$6631 ( \6724 , \6722 , \6723 );
not \U$6632 ( \6725 , \6724 );
not \U$6633 ( \6726 , \5693 );
not \U$6634 ( \6727 , \6690 );
or \U$6635 ( \6728 , \6726 , \6727 );
not \U$6636 ( \6729 , \5362 );
not \U$6637 ( \6730 , \5686 );
or \U$6638 ( \6731 , \6729 , \6730 );
or \U$6639 ( \6732 , \5410 , \5362 );
nand \U$6640 ( \6733 , \6731 , \6732 );
nand \U$6641 ( \6734 , \6733 , \5824 );
nand \U$6642 ( \6735 , \6728 , \6734 );
buf \U$6643 ( \6736 , \4692 );
and \U$6644 ( \6737 , \6736 , \6654 );
buf \U$6645 ( \6738 , \4693 );
not \U$6646 ( \6739 , \4712 );
nand \U$6647 ( \6740 , \6738 , \6739 );
nor \U$6648 ( \6741 , \6737 , \6740 );
nor \U$6649 ( \6742 , \6735 , \6741 );
not \U$6650 ( \6743 , \6742 );
nand \U$6651 ( \6744 , \6735 , \6741 );
nand \U$6652 ( \6745 , \6743 , \6744 );
nand \U$6653 ( \6746 , \6725 , \6745 );
not \U$6654 ( \6747 , \5693 );
not \U$6655 ( \6748 , \6733 );
or \U$6656 ( \6749 , \6747 , \6748 );
not \U$6657 ( \6750 , \5597 );
not \U$6658 ( \6751 , \6568 );
or \U$6659 ( \6752 , \6750 , \6751 );
or \U$6660 ( \6753 , \5410 , \5597 );
nand \U$6661 ( \6754 , \6752 , \6753 );
nand \U$6662 ( \6755 , \6754 , \5824 );
nand \U$6663 ( \6756 , \6749 , \6755 );
not \U$6664 ( \6757 , \6756 );
nand \U$6665 ( \6758 , \5851 , \5842 );
nand \U$6666 ( \6759 , \6757 , \6758 );
not \U$6667 ( \6760 , \6759 );
not \U$6668 ( \6761 , \5693 );
not \U$6669 ( \6762 , \6754 );
or \U$6670 ( \6763 , \6761 , \6762 );
nand \U$6671 ( \6764 , \5683 , \6190 );
nand \U$6672 ( \6765 , \6763 , \6764 );
nand \U$6673 ( \6766 , \6371 , \5692 );
and \U$6674 ( \6767 , \5411 , \6766 );
nand \U$6675 ( \6768 , \6765 , \6767 );
not \U$6676 ( \6769 , \6768 );
not \U$6677 ( \6770 , \6769 );
or \U$6678 ( \6771 , \6760 , \6770 );
not \U$6679 ( \6772 , \6758 );
nand \U$6680 ( \6773 , \6772 , \6756 );
nand \U$6681 ( \6774 , \6771 , \6773 );
nand \U$6682 ( \6775 , \6746 , \6774 );
not \U$6683 ( \6776 , \6745 );
nand \U$6684 ( \6777 , \6776 , \6724 );
nand \U$6685 ( \6778 , \6775 , \6777 );
not \U$6686 ( \6779 , \6778 );
not \U$6687 ( \6780 , \6707 );
xnor \U$6688 ( \6781 , \6683 , \6694 );
not \U$6689 ( \6782 , \6781 );
or \U$6690 ( \6783 , \6780 , \6782 );
or \U$6691 ( \6784 , \6781 , \6707 );
nand \U$6692 ( \6785 , \6783 , \6784 );
buf \U$6693 ( \6786 , \6744 );
nand \U$6694 ( \6787 , \6785 , \6786 );
not \U$6695 ( \6788 , \6787 );
or \U$6696 ( \6789 , \6779 , \6788 );
not \U$6697 ( \6790 , \6785 );
not \U$6698 ( \6791 , \6786 );
nand \U$6699 ( \6792 , \6790 , \6791 );
nand \U$6700 ( \6793 , \6789 , \6792 );
and \U$6701 ( \6794 , \6714 , \6793 );
nor \U$6702 ( \6795 , \6682 , \6713 );
nor \U$6703 ( \6796 , \6794 , \6795 );
not \U$6704 ( \6797 , \6584 );
nor \U$6705 ( \6798 , \6797 , \6588 );
not \U$6706 ( \6799 , \6798 );
not \U$6707 ( \6800 , \6551 );
and \U$6708 ( \6801 , \6799 , \6800 );
and \U$6709 ( \6802 , \6551 , \6798 );
nor \U$6710 ( \6803 , \6801 , \6802 );
buf \U$6711 ( \6804 , \6677 );
and \U$6712 ( \6805 , \6804 , \6660 );
and \U$6713 ( \6806 , \6673 , \6676 );
nor \U$6714 ( \6807 , \6805 , \6806 );
nor \U$6715 ( \6808 , \6803 , \6807 );
or \U$6716 ( \6809 , \6796 , \6808 );
nand \U$6717 ( \6810 , \6803 , \6807 );
nand \U$6718 ( \6811 , \6809 , \6810 );
and \U$6719 ( \6812 , \6652 , \6811 );
and \U$6720 ( \6813 , \6590 , \6651 );
or \U$6721 ( \6814 , \6812 , \6813 );
not \U$6722 ( \6815 , \5683 );
not \U$6723 ( \6816 , \6598 );
or \U$6724 ( \6817 , \6815 , \6816 );
not \U$6725 ( \6818 , \3151 );
not \U$6726 ( \6819 , \5686 );
or \U$6727 ( \6820 , \6818 , \6819 );
or \U$6728 ( \6821 , \5686 , \3151 );
nand \U$6729 ( \6822 , \6820 , \6821 );
nand \U$6730 ( \6823 , \6822 , \5693 );
nand \U$6731 ( \6824 , \6817 , \6823 );
not \U$6732 ( \6825 , \6824 );
nand \U$6733 ( \6826 , \4271 , \5838 );
nand \U$6734 ( \6827 , \6825 , \6826 );
not \U$6735 ( \6828 , \6827 );
not \U$6736 ( \6829 , \6636 );
not \U$6737 ( \6830 , \1719 );
or \U$6738 ( \6831 , \6829 , \6830 );
and \U$6739 ( \6832 , \5362 , \1726 );
not \U$6740 ( \6833 , \5362 );
and \U$6741 ( \6834 , \6833 , \5248 );
or \U$6742 ( \6835 , \6832 , \6834 );
nand \U$6743 ( \6836 , \4161 , \6835 );
nand \U$6744 ( \6837 , \6831 , \6836 );
not \U$6745 ( \6838 , \6837 );
or \U$6746 ( \6839 , \6828 , \6838 );
not \U$6747 ( \6840 , \6826 );
nand \U$6748 ( \6841 , \6840 , \6824 );
nand \U$6749 ( \6842 , \6839 , \6841 );
not \U$6750 ( \6843 , \6628 );
not \U$6751 ( \6844 , \6371 );
not \U$6752 ( \6845 , \4153 );
or \U$6753 ( \6846 , \6844 , \6845 );
nand \U$6754 ( \6847 , \6846 , \4256 );
nand \U$6755 ( \6848 , \6843 , \6847 );
nand \U$6756 ( \6849 , \4439 , \6848 );
not \U$6757 ( \6850 , \3843 );
not \U$6758 ( \6851 , \4698 );
or \U$6759 ( \6852 , \6850 , \6851 );
or \U$6760 ( \6853 , \4698 , \3843 );
nand \U$6761 ( \6854 , \6852 , \6853 );
not \U$6762 ( \6855 , \6854 );
not \U$6763 ( \6856 , \4711 );
or \U$6764 ( \6857 , \6855 , \6856 );
not \U$6765 ( \6858 , \4315 );
not \U$6766 ( \6859 , \6739 );
or \U$6767 ( \6860 , \6858 , \6859 );
or \U$6768 ( \6861 , \5546 , \4315 );
nand \U$6769 ( \6862 , \6860 , \6861 );
nand \U$6770 ( \6863 , \4696 , \6862 );
nand \U$6771 ( \6864 , \6857 , \6863 );
xor \U$6772 ( \6865 , \6849 , \6864 );
not \U$6773 ( \6866 , \3967 );
not \U$6774 ( \6867 , \6866 );
nand \U$6775 ( \6868 , \5235 , \4793 );
not \U$6776 ( \6869 , \4793 );
nand \U$6777 ( \6870 , \6869 , \5232 );
and \U$6778 ( \6871 , \6868 , \6870 );
not \U$6779 ( \6872 , \6871 );
and \U$6780 ( \6873 , \6867 , \6872 );
not \U$6781 ( \6874 , \3977 );
not \U$6782 ( \6875 , \4327 );
and \U$6783 ( \6876 , \6874 , \6875 );
and \U$6784 ( \6877 , \5235 , \4327 );
nor \U$6785 ( \6878 , \6876 , \6877 );
nor \U$6786 ( \6879 , \4374 , \6878 );
nor \U$6787 ( \6880 , \6873 , \6879 );
xor \U$6788 ( \6881 , \6865 , \6880 );
xor \U$6789 ( \6882 , \6842 , \6881 );
nand \U$6790 ( \6883 , \6600 , \6607 );
not \U$6791 ( \6884 , \6883 );
not \U$6792 ( \6885 , \6623 );
not \U$6793 ( \6886 , \6885 );
not \U$6794 ( \6887 , \3967 );
or \U$6795 ( \6888 , \6886 , \6887 );
not \U$6796 ( \6889 , \6868 );
not \U$6797 ( \6890 , \6870 );
or \U$6798 ( \6891 , \6889 , \6890 );
nand \U$6799 ( \6892 , \6891 , \4373 );
nand \U$6800 ( \6893 , \6888 , \6892 );
nor \U$6801 ( \6894 , \6884 , \6893 );
not \U$6802 ( \6895 , \5850 );
not \U$6803 ( \6896 , \6854 );
not \U$6804 ( \6897 , \6896 );
and \U$6805 ( \6898 , \6895 , \6897 );
and \U$6806 ( \6899 , \4711 , \6647 );
nor \U$6807 ( \6900 , \6898 , \6899 );
or \U$6808 ( \6901 , \6894 , \6900 );
nand \U$6809 ( \6902 , \6893 , \6884 );
nand \U$6810 ( \6903 , \6901 , \6902 );
not \U$6811 ( \6904 , \6903 );
not \U$6812 ( \6905 , \5824 );
not \U$6813 ( \6906 , \6822 );
or \U$6814 ( \6907 , \6905 , \6906 );
not \U$6815 ( \6908 , \3822 );
not \U$6816 ( \6909 , \5686 );
or \U$6817 ( \6910 , \6908 , \6909 );
or \U$6818 ( \6911 , \5410 , \3822 );
nand \U$6819 ( \6912 , \6910 , \6911 );
nand \U$6820 ( \6913 , \6912 , \5693 );
nand \U$6821 ( \6914 , \6907 , \6913 );
not \U$6822 ( \6915 , \6914 );
not \U$6823 ( \6916 , \4116 );
not \U$6824 ( \6917 , \6190 );
and \U$6825 ( \6918 , \6916 , \6917 );
not \U$6826 ( \6919 , \5837 );
and \U$6827 ( \6920 , \5221 , \6919 );
nor \U$6828 ( \6921 , \6918 , \6920 );
nor \U$6829 ( \6922 , \6921 , \5322 );
not \U$6830 ( \6923 , \5597 );
not \U$6831 ( \6924 , \4120 );
or \U$6832 ( \6925 , \6923 , \6924 );
or \U$6833 ( \6926 , \4180 , \5597 );
nand \U$6834 ( \6927 , \6925 , \6926 );
not \U$6835 ( \6928 , \4270 );
nor \U$6836 ( \6929 , \6927 , \6928 );
nor \U$6837 ( \6930 , \6922 , \6929 );
not \U$6838 ( \6931 , \6930 );
or \U$6839 ( \6932 , \6915 , \6931 );
not \U$6840 ( \6933 , \6929 );
not \U$6841 ( \6934 , \6933 );
not \U$6842 ( \6935 , \6921 );
nand \U$6843 ( \6936 , \5323 , \6935 );
not \U$6844 ( \6937 , \6936 );
or \U$6845 ( \6938 , \6934 , \6937 );
not \U$6846 ( \6939 , \6914 );
nand \U$6847 ( \6940 , \6938 , \6939 );
nand \U$6848 ( \6941 , \6932 , \6940 );
not \U$6849 ( \6942 , \6835 );
not \U$6850 ( \6943 , \4146 );
or \U$6851 ( \6944 , \6942 , \6943 );
not \U$6852 ( \6945 , \5264 );
not \U$6853 ( \6946 , \4170 );
or \U$6854 ( \6947 , \6945 , \6946 );
or \U$6855 ( \6948 , \4167 , \5264 );
nand \U$6856 ( \6949 , \6947 , \6948 );
nand \U$6857 ( \6950 , \1722 , \6949 );
nand \U$6858 ( \6951 , \6944 , \6950 );
not \U$6859 ( \6952 , \6951 );
and \U$6860 ( \6953 , \6941 , \6952 );
not \U$6861 ( \6954 , \6941 );
and \U$6862 ( \6955 , \6954 , \6951 );
nor \U$6863 ( \6956 , \6953 , \6955 );
not \U$6864 ( \6957 , \6956 );
and \U$6865 ( \6958 , \6904 , \6957 );
and \U$6866 ( \6959 , \6903 , \6956 );
nor \U$6867 ( \6960 , \6958 , \6959 );
xnor \U$6868 ( \6961 , \6882 , \6960 );
not \U$6869 ( \6962 , \6961 );
xor \U$6870 ( \6963 , \6626 , \6638 );
and \U$6871 ( \6964 , \6963 , \6649 );
and \U$6872 ( \6965 , \6626 , \6638 );
or \U$6873 ( \6966 , \6964 , \6965 );
not \U$6874 ( \6967 , \6966 );
not \U$6875 ( \6968 , \6837 );
not \U$6876 ( \6969 , \6824 );
not \U$6877 ( \6970 , \6826 );
and \U$6878 ( \6971 , \6969 , \6970 );
and \U$6879 ( \6972 , \6824 , \6826 );
nor \U$6880 ( \6973 , \6971 , \6972 );
not \U$6881 ( \6974 , \6973 );
and \U$6882 ( \6975 , \6968 , \6974 );
and \U$6883 ( \6976 , \6837 , \6973 );
nor \U$6884 ( \6977 , \6975 , \6976 );
nand \U$6885 ( \6978 , \6967 , \6977 );
not \U$6886 ( \6979 , \6978 );
not \U$6887 ( \6980 , \6900 );
xor \U$6888 ( \6981 , \6883 , \6980 );
xnor \U$6889 ( \6982 , \6981 , \6893 );
not \U$6890 ( \6983 , \6982 );
or \U$6891 ( \6984 , \6979 , \6983 );
not \U$6892 ( \6985 , \6977 );
nand \U$6893 ( \6986 , \6985 , \6966 );
nand \U$6894 ( \6987 , \6984 , \6986 );
not \U$6895 ( \6988 , \6987 );
nand \U$6896 ( \6989 , \6962 , \6988 );
xor \U$6897 ( \6990 , \6977 , \6967 );
xor \U$6898 ( \6991 , \6990 , \6982 );
not \U$6899 ( \6992 , \6991 );
xor \U$6900 ( \6993 , \6608 , \6614 );
and \U$6901 ( \6994 , \6993 , \6650 );
and \U$6902 ( \6995 , \6608 , \6614 );
or \U$6903 ( \6996 , \6994 , \6995 );
not \U$6904 ( \6997 , \6996 );
nand \U$6905 ( \6998 , \6992 , \6997 );
nand \U$6906 ( \6999 , \6814 , \6989 , \6998 );
not \U$6907 ( \7000 , \6987 );
not \U$6908 ( \7001 , \6961 );
or \U$6909 ( \7002 , \7000 , \7001 );
nand \U$6910 ( \7003 , \6991 , \6996 );
nand \U$6911 ( \7004 , \7002 , \7003 );
nand \U$6912 ( \7005 , \7004 , \6989 );
nand \U$6913 ( \7006 , \6999 , \7005 );
not \U$6914 ( \7007 , \6878 );
not \U$6915 ( \7008 , \7007 );
not \U$6916 ( \7009 , \3967 );
or \U$6917 ( \7010 , \7008 , \7009 );
not \U$6918 ( \7011 , \3843 );
not \U$6919 ( \7012 , \5235 );
or \U$6920 ( \7013 , \7011 , \7012 );
or \U$6921 ( \7014 , \3977 , \3843 );
nand \U$6922 ( \7015 , \7013 , \7014 );
nand \U$6923 ( \7016 , \4375 , \7015 );
nand \U$6924 ( \7017 , \7010 , \7016 );
not \U$6925 ( \7018 , \5362 );
not \U$6926 ( \7019 , \4360 );
or \U$6927 ( \7020 , \7018 , \7019 );
or \U$6928 ( \7021 , \4184 , \5362 );
nand \U$6929 ( \7022 , \7020 , \7021 );
not \U$6930 ( \7023 , \7022 );
not \U$6931 ( \7024 , \4271 );
or \U$6932 ( \7025 , \7023 , \7024 );
not \U$6933 ( \7026 , \6927 );
nand \U$6934 ( \7027 , \7026 , \4267 );
nand \U$6935 ( \7028 , \7025 , \7027 );
not \U$6936 ( \7029 , \6912 );
not \U$6937 ( \7030 , \5684 );
or \U$6938 ( \7031 , \7029 , \7030 );
not \U$6939 ( \7032 , \6181 );
not \U$6940 ( \7033 , \3126 );
and \U$6941 ( \7034 , \7032 , \7033 );
and \U$6942 ( \7035 , \5411 , \3126 );
nor \U$6943 ( \7036 , \7034 , \7035 );
nand \U$6944 ( \7037 , \7036 , \5693 );
nand \U$6945 ( \7038 , \7031 , \7037 );
and \U$6946 ( \7039 , \7028 , \7038 );
not \U$6947 ( \7040 , \7028 );
not \U$6948 ( \7041 , \7038 );
and \U$6949 ( \7042 , \7040 , \7041 );
nor \U$6950 ( \7043 , \7039 , \7042 );
xnor \U$6951 ( \7044 , \7017 , \7043 );
not \U$6952 ( \7045 , \6842 );
not \U$6953 ( \7046 , \6881 );
or \U$6954 ( \7047 , \7045 , \7046 );
not \U$6955 ( \7048 , \6880 );
buf \U$6956 ( \7049 , \6849 );
not \U$6957 ( \7050 , \7049 );
not \U$6958 ( \7051 , \6864 );
or \U$6959 ( \7052 , \7050 , \7051 );
or \U$6960 ( \7053 , \6864 , \7049 );
nand \U$6961 ( \7054 , \7052 , \7053 );
nand \U$6962 ( \7055 , \7048 , \7054 );
nand \U$6963 ( \7056 , \7047 , \7055 );
xor \U$6964 ( \7057 , \7044 , \7056 );
not \U$6965 ( \7058 , \6864 );
nor \U$6966 ( \7059 , \7058 , \7049 );
not \U$6967 ( \7060 , \7059 );
nand \U$6968 ( \7061 , \6941 , \6951 );
not \U$6969 ( \7062 , \6933 );
not \U$6970 ( \7063 , \6936 );
or \U$6971 ( \7064 , \7062 , \7063 );
nand \U$6972 ( \7065 , \7064 , \6914 );
and \U$6973 ( \7066 , \7061 , \7065 );
not \U$6974 ( \7067 , \7066 );
or \U$6975 ( \7068 , \7060 , \7067 );
not \U$6976 ( \7069 , \7065 );
not \U$6977 ( \7070 , \7061 );
or \U$6978 ( \7071 , \7069 , \7070 );
not \U$6979 ( \7072 , \7059 );
nand \U$6980 ( \7073 , \7071 , \7072 );
nand \U$6981 ( \7074 , \7068 , \7073 );
not \U$6982 ( \7075 , \4123 );
nand \U$6983 ( \7076 , \7075 , \5838 );
not \U$6984 ( \7077 , \7076 );
not \U$6985 ( \7078 , \7077 );
and \U$6986 ( \7079 , \4146 , \6949 );
not \U$6987 ( \7080 , \4153 );
not \U$6988 ( \7081 , \4793 );
and \U$6989 ( \7082 , \7080 , \7081 );
and \U$6990 ( \7083 , \4798 , \4793 );
nor \U$6991 ( \7084 , \7082 , \7083 );
nor \U$6992 ( \7085 , \4160 , \7084 );
nor \U$6993 ( \7086 , \7079 , \7085 );
not \U$6994 ( \7087 , \7086 );
or \U$6995 ( \7088 , \7078 , \7087 );
not \U$6996 ( \7089 , \7085 );
not \U$6997 ( \7090 , \7089 );
nand \U$6998 ( \7091 , \4146 , \6949 );
not \U$6999 ( \7092 , \7091 );
or \U$7000 ( \7093 , \7090 , \7092 );
nand \U$7001 ( \7094 , \7093 , \7076 );
nand \U$7002 ( \7095 , \7088 , \7094 );
not \U$7003 ( \7096 , \6862 );
not \U$7004 ( \7097 , \4711 );
or \U$7005 ( \7098 , \7096 , \7097 );
not \U$7006 ( \7099 , \3151 );
not \U$7007 ( \7100 , \5352 );
or \U$7008 ( \7101 , \7099 , \7100 );
or \U$7009 ( \7102 , \4698 , \3151 );
nand \U$7010 ( \7103 , \7101 , \7102 );
nand \U$7011 ( \7104 , \6121 , \7103 );
nand \U$7012 ( \7105 , \7098 , \7104 );
xor \U$7013 ( \7106 , \7095 , \7105 );
and \U$7014 ( \7107 , \7074 , \7106 );
not \U$7015 ( \7108 , \7074 );
not \U$7016 ( \7109 , \7106 );
and \U$7017 ( \7110 , \7108 , \7109 );
nor \U$7018 ( \7111 , \7107 , \7110 );
xnor \U$7019 ( \7112 , \7057 , \7111 );
not \U$7020 ( \7113 , \7112 );
xor \U$7021 ( \7114 , \6881 , \6842 );
not \U$7022 ( \7115 , \6903 );
nand \U$7023 ( \7116 , \7115 , \6956 );
and \U$7024 ( \7117 , \7114 , \7116 );
not \U$7025 ( \7118 , \6903 );
nor \U$7026 ( \7119 , \7118 , \6956 );
nor \U$7027 ( \7120 , \7117 , \7119 );
nand \U$7028 ( \7121 , \7113 , \7120 );
nand \U$7029 ( \7122 , \7006 , \7121 );
not \U$7030 ( \7123 , \7015 );
not \U$7031 ( \7124 , \4377 );
or \U$7032 ( \7125 , \7123 , \7124 );
nand \U$7033 ( \7126 , \3976 , \6426 );
nand \U$7034 ( \7127 , \7125 , \7126 );
not \U$7035 ( \7128 , \6654 );
not \U$7036 ( \7129 , \7128 );
not \U$7037 ( \7130 , \4396 );
or \U$7038 ( \7131 , \7129 , \7130 );
not \U$7039 ( \7132 , \5839 );
or \U$7040 ( \7133 , \4396 , \7132 );
nand \U$7041 ( \7134 , \7131 , \7133 );
not \U$7042 ( \7135 , \7134 );
not \U$7043 ( \7136 , \4131 );
or \U$7044 ( \7137 , \7135 , \7136 );
not \U$7045 ( \7138 , \5597 );
not \U$7046 ( \7139 , \4137 );
or \U$7047 ( \7140 , \7138 , \7139 );
or \U$7048 ( \7141 , \4396 , \5597 );
nand \U$7049 ( \7142 , \7140 , \7141 );
nand \U$7050 ( \7143 , \5287 , \7142 );
nand \U$7051 ( \7144 , \7137 , \7143 );
xor \U$7052 ( \7145 , \7127 , \7144 );
not \U$7053 ( \7146 , \4127 );
not \U$7054 ( \7147 , \4438 );
or \U$7055 ( \7148 , \7146 , \7147 );
nand \U$7056 ( \7149 , \7148 , \5839 );
buf \U$7057 ( \7150 , \4122 );
nand \U$7058 ( \7151 , \7149 , \7150 , \4140 );
not \U$7059 ( \7152 , \7151 );
not \U$7060 ( \7153 , \7103 );
not \U$7061 ( \7154 , \4711 );
or \U$7062 ( \7155 , \7153 , \7154 );
nand \U$7063 ( \7156 , \6121 , \6459 );
nand \U$7064 ( \7157 , \7155 , \7156 );
not \U$7065 ( \7158 , \7157 );
or \U$7066 ( \7159 , \7152 , \7158 );
or \U$7067 ( \7160 , \7157 , \7151 );
nand \U$7068 ( \7161 , \7159 , \7160 );
xor \U$7069 ( \7162 , \7145 , \7161 );
not \U$7070 ( \7163 , \7106 );
not \U$7071 ( \7164 , \7074 );
or \U$7072 ( \7165 , \7163 , \7164 );
not \U$7073 ( \7166 , \7065 );
not \U$7074 ( \7167 , \7061 );
or \U$7075 ( \7168 , \7166 , \7167 );
nand \U$7076 ( \7169 , \7168 , \7059 );
nand \U$7077 ( \7170 , \7165 , \7169 );
xor \U$7078 ( \7171 , \7162 , \7170 );
not \U$7079 ( \7172 , \7028 );
nand \U$7080 ( \7173 , \7172 , \7041 );
and \U$7081 ( \7174 , \7017 , \7173 );
nor \U$7082 ( \7175 , \7172 , \7041 );
nor \U$7083 ( \7176 , \7174 , \7175 );
not \U$7084 ( \7177 , \7176 );
not \U$7085 ( \7178 , \7177 );
not \U$7086 ( \7179 , \7105 );
not \U$7087 ( \7180 , \7095 );
or \U$7088 ( \7181 , \7179 , \7180 );
not \U$7089 ( \7182 , \7089 );
not \U$7090 ( \7183 , \7091 );
or \U$7091 ( \7184 , \7182 , \7183 );
nand \U$7092 ( \7185 , \7184 , \7077 );
nand \U$7093 ( \7186 , \7181 , \7185 );
not \U$7094 ( \7187 , \7186 );
not \U$7095 ( \7188 , \7187 );
or \U$7096 ( \7189 , \7178 , \7188 );
nand \U$7097 ( \7190 , \7186 , \7176 );
nand \U$7098 ( \7191 , \7189 , \7190 );
not \U$7099 ( \7192 , \5684 );
not \U$7100 ( \7193 , \7036 );
or \U$7101 ( \7194 , \7192 , \7193 );
nand \U$7102 ( \7195 , \6438 , \5693 );
nand \U$7103 ( \7196 , \7194 , \7195 );
not \U$7104 ( \7197 , \7022 );
not \U$7105 ( \7198 , \4354 );
or \U$7106 ( \7199 , \7197 , \7198 );
not \U$7107 ( \7200 , \6416 );
nand \U$7108 ( \7201 , \7200 , \4271 );
nand \U$7109 ( \7202 , \7199 , \7201 );
and \U$7110 ( \7203 , \7196 , \7202 );
not \U$7111 ( \7204 , \7196 );
not \U$7112 ( \7205 , \7202 );
and \U$7113 ( \7206 , \7204 , \7205 );
nor \U$7114 ( \7207 , \7203 , \7206 );
not \U$7115 ( \7208 , \7084 );
not \U$7116 ( \7209 , \7208 );
not \U$7117 ( \7210 , \1719 );
or \U$7118 ( \7211 , \7209 , \7210 );
nand \U$7119 ( \7212 , \1724 , \6467 );
nand \U$7120 ( \7213 , \7211 , \7212 );
not \U$7121 ( \7214 , \7213 );
and \U$7122 ( \7215 , \7207 , \7214 );
not \U$7123 ( \7216 , \7207 );
and \U$7124 ( \7217 , \7216 , \7213 );
or \U$7125 ( \7218 , \7215 , \7217 );
and \U$7126 ( \7219 , \7191 , \7218 );
not \U$7127 ( \7220 , \7191 );
not \U$7128 ( \7221 , \7218 );
and \U$7129 ( \7222 , \7220 , \7221 );
nor \U$7130 ( \7223 , \7219 , \7222 );
xnor \U$7131 ( \7224 , \7171 , \7223 );
not \U$7132 ( \7225 , \7044 );
not \U$7133 ( \7226 , \7225 );
not \U$7134 ( \7227 , \7056 );
or \U$7135 ( \7228 , \7226 , \7227 );
not \U$7136 ( \7229 , \7111 );
nand \U$7137 ( \7230 , \7228 , \7229 );
not \U$7138 ( \7231 , \7056 );
nand \U$7139 ( \7232 , \7231 , \7044 );
nand \U$7140 ( \7233 , \7230 , \7232 );
nor \U$7141 ( \7234 , \7224 , \7233 );
not \U$7142 ( \7235 , \7112 );
nor \U$7143 ( \7236 , \7235 , \7120 );
nor \U$7144 ( \7237 , \7234 , \7236 );
nand \U$7145 ( \7238 , \7122 , \7237 );
not \U$7146 ( \7239 , \7213 );
not \U$7147 ( \7240 , \7207 );
or \U$7148 ( \7241 , \7239 , \7240 );
nand \U$7149 ( \7242 , \7202 , \7196 );
nand \U$7150 ( \7243 , \7241 , \7242 );
not \U$7151 ( \7244 , \7243 );
not \U$7152 ( \7245 , \7142 );
not \U$7153 ( \7246 , \4131 );
or \U$7154 ( \7247 , \7245 , \7246 );
nand \U$7155 ( \7248 , \5287 , \6362 );
nand \U$7156 ( \7249 , \7247 , \7248 );
not \U$7157 ( \7250 , \7249 );
not \U$7158 ( \7251 , \7250 );
not \U$7159 ( \7252 , \7151 );
and \U$7160 ( \7253 , \7157 , \7252 );
not \U$7161 ( \7254 , \7253 );
or \U$7162 ( \7255 , \7251 , \7254 );
or \U$7163 ( \7256 , \7253 , \7250 );
nand \U$7164 ( \7257 , \7255 , \7256 );
not \U$7165 ( \7258 , \7257 );
or \U$7166 ( \7259 , \7244 , \7258 );
nand \U$7167 ( \7260 , \7253 , \7249 );
nand \U$7168 ( \7261 , \7259 , \7260 );
not \U$7169 ( \7262 , \7261 );
not \U$7170 ( \7263 , \6367 );
not \U$7171 ( \7264 , \7263 );
not \U$7172 ( \7265 , \6396 );
or \U$7173 ( \7266 , \7264 , \7265 );
or \U$7174 ( \7267 , \6396 , \7263 );
nand \U$7175 ( \7268 , \7266 , \7267 );
xor \U$7176 ( \7269 , \6234 , \6249 );
xor \U$7177 ( \7270 , \7269 , \6262 );
and \U$7178 ( \7271 , \7268 , \7270 );
not \U$7179 ( \7272 , \7268 );
not \U$7180 ( \7273 , \7270 );
and \U$7181 ( \7274 , \7272 , \7273 );
nor \U$7182 ( \7275 , \7271 , \7274 );
not \U$7183 ( \7276 , \7275 );
or \U$7184 ( \7277 , \7262 , \7276 );
or \U$7185 ( \7278 , \7275 , \7261 );
nand \U$7186 ( \7279 , \7277 , \7278 );
not \U$7187 ( \7280 , \7279 );
xor \U$7188 ( \7281 , \6451 , \6461 );
xor \U$7189 ( \7282 , \7281 , \6470 );
not \U$7190 ( \7283 , \7282 );
not \U$7191 ( \7284 , \6420 );
not \U$7192 ( \7285 , \6442 );
and \U$7193 ( \7286 , \7284 , \7285 );
and \U$7194 ( \7287 , \6420 , \6442 );
nor \U$7195 ( \7288 , \7286 , \7287 );
and \U$7196 ( \7289 , \6431 , \7288 );
not \U$7197 ( \7290 , \6431 );
not \U$7198 ( \7291 , \7288 );
and \U$7199 ( \7292 , \7290 , \7291 );
nor \U$7200 ( \7293 , \7289 , \7292 );
not \U$7201 ( \7294 , \7293 );
or \U$7202 ( \7295 , \7283 , \7294 );
xor \U$7203 ( \7296 , \7127 , \7144 );
and \U$7204 ( \7297 , \7296 , \7161 );
and \U$7205 ( \7298 , \7127 , \7144 );
or \U$7206 ( \7299 , \7297 , \7298 );
nand \U$7207 ( \7300 , \7295 , \7299 );
not \U$7208 ( \7301 , \7282 );
not \U$7209 ( \7302 , \7293 );
nand \U$7210 ( \7303 , \7301 , \7302 );
nand \U$7211 ( \7304 , \7300 , \7303 );
not \U$7212 ( \7305 , \7304 );
not \U$7213 ( \7306 , \6477 );
not \U$7214 ( \7307 , \6445 );
not \U$7215 ( \7308 , \7307 );
and \U$7216 ( \7309 , \7306 , \7308 );
and \U$7217 ( \7310 , \6477 , \7307 );
nor \U$7218 ( \7311 , \7309 , \7310 );
not \U$7219 ( \7312 , \7311 );
or \U$7220 ( \7313 , \7305 , \7312 );
or \U$7221 ( \7314 , \7304 , \7311 );
nand \U$7222 ( \7315 , \7313 , \7314 );
not \U$7223 ( \7316 , \7315 );
or \U$7224 ( \7317 , \7280 , \7316 );
or \U$7225 ( \7318 , \7315 , \7279 );
nand \U$7226 ( \7319 , \7317 , \7318 );
xor \U$7227 ( \7320 , \7282 , \7302 );
xnor \U$7228 ( \7321 , \7320 , \7299 );
not \U$7229 ( \7322 , \7321 );
not \U$7230 ( \7323 , \7243 );
not \U$7231 ( \7324 , \7323 );
not \U$7232 ( \7325 , \7257 );
and \U$7233 ( \7326 , \7324 , \7325 );
and \U$7234 ( \7327 , \7323 , \7257 );
nor \U$7235 ( \7328 , \7326 , \7327 );
not \U$7236 ( \7329 , \7328 );
not \U$7237 ( \7330 , \7218 );
not \U$7238 ( \7331 , \7191 );
or \U$7239 ( \7332 , \7330 , \7331 );
nand \U$7240 ( \7333 , \7186 , \7177 );
nand \U$7241 ( \7334 , \7332 , \7333 );
not \U$7242 ( \7335 , \7334 );
or \U$7243 ( \7336 , \7329 , \7335 );
or \U$7244 ( \7337 , \7334 , \7328 );
nand \U$7245 ( \7338 , \7336 , \7337 );
not \U$7246 ( \7339 , \7338 );
or \U$7247 ( \7340 , \7322 , \7339 );
not \U$7248 ( \7341 , \7328 );
nand \U$7249 ( \7342 , \7341 , \7334 );
nand \U$7250 ( \7343 , \7340 , \7342 );
nor \U$7251 ( \7344 , \7319 , \7343 );
not \U$7252 ( \7345 , \7344 );
xor \U$7253 ( \7346 , \7328 , \7334 );
xnor \U$7254 ( \7347 , \7346 , \7321 );
not \U$7255 ( \7348 , \7347 );
not \U$7256 ( \7349 , \7223 );
or \U$7257 ( \7350 , \7162 , \7170 );
not \U$7258 ( \7351 , \7350 );
or \U$7259 ( \7352 , \7349 , \7351 );
nand \U$7260 ( \7353 , \7162 , \7170 );
nand \U$7261 ( \7354 , \7352 , \7353 );
not \U$7262 ( \7355 , \7354 );
nand \U$7263 ( \7356 , \7348 , \7355 );
nand \U$7264 ( \7357 , \7224 , \7233 );
nand \U$7265 ( \7358 , \7238 , \7345 , \7356 , \7357 );
nand \U$7266 ( \7359 , \7347 , \7354 );
nand \U$7267 ( \7360 , \7343 , \7319 );
and \U$7268 ( \7361 , \7359 , \7360 );
nor \U$7269 ( \7362 , \7361 , \7344 );
and \U$7270 ( \7363 , \6298 , \6266 );
not \U$7271 ( \7364 , \6298 );
and \U$7272 ( \7365 , \7364 , \6265 );
nor \U$7273 ( \7366 , \7363 , \7365 );
and \U$7274 ( \7367 , \7366 , \6291 );
not \U$7275 ( \7368 , \7366 );
not \U$7276 ( \7369 , \6291 );
and \U$7277 ( \7370 , \7368 , \7369 );
nor \U$7278 ( \7371 , \7367 , \7370 );
not \U$7279 ( \7372 , \7273 );
not \U$7280 ( \7373 , \7268 );
not \U$7281 ( \7374 , \7373 );
or \U$7282 ( \7375 , \7372 , \7374 );
nand \U$7283 ( \7376 , \7375 , \7261 );
not \U$7284 ( \7377 , \7373 );
nand \U$7285 ( \7378 , \7377 , \7270 );
and \U$7286 ( \7379 , \7376 , \7378 );
xor \U$7287 ( \7380 , \7371 , \7379 );
xor \U$7288 ( \7381 , \6406 , \6400 );
not \U$7289 ( \7382 , \7381 );
not \U$7290 ( \7383 , \6482 );
and \U$7291 ( \7384 , \7382 , \7383 );
and \U$7292 ( \7385 , \6482 , \7381 );
nor \U$7293 ( \7386 , \7384 , \7385 );
xor \U$7294 ( \7387 , \7380 , \7386 );
not \U$7295 ( \7388 , \7311 );
not \U$7296 ( \7389 , \7388 );
not \U$7297 ( \7390 , \7279 );
not \U$7298 ( \7391 , \7390 );
or \U$7299 ( \7392 , \7389 , \7391 );
not \U$7300 ( \7393 , \7304 );
nand \U$7301 ( \7394 , \7392 , \7393 );
nand \U$7302 ( \7395 , \7279 , \7311 );
nand \U$7303 ( \7396 , \7394 , \7395 );
nor \U$7304 ( \7397 , \7387 , \7396 );
nor \U$7305 ( \7398 , \7362 , \7397 );
nand \U$7306 ( \7399 , \7358 , \7398 );
not \U$7307 ( \7400 , \7399 );
nand \U$7308 ( \7401 , \6494 , \6499 , \6497 );
not \U$7309 ( \7402 , \6491 );
not \U$7310 ( \7403 , \6352 );
not \U$7311 ( \7404 , \6487 );
or \U$7312 ( \7405 , \7403 , \7404 );
or \U$7313 ( \7406 , \6487 , \6352 );
nand \U$7314 ( \7407 , \7405 , \7406 );
not \U$7315 ( \7408 , \7407 );
or \U$7316 ( \7409 , \7402 , \7408 );
or \U$7317 ( \7410 , \7407 , \6491 );
nand \U$7318 ( \7411 , \7409 , \7410 );
xor \U$7319 ( \7412 , \7371 , \7379 );
and \U$7320 ( \7413 , \7412 , \7386 );
and \U$7321 ( \7414 , \7371 , \7379 );
or \U$7322 ( \7415 , \7413 , \7414 );
nand \U$7323 ( \7416 , \7411 , \7415 );
nand \U$7324 ( \7417 , \7387 , \7396 );
and \U$7325 ( \7418 , \7401 , \7416 , \7417 );
not \U$7326 ( \7419 , \7418 );
or \U$7327 ( \7420 , \7400 , \7419 );
not \U$7328 ( \7421 , \7411 );
not \U$7329 ( \7422 , \7415 );
nand \U$7330 ( \7423 , \7421 , \7422 );
not \U$7331 ( \7424 , \7423 );
buf \U$7332 ( \7425 , \7401 );
nand \U$7333 ( \7426 , \7424 , \7425 );
nand \U$7334 ( \7427 , \7420 , \7426 );
nor \U$7335 ( \7428 , \5502 , \6503 );
nand \U$7336 ( \7429 , \6517 , \6518 , \7427 , \7428 );
not \U$7337 ( \7430 , \5511 );
not \U$7338 ( \7431 , \5743 );
nand \U$7339 ( \7432 , \7430 , \7431 );
not \U$7340 ( \7433 , \5926 );
nand \U$7341 ( \7434 , \7433 , \5751 );
and \U$7342 ( \7435 , \7432 , \7434 );
nor \U$7343 ( \7436 , \7435 , \5745 );
and \U$7344 ( \7437 , \7436 , \5503 );
nor \U$7345 ( \7438 , \5500 , \5498 );
not \U$7346 ( \7439 , \7438 );
not \U$7347 ( \7440 , \5310 );
or \U$7348 ( \7441 , \7439 , \7440 );
or \U$7349 ( \7442 , \5204 , \5309 );
nand \U$7350 ( \7443 , \7441 , \7442 );
nor \U$7351 ( \7444 , \7437 , \7443 );
nand \U$7352 ( \7445 , \7429 , \7444 );
not \U$7353 ( \7446 , \7445 );
nand \U$7354 ( \7447 , \6516 , \7446 );
not \U$7355 ( \7448 , \7447 );
or \U$7356 ( \7449 , \5194 , \7448 );
not \U$7357 ( \7450 , \5191 );
not \U$7358 ( \7451 , \4935 );
nand \U$7359 ( \7452 , \4547 , \4844 );
or \U$7360 ( \7453 , \7451 , \7452 );
not \U$7361 ( \7454 , \4934 );
nand \U$7362 ( \7455 , \7454 , \4855 );
nand \U$7363 ( \7456 , \7453 , \7455 );
buf \U$7364 ( \7457 , \5006 );
nor \U$7365 ( \7458 , \7457 , \5010 );
nor \U$7366 ( \7459 , \7456 , \7458 );
nand \U$7367 ( \7460 , \5113 , \5155 );
not \U$7368 ( \7461 , \7460 );
nand \U$7369 ( \7462 , \7461 , \5064 , \5011 );
or \U$7370 ( \7463 , \7459 , \7462 );
not \U$7371 ( \7464 , \4948 );
not \U$7372 ( \7465 , \5061 );
or \U$7373 ( \7466 , \7464 , \7465 );
nand \U$7374 ( \7467 , \7466 , \5063 );
nand \U$7375 ( \7468 , \7467 , \5058 );
not \U$7376 ( \7469 , \7468 );
not \U$7377 ( \7470 , \7460 );
and \U$7378 ( \7471 , \7469 , \7470 );
not \U$7379 ( \7472 , \5155 );
nor \U$7380 ( \7473 , \5068 , \5112 );
not \U$7381 ( \7474 , \7473 );
or \U$7382 ( \7475 , \7472 , \7474 );
or \U$7383 ( \7476 , \5154 , \5118 );
nand \U$7384 ( \7477 , \7475 , \7476 );
nor \U$7385 ( \7478 , \7471 , \7477 );
nand \U$7386 ( \7479 , \7463 , \7478 );
and \U$7387 ( \7480 , \7450 , \7479 );
and \U$7388 ( \7481 , \5183 , \5190 );
nor \U$7389 ( \7482 , \7480 , \7481 );
nand \U$7390 ( \7483 , \7449 , \7482 );
and \U$7391 ( \7484 , \4171 , \4974 );
not \U$7392 ( \7485 , \7484 );
and \U$7393 ( \7486 , \4905 , \5164 );
and \U$7394 ( \7487 , \3833 , \4974 );
nor \U$7395 ( \7488 , \7486 , \7487 );
not \U$7396 ( \7489 , \7488 );
or \U$7397 ( \7490 , \7485 , \7489 );
or \U$7398 ( \7491 , \7488 , \7484 );
nand \U$7399 ( \7492 , \7490 , \7491 );
not \U$7400 ( \7493 , \7492 );
xor \U$7401 ( \7494 , \5160 , \5161 );
and \U$7402 ( \7495 , \7494 , \5166 );
and \U$7403 ( \7496 , \5160 , \5161 );
nor \U$7404 ( \7497 , \7495 , \7496 );
not \U$7405 ( \7498 , \7497 );
or \U$7406 ( \7499 , \7493 , \7498 );
or \U$7407 ( \7500 , \7497 , \7492 );
nand \U$7408 ( \7501 , \7499 , \7500 );
not \U$7409 ( \7502 , \7501 );
not \U$7410 ( \7503 , \5179 );
or \U$7411 ( \7504 , \7503 , \5167 );
not \U$7412 ( \7505 , \5169 );
or \U$7413 ( \7506 , \5175 , \7505 );
nand \U$7414 ( \7507 , \7504 , \7506 );
not \U$7415 ( \7508 , \7507 );
or \U$7416 ( \7509 , \7502 , \7508 );
or \U$7417 ( \7510 , \7507 , \7501 );
nand \U$7418 ( \7511 , \7509 , \7510 );
not \U$7419 ( \7512 , \7511 );
and \U$7420 ( \7513 , \7483 , \7512 );
not \U$7421 ( \7514 , \7483 );
and \U$7422 ( \7515 , \7514 , \7511 );
nor \U$7423 ( \7516 , \7513 , \7515 );
buf \U$7424 ( \7517 , \7516 );
and \U$7425 ( \7518 , \5012 , \5064 , \5114 , \5155 );
not \U$7426 ( \7519 , \7518 );
not \U$7427 ( \7520 , \7447 );
or \U$7428 ( \7521 , \7519 , \7520 );
not \U$7429 ( \7522 , \7479 );
nand \U$7430 ( \7523 , \7521 , \7522 );
nor \U$7431 ( \7524 , \7481 , \5191 );
and \U$7432 ( \7525 , \7523 , \7524 );
not \U$7433 ( \7526 , \7523 );
not \U$7434 ( \7527 , \7524 );
and \U$7435 ( \7528 , \7526 , \7527 );
nor \U$7436 ( \7529 , \7525 , \7528 );
buf \U$7437 ( \7530 , \7529 );
and \U$7438 ( \7531 , \5012 , \5064 , \5114 );
not \U$7439 ( \7532 , \7531 );
not \U$7440 ( \7533 , \5929 );
not \U$7441 ( \7534 , \6514 );
or \U$7442 ( \7535 , \7533 , \7534 );
nand \U$7443 ( \7536 , \7535 , \7446 );
not \U$7444 ( \7537 , \7536 );
or \U$7445 ( \7538 , \7532 , \7537 );
nand \U$7446 ( \7539 , \5064 , \5011 );
or \U$7447 ( \7540 , \7459 , \7539 );
nand \U$7448 ( \7541 , \7540 , \7468 );
and \U$7449 ( \7542 , \7541 , \5114 );
nor \U$7450 ( \7543 , \7542 , \7473 );
nand \U$7451 ( \7544 , \7538 , \7543 );
nand \U$7452 ( \7545 , \7476 , \5155 );
not \U$7453 ( \7546 , \7545 );
and \U$7454 ( \7547 , \7544 , \7546 );
not \U$7455 ( \7548 , \7544 );
and \U$7456 ( \7549 , \7548 , \7545 );
nor \U$7457 ( \7550 , \7547 , \7549 );
buf \U$7458 ( \7551 , \7550 );
not \U$7459 ( \7552 , \5012 );
not \U$7460 ( \7553 , \5064 );
nor \U$7461 ( \7554 , \7552 , \7553 );
not \U$7462 ( \7555 , \7554 );
not \U$7463 ( \7556 , \7536 );
or \U$7464 ( \7557 , \7555 , \7556 );
not \U$7465 ( \7558 , \7541 );
nand \U$7466 ( \7559 , \7557 , \7558 );
not \U$7467 ( \7560 , \7473 );
nand \U$7468 ( \7561 , \7560 , \5114 );
not \U$7469 ( \7562 , \7561 );
and \U$7470 ( \7563 , \7559 , \7562 );
not \U$7471 ( \7564 , \7559 );
and \U$7472 ( \7565 , \7564 , \7561 );
nor \U$7473 ( \7566 , \7563 , \7565 );
buf \U$7474 ( \7567 , \7566 );
not \U$7475 ( \7568 , \5012 );
not \U$7476 ( \7569 , \7536 );
or \U$7477 ( \7570 , \7568 , \7569 );
buf \U$7478 ( \7571 , \7456 );
and \U$7479 ( \7572 , \7571 , \5011 );
nor \U$7480 ( \7573 , \7572 , \7458 );
nand \U$7481 ( \7574 , \7570 , \7573 );
not \U$7482 ( \7575 , \7553 );
nand \U$7483 ( \7576 , \7575 , \7468 );
not \U$7484 ( \7577 , \7576 );
and \U$7485 ( \7578 , \7574 , \7577 );
not \U$7486 ( \7579 , \7574 );
and \U$7487 ( \7580 , \7579 , \7576 );
nor \U$7488 ( \7581 , \7578 , \7580 );
buf \U$7489 ( \7582 , \7581 );
not \U$7490 ( \7583 , \4845 );
nor \U$7491 ( \7584 , \7583 , \7451 );
not \U$7492 ( \7585 , \7584 );
not \U$7493 ( \7586 , \7447 );
or \U$7494 ( \7587 , \7585 , \7586 );
not \U$7495 ( \7588 , \7571 );
nand \U$7496 ( \7589 , \7587 , \7588 );
not \U$7497 ( \7590 , \7458 );
nand \U$7498 ( \7591 , \7590 , \5011 );
not \U$7499 ( \7592 , \7591 );
and \U$7500 ( \7593 , \7589 , \7592 );
not \U$7501 ( \7594 , \7589 );
and \U$7502 ( \7595 , \7594 , \7591 );
nor \U$7503 ( \7596 , \7593 , \7595 );
buf \U$7504 ( \7597 , \7596 );
not \U$7505 ( \7598 , \4845 );
not \U$7506 ( \7599 , \7536 );
or \U$7507 ( \7600 , \7598 , \7599 );
nand \U$7508 ( \7601 , \7600 , \7452 );
not \U$7509 ( \7602 , \7451 );
nand \U$7510 ( \7603 , \7602 , \7455 );
not \U$7511 ( \7604 , \7603 );
and \U$7512 ( \7605 , \7601 , \7604 );
not \U$7513 ( \7606 , \7601 );
and \U$7514 ( \7607 , \7606 , \7603 );
nor \U$7515 ( \7608 , \7605 , \7607 );
buf \U$7516 ( \7609 , \7608 );
nand \U$7517 ( \7610 , \7452 , \4845 );
xnor \U$7518 ( \7611 , \7447 , \7610 );
buf \U$7519 ( \7612 , \7611 );
buf \U$7520 ( \7613 , \5501 );
not \U$7521 ( \7614 , \7613 );
not \U$7522 ( \7615 , \5928 );
not \U$7523 ( \7616 , \7615 );
not \U$7524 ( \7617 , \6503 );
and \U$7525 ( \7618 , \7617 , \6158 , \6081 );
not \U$7526 ( \7619 , \7618 );
not \U$7527 ( \7620 , \7427 );
or \U$7528 ( \7621 , \7619 , \7620 );
nand \U$7529 ( \7622 , \7621 , \6513 );
not \U$7530 ( \7623 , \7622 );
or \U$7531 ( \7624 , \7616 , \7623 );
not \U$7532 ( \7625 , \7436 );
nand \U$7533 ( \7626 , \7624 , \7625 );
not \U$7534 ( \7627 , \7626 );
or \U$7535 ( \7628 , \7614 , \7627 );
buf \U$7536 ( \7629 , \7438 );
not \U$7537 ( \7630 , \7629 );
nand \U$7538 ( \7631 , \7628 , \7630 );
nand \U$7539 ( \7632 , \5310 , \7442 );
not \U$7540 ( \7633 , \7632 );
and \U$7541 ( \7634 , \7631 , \7633 );
not \U$7542 ( \7635 , \7631 );
and \U$7543 ( \7636 , \7635 , \7632 );
nor \U$7544 ( \7637 , \7634 , \7636 );
buf \U$7545 ( \7638 , \7637 );
not \U$7546 ( \7639 , \7629 );
nand \U$7547 ( \7640 , \7639 , \7613 );
not \U$7548 ( \7641 , \7640 );
and \U$7549 ( \7642 , \7626 , \7641 );
not \U$7550 ( \7643 , \7626 );
and \U$7551 ( \7644 , \7643 , \7640 );
nor \U$7552 ( \7645 , \7642 , \7644 );
buf \U$7553 ( \7646 , \7645 );
not \U$7554 ( \7647 , \5927 );
not \U$7555 ( \7648 , \7622 );
or \U$7556 ( \7649 , \7647 , \7648 );
nand \U$7557 ( \7650 , \7649 , \7434 );
nand \U$7558 ( \7651 , \7432 , \5746 );
not \U$7559 ( \7652 , \7651 );
and \U$7560 ( \7653 , \7650 , \7652 );
not \U$7561 ( \7654 , \7650 );
and \U$7562 ( \7655 , \7654 , \7651 );
nor \U$7563 ( \7656 , \7653 , \7655 );
buf \U$7564 ( \7657 , \7656 );
nand \U$7565 ( \7658 , \5927 , \7434 );
not \U$7566 ( \7659 , \7658 );
and \U$7567 ( \7660 , \7622 , \7659 );
not \U$7568 ( \7661 , \7622 );
and \U$7569 ( \7662 , \7661 , \7658 );
nor \U$7570 ( \7663 , \7660 , \7662 );
buf \U$7571 ( \7664 , \7663 );
not \U$7572 ( \7665 , \7617 );
and \U$7573 ( \7666 , \7401 , \7416 , \7417 );
not \U$7574 ( \7667 , \7398 );
nand \U$7575 ( \7668 , \7666 , \7667 );
buf \U$7576 ( \7669 , \7358 );
not \U$7577 ( \7670 , \7669 );
nand \U$7578 ( \7671 , \7670 , \7418 );
nand \U$7579 ( \7672 , \7668 , \7671 , \7426 );
not \U$7580 ( \7673 , \7672 );
or \U$7581 ( \7674 , \7665 , \7673 );
not \U$7582 ( \7675 , \6504 );
nand \U$7583 ( \7676 , \7674 , \7675 );
buf \U$7584 ( \7677 , \6158 );
and \U$7585 ( \7678 , \7676 , \7677 );
buf \U$7586 ( \7679 , \6506 );
nor \U$7587 ( \7680 , \7678 , \7679 );
nand \U$7588 ( \7681 , \6081 , \6511 );
and \U$7589 ( \7682 , \7680 , \7681 );
not \U$7590 ( \7683 , \7680 );
not \U$7591 ( \7684 , \7681 );
and \U$7592 ( \7685 , \7683 , \7684 );
nor \U$7593 ( \7686 , \7682 , \7685 );
buf \U$7594 ( \7687 , \7686 );
not \U$7595 ( \7688 , \7677 );
nor \U$7596 ( \7689 , \7688 , \7679 );
and \U$7597 ( \7690 , \7689 , \7676 );
not \U$7598 ( \7691 , \7689 );
not \U$7599 ( \7692 , \7676 );
and \U$7600 ( \7693 , \7691 , \7692 );
nor \U$7601 ( \7694 , \7690 , \7693 );
buf \U$7602 ( \7695 , \7694 );
nand \U$7603 ( \7696 , \7668 , \6501 , \7426 , \7671 );
nand \U$7604 ( \7697 , \6347 , \7617 );
not \U$7605 ( \7698 , \7697 );
and \U$7606 ( \7699 , \7696 , \7698 );
not \U$7607 ( \7700 , \7696 );
and \U$7608 ( \7701 , \7700 , \7697 );
nor \U$7609 ( \7702 , \7699 , \7701 );
buf \U$7610 ( \7703 , \7702 );
and \U$7611 ( \7704 , \7416 , \7417 );
nand \U$7612 ( \7705 , \7670 , \7704 );
nand \U$7613 ( \7706 , \7667 , \7704 );
buf \U$7614 ( \7707 , \7423 );
nand \U$7615 ( \7708 , \7705 , \7706 , \7707 );
nand \U$7616 ( \7709 , \6501 , \7425 );
not \U$7617 ( \7710 , \7709 );
and \U$7618 ( \7711 , \7708 , \7710 );
not \U$7619 ( \7712 , \7708 );
and \U$7620 ( \7713 , \7712 , \7709 );
nor \U$7621 ( \7714 , \7711 , \7713 );
buf \U$7622 ( \7715 , \7714 );
and \U$7623 ( \7716 , \7416 , \7707 );
not \U$7624 ( \7717 , \7417 );
not \U$7625 ( \7718 , \7362 );
nand \U$7626 ( \7719 , \7718 , \7669 );
not \U$7627 ( \7720 , \7719 );
or \U$7628 ( \7721 , \7717 , \7720 );
not \U$7629 ( \7722 , \7397 );
nand \U$7630 ( \7723 , \7721 , \7722 );
and \U$7631 ( \7724 , \7716 , \7723 );
not \U$7632 ( \7725 , \7716 );
not \U$7633 ( \7726 , \7723 );
and \U$7634 ( \7727 , \7725 , \7726 );
nor \U$7635 ( \7728 , \7724 , \7727 );
buf \U$7636 ( \7729 , \7728 );
nand \U$7637 ( \7730 , \7417 , \7722 );
not \U$7638 ( \7731 , \7730 );
and \U$7639 ( \7732 , \7719 , \7731 );
not \U$7640 ( \7733 , \7719 );
and \U$7641 ( \7734 , \7733 , \7730 );
nor \U$7642 ( \7735 , \7732 , \7734 );
buf \U$7643 ( \7736 , \7735 );
buf \U$7644 ( \7737 , \7122 );
not \U$7645 ( \7738 , \7357 );
or \U$7646 ( \7739 , \7737 , \7738 );
and \U$7647 ( \7740 , \7236 , \7357 );
nor \U$7648 ( \7741 , \7740 , \7234 );
nand \U$7649 ( \7742 , \7739 , \7741 );
and \U$7650 ( \7743 , \7742 , \7356 );
not \U$7651 ( \7744 , \7359 );
nor \U$7652 ( \7745 , \7743 , \7744 );
nand \U$7653 ( \7746 , \7345 , \7360 );
and \U$7654 ( \7747 , \7745 , \7746 );
not \U$7655 ( \7748 , \7745 );
not \U$7656 ( \7749 , \7746 );
and \U$7657 ( \7750 , \7748 , \7749 );
nor \U$7658 ( \7751 , \7747 , \7750 );
buf \U$7659 ( \7752 , \7751 );
nand \U$7660 ( \7753 , \7359 , \7356 );
not \U$7661 ( \7754 , \7753 );
and \U$7662 ( \7755 , \7742 , \7754 );
not \U$7663 ( \7756 , \7742 );
and \U$7664 ( \7757 , \7756 , \7753 );
nor \U$7665 ( \7758 , \7755 , \7757 );
buf \U$7666 ( \7759 , \7758 );
not \U$7667 ( \7760 , \7236 );
nand \U$7668 ( \7761 , \7737 , \7760 );
not \U$7669 ( \7762 , \7234 );
nand \U$7670 ( \7763 , \7762 , \7357 );
not \U$7671 ( \7764 , \7763 );
and \U$7672 ( \7765 , \7761 , \7764 );
not \U$7673 ( \7766 , \7761 );
and \U$7674 ( \7767 , \7766 , \7763 );
nor \U$7675 ( \7768 , \7765 , \7767 );
buf \U$7676 ( \7769 , \7768 );
nand \U$7677 ( \7770 , \7760 , \7121 );
not \U$7678 ( \7771 , \7006 );
and \U$7679 ( \7772 , \7770 , \7771 );
not \U$7680 ( \7773 , \7770 );
and \U$7681 ( \7774 , \7773 , \7006 );
nor \U$7682 ( \7775 , \7772 , \7774 );
buf \U$7683 ( \7776 , \7775 );
not \U$7684 ( \7777 , \6987 );
not \U$7685 ( \7778 , \6961 );
or \U$7686 ( \7779 , \7777 , \7778 );
nand \U$7687 ( \7780 , \7779 , \6989 );
and \U$7688 ( \7781 , \6814 , \6998 );
not \U$7689 ( \7782 , \7003 );
nor \U$7690 ( \7783 , \7781 , \7782 );
and \U$7691 ( \7784 , \7780 , \7783 );
not \U$7692 ( \7785 , \7780 );
not \U$7693 ( \7786 , \7783 );
and \U$7694 ( \7787 , \7785 , \7786 );
nor \U$7695 ( \7788 , \7784 , \7787 );
buf \U$7696 ( \7789 , \7788 );
nand \U$7697 ( \7790 , \6998 , \7003 );
not \U$7698 ( \7791 , \6814 );
and \U$7699 ( \7792 , \7790 , \7791 );
not \U$7700 ( \7793 , \7790 );
and \U$7701 ( \7794 , \7793 , \6814 );
nor \U$7702 ( \7795 , \7792 , \7794 );
buf \U$7703 ( \7796 , \7795 );
xor \U$7704 ( \7797 , \6590 , \6651 );
xor \U$7705 ( \7798 , \7797 , \6811 );
buf \U$7706 ( \7799 , \7798 );
not \U$7707 ( \7800 , \6808 );
nand \U$7708 ( \7801 , \7800 , \6810 );
or \U$7709 ( \7802 , \6795 , \6793 );
nand \U$7710 ( \7803 , \7802 , \6714 );
and \U$7711 ( \7804 , \7801 , \7803 );
not \U$7712 ( \7805 , \7801 );
not \U$7713 ( \7806 , \7803 );
and \U$7714 ( \7807 , \7805 , \7806 );
nor \U$7715 ( \7808 , \7804 , \7807 );
buf \U$7716 ( \7809 , \7808 );
not \U$7717 ( \7810 , \6795 );
nand \U$7718 ( \7811 , \7810 , \6714 );
buf \U$7719 ( \7812 , \6793 );
not \U$7720 ( \7813 , \7812 );
and \U$7721 ( \7814 , \7811 , \7813 );
not \U$7722 ( \7815 , \7811 );
and \U$7723 ( \7816 , \7815 , \7812 );
nor \U$7724 ( \7817 , \7814 , \7816 );
buf \U$7725 ( \7818 , \7817 );
endmodule

