//
// Conformal-LEC Version 20.10-d215 (04-Sep-2020)
//
module top(RIa139848_33,RIa138a38_3,RIa139c80_42,RIa139cf8_43,RIa139c08_41,RIa139de8_45,RIa139d70_44,RIa139e60_46,RIa139ed8_47,
        RIa139f50_48,RIa138ee8_13,RIa139398_23,RIa1398c0_34,RIa138e70_12,RIa1389c0_2,RIa139320_22,RIa139938_35,RIa138df8_11,RIa138948_1,
        RIa1392a8_21,RIa1399b0_36,RIa139aa0_38,RIa139b18_39,RIa139b90_40,RIa139410_24,RIa138ab0_4,RIa138f60_14,RIa138fd8_15,RIa138b28_5,
        RIa139488_25,RIa139050_16,RIa138ba0_6,RIa139500_26,RIa1395f0_28,RIa138c90_8,RIa139140_18,RIa139230_20,RIa138d80_10,RIa1396e0_30,
        RIa1391b8_19,RIa138d08_9,RIa139668_29,RIa1390c8_17,RIa138c18_7,RIa139578_27,RIa139a28_37,RIa1397d0_32,RIa139758_31,R_31_942aab8,
        R_32_942ab60,R_33_942ac08,R_34_942acb0,R_35_942ad58,R_36_942ae00,R_37_942aea8,R_38_942af50,R_39_942aff8,R_3a_942b0a0,R_3b_942b148,
        R_3c_942b1f0,R_3d_942b298,R_3e_942b340,R_3f_942b3e8,R_40_942b490,R_41_942b538,R_42_942b5e0,R_43_942b688,R_44_942b730);
input RIa139848_33,RIa138a38_3,RIa139c80_42,RIa139cf8_43,RIa139c08_41,RIa139de8_45,RIa139d70_44,RIa139e60_46,RIa139ed8_47,
        RIa139f50_48,RIa138ee8_13,RIa139398_23,RIa1398c0_34,RIa138e70_12,RIa1389c0_2,RIa139320_22,RIa139938_35,RIa138df8_11,RIa138948_1,
        RIa1392a8_21,RIa1399b0_36,RIa139aa0_38,RIa139b18_39,RIa139b90_40,RIa139410_24,RIa138ab0_4,RIa138f60_14,RIa138fd8_15,RIa138b28_5,
        RIa139488_25,RIa139050_16,RIa138ba0_6,RIa139500_26,RIa1395f0_28,RIa138c90_8,RIa139140_18,RIa139230_20,RIa138d80_10,RIa1396e0_30,
        RIa1391b8_19,RIa138d08_9,RIa139668_29,RIa1390c8_17,RIa138c18_7,RIa139578_27,RIa139a28_37,RIa1397d0_32,RIa139758_31;
output R_31_942aab8,R_32_942ab60,R_33_942ac08,R_34_942acb0,R_35_942ad58,R_36_942ae00,R_37_942aea8,R_38_942af50,R_39_942aff8,
        R_3a_942b0a0,R_3b_942b148,R_3c_942b1f0,R_3d_942b298,R_3e_942b340,R_3f_942b3e8,R_40_942b490,R_41_942b538,R_42_942b5e0,R_43_942b688,
        R_44_942b730;


wire \63_ZERO , \64_ONE , \65 , \66 , \67 , \68 , \69 , \70 , \71 ,
         \72 , \73 , \74 , \75 , \76 , \77 , \78 , \79 , \80 , \81 ,
         \82 , \83 , \84 , \85 , \86 , \87 , \88 , \89 , \90 , \91 ,
         \92 , \93 , \94 , \95 , \96 , \97 , \98 , \99 , \100 , \101 ,
         \102 , \103 , \104 , \105 , \106 , \107 , \108 , \109 , \110 , \111 ,
         \112 , \113 , \114 , \115 , \116 , \117 , \118 , \119 , \120 , \121 ,
         \122 , \123 , \124 , \125 , \126 , \127 , \128 , \129 , \130 , \131 ,
         \132 , \133 , \134 , \135 , \136 , \137 , \138 , \139 , \140 , \141 ,
         \142 , \143 , \144 , \145 , \146 , \147 , \148 , \149 , \150 , \151 ,
         \152 , \153 , \154 , \155 , \156 , \157 , \158 , \159 , \160 , \161 ,
         \162 , \163 , \164 , \165 , \166 , \167 , \168 , \169 , \170 , \171 ,
         \172 , \173 , \174 , \175 , \176 , \177 , \178 , \179 , \180 , \181 ,
         \182 , \183 , \184 , \185 , \186 , \187 , \188 , \189 , \190 , \191 ,
         \192 , \193 , \194 , \195 , \196 , \197 , \198 , \199 , \200 , \201 ,
         \202 , \203 , \204 , \205 , \206 , \207 , \208 , \209 , \210 , \211 ,
         \212 , \213 , \214 , \215 , \216 , \217 , \218 , \219 , \220 , \221 ,
         \222 , \223 , \224 , \225 , \226 , \227 , \228 , \229 , \230 , \231 ,
         \232 , \233 , \234 , \235 , \236 , \237 , \238 , \239 , \240 , \241 ,
         \242 , \243 , \244 , \245 , \246 , \247 , \248 , \249 , \250 , \251 ,
         \252 , \253 , \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 ,
         \262 , \263 , \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 ,
         \272 , \273 , \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 ,
         \282 , \283 , \284 , \285 , \286 , \287 , \288 , \289 , \290 , \291 ,
         \292 , \293 , \294 , \295 , \296 , \297 , \298 , \299 , \300 , \301 ,
         \302 , \303 , \304 , \305 , \306 , \307 , \308 , \309 , \310 , \311 ,
         \312 , \313 , \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321 ,
         \322 , \323 , \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331 ,
         \332 , \333 , \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 ,
         \342 , \343 , \344 , \345 , \346 , \347 , \348 , \349 , \350 , \351 ,
         \352 , \353 , \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 ,
         \362 , \363 , \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 ,
         \372 , \373 , \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 ,
         \382 , \383 , \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 ,
         \392 , \393 , \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 ,
         \402 , \403 , \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 ,
         \412 , \413 , \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 ,
         \422 , \423 , \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 ,
         \432 , \433 , \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 ,
         \442 , \443 , \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 ,
         \452 , \453 , \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 ,
         \462 , \463 , \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 ,
         \472 , \473 , \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 ,
         \482 , \483 , \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 ,
         \492 , \493 , \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 ,
         \502 , \503 , \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 ,
         \512 , \513 , \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 ,
         \522 , \523 , \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 ,
         \532 , \533 , \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 ,
         \542 , \543 , \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 ,
         \552 , \553 , \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 ,
         \562 , \563 , \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 ,
         \572 , \573 , \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 ,
         \582 , \583 , \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 ,
         \592 , \593 , \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 ,
         \602 , \603 , \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 ,
         \612 , \613 , \614 , \615 , \616 , \617 , \618 , \619 , \620 , \621 ,
         \622 , \623 , \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 ,
         \632 , \633 , \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 ,
         \642 , \643 , \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 ,
         \652 , \653 , \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 ,
         \662 , \663 , \664 , \665 , \666 , \667 , \668 , \669 , \670 , \671 ,
         \672 , \673 , \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 ,
         \682 , \683 , \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 ,
         \692 , \693 , \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 ,
         \702 , \703 , \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 ,
         \712 , \713 , \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 ,
         \722 , \723 , \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 ,
         \732 , \733 , \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 ,
         \742 , \743 , \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 ,
         \752 , \753 , \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 ,
         \762 , \763 , \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 ,
         \772 , \773 , \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 ,
         \782 , \783 , \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 ,
         \792 , \793 , \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 ,
         \802 , \803 , \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 ,
         \812 , \813 , \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 ,
         \822 , \823 , \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 ,
         \832 , \833 , \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 ,
         \842 , \843 , \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 ,
         \852 , \853 , \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 ,
         \862 , \863 , \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 ,
         \872 , \873 , \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 ,
         \882 , \883 , \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 ,
         \892 , \893 , \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 ,
         \902 , \903 , \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 ,
         \912 , \913 , \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 ,
         \922 , \923 , \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 ,
         \932 , \933 , \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 ,
         \942 , \943 , \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 ,
         \952 , \953 , \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 ,
         \962 , \963 , \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 ,
         \972 , \973 , \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 ,
         \982 , \983 , \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 ,
         \992 , \993 , \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 ,
         \1002 , \1003 , \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 ,
         \1012 , \1013 , \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 ,
         \1022 , \1023 , \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 ,
         \1032 , \1033 , \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 ,
         \1042 , \1043 , \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 ,
         \1052 , \1053 , \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 ,
         \1062 , \1063 , \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 ,
         \1072 , \1073 , \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 ,
         \1082 , \1083 , \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 ,
         \1092 , \1093 , \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 ,
         \1102 , \1103 , \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 ,
         \1112 , \1113 , \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 ,
         \1122 , \1123 , \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 ,
         \1132 , \1133 , \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 ,
         \1142 , \1143 , \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 ,
         \1152 , \1153 , \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 ,
         \1162 , \1163 , \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 ,
         \1172 , \1173 , \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 ,
         \1182 , \1183 , \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 ,
         \1192 , \1193 , \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 ,
         \1202 , \1203 , \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 ,
         \1212 , \1213 , \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 ,
         \1222 , \1223 , \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 ,
         \1232 , \1233 , \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 ,
         \1242 , \1243 , \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 ,
         \1252 , \1253 , \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 ,
         \1262 , \1263 , \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 ,
         \1272 , \1273 , \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 ,
         \1282 , \1283 , \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 ,
         \1292 , \1293 , \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 ,
         \1302 , \1303 , \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 ,
         \1312 , \1313 , \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 ,
         \1322 , \1323 , \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 ,
         \1332 , \1333 , \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 ,
         \1342 , \1343 , \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 ,
         \1352 , \1353 , \1354 , \1355 , \1356 , \1357 , \1358 , \1359 , \1360 , \1361 ,
         \1362 , \1363 , \1364 , \1365 , \1366 , \1367 , \1368 , \1369 , \1370 , \1371 ,
         \1372 , \1373 , \1374 , \1375 , \1376 , \1377 , \1378 , \1379 , \1380 , \1381 ,
         \1382 , \1383 , \1384 , \1385 , \1386 , \1387 , \1388 , \1389 , \1390 , \1391 ,
         \1392 , \1393 , \1394 , \1395 , \1396 , \1397 , \1398 , \1399 , \1400 , \1401 ,
         \1402 , \1403 , \1404 , \1405 , \1406 , \1407 ;
buf \U$labajz155 ( R_31_942aab8, \1236 );
buf \U$labajz156 ( R_32_942ab60, \1243 );
buf \U$labajz157 ( R_33_942ac08, \1271 );
buf \U$labajz158 ( R_34_942acb0, \1278 );
buf \U$labajz159 ( R_35_942ad58, \1294 );
buf \U$labajz160 ( R_36_942ae00, \1297 );
buf \U$labajz161 ( R_37_942aea8, \1311 );
buf \U$labajz162 ( R_38_942af50, \1319 );
buf \U$labajz163 ( R_39_942aff8, \1339 );
buf \U$labajz164 ( R_3a_942b0a0, \1346 );
buf \U$labajz165 ( R_3b_942b148, \1355 );
buf \U$labajz166 ( R_3c_942b1f0, \1364 );
buf \U$labajz167 ( R_3d_942b298, \1371 );
buf \U$labajz168 ( R_3e_942b340, \1378 );
buf \U$labajz169 ( R_3f_942b3e8, \1385 );
buf \U$labajz170 ( R_40_942b490, \1392 );
buf \U$labajz171 ( R_41_942b538, \1395 );
buf \U$labajz172 ( R_42_942b5e0, \1399 );
buf \U$labajz173 ( R_43_942b688, \1405 );
buf \U$labajz174 ( R_44_942b730, \1407 );
not \U$1 ( \65 , RIa138948_1);
nor \U$2 ( \66 , RIa139ed8_47, RIa139f50_48);
not \U$3 ( \67 , \66 );
or \U$4 ( \68 , \65 , \67 );
and \U$5 ( \69 , RIa138df8_11, RIa139f50_48);
and \U$6 ( \70 , RIa1392a8_21, RIa139ed8_47);
nor \U$7 ( \71 , \69 , \70 );
nand \U$8 ( \72 , \68 , \71 );
buf \U$9 ( \73 , \72 );
nand \U$10 ( \74 , RIa139848_33, \73 );
nor \U$11 ( \75 , RIa139ed8_47, RIa139f50_48);
not \U$12 ( \76 , \75 );
not \U$13 ( \77 , RIa138a38_3);
not \U$14 ( \78 , \77 );
or \U$15 ( \79 , \76 , \78 );
nand \U$16 ( \80 , RIa138ee8_13, RIa139f50_48);
not \U$17 ( \81 , RIa139398_23);
nand \U$18 ( \82 , \80 , \81 , RIa139ed8_47);
nand \U$19 ( \83 , \79 , \82 );
nor \U$20 ( \84 , RIa139ed8_47, RIa138ee8_13);
and \U$21 ( \85 , \84 , RIa139f50_48);
nor \U$22 ( \86 , \83 , \85 );
buf \U$23 ( \87 , \86 );
not \U$24 ( \88 , \87 );
not \U$25 ( \89 , \88 );
nand \U$26 ( \90 , \89 , RIa139758_31);
xor \U$27 ( \91 , \74 , \90 );
not \U$28 ( \92 , RIa1389c0_2);
nor \U$29 ( \93 , RIa139ed8_47, RIa139f50_48);
not \U$30 ( \94 , \93 );
or \U$31 ( \95 , \92 , \94 );
and \U$32 ( \96 , RIa138e70_12, RIa139f50_48);
and \U$33 ( \97 , RIa139320_22, RIa139ed8_47);
nor \U$34 ( \98 , \96 , \97 );
nand \U$35 ( \99 , \95 , \98 );
buf \U$36 ( \100 , \99 );
and \U$37 ( \101 , \100 , RIa1397d0_32);
not \U$38 ( \102 , \101 );
and \U$39 ( \103 , \91 , \102 );
and \U$40 ( \104 , \90 , \74 );
nor \U$41 ( \105 , \103 , \104 );
not \U$42 ( \106 , \105 );
nand \U$43 ( \107 , \100 , RIa139758_31);
nand \U$44 ( \108 , \73 , RIa1397d0_32);
xor \U$45 ( \109 , \107 , \108 );
and \U$46 ( \110 , \106 , \109 );
and \U$47 ( \111 , \107 , \108 );
nor \U$48 ( \112 , \110 , \111 );
and \U$49 ( \113 , \73 , RIa139758_31);
or \U$50 ( \114 , \112 , \113 );
not \U$51 ( \115 , \114 );
not \U$52 ( \116 , RIa138b28_5);
not \U$53 ( \117 , \66 );
or \U$54 ( \118 , \116 , \117 );
and \U$55 ( \119 , RIa138fd8_15, RIa139f50_48);
and \U$56 ( \120 , RIa139488_25, RIa139ed8_47);
nor \U$57 ( \121 , \119 , \120 );
nand \U$58 ( \122 , \118 , \121 );
buf \U$59 ( \123 , \122 );
nand \U$60 ( \124 , \123 , RIa1397d0_32);
not \U$61 ( \125 , \124 );
nor \U$62 ( \126 , RIa139ed8_47, RIa139f50_48);
not \U$63 ( \127 , \126 );
not \U$64 ( \128 , RIa138ba0_6);
or \U$65 ( \129 , \127 , \128 );
and \U$66 ( \130 , RIa139050_16, RIa139f50_48);
and \U$67 ( \131 , RIa139500_26, RIa139ed8_47);
nor \U$68 ( \132 , \130 , \131 );
nand \U$69 ( \133 , \129 , \132 );
buf \U$70 ( \134 , \133 );
and \U$71 ( \135 , \134 , RIa139758_31);
not \U$72 ( \136 , \135 );
or \U$73 ( \137 , \125 , \136 );
or \U$74 ( \138 , \135 , \124 );
nand \U$75 ( \139 , \137 , \138 );
nand \U$76 ( \140 , \89 , RIa1398c0_34);
xnor \U$77 ( \141 , \139 , \140 );
nand \U$78 ( \142 , \123 , RIa139848_33);
not \U$79 ( \143 , \142 );
not \U$80 ( \144 , \143 );
nand \U$81 ( \145 , \134 , RIa1397d0_32);
not \U$82 ( \146 , \145 );
not \U$83 ( \147 , \146 );
or \U$84 ( \148 , \144 , \147 );
not \U$85 ( \149 , \142 );
not \U$86 ( \150 , \145 );
or \U$87 ( \151 , \149 , \150 );
not \U$88 ( \152 , \87 );
not \U$89 ( \153 , RIa139938_35);
nor \U$90 ( \154 , \152 , \153 );
nand \U$91 ( \155 , \151 , \154 );
nand \U$92 ( \156 , \148 , \155 );
nand \U$93 ( \157 , \100 , RIa1399b0_36);
not \U$94 ( \158 , \157 );
not \U$95 ( \159 , \158 );
nand \U$96 ( \160 , \73 , RIa139a28_37);
not \U$97 ( \161 , \160 );
not \U$98 ( \162 , \161 );
or \U$99 ( \163 , \159 , \162 );
not \U$100 ( \164 , \157 );
not \U$101 ( \165 , \160 );
or \U$102 ( \166 , \164 , \165 );
not \U$103 ( \167 , RIa138ab0_4);
nor \U$104 ( \168 , RIa139ed8_47, RIa139f50_48);
not \U$105 ( \169 , \168 );
or \U$106 ( \170 , \167 , \169 );
and \U$107 ( \171 , RIa138f60_14, RIa139f50_48);
and \U$108 ( \172 , RIa139410_24, RIa139ed8_47);
nor \U$109 ( \173 , \171 , \172 );
nand \U$110 ( \174 , \170 , \173 );
buf \U$111 ( \175 , \174 );
and \U$112 ( \176 , \175 , RIa1398c0_34);
nand \U$113 ( \177 , \166 , \176 );
nand \U$114 ( \178 , \163 , \177 );
nor \U$115 ( \179 , \156 , \178 );
not \U$116 ( \180 , \179 );
nand \U$117 ( \181 , \156 , \178 );
nand \U$118 ( \182 , \180 , \181 );
nand \U$119 ( \183 , \73 , RIa1399b0_36);
not \U$120 ( \184 , \183 );
nand \U$121 ( \185 , \100 , RIa139938_35);
not \U$122 ( \186 , \185 );
not \U$123 ( \187 , \186 );
or \U$124 ( \188 , \184 , \187 );
not \U$125 ( \189 , \183 );
nand \U$126 ( \190 , \185 , \189 );
nand \U$127 ( \191 , \188 , \190 );
buf \U$128 ( \192 , \175 );
nand \U$129 ( \193 , \192 , RIa139848_33);
not \U$130 ( \194 , \193 );
and \U$131 ( \195 , \191 , \194 );
not \U$132 ( \196 , \191 );
and \U$133 ( \197 , \196 , \193 );
nor \U$134 ( \198 , \195 , \197 );
not \U$135 ( \199 , \198 );
and \U$136 ( \200 , \182 , \199 );
not \U$137 ( \201 , \182 );
and \U$138 ( \202 , \201 , \198 );
nor \U$139 ( \203 , \200 , \202 );
xor \U$140 ( \204 , \141 , \203 );
nor \U$141 ( \205 , RIa139ed8_47, RIa1390c8_17);
and \U$142 ( \206 , \205 , RIa139f50_48);
not \U$143 ( \207 , RIa138c18_7);
not \U$144 ( \208 , \207 );
not \U$145 ( \209 , \75 );
or \U$146 ( \210 , \208 , \209 );
not \U$147 ( \211 , RIa139578_27);
nand \U$148 ( \212 , RIa1390c8_17, RIa139f50_48);
nand \U$149 ( \213 , \211 , \212 , RIa139ed8_47);
nand \U$150 ( \214 , \210 , \213 );
nor \U$151 ( \215 , \206 , \214 );
buf \U$152 ( \216 , \215 );
nand \U$153 ( \217 , \216 , RIa139758_31);
not \U$154 ( \218 , \153 );
nand \U$155 ( \219 , \218 , \175 );
nand \U$156 ( \220 , \100 , RIa139a28_37);
nand \U$157 ( \221 , \219 , \220 );
nand \U$158 ( \222 , \72 , RIa139aa0_38);
nand \U$159 ( \223 , \220 , \222 );
nand \U$160 ( \224 , \219 , \222 );
nand \U$161 ( \225 , \221 , \223 , \224 );
xor \U$162 ( \226 , \217 , \225 );
not \U$163 ( \227 , \88 );
and \U$164 ( \228 , \227 , RIa1399b0_36);
not \U$165 ( \229 , \228 );
not \U$166 ( \230 , RIa138c90_8);
not \U$167 ( \231 , \168 );
or \U$168 ( \232 , \230 , \231 );
and \U$169 ( \233 , RIa139140_18, RIa139f50_48);
and \U$170 ( \234 , RIa1395f0_28, RIa139ed8_47);
nor \U$171 ( \235 , \233 , \234 );
nand \U$172 ( \236 , \232 , \235 );
nand \U$173 ( \237 , \236 , RIa139758_31);
nand \U$174 ( \238 , \123 , RIa1398c0_34);
xor \U$175 ( \239 , \237 , \238 );
and \U$176 ( \240 , \229 , \239 );
and \U$177 ( \241 , \237 , \238 );
nor \U$178 ( \242 , \240 , \241 );
not \U$179 ( \243 , \242 );
and \U$180 ( \244 , \226 , \243 );
and \U$181 ( \245 , \217 , \225 );
nor \U$182 ( \246 , \244 , \245 );
and \U$183 ( \247 , \204 , \246 );
and \U$184 ( \248 , \141 , \203 );
or \U$185 ( \249 , \247 , \248 );
not \U$186 ( \250 , \249 );
not \U$187 ( \251 , \186 );
not \U$188 ( \252 , \189 );
and \U$189 ( \253 , \251 , \252 );
and \U$190 ( \254 , \191 , \193 );
nor \U$191 ( \255 , \253 , \254 );
not \U$192 ( \256 , \73 );
not \U$193 ( \257 , \256 );
nand \U$194 ( \258 , \257 , RIa139938_35);
nand \U$195 ( \259 , \192 , RIa1397d0_32);
xor \U$196 ( \260 , \258 , \259 );
nand \U$197 ( \261 , \100 , RIa1398c0_34);
xnor \U$198 ( \262 , \260 , \261 );
xor \U$199 ( \263 , \255 , \262 );
not \U$200 ( \264 , \140 );
not \U$201 ( \265 , \139 );
or \U$202 ( \266 , \264 , \265 );
not \U$203 ( \267 , \135 );
nand \U$204 ( \268 , \267 , \124 );
nand \U$205 ( \269 , \266 , \268 );
not \U$206 ( \270 , \269 );
nand \U$207 ( \271 , \89 , RIa139848_33);
not \U$208 ( \272 , \271 );
and \U$209 ( \273 , \123 , RIa139758_31);
not \U$210 ( \274 , \273 );
and \U$211 ( \275 , \272 , \274 );
and \U$212 ( \276 , \271 , \273 );
nor \U$213 ( \277 , \275 , \276 );
not \U$214 ( \278 , \277 );
and \U$215 ( \279 , \270 , \278 );
and \U$216 ( \280 , \269 , \277 );
nor \U$217 ( \281 , \279 , \280 );
xor \U$218 ( \282 , \263 , \281 );
not \U$219 ( \283 , \179 );
and \U$220 ( \284 , \283 , \198 );
not \U$221 ( \285 , \181 );
nor \U$222 ( \286 , \284 , \285 );
and \U$223 ( \287 , \282 , \286 );
not \U$224 ( \288 , \282 );
not \U$225 ( \289 , \286 );
and \U$226 ( \290 , \288 , \289 );
nor \U$227 ( \291 , \287 , \290 );
not \U$228 ( \292 , \291 );
not \U$229 ( \293 , \292 );
or \U$230 ( \294 , \250 , \293 );
nand \U$231 ( \295 , \282 , \289 );
nand \U$232 ( \296 , \294 , \295 );
not \U$233 ( \297 , \269 );
or \U$234 ( \298 , \297 , \277 );
not \U$235 ( \299 , \271 );
or \U$236 ( \300 , \299 , \273 );
nand \U$237 ( \301 , \298 , \300 );
not \U$238 ( \302 , \301 );
nand \U$239 ( \303 , \73 , RIa1398c0_34);
nand \U$240 ( \304 , \100 , RIa139848_33);
xor \U$241 ( \305 , \303 , \304 );
nand \U$242 ( \306 , \192 , RIa139758_31);
not \U$243 ( \307 , \306 );
and \U$244 ( \308 , \305 , \307 );
not \U$245 ( \309 , \305 );
and \U$246 ( \310 , \309 , \306 );
nor \U$247 ( \311 , \308 , \310 );
not \U$248 ( \312 , \311 );
nand \U$249 ( \313 , RIa1397d0_32, \89 );
not \U$250 ( \314 , \313 );
not \U$251 ( \315 , \261 );
not \U$252 ( \316 , \260 );
or \U$253 ( \317 , \315 , \316 );
nand \U$254 ( \318 , \259 , \258 );
nand \U$255 ( \319 , \317 , \318 );
not \U$256 ( \320 , \319 );
not \U$257 ( \321 , \320 );
or \U$258 ( \322 , \314 , \321 );
not \U$259 ( \323 , \313 );
nand \U$260 ( \324 , \319 , \323 );
nand \U$261 ( \325 , \322 , \324 );
not \U$262 ( \326 , \325 );
or \U$263 ( \327 , \312 , \326 );
or \U$264 ( \328 , \325 , \311 );
nand \U$265 ( \329 , \327 , \328 );
not \U$266 ( \330 , \329 );
not \U$267 ( \331 , \330 );
or \U$268 ( \332 , \302 , \331 );
not \U$269 ( \333 , \301 );
nand \U$270 ( \334 , \333 , \329 );
nand \U$271 ( \335 , \332 , \334 );
not \U$272 ( \336 , \335 );
xor \U$273 ( \337 , \255 , \262 );
and \U$274 ( \338 , \337 , \281 );
and \U$275 ( \339 , \255 , \262 );
or \U$276 ( \340 , \338 , \339 );
not \U$277 ( \341 , \340 );
and \U$278 ( \342 , \336 , \341 );
and \U$279 ( \343 , \335 , \340 );
nor \U$280 ( \344 , \342 , \343 );
nor \U$281 ( \345 , \296 , \344 );
not \U$282 ( \346 , \345 );
not \U$283 ( \347 , \222 );
and \U$284 ( \348 , \99 , RIa139b18_39);
buf \U$285 ( \349 , \348 );
nand \U$286 ( \350 , \347 , \349 );
not \U$287 ( \351 , \350 );
not \U$288 ( \352 , \351 );
nand \U$289 ( \353 , \215 , RIa1397d0_32);
and \U$290 ( \354 , \134 , RIa139848_33);
xnor \U$291 ( \355 , \353 , \354 );
not \U$292 ( \356 , \355 );
or \U$293 ( \357 , \352 , \356 );
or \U$294 ( \358 , \355 , \351 );
nand \U$295 ( \359 , \357 , \358 );
not \U$296 ( \360 , \359 );
not \U$297 ( \361 , \239 );
not \U$298 ( \362 , \228 );
and \U$299 ( \363 , \361 , \362 );
and \U$300 ( \364 , \239 , \228 );
nor \U$301 ( \365 , \363 , \364 );
not \U$302 ( \366 , \365 );
and \U$303 ( \367 , \360 , \366 );
and \U$304 ( \368 , \359 , \365 );
nor \U$305 ( \369 , \367 , \368 );
not \U$306 ( \370 , \100 );
not \U$307 ( \371 , RIa139aa0_38);
or \U$308 ( \372 , \370 , \371 );
not \U$309 ( \373 , RIa139b18_39);
or \U$310 ( \374 , \256 , \373 );
nand \U$311 ( \375 , \372 , \374 );
and \U$312 ( \376 , \350 , \375 );
not \U$313 ( \377 , \376 );
nand \U$314 ( \378 , \216 , RIa139848_33);
not \U$315 ( \379 , \378 );
and \U$316 ( \380 , \72 , RIa139b90_40);
and \U$317 ( \381 , \348 , \380 );
not \U$318 ( \382 , \381 );
and \U$319 ( \383 , \379 , \382 );
and \U$320 ( \384 , \348 , \380 );
and \U$321 ( \385 , \378 , \384 );
nor \U$322 ( \386 , \383 , \385 );
not \U$323 ( \387 , \386 );
and \U$324 ( \388 , \377 , \387 );
not \U$325 ( \389 , \384 );
and \U$326 ( \390 , \378 , \389 );
nor \U$327 ( \391 , \388 , \390 );
or \U$328 ( \392 , \369 , \391 );
not \U$329 ( \393 , \365 );
nand \U$330 ( \394 , \393 , \359 );
nand \U$331 ( \395 , \392 , \394 );
not \U$332 ( \396 , \395 );
and \U$333 ( \397 , \122 , RIa139938_35);
and \U$334 ( \398 , \134 , RIa1398c0_34);
xor \U$335 ( \399 , \397 , \398 );
and \U$336 ( \400 , \87 , RIa139a28_37);
and \U$337 ( \401 , \399 , \400 );
and \U$338 ( \402 , \397 , \398 );
or \U$339 ( \403 , \401 , \402 );
xor \U$340 ( \404 , \222 , \220 );
xnor \U$341 ( \405 , \404 , \219 );
xor \U$342 ( \406 , \403 , \405 );
not \U$343 ( \407 , RIa138d08_9);
nand \U$344 ( \408 , \407 , \93 );
not \U$345 ( \409 , RIa139ed8_47);
not \U$346 ( \410 , RIa1391b8_19);
nand \U$347 ( \411 , \409 , \410 , RIa139f50_48);
not \U$348 ( \412 , RIa139668_29);
nand \U$349 ( \413 , RIa1391b8_19, RIa139f50_48);
nand \U$350 ( \414 , \412 , \413 , RIa139ed8_47);
nand \U$351 ( \415 , \408 , \411 , \414 );
not \U$352 ( \416 , \415 );
nand \U$353 ( \417 , \416 , RIa139758_31);
and \U$354 ( \418 , \174 , RIa1399b0_36);
and \U$355 ( \419 , \236 , RIa1397d0_32);
nor \U$356 ( \420 , \418 , \419 );
or \U$357 ( \421 , \417 , \420 );
nand \U$358 ( \422 , \418 , \419 );
nand \U$359 ( \423 , \421 , \422 );
and \U$360 ( \424 , \406 , \423 );
and \U$361 ( \425 , \403 , \405 );
or \U$362 ( \426 , \424 , \425 );
not \U$363 ( \427 , \426 );
not \U$364 ( \428 , \427 );
not \U$365 ( \429 , \242 );
not \U$366 ( \430 , \226 );
or \U$367 ( \431 , \429 , \430 );
or \U$368 ( \432 , \242 , \226 );
nand \U$369 ( \433 , \431 , \432 );
not \U$370 ( \434 , \433 );
not \U$371 ( \435 , \434 );
or \U$372 ( \436 , \428 , \435 );
nand \U$373 ( \437 , \433 , \426 );
nand \U$374 ( \438 , \436 , \437 );
not \U$375 ( \439 , \438 );
or \U$376 ( \440 , \396 , \439 );
nand \U$377 ( \441 , \433 , \427 );
nand \U$378 ( \442 , \440 , \441 );
not \U$379 ( \443 , \442 );
xor \U$380 ( \444 , \141 , \203 );
xor \U$381 ( \445 , \444 , \246 );
not \U$382 ( \446 , \445 );
xor \U$383 ( \447 , \158 , \161 );
xor \U$384 ( \448 , \447 , \176 );
not \U$385 ( \449 , \448 );
xor \U$386 ( \450 , \146 , \143 );
xnor \U$387 ( \451 , \450 , \154 );
not \U$388 ( \452 , \451 );
not \U$389 ( \453 , \452 );
or \U$390 ( \454 , \449 , \453 );
not \U$391 ( \455 , \355 );
not \U$392 ( \456 , \350 );
or \U$393 ( \457 , \455 , \456 );
not \U$394 ( \458 , \354 );
nand \U$395 ( \459 , \458 , \353 );
nand \U$396 ( \460 , \457 , \459 );
nand \U$397 ( \461 , \454 , \460 );
not \U$398 ( \462 , \448 );
nand \U$399 ( \463 , \462 , \451 );
and \U$400 ( \464 , \461 , \463 );
not \U$401 ( \465 , \464 );
nand \U$402 ( \466 , \446 , \465 );
nand \U$403 ( \467 , \443 , \466 );
nand \U$404 ( \468 , \445 , \464 );
nand \U$405 ( \469 , \467 , \468 );
not \U$406 ( \470 , \469 );
not \U$407 ( \471 , \249 );
not \U$408 ( \472 , \471 );
not \U$409 ( \473 , \292 );
or \U$410 ( \474 , \472 , \473 );
nand \U$411 ( \475 , \291 , \249 );
nand \U$412 ( \476 , \474 , \475 );
not \U$413 ( \477 , \476 );
nand \U$414 ( \478 , \470 , \477 );
nand \U$415 ( \479 , \346 , \478 );
not \U$416 ( \480 , \340 );
not \U$417 ( \481 , \480 );
not \U$418 ( \482 , \335 );
or \U$419 ( \483 , \481 , \482 );
not \U$420 ( \484 , \330 );
nand \U$421 ( \485 , \484 , \301 );
nand \U$422 ( \486 , \483 , \485 );
not \U$423 ( \487 , \91 );
not \U$424 ( \488 , \101 );
and \U$425 ( \489 , \487 , \488 );
and \U$426 ( \490 , \91 , \101 );
nor \U$427 ( \491 , \489 , \490 );
and \U$428 ( \492 , \305 , \306 );
and \U$429 ( \493 , \304 , \303 );
nor \U$430 ( \494 , \492 , \493 );
xnor \U$431 ( \495 , \491 , \494 );
not \U$432 ( \496 , \320 );
not \U$433 ( \497 , \323 );
and \U$434 ( \498 , \496 , \497 );
not \U$435 ( \499 , \311 );
and \U$436 ( \500 , \325 , \499 );
nor \U$437 ( \501 , \498 , \500 );
xor \U$438 ( \502 , \495 , \501 );
nand \U$439 ( \503 , \486 , \502 );
or \U$440 ( \504 , \501 , \495 );
or \U$441 ( \505 , \491 , \494 );
nand \U$442 ( \506 , \504 , \505 );
not \U$443 ( \507 , \109 );
not \U$444 ( \508 , \105 );
or \U$445 ( \509 , \507 , \508 );
or \U$446 ( \510 , \105 , \109 );
nand \U$447 ( \511 , \509 , \510 );
nand \U$448 ( \512 , \506 , \511 );
nand \U$449 ( \513 , \503 , \512 );
nor \U$450 ( \514 , \479 , \513 );
not \U$451 ( \515 , \514 );
and \U$452 ( \516 , \123 , RIa139a28_37);
not \U$453 ( \517 , \516 );
not \U$454 ( \518 , \415 );
and \U$455 ( \519 , \518 , RIa139848_33);
not \U$456 ( \520 , \519 );
or \U$457 ( \521 , \517 , \520 );
not \U$458 ( \522 , RIa138d80_10);
not \U$459 ( \523 , \168 );
or \U$460 ( \524 , \522 , \523 );
and \U$461 ( \525 , RIa139230_20, RIa139f50_48);
and \U$462 ( \526 , RIa1396e0_30, RIa139ed8_47);
nor \U$463 ( \527 , \525 , \526 );
nand \U$464 ( \528 , \524 , \527 );
buf \U$465 ( \529 , \528 );
nand \U$466 ( \530 , \529 , RIa1397d0_32);
nand \U$467 ( \531 , \521 , \530 );
not \U$468 ( \532 , \516 );
not \U$469 ( \533 , \519 );
nand \U$470 ( \534 , \532 , \533 );
and \U$471 ( \535 , \531 , \534 );
not \U$472 ( \536 , \535 );
and \U$473 ( \537 , \215 , RIa139938_35);
not \U$474 ( \538 , \537 );
not \U$475 ( \539 , RIa139aa0_38);
not \U$476 ( \540 , \175 );
or \U$477 ( \541 , \539 , \540 );
nand \U$478 ( \542 , \134 , RIa1399b0_36);
nand \U$479 ( \543 , \541 , \542 );
not \U$480 ( \544 , \543 );
or \U$481 ( \545 , \538 , \544 );
and \U$482 ( \546 , \134 , RIa139aa0_38);
nand \U$483 ( \547 , \418 , \546 );
nand \U$484 ( \548 , \545 , \547 );
not \U$485 ( \549 , \548 );
nand \U$486 ( \550 , \87 , RIa139b90_40);
not \U$487 ( \551 , \550 );
nand \U$488 ( \552 , \551 , \349 );
not \U$489 ( \553 , \552 );
and \U$490 ( \554 , \549 , \553 );
and \U$491 ( \555 , \548 , \552 );
nor \U$492 ( \556 , \554 , \555 );
nor \U$493 ( \557 , \536 , \556 );
not \U$494 ( \558 , \557 );
and \U$495 ( \559 , \216 , RIa1398c0_34);
and \U$496 ( \560 , \134 , RIa139938_35);
and \U$497 ( \561 , \559 , \560 );
not \U$498 ( \562 , \559 );
not \U$499 ( \563 , \560 );
and \U$500 ( \564 , \562 , \563 );
nor \U$501 ( \565 , \561 , \564 );
not \U$502 ( \566 , \565 );
nor \U$503 ( \567 , \348 , \380 );
or \U$504 ( \568 , \567 , \381 );
not \U$505 ( \569 , \568 );
not \U$506 ( \570 , \569 );
and \U$507 ( \571 , \566 , \570 );
and \U$508 ( \572 , \565 , \569 );
nor \U$509 ( \573 , \571 , \572 );
not \U$510 ( \574 , \535 );
nand \U$511 ( \575 , \556 , \574 );
nand \U$512 ( \576 , \558 , \573 , \575 );
and \U$513 ( \577 , \122 , RIa139aa0_38);
and \U$514 ( \578 , \236 , RIa139938_35);
xor \U$515 ( \579 , \577 , \578 );
and \U$516 ( \580 , \518 , RIa1398c0_34);
and \U$517 ( \581 , \579 , \580 );
and \U$518 ( \582 , \577 , \578 );
or \U$519 ( \583 , \581 , \582 );
not \U$520 ( \584 , \583 );
not \U$521 ( \585 , \584 );
not \U$522 ( \586 , RIa139848_33);
not \U$523 ( \587 , \529 );
or \U$524 ( \588 , \586 , \587 );
nand \U$525 ( \589 , \134 , RIa139a28_37);
nand \U$526 ( \590 , \588 , \589 );
not \U$527 ( \591 , \590 );
and \U$528 ( \592 , \216 , RIa1399b0_36);
not \U$529 ( \593 , \592 );
or \U$530 ( \594 , \591 , \593 );
and \U$531 ( \595 , \528 , RIa139a28_37);
nand \U$532 ( \596 , \595 , \354 );
nand \U$533 ( \597 , \594 , \596 );
not \U$534 ( \598 , \597 );
not \U$535 ( \599 , \598 );
or \U$536 ( \600 , \585 , \599 );
or \U$537 ( \601 , \584 , \598 );
buf \U$538 ( \602 , \543 );
nand \U$539 ( \603 , \547 , \602 );
buf \U$540 ( \604 , \537 );
and \U$541 ( \605 , \603 , \604 );
not \U$542 ( \606 , \603 );
not \U$543 ( \607 , \604 );
and \U$544 ( \608 , \606 , \607 );
nor \U$545 ( \609 , \605 , \608 );
nand \U$546 ( \610 , \601 , \609 );
nand \U$547 ( \611 , \600 , \610 );
and \U$548 ( \612 , \576 , \611 );
not \U$549 ( \613 , \557 );
and \U$550 ( \614 , \575 , \613 );
nor \U$551 ( \615 , \614 , \573 );
nor \U$552 ( \616 , \612 , \615 );
not \U$553 ( \617 , \616 );
not \U$554 ( \618 , \556 );
not \U$555 ( \619 , \535 );
and \U$556 ( \620 , \618 , \619 );
not \U$557 ( \621 , \552 );
nor \U$558 ( \622 , \621 , \548 );
nor \U$559 ( \623 , \620 , \622 );
not \U$560 ( \624 , \623 );
not \U$561 ( \625 , \422 );
nor \U$562 ( \626 , \625 , \420 );
xor \U$563 ( \627 , \626 , \417 );
not \U$564 ( \628 , \568 );
not \U$565 ( \629 , \565 );
or \U$566 ( \630 , \628 , \629 );
not \U$567 ( \631 , \559 );
nand \U$568 ( \632 , \631 , \563 );
nand \U$569 ( \633 , \630 , \632 );
xor \U$570 ( \634 , \627 , \633 );
not \U$571 ( \635 , \634 );
and \U$572 ( \636 , \624 , \635 );
and \U$573 ( \637 , \623 , \634 );
nor \U$574 ( \638 , \636 , \637 );
not \U$575 ( \639 , \638 );
not \U$576 ( \640 , \639 );
or \U$577 ( \641 , \617 , \640 );
not \U$578 ( \642 , \616 );
nand \U$579 ( \643 , \642 , \638 );
nand \U$580 ( \644 , \641 , \643 );
not \U$581 ( \645 , \386 );
and \U$582 ( \646 , \376 , \645 );
not \U$583 ( \647 , \376 );
and \U$584 ( \648 , \647 , \386 );
nor \U$585 ( \649 , \646 , \648 );
nand \U$586 ( \650 , \236 , RIa139848_33);
and \U$587 ( \651 , \174 , RIa139a28_37);
and \U$588 ( \652 , \650 , \651 );
not \U$589 ( \653 , \650 );
not \U$590 ( \654 , \651 );
and \U$591 ( \655 , \653 , \654 );
nor \U$592 ( \656 , \652 , \655 );
nand \U$593 ( \657 , \416 , RIa1397d0_32);
xor \U$594 ( \658 , \656 , \657 );
not \U$595 ( \659 , \658 );
nand \U$596 ( \660 , \122 , RIa1399b0_36);
nand \U$597 ( \661 , \528 , RIa139758_31);
xor \U$598 ( \662 , \660 , \661 );
nand \U$599 ( \663 , \87 , RIa139aa0_38);
xor \U$600 ( \664 , \662 , \663 );
nand \U$601 ( \665 , \659 , \664 );
not \U$602 ( \666 , \665 );
and \U$603 ( \667 , \175 , RIa139b18_39);
not \U$604 ( \668 , \667 );
nor \U$605 ( \669 , \668 , \550 );
not \U$606 ( \670 , \669 );
and \U$607 ( \671 , \236 , RIa1398c0_34);
not \U$608 ( \672 , \671 );
and \U$609 ( \673 , \86 , RIa139b18_39);
nand \U$610 ( \674 , \100 , RIa139b90_40);
xor \U$611 ( \675 , \673 , \674 );
not \U$612 ( \676 , \675 );
or \U$613 ( \677 , \672 , \676 );
or \U$614 ( \678 , \675 , \671 );
nand \U$615 ( \679 , \677 , \678 );
not \U$616 ( \680 , \679 );
or \U$617 ( \681 , \670 , \680 );
not \U$618 ( \682 , \675 );
nand \U$619 ( \683 , \682 , \671 );
nand \U$620 ( \684 , \681 , \683 );
not \U$621 ( \685 , \684 );
or \U$622 ( \686 , \666 , \685 );
not \U$623 ( \687 , \664 );
nand \U$624 ( \688 , \687 , \658 );
nand \U$625 ( \689 , \686 , \688 );
xor \U$626 ( \690 , \649 , \689 );
xor \U$627 ( \691 , \660 , \661 );
and \U$628 ( \692 , \691 , \663 );
and \U$629 ( \693 , \660 , \661 );
or \U$630 ( \694 , \692 , \693 );
not \U$631 ( \695 , \694 );
xor \U$632 ( \696 , \397 , \398 );
xor \U$633 ( \697 , \696 , \400 );
not \U$634 ( \698 , \697 );
or \U$635 ( \699 , \695 , \698 );
or \U$636 ( \700 , \694 , \697 );
nand \U$637 ( \701 , \699 , \700 );
buf \U$638 ( \702 , \650 );
or \U$639 ( \703 , \657 , \702 );
nand \U$640 ( \704 , \703 , \654 );
nand \U$641 ( \705 , \657 , \702 );
nand \U$642 ( \706 , \704 , \705 );
and \U$643 ( \707 , \701 , \706 );
not \U$644 ( \708 , \701 );
not \U$645 ( \709 , \706 );
and \U$646 ( \710 , \708 , \709 );
or \U$647 ( \711 , \707 , \710 );
xor \U$648 ( \712 , \690 , \711 );
not \U$649 ( \713 , \712 );
and \U$650 ( \714 , \644 , \713 );
not \U$651 ( \715 , \644 );
and \U$652 ( \716 , \715 , \712 );
nor \U$653 ( \717 , \714 , \716 );
not \U$654 ( \718 , \717 );
not \U$655 ( \719 , \658 );
not \U$656 ( \720 , \664 );
and \U$657 ( \721 , \719 , \720 );
and \U$658 ( \722 , \658 , \664 );
nor \U$659 ( \723 , \721 , \722 );
xor \U$660 ( \724 , \723 , \684 );
not \U$661 ( \725 , \724 );
not \U$662 ( \726 , \725 );
buf \U$663 ( \727 , \546 );
not \U$664 ( \728 , \727 );
not \U$665 ( \729 , RIa139a28_37);
not \U$666 ( \730 , \216 );
or \U$667 ( \731 , \729 , \730 );
buf \U$668 ( \732 , \236 );
nand \U$669 ( \733 , \732 , RIa1399b0_36);
nand \U$670 ( \734 , \731 , \733 );
not \U$671 ( \735 , \734 );
or \U$672 ( \736 , \728 , \735 );
nand \U$673 ( \737 , \732 , RIa139a28_37);
not \U$674 ( \738 , \737 );
nand \U$675 ( \739 , \738 , \592 );
nand \U$676 ( \740 , \736 , \739 );
not \U$677 ( \741 , \740 );
not \U$678 ( \742 , \550 );
not \U$679 ( \743 , \667 );
and \U$680 ( \744 , \742 , \743 );
and \U$681 ( \745 , \550 , \667 );
nor \U$682 ( \746 , \744 , \745 );
not \U$683 ( \747 , \746 );
and \U$684 ( \748 , \123 , RIa139b90_40);
nand \U$685 ( \749 , \667 , \748 );
not \U$686 ( \750 , \749 );
not \U$687 ( \751 , \750 );
or \U$688 ( \752 , \747 , \751 );
or \U$689 ( \753 , \746 , \750 );
nand \U$690 ( \754 , \752 , \753 );
not \U$691 ( \755 , \754 );
or \U$692 ( \756 , \741 , \755 );
not \U$693 ( \757 , \746 );
nand \U$694 ( \758 , \757 , \750 );
nand \U$695 ( \759 , \756 , \758 );
buf \U$696 ( \760 , \519 );
not \U$697 ( \761 , \760 );
xnor \U$698 ( \762 , \516 , \530 );
not \U$699 ( \763 , \762 );
or \U$700 ( \764 , \761 , \763 );
or \U$701 ( \765 , \760 , \762 );
nand \U$702 ( \766 , \764 , \765 );
not \U$703 ( \767 , \766 );
or \U$704 ( \768 , \759 , \767 );
xor \U$705 ( \769 , \669 , \679 );
nand \U$706 ( \770 , \768 , \769 );
nand \U$707 ( \771 , \759 , \767 );
nand \U$708 ( \772 , \770 , \771 );
not \U$709 ( \773 , \772 );
or \U$710 ( \774 , \726 , \773 );
xor \U$711 ( \775 , \556 , \611 );
not \U$712 ( \776 , \574 );
not \U$713 ( \777 , \573 );
or \U$714 ( \778 , \776 , \777 );
or \U$715 ( \779 , \574 , \573 );
nand \U$716 ( \780 , \778 , \779 );
xor \U$717 ( \781 , \775 , \780 );
not \U$718 ( \782 , \781 );
nand \U$719 ( \783 , \774 , \782 );
or \U$720 ( \784 , \772 , \725 );
nand \U$721 ( \785 , \783 , \784 );
not \U$722 ( \786 , \785 );
nand \U$723 ( \787 , \718 , \786 );
not \U$724 ( \788 , \787 );
not \U$725 ( \789 , \623 );
and \U$726 ( \790 , \789 , \634 );
and \U$727 ( \791 , \627 , \633 );
nor \U$728 ( \792 , \790 , \791 );
not \U$729 ( \793 , \792 );
xor \U$730 ( \794 , \403 , \405 );
xor \U$731 ( \795 , \794 , \423 );
not \U$732 ( \796 , \795 );
not \U$733 ( \797 , \796 );
not \U$734 ( \798 , \706 );
not \U$735 ( \799 , \701 );
or \U$736 ( \800 , \798 , \799 );
not \U$737 ( \801 , \697 );
nand \U$738 ( \802 , \801 , \694 );
nand \U$739 ( \803 , \800 , \802 );
not \U$740 ( \804 , \803 );
not \U$741 ( \805 , \804 );
or \U$742 ( \806 , \797 , \805 );
nand \U$743 ( \807 , \803 , \795 );
nand \U$744 ( \808 , \806 , \807 );
not \U$745 ( \809 , \808 );
and \U$746 ( \810 , \793 , \809 );
and \U$747 ( \811 , \792 , \808 );
nor \U$748 ( \812 , \810 , \811 );
not \U$749 ( \813 , \812 );
xor \U$750 ( \814 , \649 , \689 );
and \U$751 ( \815 , \814 , \711 );
and \U$752 ( \816 , \649 , \689 );
or \U$753 ( \817 , \815 , \816 );
not \U$754 ( \818 , \391 );
and \U$755 ( \819 , \369 , \818 );
not \U$756 ( \820 , \369 );
and \U$757 ( \821 , \820 , \391 );
nor \U$758 ( \822 , \819 , \821 );
not \U$759 ( \823 , \822 );
and \U$760 ( \824 , \817 , \823 );
not \U$761 ( \825 , \817 );
and \U$762 ( \826 , \825 , \822 );
nor \U$763 ( \827 , \824 , \826 );
not \U$764 ( \828 , \827 );
or \U$765 ( \829 , \813 , \828 );
or \U$766 ( \830 , \827 , \812 );
nand \U$767 ( \831 , \829 , \830 );
not \U$768 ( \832 , \712 );
not \U$769 ( \833 , \616 );
nand \U$770 ( \834 , \833 , \639 );
not \U$771 ( \835 , \834 );
or \U$772 ( \836 , \832 , \835 );
nand \U$773 ( \837 , \638 , \616 );
nand \U$774 ( \838 , \836 , \837 );
nand \U$775 ( \839 , \831 , \838 );
not \U$776 ( \840 , \839 );
or \U$777 ( \841 , \788 , \840 );
and \U$778 ( \842 , \827 , \812 );
nor \U$779 ( \843 , \842 , \838 );
not \U$780 ( \844 , \827 );
not \U$781 ( \845 , \812 );
nand \U$782 ( \846 , \844 , \845 );
nand \U$783 ( \847 , \843 , \846 );
nand \U$784 ( \848 , \841 , \847 );
not \U$785 ( \849 , \823 );
not \U$786 ( \850 , \817 );
not \U$787 ( \851 , \850 );
or \U$788 ( \852 , \849 , \851 );
nand \U$789 ( \853 , \852 , \846 );
and \U$790 ( \854 , \448 , \451 );
not \U$791 ( \855 , \448 );
and \U$792 ( \856 , \855 , \452 );
nor \U$793 ( \857 , \854 , \856 );
not \U$794 ( \858 , \460 );
xor \U$795 ( \859 , \857 , \858 );
not \U$796 ( \860 , \395 );
not \U$797 ( \861 , \438 );
not \U$798 ( \862 , \861 );
or \U$799 ( \863 , \860 , \862 );
not \U$800 ( \864 , \395 );
nand \U$801 ( \865 , \864 , \438 );
nand \U$802 ( \866 , \863 , \865 );
xor \U$803 ( \867 , \859 , \866 );
not \U$804 ( \868 , \792 );
not \U$805 ( \869 , \868 );
not \U$806 ( \870 , \808 );
or \U$807 ( \871 , \869 , \870 );
not \U$808 ( \872 , \804 );
nand \U$809 ( \873 , \872 , \796 );
nand \U$810 ( \874 , \871 , \873 );
xor \U$811 ( \875 , \867 , \874 );
nand \U$812 ( \876 , \853 , \875 );
xor \U$813 ( \877 , \464 , \445 );
xor \U$814 ( \878 , \877 , \442 );
xor \U$815 ( \879 , \859 , \866 );
and \U$816 ( \880 , \879 , \874 );
and \U$817 ( \881 , \859 , \866 );
or \U$818 ( \882 , \880 , \881 );
nand \U$819 ( \883 , \878 , \882 );
nand \U$820 ( \884 , \876 , \883 );
nor \U$821 ( \885 , \848 , \884 );
nor \U$822 ( \886 , \853 , \875 );
nand \U$823 ( \887 , \886 , \883 );
not \U$824 ( \888 , \882 );
not \U$825 ( \889 , \878 );
nand \U$826 ( \890 , \888 , \889 );
nand \U$827 ( \891 , \887 , \890 );
nor \U$828 ( \892 , \885 , \891 );
nand \U$829 ( \893 , \215 , RIa139b18_39);
nand \U$830 ( \894 , \134 , RIa139b90_40);
or \U$831 ( \895 , \893 , \894 );
and \U$832 ( \896 , \529 , RIa139938_35);
and \U$833 ( \897 , \895 , \896 );
not \U$834 ( \898 , \895 );
not \U$835 ( \899 , \896 );
and \U$836 ( \900 , \898 , \899 );
nor \U$837 ( \901 , \897 , \900 );
not \U$838 ( \902 , \901 );
and \U$839 ( \903 , \134 , RIa139b18_39);
xor \U$840 ( \904 , \903 , \748 );
not \U$841 ( \905 , \904 );
and \U$842 ( \906 , \902 , \905 );
and \U$843 ( \907 , \895 , \899 );
nor \U$844 ( \908 , \906 , \907 );
not \U$845 ( \909 , \908 );
nand \U$846 ( \910 , \580 , \896 );
not \U$847 ( \911 , RIa139938_35);
not \U$848 ( \912 , \416 );
not \U$849 ( \913 , \912 );
not \U$850 ( \914 , \913 );
or \U$851 ( \915 , \911 , \914 );
buf \U$852 ( \916 , \529 );
nand \U$853 ( \917 , \916 , RIa1398c0_34);
nand \U$854 ( \918 , \915 , \917 );
nand \U$855 ( \919 , \910 , \918 );
and \U$856 ( \920 , \903 , \748 );
xor \U$857 ( \921 , \919 , \920 );
not \U$858 ( \922 , \921 );
or \U$859 ( \923 , \909 , \922 );
or \U$860 ( \924 , \908 , \921 );
nand \U$861 ( \925 , \923 , \924 );
not \U$862 ( \926 , \925 );
not \U$863 ( \927 , \926 );
and \U$864 ( \928 , RIa139b18_39, \123 );
and \U$865 ( \929 , \192 , RIa139b90_40);
nor \U$866 ( \930 , \928 , \929 );
nor \U$867 ( \931 , \750 , \930 );
not \U$868 ( \932 , \931 );
not \U$869 ( \933 , \737 );
nand \U$870 ( \934 , \416 , RIa1399b0_36);
not \U$871 ( \935 , \934 );
and \U$872 ( \936 , \215 , RIa139aa0_38);
not \U$873 ( \937 , \936 );
or \U$874 ( \938 , \935 , \937 );
or \U$875 ( \939 , \936 , \934 );
nand \U$876 ( \940 , \938 , \939 );
not \U$877 ( \941 , \940 );
or \U$878 ( \942 , \933 , \941 );
not \U$879 ( \943 , \936 );
nand \U$880 ( \944 , \943 , \934 );
nand \U$881 ( \945 , \942 , \944 );
not \U$882 ( \946 , \945 );
or \U$883 ( \947 , \932 , \946 );
or \U$884 ( \948 , \945 , \931 );
nand \U$885 ( \949 , \947 , \948 );
not \U$886 ( \950 , \949 );
nand \U$887 ( \951 , \739 , \734 );
not \U$888 ( \952 , \727 );
and \U$889 ( \953 , \951 , \952 );
not \U$890 ( \954 , \951 );
and \U$891 ( \955 , \954 , \727 );
nor \U$892 ( \956 , \953 , \955 );
not \U$893 ( \957 , \956 );
and \U$894 ( \958 , \950 , \957 );
and \U$895 ( \959 , \949 , \956 );
nor \U$896 ( \960 , \958 , \959 );
not \U$897 ( \961 , \960 );
not \U$898 ( \962 , \961 );
or \U$899 ( \963 , \927 , \962 );
nand \U$900 ( \964 , \960 , \925 );
nand \U$901 ( \965 , \963 , \964 );
xnor \U$902 ( \966 , \904 , \901 );
not \U$903 ( \967 , \966 );
not \U$904 ( \968 , \967 );
nand \U$905 ( \969 , \913 , RIa139a28_37);
not \U$906 ( \970 , \969 );
and \U$907 ( \971 , \528 , RIa1399b0_36);
not \U$908 ( \972 , \971 );
not \U$909 ( \973 , \972 );
and \U$910 ( \974 , \236 , RIa139aa0_38);
not \U$911 ( \975 , \974 );
or \U$912 ( \976 , \973 , \975 );
not \U$913 ( \977 , \974 );
nand \U$914 ( \978 , \977 , \971 );
nand \U$915 ( \979 , \976 , \978 );
not \U$916 ( \980 , \979 );
or \U$917 ( \981 , \970 , \980 );
nand \U$918 ( \982 , \977 , \972 );
nand \U$919 ( \983 , \981 , \982 );
not \U$920 ( \984 , \983 );
not \U$921 ( \985 , \984 );
not \U$922 ( \986 , \737 );
not \U$923 ( \987 , \940 );
not \U$924 ( \988 , \987 );
or \U$925 ( \989 , \986 , \988 );
not \U$926 ( \990 , \737 );
nand \U$927 ( \991 , \990 , \940 );
nand \U$928 ( \992 , \989 , \991 );
not \U$929 ( \993 , \992 );
or \U$930 ( \994 , \985 , \993 );
or \U$931 ( \995 , \984 , \992 );
nand \U$932 ( \996 , \994 , \995 );
not \U$933 ( \997 , \996 );
or \U$934 ( \998 , \968 , \997 );
not \U$935 ( \999 , \984 );
nand \U$936 ( \1000 , \999 , \992 );
nand \U$937 ( \1001 , \998 , \1000 );
nand \U$938 ( \1002 , \965 , \1001 );
not \U$939 ( \1003 , \1002 );
nand \U$940 ( \1004 , \732 , RIa139b90_40);
nand \U$941 ( \1005 , \529 , RIa139aa0_38);
nor \U$942 ( \1006 , \1004 , \1005 );
xnor \U$943 ( \1007 , \1004 , \1005 );
not \U$944 ( \1008 , \912 );
nand \U$945 ( \1009 , \1008 , RIa139b18_39);
or \U$946 ( \1010 , \1007 , \1009 );
nand \U$947 ( \1011 , \529 , RIa139b90_40);
nor \U$948 ( \1012 , \1011 , \373 );
nand \U$949 ( \1013 , \1008 , \1012 );
nand \U$950 ( \1014 , \1010 , \1013 );
xor \U$951 ( \1015 , \1006 , \1014 );
nand \U$952 ( \1016 , \416 , RIa139aa0_38);
not \U$953 ( \1017 , \1016 );
not \U$954 ( \1018 , \595 );
and \U$955 ( \1019 , \1017 , \1018 );
and \U$956 ( \1020 , \1016 , \595 );
nor \U$957 ( \1021 , \1019 , \1020 );
nand \U$958 ( \1022 , \216 , RIa139b90_40);
not \U$959 ( \1023 , \1022 );
nand \U$960 ( \1024 , \732 , RIa139b18_39);
not \U$961 ( \1025 , \1024 );
and \U$962 ( \1026 , \1023 , \1025 );
and \U$963 ( \1027 , \1022 , \1024 );
nor \U$964 ( \1028 , \1026 , \1027 );
not \U$965 ( \1029 , \1028 );
and \U$966 ( \1030 , \1021 , \1029 );
not \U$967 ( \1031 , \1021 );
and \U$968 ( \1032 , \1031 , \1028 );
nor \U$969 ( \1033 , \1030 , \1032 );
and \U$970 ( \1034 , \1015 , \1033 );
and \U$971 ( \1035 , \1006 , \1014 );
or \U$972 ( \1036 , \1034 , \1035 );
xnor \U$973 ( \1037 , \979 , \969 );
not \U$974 ( \1038 , \1037 );
not \U$975 ( \1039 , \895 );
and \U$976 ( \1040 , \893 , \894 );
nor \U$977 ( \1041 , \1039 , \1040 );
not \U$978 ( \1042 , \1022 );
not \U$979 ( \1043 , \1024 );
nand \U$980 ( \1044 , \1042 , \1043 );
not \U$981 ( \1045 , \1044 );
and \U$982 ( \1046 , \1041 , \1045 );
not \U$983 ( \1047 , \1041 );
and \U$984 ( \1048 , \1047 , \1044 );
nor \U$985 ( \1049 , \1046 , \1048 );
not \U$986 ( \1050 , \1049 );
or \U$987 ( \1051 , \1038 , \1050 );
or \U$988 ( \1052 , \1037 , \1049 );
nand \U$989 ( \1053 , \1051 , \1052 );
not \U$990 ( \1054 , \595 );
not \U$991 ( \1055 , \1054 );
not \U$992 ( \1056 , \1016 );
or \U$993 ( \1057 , \1055 , \1056 );
or \U$994 ( \1058 , \1016 , \1054 );
nand \U$995 ( \1059 , \1058 , \1029 );
nand \U$996 ( \1060 , \1057 , \1059 );
nand \U$997 ( \1061 , \1053 , \1060 );
nand \U$998 ( \1062 , \1036 , \1061 );
not \U$999 ( \1063 , \1053 );
not \U$1000 ( \1064 , \1060 );
nand \U$1001 ( \1065 , \1063 , \1064 );
nand \U$1002 ( \1066 , \1062 , \1065 );
not \U$1003 ( \1067 , \1066 );
not \U$1004 ( \1068 , \966 );
not \U$1005 ( \1069 , \1068 );
not \U$1006 ( \1070 , \996 );
not \U$1007 ( \1071 , \1070 );
or \U$1008 ( \1072 , \1069 , \1071 );
nand \U$1009 ( \1073 , \996 , \966 );
nand \U$1010 ( \1074 , \1072 , \1073 );
not \U$1011 ( \1075 , \1037 );
not \U$1012 ( \1076 , \1075 );
not \U$1013 ( \1077 , \1049 );
or \U$1014 ( \1078 , \1076 , \1077 );
not \U$1015 ( \1079 , \1041 );
nand \U$1016 ( \1080 , \1079 , \1044 );
nand \U$1017 ( \1081 , \1078 , \1080 );
nand \U$1018 ( \1082 , \1074 , \1081 );
not \U$1019 ( \1083 , \1082 );
or \U$1020 ( \1084 , \1067 , \1083 );
not \U$1021 ( \1085 , \1074 );
not \U$1022 ( \1086 , \1081 );
nand \U$1023 ( \1087 , \1085 , \1086 );
nand \U$1024 ( \1088 , \1084 , \1087 );
not \U$1025 ( \1089 , \1088 );
or \U$1026 ( \1090 , \1003 , \1089 );
not \U$1027 ( \1091 , \965 );
not \U$1028 ( \1092 , \1001 );
nand \U$1029 ( \1093 , \1091 , \1092 );
nand \U$1030 ( \1094 , \1090 , \1093 );
not \U$1031 ( \1095 , \740 );
and \U$1032 ( \1096 , \754 , \1095 );
not \U$1033 ( \1097 , \754 );
and \U$1034 ( \1098 , \1097 , \740 );
nor \U$1035 ( \1099 , \1096 , \1098 );
xor \U$1036 ( \1100 , \577 , \578 );
xor \U$1037 ( \1101 , \1100 , \580 );
not \U$1038 ( \1102 , \1101 );
not \U$1039 ( \1103 , \1102 );
nand \U$1040 ( \1104 , \596 , \590 );
and \U$1041 ( \1105 , \1104 , \592 );
not \U$1042 ( \1106 , \1104 );
not \U$1043 ( \1107 , \592 );
and \U$1044 ( \1108 , \1106 , \1107 );
nor \U$1045 ( \1109 , \1105 , \1108 );
not \U$1046 ( \1110 , \1109 );
not \U$1047 ( \1111 , \1110 );
or \U$1048 ( \1112 , \1103 , \1111 );
nand \U$1049 ( \1113 , \1109 , \1101 );
nand \U$1050 ( \1114 , \1112 , \1113 );
not \U$1051 ( \1115 , \918 );
not \U$1052 ( \1116 , \920 );
or \U$1053 ( \1117 , \1115 , \1116 );
nand \U$1054 ( \1118 , \1117 , \910 );
not \U$1055 ( \1119 , \1118 );
and \U$1056 ( \1120 , \1114 , \1119 );
not \U$1057 ( \1121 , \1114 );
and \U$1058 ( \1122 , \1121 , \1118 );
nor \U$1059 ( \1123 , \1120 , \1122 );
xor \U$1060 ( \1124 , \1099 , \1123 );
not \U$1061 ( \1125 , \956 );
not \U$1062 ( \1126 , \1125 );
not \U$1063 ( \1127 , \949 );
or \U$1064 ( \1128 , \1126 , \1127 );
not \U$1065 ( \1129 , \931 );
nand \U$1066 ( \1130 , \1129 , \945 );
nand \U$1067 ( \1131 , \1128 , \1130 );
xor \U$1068 ( \1132 , \1124 , \1131 );
not \U$1069 ( \1133 , \1132 );
not \U$1070 ( \1134 , \925 );
not \U$1071 ( \1135 , \961 );
or \U$1072 ( \1136 , \1134 , \1135 );
not \U$1073 ( \1137 , \908 );
nand \U$1074 ( \1138 , \1137 , \921 );
nand \U$1075 ( \1139 , \1136 , \1138 );
not \U$1076 ( \1140 , \1139 );
nand \U$1077 ( \1141 , \1133 , \1140 );
not \U$1078 ( \1142 , \1141 );
or \U$1079 ( \1143 , \1094 , \1142 );
and \U$1080 ( \1144 , \583 , \597 );
not \U$1081 ( \1145 , \583 );
and \U$1082 ( \1146 , \1145 , \598 );
nor \U$1083 ( \1147 , \1144 , \1146 );
not \U$1084 ( \1148 , \609 );
xnor \U$1085 ( \1149 , \1147 , \1148 );
not \U$1086 ( \1150 , \1149 );
not \U$1087 ( \1151 , \1102 );
not \U$1088 ( \1152 , \1109 );
or \U$1089 ( \1153 , \1151 , \1152 );
nand \U$1090 ( \1154 , \1153 , \1118 );
nand \U$1091 ( \1155 , \1110 , \1101 );
nand \U$1092 ( \1156 , \1154 , \1155 );
not \U$1093 ( \1157 , \1156 );
and \U$1094 ( \1158 , \1150 , \1157 );
and \U$1095 ( \1159 , \1149 , \1156 );
nor \U$1096 ( \1160 , \1158 , \1159 );
not \U$1097 ( \1161 , \1160 );
not \U$1098 ( \1162 , \759 );
not \U$1099 ( \1163 , \1162 );
not \U$1100 ( \1164 , \766 );
not \U$1101 ( \1165 , \769 );
or \U$1102 ( \1166 , \1164 , \1165 );
or \U$1103 ( \1167 , \769 , \766 );
nand \U$1104 ( \1168 , \1166 , \1167 );
not \U$1105 ( \1169 , \1168 );
or \U$1106 ( \1170 , \1163 , \1169 );
or \U$1107 ( \1171 , \1168 , \1162 );
nand \U$1108 ( \1172 , \1170 , \1171 );
not \U$1109 ( \1173 , \1172 );
and \U$1110 ( \1174 , \1161 , \1173 );
and \U$1111 ( \1175 , \1160 , \1172 );
nor \U$1112 ( \1176 , \1174 , \1175 );
xor \U$1113 ( \1177 , \1099 , \1123 );
and \U$1114 ( \1178 , \1177 , \1131 );
and \U$1115 ( \1179 , \1099 , \1123 );
or \U$1116 ( \1180 , \1178 , \1179 );
nand \U$1117 ( \1181 , \1176 , \1180 );
nand \U$1118 ( \1182 , \1132 , \1139 );
and \U$1119 ( \1183 , \1181 , \1182 );
nand \U$1120 ( \1184 , \1143 , \1183 );
xor \U$1121 ( \1185 , \724 , \772 );
xnor \U$1122 ( \1186 , \1185 , \781 );
not \U$1123 ( \1187 , \1172 );
not \U$1124 ( \1188 , \1160 );
not \U$1125 ( \1189 , \1188 );
or \U$1126 ( \1190 , \1187 , \1189 );
not \U$1127 ( \1191 , \1149 );
nand \U$1128 ( \1192 , \1191 , \1156 );
nand \U$1129 ( \1193 , \1190 , \1192 );
nand \U$1130 ( \1194 , \1186 , \1193 );
not \U$1131 ( \1195 , \1176 );
not \U$1132 ( \1196 , \1180 );
nand \U$1133 ( \1197 , \1195 , \1196 );
nand \U$1134 ( \1198 , \1194 , \1197 );
not \U$1135 ( \1199 , \1198 );
nand \U$1136 ( \1200 , \1184 , \1199 );
nand \U$1137 ( \1201 , \843 , \846 );
not \U$1138 ( \1202 , \1201 );
not \U$1139 ( \1203 , \1186 );
not \U$1140 ( \1204 , \1193 );
nand \U$1141 ( \1205 , \1203 , \1204 );
nand \U$1142 ( \1206 , \717 , \785 );
nand \U$1143 ( \1207 , \1205 , \1206 );
nor \U$1144 ( \1208 , \1202 , \1207 );
nand \U$1145 ( \1209 , \1200 , \1208 );
not \U$1146 ( \1210 , \1209 );
not \U$1147 ( \1211 , \884 );
nand \U$1148 ( \1212 , \1210 , \1211 );
nand \U$1149 ( \1213 , \892 , \1212 );
not \U$1150 ( \1214 , \1213 );
or \U$1151 ( \1215 , \515 , \1214 );
not \U$1152 ( \1216 , \503 );
nor \U$1153 ( \1217 , \1216 , \345 );
not \U$1154 ( \1218 , \1217 );
not \U$1155 ( \1219 , \344 );
not \U$1156 ( \1220 , \296 );
or \U$1157 ( \1221 , \1219 , \1220 );
nand \U$1158 ( \1222 , \469 , \476 );
nand \U$1159 ( \1223 , \1221 , \1222 );
not \U$1160 ( \1224 , \1223 );
or \U$1161 ( \1225 , \1218 , \1224 );
or \U$1162 ( \1226 , \486 , \502 );
nand \U$1163 ( \1227 , \1225 , \1226 );
and \U$1164 ( \1228 , \1227 , \512 );
nor \U$1165 ( \1229 , \506 , \511 );
nor \U$1166 ( \1230 , \1228 , \1229 );
nand \U$1167 ( \1231 , \1215 , \1230 );
not \U$1168 ( \1232 , \1231 );
or \U$1169 ( \1233 , \115 , \1232 );
nand \U$1170 ( \1234 , \112 , \113 );
nand \U$1171 ( \1235 , \1233 , \1234 );
buf \U$1172 ( \1236 , \1235 );
nand \U$1173 ( \1237 , \1234 , \114 );
not \U$1174 ( \1238 , \1237 );
not \U$1175 ( \1239 , \1231 );
or \U$1176 ( \1240 , \1238 , \1239 );
or \U$1177 ( \1241 , \1231 , \1237 );
nand \U$1178 ( \1242 , \1240 , \1241 );
buf \U$1179 ( \1243 , \1242 );
not \U$1180 ( \1244 , \503 );
nor \U$1181 ( \1245 , \479 , \884 );
not \U$1182 ( \1246 , \1245 );
nand \U$1183 ( \1247 , \848 , \1209 );
not \U$1184 ( \1248 , \1247 );
or \U$1185 ( \1249 , \1246 , \1248 );
and \U$1186 ( \1250 , \888 , \889 );
nor \U$1187 ( \1251 , \1250 , \1223 );
not \U$1188 ( \1252 , \1251 );
not \U$1189 ( \1253 , \887 );
or \U$1190 ( \1254 , \1252 , \1253 );
not \U$1191 ( \1255 , \1223 );
not \U$1192 ( \1256 , \478 );
and \U$1193 ( \1257 , \1255 , \1256 );
nor \U$1194 ( \1258 , \1257 , \345 );
nand \U$1195 ( \1259 , \1254 , \1258 );
nand \U$1196 ( \1260 , \1249 , \1259 );
not \U$1197 ( \1261 , \1260 );
or \U$1198 ( \1262 , \1244 , \1261 );
nand \U$1199 ( \1263 , \1262 , \1226 );
not \U$1200 ( \1264 , \1229 );
nand \U$1201 ( \1265 , \1264 , \512 );
not \U$1202 ( \1266 , \1265 );
and \U$1203 ( \1267 , \1263 , \1266 );
not \U$1204 ( \1268 , \1263 );
and \U$1205 ( \1269 , \1268 , \1265 );
nor \U$1206 ( \1270 , \1267 , \1269 );
buf \U$1207 ( \1271 , \1270 );
nand \U$1208 ( \1272 , \1226 , \503 );
not \U$1209 ( \1273 , \1272 );
and \U$1210 ( \1274 , \1260 , \1273 );
not \U$1211 ( \1275 , \1260 );
and \U$1212 ( \1276 , \1275 , \1272 );
nor \U$1213 ( \1277 , \1274 , \1276 );
buf \U$1214 ( \1278 , \1277 );
buf \U$1215 ( \1279 , \478 );
not \U$1216 ( \1280 , \1279 );
not \U$1217 ( \1281 , \1213 );
or \U$1218 ( \1282 , \1280 , \1281 );
nand \U$1219 ( \1283 , \1282 , \1222 );
and \U$1220 ( \1284 , \344 , \296 );
not \U$1221 ( \1285 , \344 );
not \U$1222 ( \1286 , \296 );
and \U$1223 ( \1287 , \1285 , \1286 );
nor \U$1224 ( \1288 , \1284 , \1287 );
and \U$1225 ( \1289 , \1283 , \1288 );
not \U$1226 ( \1290 , \1283 );
not \U$1227 ( \1291 , \1288 );
and \U$1228 ( \1292 , \1290 , \1291 );
nor \U$1229 ( \1293 , \1289 , \1292 );
buf \U$1230 ( \1294 , \1293 );
nand \U$1231 ( \1295 , \1279 , \1222 );
xnor \U$1232 ( \1296 , \1295 , \1213 );
buf \U$1233 ( \1297 , \1296 );
buf \U$1234 ( \1298 , \876 );
not \U$1235 ( \1299 , \1298 );
not \U$1236 ( \1300 , \1247 );
or \U$1237 ( \1301 , \1299 , \1300 );
buf \U$1238 ( \1302 , \886 );
not \U$1239 ( \1303 , \1302 );
nand \U$1240 ( \1304 , \1301 , \1303 );
nand \U$1241 ( \1305 , \883 , \890 );
not \U$1242 ( \1306 , \1305 );
and \U$1243 ( \1307 , \1304 , \1306 );
not \U$1244 ( \1308 , \1304 );
and \U$1245 ( \1309 , \1308 , \1305 );
nor \U$1246 ( \1310 , \1307 , \1309 );
buf \U$1247 ( \1311 , \1310 );
not \U$1248 ( \1312 , \1302 );
nand \U$1249 ( \1313 , \1312 , \1298 );
not \U$1250 ( \1314 , \1313 );
and \U$1251 ( \1315 , \1247 , \1314 );
not \U$1252 ( \1316 , \1247 );
and \U$1253 ( \1317 , \1316 , \1313 );
nor \U$1254 ( \1318 , \1315 , \1317 );
buf \U$1255 ( \1319 , \1318 );
not \U$1256 ( \1320 , \1184 );
not \U$1257 ( \1321 , \1199 );
or \U$1258 ( \1322 , \1320 , \1321 );
nand \U$1259 ( \1323 , \1204 , \1203 );
nand \U$1260 ( \1324 , \1322 , \1323 );
not \U$1261 ( \1325 , \1324 );
buf \U$1262 ( \1326 , \1206 );
not \U$1263 ( \1327 , \1326 );
not \U$1264 ( \1328 , \1327 );
and \U$1265 ( \1329 , \1325 , \1328 );
buf \U$1266 ( \1330 , \787 );
not \U$1267 ( \1331 , \1330 );
nor \U$1268 ( \1332 , \1329 , \1331 );
nand \U$1269 ( \1333 , \847 , \839 );
and \U$1270 ( \1334 , \1332 , \1333 );
not \U$1271 ( \1335 , \1332 );
not \U$1272 ( \1336 , \1333 );
and \U$1273 ( \1337 , \1335 , \1336 );
nor \U$1274 ( \1338 , \1334 , \1337 );
buf \U$1275 ( \1339 , \1338 );
nand \U$1276 ( \1340 , \1330 , \1326 );
and \U$1277 ( \1341 , \1324 , \1340 );
not \U$1278 ( \1342 , \1324 );
not \U$1279 ( \1343 , \1340 );
and \U$1280 ( \1344 , \1342 , \1343 );
nor \U$1281 ( \1345 , \1341 , \1344 );
buf \U$1282 ( \1346 , \1345 );
buf \U$1283 ( \1347 , \1184 );
nand \U$1284 ( \1348 , \1347 , \1197 );
nand \U$1285 ( \1349 , \1323 , \1194 );
not \U$1286 ( \1350 , \1349 );
and \U$1287 ( \1351 , \1348 , \1350 );
not \U$1288 ( \1352 , \1348 );
and \U$1289 ( \1353 , \1352 , \1349 );
nor \U$1290 ( \1354 , \1351 , \1353 );
buf \U$1291 ( \1355 , \1354 );
and \U$1292 ( \1356 , \1094 , \1182 );
nor \U$1293 ( \1357 , \1356 , \1142 );
nand \U$1294 ( \1358 , \1181 , \1197 );
and \U$1295 ( \1359 , \1357 , \1358 );
not \U$1296 ( \1360 , \1357 );
not \U$1297 ( \1361 , \1358 );
and \U$1298 ( \1362 , \1360 , \1361 );
nor \U$1299 ( \1363 , \1359 , \1362 );
buf \U$1300 ( \1364 , \1363 );
nand \U$1301 ( \1365 , \1141 , \1182 );
not \U$1302 ( \1366 , \1094 );
and \U$1303 ( \1367 , \1365 , \1366 );
not \U$1304 ( \1368 , \1365 );
and \U$1305 ( \1369 , \1368 , \1094 );
nor \U$1306 ( \1370 , \1367 , \1369 );
buf \U$1307 ( \1371 , \1370 );
and \U$1308 ( \1372 , \1002 , \1093 );
and \U$1309 ( \1373 , \1372 , \1088 );
not \U$1310 ( \1374 , \1372 );
not \U$1311 ( \1375 , \1088 );
and \U$1312 ( \1376 , \1374 , \1375 );
nor \U$1313 ( \1377 , \1373 , \1376 );
buf \U$1314 ( \1378 , \1377 );
and \U$1315 ( \1379 , \1082 , \1087 );
and \U$1316 ( \1380 , \1379 , \1066 );
not \U$1317 ( \1381 , \1379 );
not \U$1318 ( \1382 , \1066 );
and \U$1319 ( \1383 , \1381 , \1382 );
nor \U$1320 ( \1384 , \1380 , \1383 );
buf \U$1321 ( \1385 , \1384 );
nand \U$1322 ( \1386 , \1065 , \1061 );
not \U$1323 ( \1387 , \1036 );
and \U$1324 ( \1388 , \1386 , \1387 );
not \U$1325 ( \1389 , \1386 );
and \U$1326 ( \1390 , \1389 , \1036 );
nor \U$1327 ( \1391 , \1388 , \1390 );
buf \U$1328 ( \1392 , \1391 );
xor \U$1329 ( \1393 , \1006 , \1014 );
xor \U$1330 ( \1394 , \1393 , \1033 );
buf \U$1331 ( \1395 , \1394 );
not \U$1332 ( \1396 , \1009 );
nand \U$1333 ( \1397 , \1396 , \1013 );
xor \U$1334 ( \1398 , \1397 , \1007 );
buf \U$1335 ( \1399 , \1398 );
not \U$1336 ( \1400 , \1013 );
and \U$1337 ( \1401 , \913 , RIa139b90_40);
and \U$1338 ( \1402 , \916 , RIa139b18_39);
nor \U$1339 ( \1403 , \1401 , \1402 );
nor \U$1340 ( \1404 , \1400 , \1403 );
buf \U$1341 ( \1405 , \1404 );
not \U$1342 ( \1406 , \1011 );
buf \U$1343 ( \1407 , \1406 );
endmodule

