//
// Conformal-LEC Version 20.10-d215 (04-Sep-2020)
//
module top(RIa148a08_33,RIa147bf8_3,RIa148e40_42,RIa148eb8_43,RIa148dc8_41,RIa148fa8_45,RIa148f30_44,RIa149020_46,RIa149098_47,
        RIa149110_48,RIa1480a8_13,RIa148558_23,RIa148a80_34,RIa148030_12,RIa147b80_2,RIa1484e0_22,RIa148af8_35,RIa147fb8_11,RIa147b08_1,
        RIa148468_21,RIa148b70_36,RIa148c60_38,RIa148cd8_39,RIa148d50_40,RIa1485d0_24,RIa147c70_4,RIa148120_14,RIa148198_15,RIa147ce8_5,
        RIa148648_25,RIa148210_16,RIa147d60_6,RIa1486c0_26,RIa1487b0_28,RIa147e50_8,RIa148300_18,RIa1483f0_20,RIa147f40_10,RIa1488a0_30,
        RIa148378_19,RIa147ec8_9,RIa148828_29,RIa148288_17,RIa147dd8_7,RIa148738_27,RIa148be8_37,RIa148990_32,RIa148918_31,R_31_942fc58,
        R_32_942fd00,R_33_942fda8,R_34_942fe50,R_35_942fef8,R_36_942ffa0,R_37_9430048,R_38_94300f0,R_39_9430198,R_3a_9430240,R_3b_94302e8,
        R_3c_9430390);
input RIa148a08_33,RIa147bf8_3,RIa148e40_42,RIa148eb8_43,RIa148dc8_41,RIa148fa8_45,RIa148f30_44,RIa149020_46,RIa149098_47,
        RIa149110_48,RIa1480a8_13,RIa148558_23,RIa148a80_34,RIa148030_12,RIa147b80_2,RIa1484e0_22,RIa148af8_35,RIa147fb8_11,RIa147b08_1,
        RIa148468_21,RIa148b70_36,RIa148c60_38,RIa148cd8_39,RIa148d50_40,RIa1485d0_24,RIa147c70_4,RIa148120_14,RIa148198_15,RIa147ce8_5,
        RIa148648_25,RIa148210_16,RIa147d60_6,RIa1486c0_26,RIa1487b0_28,RIa147e50_8,RIa148300_18,RIa1483f0_20,RIa147f40_10,RIa1488a0_30,
        RIa148378_19,RIa147ec8_9,RIa148828_29,RIa148288_17,RIa147dd8_7,RIa148738_27,RIa148be8_37,RIa148990_32,RIa148918_31;
output R_31_942fc58,R_32_942fd00,R_33_942fda8,R_34_942fe50,R_35_942fef8,R_36_942ffa0,R_37_9430048,R_38_94300f0,R_39_9430198,
        R_3a_9430240,R_3b_94302e8,R_3c_9430390;

wire \55_ZERO , \56_ONE , \57 , \58 , \59 , \60 , \61 , \62 , \63 ,
         \64 , \65 , \66 , \67 , \68 , \69 , \70 , \71 , \72 , \73 ,
         \74 , \75 , \76 , \77 , \78 , \79 , \80 , \81 , \82 , \83 ,
         \84 , \85 , \86 , \87 , \88 , \89 , \90 , \91 , \92 , \93 ,
         \94 , \95 , \96 , \97 , \98 , \99 , \100 , \101 , \102 , \103 ,
         \104 , \105 , \106 , \107 , \108 , \109 , \110 , \111 , \112 , \113 ,
         \114 , \115 , \116 , \117 , \118 , \119 , \120 , \121 , \122 , \123 ,
         \124 , \125 , \126 , \127 , \128 , \129 , \130 , \131 , \132 , \133 ,
         \134 , \135 , \136 , \137 , \138 , \139 , \140 , \141 , \142 , \143 ,
         \144 , \145 , \146 , \147 , \148 , \149 , \150 , \151 , \152 , \153 ,
         \154 , \155 , \156 , \157 , \158 , \159 , \160 , \161 , \162 , \163 ,
         \164 , \165 , \166 , \167 , \168 , \169 , \170 , \171 , \172 , \173 ,
         \174 , \175 , \176 , \177 , \178 , \179 , \180 , \181 , \182 , \183 ,
         \184 , \185 , \186 , \187 , \188 , \189 , \190 , \191 , \192 , \193 ,
         \194 , \195 , \196 , \197 , \198 , \199 , \200 , \201 , \202 , \203 ,
         \204 , \205 , \206 , \207 , \208 , \209 , \210 , \211 , \212 , \213 ,
         \214 , \215 , \216 , \217 , \218 , \219 , \220 , \221 , \222 , \223 ,
         \224 , \225 , \226 , \227 , \228 , \229 , \230 , \231 , \232 , \233 ,
         \234 , \235 , \236 , \237 , \238 , \239 , \240 , \241 , \242 , \243 ,
         \244 , \245 , \246 , \247 , \248 , \249 , \250 , \251 , \252 , \253 ,
         \254 , \255 , \256 , \257 , \258 , \259 , \260 , \261 , \262 , \263 ,
         \264 , \265 , \266 , \267 , \268 , \269 , \270 , \271 , \272 , \273 ,
         \274 , \275 , \276 , \277 , \278 , \279 , \280 , \281 , \282 , \283 ,
         \284 , \285 , \286 , \287 , \288 , \289 , \290 , \291 , \292 , \293 ,
         \294 , \295 , \296 , \297 , \298 , \299 , \300 , \301 , \302 , \303 ,
         \304 , \305 , \306 , \307 , \308 , \309 , \310 , \311 , \312 , \313 ,
         \314 , \315 , \316 , \317 , \318 , \319 , \320 , \321 , \322 , \323 ,
         \324 , \325 , \326 , \327 , \328 , \329 , \330 , \331 , \332 , \333 ,
         \334 , \335 , \336 , \337 , \338 , \339 , \340 , \341 , \342 , \343 ,
         \344 , \345 , \346 , \347 , \348 , \349 , \350 , \351 , \352 , \353 ,
         \354 , \355 , \356 , \357 , \358 , \359 , \360 , \361 , \362 , \363 ,
         \364 , \365 , \366 , \367 , \368 , \369 , \370 , \371 , \372 , \373 ,
         \374 , \375 , \376 , \377 , \378 , \379 , \380 , \381 , \382 , \383 ,
         \384 , \385 , \386 , \387 , \388 , \389 , \390 , \391 , \392 , \393 ,
         \394 , \395 , \396 , \397 , \398 , \399 , \400 , \401 , \402 , \403 ,
         \404 , \405 , \406 , \407 , \408 , \409 , \410 , \411 , \412 , \413 ,
         \414 , \415 , \416 , \417 , \418 , \419 , \420 , \421 , \422 , \423 ,
         \424 , \425 , \426 , \427 , \428 , \429 , \430 , \431 , \432 , \433 ,
         \434 , \435 , \436 , \437 , \438 , \439 , \440 , \441 , \442 , \443 ,
         \444 , \445 , \446 , \447 , \448 , \449 , \450 , \451 , \452 , \453 ,
         \454 , \455 , \456 , \457 , \458 , \459 , \460 , \461 , \462 , \463 ,
         \464 , \465 , \466 , \467 , \468 , \469 , \470 , \471 , \472 , \473 ,
         \474 , \475 , \476 , \477 , \478 , \479 , \480 , \481 , \482 , \483 ,
         \484 , \485 , \486 , \487 , \488 , \489 , \490 , \491 , \492 , \493 ,
         \494 , \495 , \496 , \497 , \498 , \499 , \500 , \501 , \502 , \503 ,
         \504 , \505 , \506 , \507 , \508 , \509 , \510 , \511 , \512 , \513 ,
         \514 , \515 , \516 , \517 , \518 , \519 , \520 , \521 , \522 , \523 ,
         \524 , \525 , \526 , \527 , \528 , \529 , \530 , \531 , \532 , \533 ,
         \534 , \535 , \536 , \537 , \538 , \539 , \540 , \541 , \542 , \543 ,
         \544 , \545 , \546 , \547 , \548 , \549 , \550 , \551 , \552 , \553 ,
         \554 , \555 , \556 , \557 , \558 , \559 , \560 , \561 , \562 , \563 ,
         \564 , \565 , \566 , \567 , \568 , \569 , \570 , \571 , \572 , \573 ,
         \574 , \575 , \576 , \577 , \578 , \579 , \580 , \581 , \582 , \583 ,
         \584 , \585 , \586 , \587 , \588 , \589 , \590 , \591 , \592 , \593 ,
         \594 , \595 , \596 , \597 , \598 , \599 , \600 , \601 , \602 , \603 ,
         \604 , \605 , \606 , \607 , \608 , \609 , \610 , \611 , \612 , \613 ,
         \614 , \615 , \616 , \617 , \618 , \619 , \620 , \621 , \622 , \623 ,
         \624 , \625 , \626 , \627 , \628 , \629 , \630 , \631 , \632 , \633 ,
         \634 , \635 , \636 , \637 , \638 , \639 , \640 , \641 , \642 , \643 ,
         \644 , \645 , \646 , \647 , \648 , \649 , \650 , \651 , \652 , \653 ,
         \654 , \655 , \656 , \657 , \658 , \659 , \660 , \661 , \662 , \663 ,
         \664 , \665 , \666 , \667 , \668 , \669 , \670 , \671 , \672 , \673 ,
         \674 , \675 , \676 , \677 , \678 , \679 , \680 , \681 , \682 , \683 ,
         \684 , \685 , \686 , \687 , \688 , \689 , \690 , \691 , \692 , \693 ,
         \694 , \695 , \696 , \697 , \698 , \699 , \700 , \701 , \702 , \703 ,
         \704 , \705 , \706 , \707 , \708 , \709 , \710 , \711 , \712 , \713 ,
         \714 , \715 , \716 , \717 , \718 , \719 , \720 , \721 , \722 , \723 ,
         \724 , \725 , \726 , \727 , \728 , \729 , \730 , \731 , \732 , \733 ,
         \734 , \735 , \736 , \737 , \738 , \739 , \740 , \741 , \742 , \743 ,
         \744 , \745 , \746 , \747 , \748 , \749 , \750 , \751 , \752 , \753 ,
         \754 , \755 , \756 , \757 , \758 , \759 , \760 , \761 , \762 , \763 ,
         \764 , \765 , \766 , \767 , \768 , \769 , \770 , \771 , \772 , \773 ,
         \774 , \775 , \776 , \777 , \778 , \779 , \780 , \781 , \782 , \783 ,
         \784 , \785 , \786 , \787 , \788 , \789 , \790 , \791 , \792 , \793 ,
         \794 , \795 , \796 , \797 , \798 , \799 , \800 , \801 , \802 , \803 ,
         \804 , \805 , \806 , \807 , \808 , \809 , \810 , \811 , \812 , \813 ,
         \814 , \815 , \816 , \817 , \818 , \819 , \820 , \821 , \822 , \823 ,
         \824 , \825 , \826 , \827 , \828 , \829 , \830 , \831 , \832 , \833 ,
         \834 , \835 , \836 , \837 , \838 , \839 , \840 , \841 , \842 , \843 ,
         \844 , \845 , \846 , \847 , \848 , \849 , \850 , \851 , \852 , \853 ,
         \854 , \855 , \856 , \857 , \858 , \859 , \860 , \861 , \862 , \863 ,
         \864 , \865 , \866 , \867 , \868 , \869 , \870 , \871 , \872 , \873 ,
         \874 , \875 , \876 , \877 , \878 , \879 , \880 , \881 , \882 , \883 ,
         \884 , \885 , \886 , \887 , \888 , \889 , \890 , \891 , \892 , \893 ,
         \894 , \895 , \896 , \897 , \898 , \899 , \900 , \901 , \902 , \903 ,
         \904 , \905 , \906 , \907 , \908 , \909 , \910 , \911 , \912 , \913 ,
         \914 , \915 , \916 , \917 , \918 , \919 , \920 , \921 , \922 , \923 ,
         \924 , \925 , \926 , \927 , \928 , \929 , \930 , \931 , \932 , \933 ,
         \934 , \935 , \936 , \937 , \938 , \939 , \940 , \941 , \942 , \943 ,
         \944 , \945 , \946 , \947 , \948 , \949 , \950 , \951 , \952 , \953 ,
         \954 , \955 , \956 , \957 , \958 , \959 , \960 , \961 , \962 , \963 ,
         \964 , \965 , \966 , \967 , \968 , \969 , \970 , \971 , \972 , \973 ,
         \974 , \975 , \976 , \977 , \978 , \979 , \980 , \981 , \982 , \983 ,
         \984 , \985 , \986 , \987 , \988 , \989 , \990 , \991 , \992 , \993 ,
         \994 , \995 , \996 , \997 , \998 , \999 , \1000 , \1001 , \1002 , \1003 ,
         \1004 , \1005 , \1006 , \1007 , \1008 , \1009 , \1010 , \1011 , \1012 , \1013 ,
         \1014 , \1015 , \1016 , \1017 , \1018 , \1019 , \1020 , \1021 , \1022 , \1023 ,
         \1024 , \1025 , \1026 , \1027 , \1028 , \1029 , \1030 , \1031 , \1032 , \1033 ,
         \1034 , \1035 , \1036 , \1037 , \1038 , \1039 , \1040 , \1041 , \1042 , \1043 ,
         \1044 , \1045 , \1046 , \1047 , \1048 , \1049 , \1050 , \1051 , \1052 , \1053 ,
         \1054 , \1055 , \1056 , \1057 , \1058 , \1059 , \1060 , \1061 , \1062 , \1063 ,
         \1064 , \1065 , \1066 , \1067 , \1068 , \1069 , \1070 , \1071 , \1072 , \1073 ,
         \1074 , \1075 , \1076 , \1077 , \1078 , \1079 , \1080 , \1081 , \1082 , \1083 ,
         \1084 , \1085 , \1086 , \1087 , \1088 , \1089 , \1090 , \1091 , \1092 , \1093 ,
         \1094 , \1095 , \1096 , \1097 , \1098 , \1099 , \1100 , \1101 , \1102 , \1103 ,
         \1104 , \1105 , \1106 , \1107 , \1108 , \1109 , \1110 , \1111 , \1112 , \1113 ,
         \1114 , \1115 , \1116 , \1117 , \1118 , \1119 , \1120 , \1121 , \1122 , \1123 ,
         \1124 , \1125 , \1126 , \1127 , \1128 , \1129 , \1130 , \1131 , \1132 , \1133 ,
         \1134 , \1135 , \1136 , \1137 , \1138 , \1139 , \1140 , \1141 , \1142 , \1143 ,
         \1144 , \1145 , \1146 , \1147 , \1148 , \1149 , \1150 , \1151 , \1152 , \1153 ,
         \1154 , \1155 , \1156 , \1157 , \1158 , \1159 , \1160 , \1161 , \1162 , \1163 ,
         \1164 , \1165 , \1166 , \1167 , \1168 , \1169 , \1170 , \1171 , \1172 , \1173 ,
         \1174 , \1175 , \1176 , \1177 , \1178 , \1179 , \1180 , \1181 , \1182 , \1183 ,
         \1184 , \1185 , \1186 , \1187 , \1188 , \1189 , \1190 , \1191 , \1192 , \1193 ,
         \1194 , \1195 , \1196 , \1197 , \1198 , \1199 , \1200 , \1201 , \1202 , \1203 ,
         \1204 , \1205 , \1206 , \1207 , \1208 , \1209 , \1210 , \1211 , \1212 , \1213 ,
         \1214 , \1215 , \1216 , \1217 , \1218 , \1219 , \1220 , \1221 , \1222 , \1223 ,
         \1224 , \1225 , \1226 , \1227 , \1228 , \1229 , \1230 , \1231 , \1232 , \1233 ,
         \1234 , \1235 , \1236 , \1237 , \1238 , \1239 , \1240 , \1241 , \1242 , \1243 ,
         \1244 , \1245 , \1246 , \1247 , \1248 , \1249 , \1250 , \1251 , \1252 , \1253 ,
         \1254 , \1255 , \1256 , \1257 , \1258 , \1259 , \1260 , \1261 , \1262 , \1263 ,
         \1264 , \1265 , \1266 , \1267 , \1268 , \1269 , \1270 , \1271 , \1272 , \1273 ,
         \1274 , \1275 , \1276 , \1277 , \1278 , \1279 , \1280 , \1281 , \1282 , \1283 ,
         \1284 , \1285 , \1286 , \1287 , \1288 , \1289 , \1290 , \1291 , \1292 , \1293 ,
         \1294 , \1295 , \1296 , \1297 , \1298 , \1299 , \1300 , \1301 , \1302 , \1303 ,
         \1304 , \1305 , \1306 , \1307 , \1308 , \1309 , \1310 , \1311 , \1312 , \1313 ,
         \1314 , \1315 , \1316 , \1317 , \1318 , \1319 , \1320 , \1321 , \1322 , \1323 ,
         \1324 , \1325 , \1326 , \1327 , \1328 , \1329 , \1330 , \1331 , \1332 , \1333 ,
         \1334 , \1335 , \1336 , \1337 , \1338 , \1339 , \1340 , \1341 , \1342 , \1343 ,
         \1344 , \1345 , \1346 , \1347 , \1348 , \1349 , \1350 , \1351 , \1352 , \1353 ,
         \1354 , \1355 , \1356 ;
buf \U$labajz149 ( R_31_942fc58, \1228 );
buf \U$labajz150 ( R_32_942fd00, \1235 );
buf \U$labajz151 ( R_33_942fda8, \1263 );
buf \U$labajz152 ( R_34_942fe50, \1270 );
buf \U$labajz153 ( R_35_942fef8, \1286 );
buf \U$labajz154 ( R_36_942ffa0, \1289 );
buf \U$labajz155 ( R_37_9430048, \1303 );
buf \U$labajz156 ( R_38_94300f0, \1311 );
buf \U$labajz157 ( R_39_9430198, \1331 );
buf \U$labajz158 ( R_3a_9430240, \1338 );
buf \U$labajz159 ( R_3b_94302e8, \1347 );
buf \U$labajz160 ( R_3c_9430390, \1356 );
not \U$1 ( \57 , RIa147b08_1);
nor \U$2 ( \58 , RIa149098_47, RIa149110_48);
not \U$3 ( \59 , \58 );
or \U$4 ( \60 , \57 , \59 );
and \U$5 ( \61 , RIa147fb8_11, RIa149110_48);
and \U$6 ( \62 , RIa148468_21, RIa149098_47);
nor \U$7 ( \63 , \61 , \62 );
nand \U$8 ( \64 , \60 , \63 );
buf \U$9 ( \65 , \64 );
nand \U$10 ( \66 , RIa148a08_33, \65 );
nor \U$11 ( \67 , RIa149098_47, RIa149110_48);
not \U$12 ( \68 , \67 );
not \U$13 ( \69 , RIa147bf8_3);
not \U$14 ( \70 , \69 );
or \U$15 ( \71 , \68 , \70 );
nand \U$16 ( \72 , RIa1480a8_13, RIa149110_48);
not \U$17 ( \73 , RIa148558_23);
nand \U$18 ( \74 , \72 , \73 , RIa149098_47);
nand \U$19 ( \75 , \71 , \74 );
nor \U$20 ( \76 , RIa149098_47, RIa1480a8_13);
and \U$21 ( \77 , \76 , RIa149110_48);
nor \U$22 ( \78 , \75 , \77 );
buf \U$23 ( \79 , \78 );
not \U$24 ( \80 , \79 );
not \U$25 ( \81 , \80 );
nand \U$26 ( \82 , \81 , RIa148918_31);
xor \U$27 ( \83 , \66 , \82 );
not \U$28 ( \84 , RIa147b80_2);
nor \U$29 ( \85 , RIa149098_47, RIa149110_48);
not \U$30 ( \86 , \85 );
or \U$31 ( \87 , \84 , \86 );
and \U$32 ( \88 , RIa148030_12, RIa149110_48);
and \U$33 ( \89 , RIa1484e0_22, RIa149098_47);
nor \U$34 ( \90 , \88 , \89 );
nand \U$35 ( \91 , \87 , \90 );
buf \U$36 ( \92 , \91 );
and \U$37 ( \93 , \92 , RIa148990_32);
not \U$38 ( \94 , \93 );
and \U$39 ( \95 , \83 , \94 );
and \U$40 ( \96 , \82 , \66 );
nor \U$41 ( \97 , \95 , \96 );
not \U$42 ( \98 , \97 );
nand \U$43 ( \99 , \92 , RIa148918_31);
nand \U$44 ( \100 , \65 , RIa148990_32);
xor \U$45 ( \101 , \99 , \100 );
and \U$46 ( \102 , \98 , \101 );
and \U$47 ( \103 , \99 , \100 );
nor \U$48 ( \104 , \102 , \103 );
and \U$49 ( \105 , \65 , RIa148918_31);
or \U$50 ( \106 , \104 , \105 );
not \U$51 ( \107 , \106 );
not \U$52 ( \108 , RIa147ce8_5);
not \U$53 ( \109 , \58 );
or \U$54 ( \110 , \108 , \109 );
and \U$55 ( \111 , RIa148198_15, RIa149110_48);
and \U$56 ( \112 , RIa148648_25, RIa149098_47);
nor \U$57 ( \113 , \111 , \112 );
nand \U$58 ( \114 , \110 , \113 );
buf \U$59 ( \115 , \114 );
nand \U$60 ( \116 , \115 , RIa148990_32);
not \U$61 ( \117 , \116 );
nor \U$62 ( \118 , RIa149098_47, RIa149110_48);
not \U$63 ( \119 , \118 );
not \U$64 ( \120 , RIa147d60_6);
or \U$65 ( \121 , \119 , \120 );
and \U$66 ( \122 , RIa148210_16, RIa149110_48);
and \U$67 ( \123 , RIa1486c0_26, RIa149098_47);
nor \U$68 ( \124 , \122 , \123 );
nand \U$69 ( \125 , \121 , \124 );
buf \U$70 ( \126 , \125 );
and \U$71 ( \127 , \126 , RIa148918_31);
not \U$72 ( \128 , \127 );
or \U$73 ( \129 , \117 , \128 );
or \U$74 ( \130 , \127 , \116 );
nand \U$75 ( \131 , \129 , \130 );
nand \U$76 ( \132 , \81 , RIa148a80_34);
xnor \U$77 ( \133 , \131 , \132 );
nand \U$78 ( \134 , \115 , RIa148a08_33);
not \U$79 ( \135 , \134 );
not \U$80 ( \136 , \135 );
nand \U$81 ( \137 , \126 , RIa148990_32);
not \U$82 ( \138 , \137 );
not \U$83 ( \139 , \138 );
or \U$84 ( \140 , \136 , \139 );
not \U$85 ( \141 , \134 );
not \U$86 ( \142 , \137 );
or \U$87 ( \143 , \141 , \142 );
not \U$88 ( \144 , \79 );
not \U$89 ( \145 , RIa148af8_35);
nor \U$90 ( \146 , \144 , \145 );
nand \U$91 ( \147 , \143 , \146 );
nand \U$92 ( \148 , \140 , \147 );
nand \U$93 ( \149 , \92 , RIa148b70_36);
not \U$94 ( \150 , \149 );
not \U$95 ( \151 , \150 );
nand \U$96 ( \152 , \65 , RIa148be8_37);
not \U$97 ( \153 , \152 );
not \U$98 ( \154 , \153 );
or \U$99 ( \155 , \151 , \154 );
not \U$100 ( \156 , \149 );
not \U$101 ( \157 , \152 );
or \U$102 ( \158 , \156 , \157 );
not \U$103 ( \159 , RIa147c70_4);
nor \U$104 ( \160 , RIa149098_47, RIa149110_48);
not \U$105 ( \161 , \160 );
or \U$106 ( \162 , \159 , \161 );
and \U$107 ( \163 , RIa148120_14, RIa149110_48);
and \U$108 ( \164 , RIa1485d0_24, RIa149098_47);
nor \U$109 ( \165 , \163 , \164 );
nand \U$110 ( \166 , \162 , \165 );
buf \U$111 ( \167 , \166 );
and \U$112 ( \168 , \167 , RIa148a80_34);
nand \U$113 ( \169 , \158 , \168 );
nand \U$114 ( \170 , \155 , \169 );
nor \U$115 ( \171 , \148 , \170 );
not \U$116 ( \172 , \171 );
nand \U$117 ( \173 , \148 , \170 );
nand \U$118 ( \174 , \172 , \173 );
nand \U$119 ( \175 , \65 , RIa148b70_36);
not \U$120 ( \176 , \175 );
nand \U$121 ( \177 , \92 , RIa148af8_35);
not \U$122 ( \178 , \177 );
not \U$123 ( \179 , \178 );
or \U$124 ( \180 , \176 , \179 );
not \U$125 ( \181 , \175 );
nand \U$126 ( \182 , \177 , \181 );
nand \U$127 ( \183 , \180 , \182 );
buf \U$128 ( \184 , \167 );
nand \U$129 ( \185 , \184 , RIa148a08_33);
not \U$130 ( \186 , \185 );
and \U$131 ( \187 , \183 , \186 );
not \U$132 ( \188 , \183 );
and \U$133 ( \189 , \188 , \185 );
nor \U$134 ( \190 , \187 , \189 );
not \U$135 ( \191 , \190 );
and \U$136 ( \192 , \174 , \191 );
not \U$137 ( \193 , \174 );
and \U$138 ( \194 , \193 , \190 );
nor \U$139 ( \195 , \192 , \194 );
xor \U$140 ( \196 , \133 , \195 );
nor \U$141 ( \197 , RIa149098_47, RIa148288_17);
and \U$142 ( \198 , \197 , RIa149110_48);
not \U$143 ( \199 , RIa147dd8_7);
not \U$144 ( \200 , \199 );
not \U$145 ( \201 , \67 );
or \U$146 ( \202 , \200 , \201 );
not \U$147 ( \203 , RIa148738_27);
nand \U$148 ( \204 , RIa148288_17, RIa149110_48);
nand \U$149 ( \205 , \203 , \204 , RIa149098_47);
nand \U$150 ( \206 , \202 , \205 );
nor \U$151 ( \207 , \198 , \206 );
buf \U$152 ( \208 , \207 );
nand \U$153 ( \209 , \208 , RIa148918_31);
not \U$154 ( \210 , \145 );
nand \U$155 ( \211 , \210 , \167 );
nand \U$156 ( \212 , \92 , RIa148be8_37);
nand \U$157 ( \213 , \211 , \212 );
nand \U$158 ( \214 , \64 , RIa148c60_38);
nand \U$159 ( \215 , \212 , \214 );
nand \U$160 ( \216 , \211 , \214 );
nand \U$161 ( \217 , \213 , \215 , \216 );
xor \U$162 ( \218 , \209 , \217 );
not \U$163 ( \219 , \80 );
and \U$164 ( \220 , \219 , RIa148b70_36);
not \U$165 ( \221 , \220 );
not \U$166 ( \222 , RIa147e50_8);
not \U$167 ( \223 , \160 );
or \U$168 ( \224 , \222 , \223 );
and \U$169 ( \225 , RIa148300_18, RIa149110_48);
and \U$170 ( \226 , RIa1487b0_28, RIa149098_47);
nor \U$171 ( \227 , \225 , \226 );
nand \U$172 ( \228 , \224 , \227 );
nand \U$173 ( \229 , \228 , RIa148918_31);
nand \U$174 ( \230 , \115 , RIa148a80_34);
xor \U$175 ( \231 , \229 , \230 );
and \U$176 ( \232 , \221 , \231 );
and \U$177 ( \233 , \229 , \230 );
nor \U$178 ( \234 , \232 , \233 );
not \U$179 ( \235 , \234 );
and \U$180 ( \236 , \218 , \235 );
and \U$181 ( \237 , \209 , \217 );
nor \U$182 ( \238 , \236 , \237 );
and \U$183 ( \239 , \196 , \238 );
and \U$184 ( \240 , \133 , \195 );
or \U$185 ( \241 , \239 , \240 );
not \U$186 ( \242 , \241 );
not \U$187 ( \243 , \178 );
not \U$188 ( \244 , \181 );
and \U$189 ( \245 , \243 , \244 );
and \U$190 ( \246 , \183 , \185 );
nor \U$191 ( \247 , \245 , \246 );
not \U$192 ( \248 , \65 );
not \U$193 ( \249 , \248 );
nand \U$194 ( \250 , \249 , RIa148af8_35);
nand \U$195 ( \251 , \184 , RIa148990_32);
xor \U$196 ( \252 , \250 , \251 );
nand \U$197 ( \253 , \92 , RIa148a80_34);
xnor \U$198 ( \254 , \252 , \253 );
xor \U$199 ( \255 , \247 , \254 );
not \U$200 ( \256 , \132 );
not \U$201 ( \257 , \131 );
or \U$202 ( \258 , \256 , \257 );
not \U$203 ( \259 , \127 );
nand \U$204 ( \260 , \259 , \116 );
nand \U$205 ( \261 , \258 , \260 );
not \U$206 ( \262 , \261 );
nand \U$207 ( \263 , \81 , RIa148a08_33);
not \U$208 ( \264 , \263 );
and \U$209 ( \265 , \115 , RIa148918_31);
not \U$210 ( \266 , \265 );
and \U$211 ( \267 , \264 , \266 );
and \U$212 ( \268 , \263 , \265 );
nor \U$213 ( \269 , \267 , \268 );
not \U$214 ( \270 , \269 );
and \U$215 ( \271 , \262 , \270 );
and \U$216 ( \272 , \261 , \269 );
nor \U$217 ( \273 , \271 , \272 );
xor \U$218 ( \274 , \255 , \273 );
not \U$219 ( \275 , \171 );
and \U$220 ( \276 , \275 , \190 );
not \U$221 ( \277 , \173 );
nor \U$222 ( \278 , \276 , \277 );
and \U$223 ( \279 , \274 , \278 );
not \U$224 ( \280 , \274 );
not \U$225 ( \281 , \278 );
and \U$226 ( \282 , \280 , \281 );
nor \U$227 ( \283 , \279 , \282 );
not \U$228 ( \284 , \283 );
not \U$229 ( \285 , \284 );
or \U$230 ( \286 , \242 , \285 );
nand \U$231 ( \287 , \274 , \281 );
nand \U$232 ( \288 , \286 , \287 );
not \U$233 ( \289 , \261 );
or \U$234 ( \290 , \289 , \269 );
not \U$235 ( \291 , \263 );
or \U$236 ( \292 , \291 , \265 );
nand \U$237 ( \293 , \290 , \292 );
not \U$238 ( \294 , \293 );
nand \U$239 ( \295 , \65 , RIa148a80_34);
nand \U$240 ( \296 , \92 , RIa148a08_33);
xor \U$241 ( \297 , \295 , \296 );
nand \U$242 ( \298 , \184 , RIa148918_31);
not \U$243 ( \299 , \298 );
and \U$244 ( \300 , \297 , \299 );
not \U$245 ( \301 , \297 );
and \U$246 ( \302 , \301 , \298 );
nor \U$247 ( \303 , \300 , \302 );
not \U$248 ( \304 , \303 );
nand \U$249 ( \305 , RIa148990_32, \81 );
not \U$250 ( \306 , \305 );
not \U$251 ( \307 , \253 );
not \U$252 ( \308 , \252 );
or \U$253 ( \309 , \307 , \308 );
nand \U$254 ( \310 , \251 , \250 );
nand \U$255 ( \311 , \309 , \310 );
not \U$256 ( \312 , \311 );
not \U$257 ( \313 , \312 );
or \U$258 ( \314 , \306 , \313 );
not \U$259 ( \315 , \305 );
nand \U$260 ( \316 , \311 , \315 );
nand \U$261 ( \317 , \314 , \316 );
not \U$262 ( \318 , \317 );
or \U$263 ( \319 , \304 , \318 );
or \U$264 ( \320 , \317 , \303 );
nand \U$265 ( \321 , \319 , \320 );
not \U$266 ( \322 , \321 );
not \U$267 ( \323 , \322 );
or \U$268 ( \324 , \294 , \323 );
not \U$269 ( \325 , \293 );
nand \U$270 ( \326 , \325 , \321 );
nand \U$271 ( \327 , \324 , \326 );
not \U$272 ( \328 , \327 );
xor \U$273 ( \329 , \247 , \254 );
and \U$274 ( \330 , \329 , \273 );
and \U$275 ( \331 , \247 , \254 );
or \U$276 ( \332 , \330 , \331 );
not \U$277 ( \333 , \332 );
and \U$278 ( \334 , \328 , \333 );
and \U$279 ( \335 , \327 , \332 );
nor \U$280 ( \336 , \334 , \335 );
nor \U$281 ( \337 , \288 , \336 );
not \U$282 ( \338 , \337 );
not \U$283 ( \339 , \214 );
and \U$284 ( \340 , \91 , RIa148cd8_39);
buf \U$285 ( \341 , \340 );
nand \U$286 ( \342 , \339 , \341 );
not \U$287 ( \343 , \342 );
not \U$288 ( \344 , \343 );
nand \U$289 ( \345 , \207 , RIa148990_32);
and \U$290 ( \346 , \126 , RIa148a08_33);
xnor \U$291 ( \347 , \345 , \346 );
not \U$292 ( \348 , \347 );
or \U$293 ( \349 , \344 , \348 );
or \U$294 ( \350 , \347 , \343 );
nand \U$295 ( \351 , \349 , \350 );
not \U$296 ( \352 , \351 );
not \U$297 ( \353 , \231 );
not \U$298 ( \354 , \220 );
and \U$299 ( \355 , \353 , \354 );
and \U$300 ( \356 , \231 , \220 );
nor \U$301 ( \357 , \355 , \356 );
not \U$302 ( \358 , \357 );
and \U$303 ( \359 , \352 , \358 );
and \U$304 ( \360 , \351 , \357 );
nor \U$305 ( \361 , \359 , \360 );
not \U$306 ( \362 , \92 );
not \U$307 ( \363 , RIa148c60_38);
or \U$308 ( \364 , \362 , \363 );
not \U$309 ( \365 , RIa148cd8_39);
or \U$310 ( \366 , \248 , \365 );
nand \U$311 ( \367 , \364 , \366 );
and \U$312 ( \368 , \342 , \367 );
not \U$313 ( \369 , \368 );
nand \U$314 ( \370 , \208 , RIa148a08_33);
not \U$315 ( \371 , \370 );
and \U$316 ( \372 , \64 , RIa148d50_40);
and \U$317 ( \373 , \340 , \372 );
not \U$318 ( \374 , \373 );
and \U$319 ( \375 , \371 , \374 );
and \U$320 ( \376 , \340 , \372 );
and \U$321 ( \377 , \370 , \376 );
nor \U$322 ( \378 , \375 , \377 );
not \U$323 ( \379 , \378 );
and \U$324 ( \380 , \369 , \379 );
not \U$325 ( \381 , \376 );
and \U$326 ( \382 , \370 , \381 );
nor \U$327 ( \383 , \380 , \382 );
or \U$328 ( \384 , \361 , \383 );
not \U$329 ( \385 , \357 );
nand \U$330 ( \386 , \385 , \351 );
nand \U$331 ( \387 , \384 , \386 );
not \U$332 ( \388 , \387 );
and \U$333 ( \389 , \114 , RIa148af8_35);
and \U$334 ( \390 , \126 , RIa148a80_34);
xor \U$335 ( \391 , \389 , \390 );
and \U$336 ( \392 , \79 , RIa148be8_37);
and \U$337 ( \393 , \391 , \392 );
and \U$338 ( \394 , \389 , \390 );
or \U$339 ( \395 , \393 , \394 );
xor \U$340 ( \396 , \214 , \212 );
xnor \U$341 ( \397 , \396 , \211 );
xor \U$342 ( \398 , \395 , \397 );
not \U$343 ( \399 , RIa147ec8_9);
nand \U$344 ( \400 , \399 , \85 );
not \U$345 ( \401 , RIa149098_47);
not \U$346 ( \402 , RIa148378_19);
nand \U$347 ( \403 , \401 , \402 , RIa149110_48);
not \U$348 ( \404 , RIa148828_29);
nand \U$349 ( \405 , RIa148378_19, RIa149110_48);
nand \U$350 ( \406 , \404 , \405 , RIa149098_47);
nand \U$351 ( \407 , \400 , \403 , \406 );
not \U$352 ( \408 , \407 );
nand \U$353 ( \409 , \408 , RIa148918_31);
and \U$354 ( \410 , \166 , RIa148b70_36);
and \U$355 ( \411 , \228 , RIa148990_32);
nor \U$356 ( \412 , \410 , \411 );
or \U$357 ( \413 , \409 , \412 );
nand \U$358 ( \414 , \410 , \411 );
nand \U$359 ( \415 , \413 , \414 );
and \U$360 ( \416 , \398 , \415 );
and \U$361 ( \417 , \395 , \397 );
or \U$362 ( \418 , \416 , \417 );
not \U$363 ( \419 , \418 );
not \U$364 ( \420 , \419 );
not \U$365 ( \421 , \234 );
not \U$366 ( \422 , \218 );
or \U$367 ( \423 , \421 , \422 );
or \U$368 ( \424 , \234 , \218 );
nand \U$369 ( \425 , \423 , \424 );
not \U$370 ( \426 , \425 );
not \U$371 ( \427 , \426 );
or \U$372 ( \428 , \420 , \427 );
nand \U$373 ( \429 , \425 , \418 );
nand \U$374 ( \430 , \428 , \429 );
not \U$375 ( \431 , \430 );
or \U$376 ( \432 , \388 , \431 );
nand \U$377 ( \433 , \425 , \419 );
nand \U$378 ( \434 , \432 , \433 );
not \U$379 ( \435 , \434 );
xor \U$380 ( \436 , \133 , \195 );
xor \U$381 ( \437 , \436 , \238 );
not \U$382 ( \438 , \437 );
xor \U$383 ( \439 , \150 , \153 );
xor \U$384 ( \440 , \439 , \168 );
not \U$385 ( \441 , \440 );
xor \U$386 ( \442 , \138 , \135 );
xnor \U$387 ( \443 , \442 , \146 );
not \U$388 ( \444 , \443 );
not \U$389 ( \445 , \444 );
or \U$390 ( \446 , \441 , \445 );
not \U$391 ( \447 , \347 );
not \U$392 ( \448 , \342 );
or \U$393 ( \449 , \447 , \448 );
not \U$394 ( \450 , \346 );
nand \U$395 ( \451 , \450 , \345 );
nand \U$396 ( \452 , \449 , \451 );
nand \U$397 ( \453 , \446 , \452 );
not \U$398 ( \454 , \440 );
nand \U$399 ( \455 , \454 , \443 );
and \U$400 ( \456 , \453 , \455 );
not \U$401 ( \457 , \456 );
nand \U$402 ( \458 , \438 , \457 );
nand \U$403 ( \459 , \435 , \458 );
nand \U$404 ( \460 , \437 , \456 );
nand \U$405 ( \461 , \459 , \460 );
not \U$406 ( \462 , \461 );
not \U$407 ( \463 , \241 );
not \U$408 ( \464 , \463 );
not \U$409 ( \465 , \284 );
or \U$410 ( \466 , \464 , \465 );
nand \U$411 ( \467 , \283 , \241 );
nand \U$412 ( \468 , \466 , \467 );
not \U$413 ( \469 , \468 );
nand \U$414 ( \470 , \462 , \469 );
nand \U$415 ( \471 , \338 , \470 );
not \U$416 ( \472 , \332 );
not \U$417 ( \473 , \472 );
not \U$418 ( \474 , \327 );
or \U$419 ( \475 , \473 , \474 );
not \U$420 ( \476 , \322 );
nand \U$421 ( \477 , \476 , \293 );
nand \U$422 ( \478 , \475 , \477 );
not \U$423 ( \479 , \83 );
not \U$424 ( \480 , \93 );
and \U$425 ( \481 , \479 , \480 );
and \U$426 ( \482 , \83 , \93 );
nor \U$427 ( \483 , \481 , \482 );
and \U$428 ( \484 , \297 , \298 );
and \U$429 ( \485 , \296 , \295 );
nor \U$430 ( \486 , \484 , \485 );
xnor \U$431 ( \487 , \483 , \486 );
not \U$432 ( \488 , \312 );
not \U$433 ( \489 , \315 );
and \U$434 ( \490 , \488 , \489 );
not \U$435 ( \491 , \303 );
and \U$436 ( \492 , \317 , \491 );
nor \U$437 ( \493 , \490 , \492 );
xor \U$438 ( \494 , \487 , \493 );
nand \U$439 ( \495 , \478 , \494 );
or \U$440 ( \496 , \493 , \487 );
or \U$441 ( \497 , \483 , \486 );
nand \U$442 ( \498 , \496 , \497 );
not \U$443 ( \499 , \101 );
not \U$444 ( \500 , \97 );
or \U$445 ( \501 , \499 , \500 );
or \U$446 ( \502 , \97 , \101 );
nand \U$447 ( \503 , \501 , \502 );
nand \U$448 ( \504 , \498 , \503 );
nand \U$449 ( \505 , \495 , \504 );
nor \U$450 ( \506 , \471 , \505 );
not \U$451 ( \507 , \506 );
and \U$452 ( \508 , \115 , RIa148be8_37);
not \U$453 ( \509 , \508 );
not \U$454 ( \510 , \407 );
and \U$455 ( \511 , \510 , RIa148a08_33);
not \U$456 ( \512 , \511 );
or \U$457 ( \513 , \509 , \512 );
not \U$458 ( \514 , RIa147f40_10);
not \U$459 ( \515 , \160 );
or \U$460 ( \516 , \514 , \515 );
and \U$461 ( \517 , RIa1483f0_20, RIa149110_48);
and \U$462 ( \518 , RIa1488a0_30, RIa149098_47);
nor \U$463 ( \519 , \517 , \518 );
nand \U$464 ( \520 , \516 , \519 );
buf \U$465 ( \521 , \520 );
nand \U$466 ( \522 , \521 , RIa148990_32);
nand \U$467 ( \523 , \513 , \522 );
not \U$468 ( \524 , \508 );
not \U$469 ( \525 , \511 );
nand \U$470 ( \526 , \524 , \525 );
and \U$471 ( \527 , \523 , \526 );
not \U$472 ( \528 , \527 );
and \U$473 ( \529 , \207 , RIa148af8_35);
not \U$474 ( \530 , \529 );
not \U$475 ( \531 , RIa148c60_38);
not \U$476 ( \532 , \167 );
or \U$477 ( \533 , \531 , \532 );
nand \U$478 ( \534 , \126 , RIa148b70_36);
nand \U$479 ( \535 , \533 , \534 );
not \U$480 ( \536 , \535 );
or \U$481 ( \537 , \530 , \536 );
and \U$482 ( \538 , \126 , RIa148c60_38);
nand \U$483 ( \539 , \410 , \538 );
nand \U$484 ( \540 , \537 , \539 );
not \U$485 ( \541 , \540 );
nand \U$486 ( \542 , \79 , RIa148d50_40);
not \U$487 ( \543 , \542 );
nand \U$488 ( \544 , \543 , \341 );
not \U$489 ( \545 , \544 );
and \U$490 ( \546 , \541 , \545 );
and \U$491 ( \547 , \540 , \544 );
nor \U$492 ( \548 , \546 , \547 );
nor \U$493 ( \549 , \528 , \548 );
not \U$494 ( \550 , \549 );
and \U$495 ( \551 , \208 , RIa148a80_34);
and \U$496 ( \552 , \126 , RIa148af8_35);
and \U$497 ( \553 , \551 , \552 );
not \U$498 ( \554 , \551 );
not \U$499 ( \555 , \552 );
and \U$500 ( \556 , \554 , \555 );
nor \U$501 ( \557 , \553 , \556 );
not \U$502 ( \558 , \557 );
nor \U$503 ( \559 , \340 , \372 );
or \U$504 ( \560 , \559 , \373 );
not \U$505 ( \561 , \560 );
not \U$506 ( \562 , \561 );
and \U$507 ( \563 , \558 , \562 );
and \U$508 ( \564 , \557 , \561 );
nor \U$509 ( \565 , \563 , \564 );
not \U$510 ( \566 , \527 );
nand \U$511 ( \567 , \548 , \566 );
nand \U$512 ( \568 , \550 , \565 , \567 );
and \U$513 ( \569 , \114 , RIa148c60_38);
and \U$514 ( \570 , \228 , RIa148af8_35);
xor \U$515 ( \571 , \569 , \570 );
and \U$516 ( \572 , \510 , RIa148a80_34);
and \U$517 ( \573 , \571 , \572 );
and \U$518 ( \574 , \569 , \570 );
or \U$519 ( \575 , \573 , \574 );
not \U$520 ( \576 , \575 );
not \U$521 ( \577 , \576 );
not \U$522 ( \578 , RIa148a08_33);
not \U$523 ( \579 , \521 );
or \U$524 ( \580 , \578 , \579 );
nand \U$525 ( \581 , \126 , RIa148be8_37);
nand \U$526 ( \582 , \580 , \581 );
not \U$527 ( \583 , \582 );
and \U$528 ( \584 , \208 , RIa148b70_36);
not \U$529 ( \585 , \584 );
or \U$530 ( \586 , \583 , \585 );
and \U$531 ( \587 , \520 , RIa148be8_37);
nand \U$532 ( \588 , \587 , \346 );
nand \U$533 ( \589 , \586 , \588 );
not \U$534 ( \590 , \589 );
not \U$535 ( \591 , \590 );
or \U$536 ( \592 , \577 , \591 );
or \U$537 ( \593 , \576 , \590 );
buf \U$538 ( \594 , \535 );
nand \U$539 ( \595 , \539 , \594 );
buf \U$540 ( \596 , \529 );
and \U$541 ( \597 , \595 , \596 );
not \U$542 ( \598 , \595 );
not \U$543 ( \599 , \596 );
and \U$544 ( \600 , \598 , \599 );
nor \U$545 ( \601 , \597 , \600 );
nand \U$546 ( \602 , \593 , \601 );
nand \U$547 ( \603 , \592 , \602 );
and \U$548 ( \604 , \568 , \603 );
not \U$549 ( \605 , \549 );
and \U$550 ( \606 , \567 , \605 );
nor \U$551 ( \607 , \606 , \565 );
nor \U$552 ( \608 , \604 , \607 );
not \U$553 ( \609 , \608 );
not \U$554 ( \610 , \548 );
not \U$555 ( \611 , \527 );
and \U$556 ( \612 , \610 , \611 );
not \U$557 ( \613 , \544 );
nor \U$558 ( \614 , \613 , \540 );
nor \U$559 ( \615 , \612 , \614 );
not \U$560 ( \616 , \615 );
not \U$561 ( \617 , \414 );
nor \U$562 ( \618 , \617 , \412 );
xor \U$563 ( \619 , \618 , \409 );
not \U$564 ( \620 , \560 );
not \U$565 ( \621 , \557 );
or \U$566 ( \622 , \620 , \621 );
not \U$567 ( \623 , \551 );
nand \U$568 ( \624 , \623 , \555 );
nand \U$569 ( \625 , \622 , \624 );
xor \U$570 ( \626 , \619 , \625 );
not \U$571 ( \627 , \626 );
and \U$572 ( \628 , \616 , \627 );
and \U$573 ( \629 , \615 , \626 );
nor \U$574 ( \630 , \628 , \629 );
not \U$575 ( \631 , \630 );
not \U$576 ( \632 , \631 );
or \U$577 ( \633 , \609 , \632 );
not \U$578 ( \634 , \608 );
nand \U$579 ( \635 , \634 , \630 );
nand \U$580 ( \636 , \633 , \635 );
not \U$581 ( \637 , \378 );
and \U$582 ( \638 , \368 , \637 );
not \U$583 ( \639 , \368 );
and \U$584 ( \640 , \639 , \378 );
nor \U$585 ( \641 , \638 , \640 );
nand \U$586 ( \642 , \228 , RIa148a08_33);
and \U$587 ( \643 , \166 , RIa148be8_37);
and \U$588 ( \644 , \642 , \643 );
not \U$589 ( \645 , \642 );
not \U$590 ( \646 , \643 );
and \U$591 ( \647 , \645 , \646 );
nor \U$592 ( \648 , \644 , \647 );
nand \U$593 ( \649 , \408 , RIa148990_32);
xor \U$594 ( \650 , \648 , \649 );
not \U$595 ( \651 , \650 );
nand \U$596 ( \652 , \114 , RIa148b70_36);
nand \U$597 ( \653 , \520 , RIa148918_31);
xor \U$598 ( \654 , \652 , \653 );
nand \U$599 ( \655 , \79 , RIa148c60_38);
xor \U$600 ( \656 , \654 , \655 );
nand \U$601 ( \657 , \651 , \656 );
not \U$602 ( \658 , \657 );
and \U$603 ( \659 , \167 , RIa148cd8_39);
not \U$604 ( \660 , \659 );
nor \U$605 ( \661 , \660 , \542 );
not \U$606 ( \662 , \661 );
and \U$607 ( \663 , \228 , RIa148a80_34);
not \U$608 ( \664 , \663 );
and \U$609 ( \665 , \78 , RIa148cd8_39);
nand \U$610 ( \666 , \92 , RIa148d50_40);
xor \U$611 ( \667 , \665 , \666 );
not \U$612 ( \668 , \667 );
or \U$613 ( \669 , \664 , \668 );
or \U$614 ( \670 , \667 , \663 );
nand \U$615 ( \671 , \669 , \670 );
not \U$616 ( \672 , \671 );
or \U$617 ( \673 , \662 , \672 );
not \U$618 ( \674 , \667 );
nand \U$619 ( \675 , \674 , \663 );
nand \U$620 ( \676 , \673 , \675 );
not \U$621 ( \677 , \676 );
or \U$622 ( \678 , \658 , \677 );
not \U$623 ( \679 , \656 );
nand \U$624 ( \680 , \679 , \650 );
nand \U$625 ( \681 , \678 , \680 );
xor \U$626 ( \682 , \641 , \681 );
xor \U$627 ( \683 , \652 , \653 );
and \U$628 ( \684 , \683 , \655 );
and \U$629 ( \685 , \652 , \653 );
or \U$630 ( \686 , \684 , \685 );
not \U$631 ( \687 , \686 );
xor \U$632 ( \688 , \389 , \390 );
xor \U$633 ( \689 , \688 , \392 );
not \U$634 ( \690 , \689 );
or \U$635 ( \691 , \687 , \690 );
or \U$636 ( \692 , \686 , \689 );
nand \U$637 ( \693 , \691 , \692 );
buf \U$638 ( \694 , \642 );
or \U$639 ( \695 , \649 , \694 );
nand \U$640 ( \696 , \695 , \646 );
nand \U$641 ( \697 , \649 , \694 );
nand \U$642 ( \698 , \696 , \697 );
and \U$643 ( \699 , \693 , \698 );
not \U$644 ( \700 , \693 );
not \U$645 ( \701 , \698 );
and \U$646 ( \702 , \700 , \701 );
or \U$647 ( \703 , \699 , \702 );
xor \U$648 ( \704 , \682 , \703 );
not \U$649 ( \705 , \704 );
and \U$650 ( \706 , \636 , \705 );
not \U$651 ( \707 , \636 );
and \U$652 ( \708 , \707 , \704 );
nor \U$653 ( \709 , \706 , \708 );
not \U$654 ( \710 , \709 );
not \U$655 ( \711 , \650 );
not \U$656 ( \712 , \656 );
and \U$657 ( \713 , \711 , \712 );
and \U$658 ( \714 , \650 , \656 );
nor \U$659 ( \715 , \713 , \714 );
xor \U$660 ( \716 , \715 , \676 );
not \U$661 ( \717 , \716 );
not \U$662 ( \718 , \717 );
buf \U$663 ( \719 , \538 );
not \U$664 ( \720 , \719 );
not \U$665 ( \721 , RIa148be8_37);
not \U$666 ( \722 , \208 );
or \U$667 ( \723 , \721 , \722 );
buf \U$668 ( \724 , \228 );
nand \U$669 ( \725 , \724 , RIa148b70_36);
nand \U$670 ( \726 , \723 , \725 );
not \U$671 ( \727 , \726 );
or \U$672 ( \728 , \720 , \727 );
nand \U$673 ( \729 , \724 , RIa148be8_37);
not \U$674 ( \730 , \729 );
nand \U$675 ( \731 , \730 , \584 );
nand \U$676 ( \732 , \728 , \731 );
not \U$677 ( \733 , \732 );
not \U$678 ( \734 , \542 );
not \U$679 ( \735 , \659 );
and \U$680 ( \736 , \734 , \735 );
and \U$681 ( \737 , \542 , \659 );
nor \U$682 ( \738 , \736 , \737 );
not \U$683 ( \739 , \738 );
and \U$684 ( \740 , \115 , RIa148d50_40);
nand \U$685 ( \741 , \659 , \740 );
not \U$686 ( \742 , \741 );
not \U$687 ( \743 , \742 );
or \U$688 ( \744 , \739 , \743 );
or \U$689 ( \745 , \738 , \742 );
nand \U$690 ( \746 , \744 , \745 );
not \U$691 ( \747 , \746 );
or \U$692 ( \748 , \733 , \747 );
not \U$693 ( \749 , \738 );
nand \U$694 ( \750 , \749 , \742 );
nand \U$695 ( \751 , \748 , \750 );
buf \U$696 ( \752 , \511 );
not \U$697 ( \753 , \752 );
xnor \U$698 ( \754 , \508 , \522 );
not \U$699 ( \755 , \754 );
or \U$700 ( \756 , \753 , \755 );
or \U$701 ( \757 , \752 , \754 );
nand \U$702 ( \758 , \756 , \757 );
not \U$703 ( \759 , \758 );
or \U$704 ( \760 , \751 , \759 );
xor \U$705 ( \761 , \661 , \671 );
nand \U$706 ( \762 , \760 , \761 );
nand \U$707 ( \763 , \751 , \759 );
nand \U$708 ( \764 , \762 , \763 );
not \U$709 ( \765 , \764 );
or \U$710 ( \766 , \718 , \765 );
xor \U$711 ( \767 , \548 , \603 );
not \U$712 ( \768 , \566 );
not \U$713 ( \769 , \565 );
or \U$714 ( \770 , \768 , \769 );
or \U$715 ( \771 , \566 , \565 );
nand \U$716 ( \772 , \770 , \771 );
xor \U$717 ( \773 , \767 , \772 );
not \U$718 ( \774 , \773 );
nand \U$719 ( \775 , \766 , \774 );
or \U$720 ( \776 , \764 , \717 );
nand \U$721 ( \777 , \775 , \776 );
not \U$722 ( \778 , \777 );
nand \U$723 ( \779 , \710 , \778 );
not \U$724 ( \780 , \779 );
not \U$725 ( \781 , \615 );
and \U$726 ( \782 , \781 , \626 );
and \U$727 ( \783 , \619 , \625 );
nor \U$728 ( \784 , \782 , \783 );
not \U$729 ( \785 , \784 );
xor \U$730 ( \786 , \395 , \397 );
xor \U$731 ( \787 , \786 , \415 );
not \U$732 ( \788 , \787 );
not \U$733 ( \789 , \788 );
not \U$734 ( \790 , \698 );
not \U$735 ( \791 , \693 );
or \U$736 ( \792 , \790 , \791 );
not \U$737 ( \793 , \689 );
nand \U$738 ( \794 , \793 , \686 );
nand \U$739 ( \795 , \792 , \794 );
not \U$740 ( \796 , \795 );
not \U$741 ( \797 , \796 );
or \U$742 ( \798 , \789 , \797 );
nand \U$743 ( \799 , \795 , \787 );
nand \U$744 ( \800 , \798 , \799 );
not \U$745 ( \801 , \800 );
and \U$746 ( \802 , \785 , \801 );
and \U$747 ( \803 , \784 , \800 );
nor \U$748 ( \804 , \802 , \803 );
not \U$749 ( \805 , \804 );
xor \U$750 ( \806 , \641 , \681 );
and \U$751 ( \807 , \806 , \703 );
and \U$752 ( \808 , \641 , \681 );
or \U$753 ( \809 , \807 , \808 );
not \U$754 ( \810 , \383 );
and \U$755 ( \811 , \361 , \810 );
not \U$756 ( \812 , \361 );
and \U$757 ( \813 , \812 , \383 );
nor \U$758 ( \814 , \811 , \813 );
not \U$759 ( \815 , \814 );
and \U$760 ( \816 , \809 , \815 );
not \U$761 ( \817 , \809 );
and \U$762 ( \818 , \817 , \814 );
nor \U$763 ( \819 , \816 , \818 );
not \U$764 ( \820 , \819 );
or \U$765 ( \821 , \805 , \820 );
or \U$766 ( \822 , \819 , \804 );
nand \U$767 ( \823 , \821 , \822 );
not \U$768 ( \824 , \704 );
not \U$769 ( \825 , \608 );
nand \U$770 ( \826 , \825 , \631 );
not \U$771 ( \827 , \826 );
or \U$772 ( \828 , \824 , \827 );
nand \U$773 ( \829 , \630 , \608 );
nand \U$774 ( \830 , \828 , \829 );
nand \U$775 ( \831 , \823 , \830 );
not \U$776 ( \832 , \831 );
or \U$777 ( \833 , \780 , \832 );
and \U$778 ( \834 , \819 , \804 );
nor \U$779 ( \835 , \834 , \830 );
not \U$780 ( \836 , \819 );
not \U$781 ( \837 , \804 );
nand \U$782 ( \838 , \836 , \837 );
nand \U$783 ( \839 , \835 , \838 );
nand \U$784 ( \840 , \833 , \839 );
not \U$785 ( \841 , \815 );
not \U$786 ( \842 , \809 );
not \U$787 ( \843 , \842 );
or \U$788 ( \844 , \841 , \843 );
nand \U$789 ( \845 , \844 , \838 );
and \U$790 ( \846 , \440 , \443 );
not \U$791 ( \847 , \440 );
and \U$792 ( \848 , \847 , \444 );
nor \U$793 ( \849 , \846 , \848 );
not \U$794 ( \850 , \452 );
xor \U$795 ( \851 , \849 , \850 );
not \U$796 ( \852 , \387 );
not \U$797 ( \853 , \430 );
not \U$798 ( \854 , \853 );
or \U$799 ( \855 , \852 , \854 );
not \U$800 ( \856 , \387 );
nand \U$801 ( \857 , \856 , \430 );
nand \U$802 ( \858 , \855 , \857 );
xor \U$803 ( \859 , \851 , \858 );
not \U$804 ( \860 , \784 );
not \U$805 ( \861 , \860 );
not \U$806 ( \862 , \800 );
or \U$807 ( \863 , \861 , \862 );
not \U$808 ( \864 , \796 );
nand \U$809 ( \865 , \864 , \788 );
nand \U$810 ( \866 , \863 , \865 );
xor \U$811 ( \867 , \859 , \866 );
nand \U$812 ( \868 , \845 , \867 );
xor \U$813 ( \869 , \456 , \437 );
xor \U$814 ( \870 , \869 , \434 );
xor \U$815 ( \871 , \851 , \858 );
and \U$816 ( \872 , \871 , \866 );
and \U$817 ( \873 , \851 , \858 );
or \U$818 ( \874 , \872 , \873 );
nand \U$819 ( \875 , \870 , \874 );
nand \U$820 ( \876 , \868 , \875 );
nor \U$821 ( \877 , \840 , \876 );
nor \U$822 ( \878 , \845 , \867 );
nand \U$823 ( \879 , \878 , \875 );
not \U$824 ( \880 , \874 );
not \U$825 ( \881 , \870 );
nand \U$826 ( \882 , \880 , \881 );
nand \U$827 ( \883 , \879 , \882 );
nor \U$828 ( \884 , \877 , \883 );
nand \U$829 ( \885 , \207 , RIa148cd8_39);
nand \U$830 ( \886 , \126 , RIa148d50_40);
or \U$831 ( \887 , \885 , \886 );
and \U$832 ( \888 , \521 , RIa148af8_35);
and \U$833 ( \889 , \887 , \888 );
not \U$834 ( \890 , \887 );
not \U$835 ( \891 , \888 );
and \U$836 ( \892 , \890 , \891 );
nor \U$837 ( \893 , \889 , \892 );
not \U$838 ( \894 , \893 );
and \U$839 ( \895 , \126 , RIa148cd8_39);
xor \U$840 ( \896 , \895 , \740 );
not \U$841 ( \897 , \896 );
and \U$842 ( \898 , \894 , \897 );
and \U$843 ( \899 , \887 , \891 );
nor \U$844 ( \900 , \898 , \899 );
not \U$845 ( \901 , \900 );
nand \U$846 ( \902 , \572 , \888 );
not \U$847 ( \903 , RIa148af8_35);
not \U$848 ( \904 , \408 );
not \U$849 ( \905 , \904 );
not \U$850 ( \906 , \905 );
or \U$851 ( \907 , \903 , \906 );
buf \U$852 ( \908 , \521 );
nand \U$853 ( \909 , \908 , RIa148a80_34);
nand \U$854 ( \910 , \907 , \909 );
nand \U$855 ( \911 , \902 , \910 );
and \U$856 ( \912 , \895 , \740 );
xor \U$857 ( \913 , \911 , \912 );
not \U$858 ( \914 , \913 );
or \U$859 ( \915 , \901 , \914 );
or \U$860 ( \916 , \900 , \913 );
nand \U$861 ( \917 , \915 , \916 );
not \U$862 ( \918 , \917 );
not \U$863 ( \919 , \918 );
and \U$864 ( \920 , RIa148cd8_39, \115 );
and \U$865 ( \921 , \184 , RIa148d50_40);
nor \U$866 ( \922 , \920 , \921 );
nor \U$867 ( \923 , \742 , \922 );
not \U$868 ( \924 , \923 );
not \U$869 ( \925 , \729 );
nand \U$870 ( \926 , \408 , RIa148b70_36);
not \U$871 ( \927 , \926 );
and \U$872 ( \928 , \207 , RIa148c60_38);
not \U$873 ( \929 , \928 );
or \U$874 ( \930 , \927 , \929 );
or \U$875 ( \931 , \928 , \926 );
nand \U$876 ( \932 , \930 , \931 );
not \U$877 ( \933 , \932 );
or \U$878 ( \934 , \925 , \933 );
not \U$879 ( \935 , \928 );
nand \U$880 ( \936 , \935 , \926 );
nand \U$881 ( \937 , \934 , \936 );
not \U$882 ( \938 , \937 );
or \U$883 ( \939 , \924 , \938 );
or \U$884 ( \940 , \937 , \923 );
nand \U$885 ( \941 , \939 , \940 );
not \U$886 ( \942 , \941 );
nand \U$887 ( \943 , \731 , \726 );
not \U$888 ( \944 , \719 );
and \U$889 ( \945 , \943 , \944 );
not \U$890 ( \946 , \943 );
and \U$891 ( \947 , \946 , \719 );
nor \U$892 ( \948 , \945 , \947 );
not \U$893 ( \949 , \948 );
and \U$894 ( \950 , \942 , \949 );
and \U$895 ( \951 , \941 , \948 );
nor \U$896 ( \952 , \950 , \951 );
not \U$897 ( \953 , \952 );
not \U$898 ( \954 , \953 );
or \U$899 ( \955 , \919 , \954 );
nand \U$900 ( \956 , \952 , \917 );
nand \U$901 ( \957 , \955 , \956 );
xnor \U$902 ( \958 , \896 , \893 );
not \U$903 ( \959 , \958 );
not \U$904 ( \960 , \959 );
nand \U$905 ( \961 , \905 , RIa148be8_37);
not \U$906 ( \962 , \961 );
and \U$907 ( \963 , \520 , RIa148b70_36);
not \U$908 ( \964 , \963 );
not \U$909 ( \965 , \964 );
and \U$910 ( \966 , \228 , RIa148c60_38);
not \U$911 ( \967 , \966 );
or \U$912 ( \968 , \965 , \967 );
not \U$913 ( \969 , \966 );
nand \U$914 ( \970 , \969 , \963 );
nand \U$915 ( \971 , \968 , \970 );
not \U$916 ( \972 , \971 );
or \U$917 ( \973 , \962 , \972 );
nand \U$918 ( \974 , \969 , \964 );
nand \U$919 ( \975 , \973 , \974 );
not \U$920 ( \976 , \975 );
not \U$921 ( \977 , \976 );
not \U$922 ( \978 , \729 );
not \U$923 ( \979 , \932 );
not \U$924 ( \980 , \979 );
or \U$925 ( \981 , \978 , \980 );
not \U$926 ( \982 , \729 );
nand \U$927 ( \983 , \982 , \932 );
nand \U$928 ( \984 , \981 , \983 );
not \U$929 ( \985 , \984 );
or \U$930 ( \986 , \977 , \985 );
or \U$931 ( \987 , \976 , \984 );
nand \U$932 ( \988 , \986 , \987 );
not \U$933 ( \989 , \988 );
or \U$934 ( \990 , \960 , \989 );
not \U$935 ( \991 , \976 );
nand \U$936 ( \992 , \991 , \984 );
nand \U$937 ( \993 , \990 , \992 );
nand \U$938 ( \994 , \957 , \993 );
not \U$939 ( \995 , \994 );
nand \U$940 ( \996 , \724 , RIa148d50_40);
nand \U$941 ( \997 , \521 , RIa148c60_38);
nor \U$942 ( \998 , \996 , \997 );
xnor \U$943 ( \999 , \996 , \997 );
not \U$944 ( \1000 , \904 );
nand \U$945 ( \1001 , \1000 , RIa148cd8_39);
or \U$946 ( \1002 , \999 , \1001 );
nand \U$947 ( \1003 , \521 , RIa148d50_40);
nor \U$948 ( \1004 , \1003 , \365 );
nand \U$949 ( \1005 , \1000 , \1004 );
nand \U$950 ( \1006 , \1002 , \1005 );
xor \U$951 ( \1007 , \998 , \1006 );
nand \U$952 ( \1008 , \408 , RIa148c60_38);
not \U$953 ( \1009 , \1008 );
not \U$954 ( \1010 , \587 );
and \U$955 ( \1011 , \1009 , \1010 );
and \U$956 ( \1012 , \1008 , \587 );
nor \U$957 ( \1013 , \1011 , \1012 );
nand \U$958 ( \1014 , \208 , RIa148d50_40);
not \U$959 ( \1015 , \1014 );
nand \U$960 ( \1016 , \724 , RIa148cd8_39);
not \U$961 ( \1017 , \1016 );
and \U$962 ( \1018 , \1015 , \1017 );
and \U$963 ( \1019 , \1014 , \1016 );
nor \U$964 ( \1020 , \1018 , \1019 );
not \U$965 ( \1021 , \1020 );
and \U$966 ( \1022 , \1013 , \1021 );
not \U$967 ( \1023 , \1013 );
and \U$968 ( \1024 , \1023 , \1020 );
nor \U$969 ( \1025 , \1022 , \1024 );
and \U$970 ( \1026 , \1007 , \1025 );
and \U$971 ( \1027 , \998 , \1006 );
or \U$972 ( \1028 , \1026 , \1027 );
xnor \U$973 ( \1029 , \971 , \961 );
not \U$974 ( \1030 , \1029 );
not \U$975 ( \1031 , \887 );
and \U$976 ( \1032 , \885 , \886 );
nor \U$977 ( \1033 , \1031 , \1032 );
not \U$978 ( \1034 , \1014 );
not \U$979 ( \1035 , \1016 );
nand \U$980 ( \1036 , \1034 , \1035 );
not \U$981 ( \1037 , \1036 );
and \U$982 ( \1038 , \1033 , \1037 );
not \U$983 ( \1039 , \1033 );
and \U$984 ( \1040 , \1039 , \1036 );
nor \U$985 ( \1041 , \1038 , \1040 );
not \U$986 ( \1042 , \1041 );
or \U$987 ( \1043 , \1030 , \1042 );
or \U$988 ( \1044 , \1029 , \1041 );
nand \U$989 ( \1045 , \1043 , \1044 );
not \U$990 ( \1046 , \587 );
not \U$991 ( \1047 , \1046 );
not \U$992 ( \1048 , \1008 );
or \U$993 ( \1049 , \1047 , \1048 );
or \U$994 ( \1050 , \1008 , \1046 );
nand \U$995 ( \1051 , \1050 , \1021 );
nand \U$996 ( \1052 , \1049 , \1051 );
nand \U$997 ( \1053 , \1045 , \1052 );
nand \U$998 ( \1054 , \1028 , \1053 );
not \U$999 ( \1055 , \1045 );
not \U$1000 ( \1056 , \1052 );
nand \U$1001 ( \1057 , \1055 , \1056 );
nand \U$1002 ( \1058 , \1054 , \1057 );
not \U$1003 ( \1059 , \1058 );
not \U$1004 ( \1060 , \958 );
not \U$1005 ( \1061 , \1060 );
not \U$1006 ( \1062 , \988 );
not \U$1007 ( \1063 , \1062 );
or \U$1008 ( \1064 , \1061 , \1063 );
nand \U$1009 ( \1065 , \988 , \958 );
nand \U$1010 ( \1066 , \1064 , \1065 );
not \U$1011 ( \1067 , \1029 );
not \U$1012 ( \1068 , \1067 );
not \U$1013 ( \1069 , \1041 );
or \U$1014 ( \1070 , \1068 , \1069 );
not \U$1015 ( \1071 , \1033 );
nand \U$1016 ( \1072 , \1071 , \1036 );
nand \U$1017 ( \1073 , \1070 , \1072 );
nand \U$1018 ( \1074 , \1066 , \1073 );
not \U$1019 ( \1075 , \1074 );
or \U$1020 ( \1076 , \1059 , \1075 );
not \U$1021 ( \1077 , \1066 );
not \U$1022 ( \1078 , \1073 );
nand \U$1023 ( \1079 , \1077 , \1078 );
nand \U$1024 ( \1080 , \1076 , \1079 );
not \U$1025 ( \1081 , \1080 );
or \U$1026 ( \1082 , \995 , \1081 );
not \U$1027 ( \1083 , \957 );
not \U$1028 ( \1084 , \993 );
nand \U$1029 ( \1085 , \1083 , \1084 );
nand \U$1030 ( \1086 , \1082 , \1085 );
not \U$1031 ( \1087 , \732 );
and \U$1032 ( \1088 , \746 , \1087 );
not \U$1033 ( \1089 , \746 );
and \U$1034 ( \1090 , \1089 , \732 );
nor \U$1035 ( \1091 , \1088 , \1090 );
xor \U$1036 ( \1092 , \569 , \570 );
xor \U$1037 ( \1093 , \1092 , \572 );
not \U$1038 ( \1094 , \1093 );
not \U$1039 ( \1095 , \1094 );
nand \U$1040 ( \1096 , \588 , \582 );
and \U$1041 ( \1097 , \1096 , \584 );
not \U$1042 ( \1098 , \1096 );
not \U$1043 ( \1099 , \584 );
and \U$1044 ( \1100 , \1098 , \1099 );
nor \U$1045 ( \1101 , \1097 , \1100 );
not \U$1046 ( \1102 , \1101 );
not \U$1047 ( \1103 , \1102 );
or \U$1048 ( \1104 , \1095 , \1103 );
nand \U$1049 ( \1105 , \1101 , \1093 );
nand \U$1050 ( \1106 , \1104 , \1105 );
not \U$1051 ( \1107 , \910 );
not \U$1052 ( \1108 , \912 );
or \U$1053 ( \1109 , \1107 , \1108 );
nand \U$1054 ( \1110 , \1109 , \902 );
not \U$1055 ( \1111 , \1110 );
and \U$1056 ( \1112 , \1106 , \1111 );
not \U$1057 ( \1113 , \1106 );
and \U$1058 ( \1114 , \1113 , \1110 );
nor \U$1059 ( \1115 , \1112 , \1114 );
xor \U$1060 ( \1116 , \1091 , \1115 );
not \U$1061 ( \1117 , \948 );
not \U$1062 ( \1118 , \1117 );
not \U$1063 ( \1119 , \941 );
or \U$1064 ( \1120 , \1118 , \1119 );
not \U$1065 ( \1121 , \923 );
nand \U$1066 ( \1122 , \1121 , \937 );
nand \U$1067 ( \1123 , \1120 , \1122 );
xor \U$1068 ( \1124 , \1116 , \1123 );
not \U$1069 ( \1125 , \1124 );
not \U$1070 ( \1126 , \917 );
not \U$1071 ( \1127 , \953 );
or \U$1072 ( \1128 , \1126 , \1127 );
not \U$1073 ( \1129 , \900 );
nand \U$1074 ( \1130 , \1129 , \913 );
nand \U$1075 ( \1131 , \1128 , \1130 );
not \U$1076 ( \1132 , \1131 );
nand \U$1077 ( \1133 , \1125 , \1132 );
not \U$1078 ( \1134 , \1133 );
or \U$1079 ( \1135 , \1086 , \1134 );
and \U$1080 ( \1136 , \575 , \589 );
not \U$1081 ( \1137 , \575 );
and \U$1082 ( \1138 , \1137 , \590 );
nor \U$1083 ( \1139 , \1136 , \1138 );
not \U$1084 ( \1140 , \601 );
xnor \U$1085 ( \1141 , \1139 , \1140 );
not \U$1086 ( \1142 , \1141 );
not \U$1087 ( \1143 , \1094 );
not \U$1088 ( \1144 , \1101 );
or \U$1089 ( \1145 , \1143 , \1144 );
nand \U$1090 ( \1146 , \1145 , \1110 );
nand \U$1091 ( \1147 , \1102 , \1093 );
nand \U$1092 ( \1148 , \1146 , \1147 );
not \U$1093 ( \1149 , \1148 );
and \U$1094 ( \1150 , \1142 , \1149 );
and \U$1095 ( \1151 , \1141 , \1148 );
nor \U$1096 ( \1152 , \1150 , \1151 );
not \U$1097 ( \1153 , \1152 );
not \U$1098 ( \1154 , \751 );
not \U$1099 ( \1155 , \1154 );
not \U$1100 ( \1156 , \758 );
not \U$1101 ( \1157 , \761 );
or \U$1102 ( \1158 , \1156 , \1157 );
or \U$1103 ( \1159 , \761 , \758 );
nand \U$1104 ( \1160 , \1158 , \1159 );
not \U$1105 ( \1161 , \1160 );
or \U$1106 ( \1162 , \1155 , \1161 );
or \U$1107 ( \1163 , \1160 , \1154 );
nand \U$1108 ( \1164 , \1162 , \1163 );
not \U$1109 ( \1165 , \1164 );
and \U$1110 ( \1166 , \1153 , \1165 );
and \U$1111 ( \1167 , \1152 , \1164 );
nor \U$1112 ( \1168 , \1166 , \1167 );
xor \U$1113 ( \1169 , \1091 , \1115 );
and \U$1114 ( \1170 , \1169 , \1123 );
and \U$1115 ( \1171 , \1091 , \1115 );
or \U$1116 ( \1172 , \1170 , \1171 );
nand \U$1117 ( \1173 , \1168 , \1172 );
nand \U$1118 ( \1174 , \1124 , \1131 );
and \U$1119 ( \1175 , \1173 , \1174 );
nand \U$1120 ( \1176 , \1135 , \1175 );
xor \U$1121 ( \1177 , \716 , \764 );
xnor \U$1122 ( \1178 , \1177 , \773 );
not \U$1123 ( \1179 , \1164 );
not \U$1124 ( \1180 , \1152 );
not \U$1125 ( \1181 , \1180 );
or \U$1126 ( \1182 , \1179 , \1181 );
not \U$1127 ( \1183 , \1141 );
nand \U$1128 ( \1184 , \1183 , \1148 );
nand \U$1129 ( \1185 , \1182 , \1184 );
nand \U$1130 ( \1186 , \1178 , \1185 );
not \U$1131 ( \1187 , \1168 );
not \U$1132 ( \1188 , \1172 );
nand \U$1133 ( \1189 , \1187 , \1188 );
nand \U$1134 ( \1190 , \1186 , \1189 );
not \U$1135 ( \1191 , \1190 );
nand \U$1136 ( \1192 , \1176 , \1191 );
nand \U$1137 ( \1193 , \835 , \838 );
not \U$1138 ( \1194 , \1193 );
not \U$1139 ( \1195 , \1178 );
not \U$1140 ( \1196 , \1185 );
nand \U$1141 ( \1197 , \1195 , \1196 );
nand \U$1142 ( \1198 , \709 , \777 );
nand \U$1143 ( \1199 , \1197 , \1198 );
nor \U$1144 ( \1200 , \1194 , \1199 );
nand \U$1145 ( \1201 , \1192 , \1200 );
not \U$1146 ( \1202 , \1201 );
not \U$1147 ( \1203 , \876 );
nand \U$1148 ( \1204 , \1202 , \1203 );
nand \U$1149 ( \1205 , \884 , \1204 );
not \U$1150 ( \1206 , \1205 );
or \U$1151 ( \1207 , \507 , \1206 );
not \U$1152 ( \1208 , \495 );
nor \U$1153 ( \1209 , \1208 , \337 );
not \U$1154 ( \1210 , \1209 );
not \U$1155 ( \1211 , \336 );
not \U$1156 ( \1212 , \288 );
or \U$1157 ( \1213 , \1211 , \1212 );
nand \U$1158 ( \1214 , \461 , \468 );
nand \U$1159 ( \1215 , \1213 , \1214 );
not \U$1160 ( \1216 , \1215 );
or \U$1161 ( \1217 , \1210 , \1216 );
or \U$1162 ( \1218 , \478 , \494 );
nand \U$1163 ( \1219 , \1217 , \1218 );
and \U$1164 ( \1220 , \1219 , \504 );
nor \U$1165 ( \1221 , \498 , \503 );
nor \U$1166 ( \1222 , \1220 , \1221 );
nand \U$1167 ( \1223 , \1207 , \1222 );
not \U$1168 ( \1224 , \1223 );
or \U$1169 ( \1225 , \107 , \1224 );
nand \U$1170 ( \1226 , \104 , \105 );
nand \U$1171 ( \1227 , \1225 , \1226 );
buf \U$1172 ( \1228 , \1227 );
nand \U$1173 ( \1229 , \1226 , \106 );
not \U$1174 ( \1230 , \1229 );
not \U$1175 ( \1231 , \1223 );
or \U$1176 ( \1232 , \1230 , \1231 );
or \U$1177 ( \1233 , \1223 , \1229 );
nand \U$1178 ( \1234 , \1232 , \1233 );
buf \U$1179 ( \1235 , \1234 );
not \U$1180 ( \1236 , \495 );
nor \U$1181 ( \1237 , \471 , \876 );
not \U$1182 ( \1238 , \1237 );
nand \U$1183 ( \1239 , \840 , \1201 );
not \U$1184 ( \1240 , \1239 );
or \U$1185 ( \1241 , \1238 , \1240 );
and \U$1186 ( \1242 , \880 , \881 );
nor \U$1187 ( \1243 , \1242 , \1215 );
not \U$1188 ( \1244 , \1243 );
not \U$1189 ( \1245 , \879 );
or \U$1190 ( \1246 , \1244 , \1245 );
not \U$1191 ( \1247 , \1215 );
not \U$1192 ( \1248 , \470 );
and \U$1193 ( \1249 , \1247 , \1248 );
nor \U$1194 ( \1250 , \1249 , \337 );
nand \U$1195 ( \1251 , \1246 , \1250 );
nand \U$1196 ( \1252 , \1241 , \1251 );
not \U$1197 ( \1253 , \1252 );
or \U$1198 ( \1254 , \1236 , \1253 );
nand \U$1199 ( \1255 , \1254 , \1218 );
not \U$1200 ( \1256 , \1221 );
nand \U$1201 ( \1257 , \1256 , \504 );
not \U$1202 ( \1258 , \1257 );
and \U$1203 ( \1259 , \1255 , \1258 );
not \U$1204 ( \1260 , \1255 );
and \U$1205 ( \1261 , \1260 , \1257 );
nor \U$1206 ( \1262 , \1259 , \1261 );
buf \U$1207 ( \1263 , \1262 );
nand \U$1208 ( \1264 , \1218 , \495 );
not \U$1209 ( \1265 , \1264 );
and \U$1210 ( \1266 , \1252 , \1265 );
not \U$1211 ( \1267 , \1252 );
and \U$1212 ( \1268 , \1267 , \1264 );
nor \U$1213 ( \1269 , \1266 , \1268 );
buf \U$1214 ( \1270 , \1269 );
buf \U$1215 ( \1271 , \470 );
not \U$1216 ( \1272 , \1271 );
not \U$1217 ( \1273 , \1205 );
or \U$1218 ( \1274 , \1272 , \1273 );
nand \U$1219 ( \1275 , \1274 , \1214 );
and \U$1220 ( \1276 , \336 , \288 );
not \U$1221 ( \1277 , \336 );
not \U$1222 ( \1278 , \288 );
and \U$1223 ( \1279 , \1277 , \1278 );
nor \U$1224 ( \1280 , \1276 , \1279 );
and \U$1225 ( \1281 , \1275 , \1280 );
not \U$1226 ( \1282 , \1275 );
not \U$1227 ( \1283 , \1280 );
and \U$1228 ( \1284 , \1282 , \1283 );
nor \U$1229 ( \1285 , \1281 , \1284 );
buf \U$1230 ( \1286 , \1285 );
nand \U$1231 ( \1287 , \1271 , \1214 );
xnor \U$1232 ( \1288 , \1287 , \1205 );
buf \U$1233 ( \1289 , \1288 );
buf \U$1234 ( \1290 , \868 );
not \U$1235 ( \1291 , \1290 );
not \U$1236 ( \1292 , \1239 );
or \U$1237 ( \1293 , \1291 , \1292 );
buf \U$1238 ( \1294 , \878 );
not \U$1239 ( \1295 , \1294 );
nand \U$1240 ( \1296 , \1293 , \1295 );
nand \U$1241 ( \1297 , \875 , \882 );
not \U$1242 ( \1298 , \1297 );
and \U$1243 ( \1299 , \1296 , \1298 );
not \U$1244 ( \1300 , \1296 );
and \U$1245 ( \1301 , \1300 , \1297 );
nor \U$1246 ( \1302 , \1299 , \1301 );
buf \U$1247 ( \1303 , \1302 );
not \U$1248 ( \1304 , \1294 );
nand \U$1249 ( \1305 , \1304 , \1290 );
not \U$1250 ( \1306 , \1305 );
and \U$1251 ( \1307 , \1239 , \1306 );
not \U$1252 ( \1308 , \1239 );
and \U$1253 ( \1309 , \1308 , \1305 );
nor \U$1254 ( \1310 , \1307 , \1309 );
buf \U$1255 ( \1311 , \1310 );
not \U$1256 ( \1312 , \1176 );
not \U$1257 ( \1313 , \1191 );
or \U$1258 ( \1314 , \1312 , \1313 );
nand \U$1259 ( \1315 , \1196 , \1195 );
nand \U$1260 ( \1316 , \1314 , \1315 );
not \U$1261 ( \1317 , \1316 );
buf \U$1262 ( \1318 , \1198 );
not \U$1263 ( \1319 , \1318 );
not \U$1264 ( \1320 , \1319 );
and \U$1265 ( \1321 , \1317 , \1320 );
buf \U$1266 ( \1322 , \779 );
not \U$1267 ( \1323 , \1322 );
nor \U$1268 ( \1324 , \1321 , \1323 );
nand \U$1269 ( \1325 , \839 , \831 );
and \U$1270 ( \1326 , \1324 , \1325 );
not \U$1271 ( \1327 , \1324 );
not \U$1272 ( \1328 , \1325 );
and \U$1273 ( \1329 , \1327 , \1328 );
nor \U$1274 ( \1330 , \1326 , \1329 );
buf \U$1275 ( \1331 , \1330 );
nand \U$1276 ( \1332 , \1322 , \1318 );
and \U$1277 ( \1333 , \1316 , \1332 );
not \U$1278 ( \1334 , \1316 );
not \U$1279 ( \1335 , \1332 );
and \U$1280 ( \1336 , \1334 , \1335 );
nor \U$1281 ( \1337 , \1333 , \1336 );
buf \U$1282 ( \1338 , \1337 );
buf \U$1283 ( \1339 , \1176 );
nand \U$1284 ( \1340 , \1339 , \1189 );
nand \U$1285 ( \1341 , \1315 , \1186 );
not \U$1286 ( \1342 , \1341 );
and \U$1287 ( \1343 , \1340 , \1342 );
not \U$1288 ( \1344 , \1340 );
and \U$1289 ( \1345 , \1344 , \1341 );
nor \U$1290 ( \1346 , \1343 , \1345 );
buf \U$1291 ( \1347 , \1346 );
and \U$1292 ( \1348 , \1086 , \1174 );
nor \U$1293 ( \1349 , \1348 , \1134 );
nand \U$1294 ( \1350 , \1173 , \1189 );
and \U$1295 ( \1351 , \1349 , \1350 );
not \U$1296 ( \1352 , \1349 );
not \U$1297 ( \1353 , \1350 );
and \U$1298 ( \1354 , \1352 , \1353 );
nor \U$1299 ( \1355 , \1351 , \1354 );
buf \U$1300 ( \1356 , \1355 );
endmodule

